module tt_um_algofoogle_raybox_zero (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire net2202;
 wire net844;
 wire \hpos[0] ;
 wire \hpos[1] ;
 wire \hpos[2] ;
 wire \hpos[3] ;
 wire \hpos[4] ;
 wire \hpos[5] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync_n;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.h[0] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.debug_overlay.vpos[0] ;
 wire \rbzero.debug_overlay.vpos[1] ;
 wire \rbzero.debug_overlay.vpos[2] ;
 wire \rbzero.debug_overlay.vpos[3] ;
 wire \rbzero.debug_overlay.vpos[4] ;
 wire \rbzero.debug_overlay.vpos[5] ;
 wire \rbzero.debug_overlay.vpos[6] ;
 wire \rbzero.debug_overlay.vpos[7] ;
 wire \rbzero.debug_overlay.vpos[8] ;
 wire \rbzero.debug_overlay.vpos[9] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.i_col[0] ;
 wire \rbzero.map_rom.i_col[1] ;
 wire \rbzero.map_rom.i_col[2] ;
 wire \rbzero.map_rom.i_col[3] ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[0] ;
 wire \rbzero.map_rom.i_row[1] ;
 wire \rbzero.map_rom.i_row[2] ;
 wire \rbzero.map_rom.i_row[3] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.o_tex_csb ;
 wire \rbzero.o_tex_out0 ;
 wire clknet_leaf_0_clk;
 wire \rbzero.o_vinf ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.rgb[0] ;
 wire \rbzero.rgb[1] ;
 wire \rbzero.rgb[2] ;
 wire \rbzero.rgb[3] ;
 wire \rbzero.rgb[4] ;
 wire \rbzero.rgb[5] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.buf_floor[0] ;
 wire \rbzero.spi_registers.buf_floor[1] ;
 wire \rbzero.spi_registers.buf_floor[2] ;
 wire \rbzero.spi_registers.buf_floor[3] ;
 wire \rbzero.spi_registers.buf_floor[4] ;
 wire \rbzero.spi_registers.buf_floor[5] ;
 wire \rbzero.spi_registers.buf_leak[0] ;
 wire \rbzero.spi_registers.buf_leak[1] ;
 wire \rbzero.spi_registers.buf_leak[2] ;
 wire \rbzero.spi_registers.buf_leak[3] ;
 wire \rbzero.spi_registers.buf_leak[4] ;
 wire \rbzero.spi_registers.buf_leak[5] ;
 wire \rbzero.spi_registers.buf_mapdx[0] ;
 wire \rbzero.spi_registers.buf_mapdx[1] ;
 wire \rbzero.spi_registers.buf_mapdx[2] ;
 wire \rbzero.spi_registers.buf_mapdx[3] ;
 wire \rbzero.spi_registers.buf_mapdx[4] ;
 wire \rbzero.spi_registers.buf_mapdxw[0] ;
 wire \rbzero.spi_registers.buf_mapdxw[1] ;
 wire \rbzero.spi_registers.buf_mapdy[0] ;
 wire \rbzero.spi_registers.buf_mapdy[1] ;
 wire \rbzero.spi_registers.buf_mapdy[2] ;
 wire \rbzero.spi_registers.buf_mapdy[3] ;
 wire \rbzero.spi_registers.buf_mapdy[4] ;
 wire \rbzero.spi_registers.buf_mapdyw[0] ;
 wire \rbzero.spi_registers.buf_mapdyw[1] ;
 wire \rbzero.spi_registers.buf_otherx[0] ;
 wire \rbzero.spi_registers.buf_otherx[1] ;
 wire \rbzero.spi_registers.buf_otherx[2] ;
 wire \rbzero.spi_registers.buf_otherx[3] ;
 wire \rbzero.spi_registers.buf_otherx[4] ;
 wire \rbzero.spi_registers.buf_othery[0] ;
 wire \rbzero.spi_registers.buf_othery[1] ;
 wire \rbzero.spi_registers.buf_othery[2] ;
 wire \rbzero.spi_registers.buf_othery[3] ;
 wire \rbzero.spi_registers.buf_othery[4] ;
 wire \rbzero.spi_registers.buf_sky[0] ;
 wire \rbzero.spi_registers.buf_sky[1] ;
 wire \rbzero.spi_registers.buf_sky[2] ;
 wire \rbzero.spi_registers.buf_sky[3] ;
 wire \rbzero.spi_registers.buf_sky[4] ;
 wire \rbzero.spi_registers.buf_sky[5] ;
 wire \rbzero.spi_registers.buf_texadd0[0] ;
 wire \rbzero.spi_registers.buf_texadd0[10] ;
 wire \rbzero.spi_registers.buf_texadd0[11] ;
 wire \rbzero.spi_registers.buf_texadd0[12] ;
 wire \rbzero.spi_registers.buf_texadd0[13] ;
 wire \rbzero.spi_registers.buf_texadd0[14] ;
 wire \rbzero.spi_registers.buf_texadd0[15] ;
 wire \rbzero.spi_registers.buf_texadd0[16] ;
 wire \rbzero.spi_registers.buf_texadd0[17] ;
 wire \rbzero.spi_registers.buf_texadd0[18] ;
 wire \rbzero.spi_registers.buf_texadd0[19] ;
 wire \rbzero.spi_registers.buf_texadd0[1] ;
 wire \rbzero.spi_registers.buf_texadd0[20] ;
 wire \rbzero.spi_registers.buf_texadd0[21] ;
 wire \rbzero.spi_registers.buf_texadd0[22] ;
 wire \rbzero.spi_registers.buf_texadd0[23] ;
 wire \rbzero.spi_registers.buf_texadd0[2] ;
 wire \rbzero.spi_registers.buf_texadd0[3] ;
 wire \rbzero.spi_registers.buf_texadd0[4] ;
 wire \rbzero.spi_registers.buf_texadd0[5] ;
 wire \rbzero.spi_registers.buf_texadd0[6] ;
 wire \rbzero.spi_registers.buf_texadd0[7] ;
 wire \rbzero.spi_registers.buf_texadd0[8] ;
 wire \rbzero.spi_registers.buf_texadd0[9] ;
 wire \rbzero.spi_registers.buf_texadd1[0] ;
 wire \rbzero.spi_registers.buf_texadd1[10] ;
 wire \rbzero.spi_registers.buf_texadd1[11] ;
 wire \rbzero.spi_registers.buf_texadd1[12] ;
 wire \rbzero.spi_registers.buf_texadd1[13] ;
 wire \rbzero.spi_registers.buf_texadd1[14] ;
 wire \rbzero.spi_registers.buf_texadd1[15] ;
 wire \rbzero.spi_registers.buf_texadd1[16] ;
 wire \rbzero.spi_registers.buf_texadd1[17] ;
 wire \rbzero.spi_registers.buf_texadd1[18] ;
 wire \rbzero.spi_registers.buf_texadd1[19] ;
 wire \rbzero.spi_registers.buf_texadd1[1] ;
 wire \rbzero.spi_registers.buf_texadd1[20] ;
 wire \rbzero.spi_registers.buf_texadd1[21] ;
 wire \rbzero.spi_registers.buf_texadd1[22] ;
 wire \rbzero.spi_registers.buf_texadd1[23] ;
 wire \rbzero.spi_registers.buf_texadd1[2] ;
 wire \rbzero.spi_registers.buf_texadd1[3] ;
 wire \rbzero.spi_registers.buf_texadd1[4] ;
 wire \rbzero.spi_registers.buf_texadd1[5] ;
 wire \rbzero.spi_registers.buf_texadd1[6] ;
 wire \rbzero.spi_registers.buf_texadd1[7] ;
 wire \rbzero.spi_registers.buf_texadd1[8] ;
 wire \rbzero.spi_registers.buf_texadd1[9] ;
 wire \rbzero.spi_registers.buf_texadd2[0] ;
 wire \rbzero.spi_registers.buf_texadd2[10] ;
 wire \rbzero.spi_registers.buf_texadd2[11] ;
 wire \rbzero.spi_registers.buf_texadd2[12] ;
 wire \rbzero.spi_registers.buf_texadd2[13] ;
 wire \rbzero.spi_registers.buf_texadd2[14] ;
 wire \rbzero.spi_registers.buf_texadd2[15] ;
 wire \rbzero.spi_registers.buf_texadd2[16] ;
 wire \rbzero.spi_registers.buf_texadd2[17] ;
 wire \rbzero.spi_registers.buf_texadd2[18] ;
 wire \rbzero.spi_registers.buf_texadd2[19] ;
 wire \rbzero.spi_registers.buf_texadd2[1] ;
 wire \rbzero.spi_registers.buf_texadd2[20] ;
 wire \rbzero.spi_registers.buf_texadd2[21] ;
 wire \rbzero.spi_registers.buf_texadd2[22] ;
 wire \rbzero.spi_registers.buf_texadd2[23] ;
 wire \rbzero.spi_registers.buf_texadd2[2] ;
 wire \rbzero.spi_registers.buf_texadd2[3] ;
 wire \rbzero.spi_registers.buf_texadd2[4] ;
 wire \rbzero.spi_registers.buf_texadd2[5] ;
 wire \rbzero.spi_registers.buf_texadd2[6] ;
 wire \rbzero.spi_registers.buf_texadd2[7] ;
 wire \rbzero.spi_registers.buf_texadd2[8] ;
 wire \rbzero.spi_registers.buf_texadd2[9] ;
 wire \rbzero.spi_registers.buf_texadd3[0] ;
 wire \rbzero.spi_registers.buf_texadd3[10] ;
 wire \rbzero.spi_registers.buf_texadd3[11] ;
 wire \rbzero.spi_registers.buf_texadd3[12] ;
 wire \rbzero.spi_registers.buf_texadd3[13] ;
 wire \rbzero.spi_registers.buf_texadd3[14] ;
 wire \rbzero.spi_registers.buf_texadd3[15] ;
 wire \rbzero.spi_registers.buf_texadd3[16] ;
 wire \rbzero.spi_registers.buf_texadd3[17] ;
 wire \rbzero.spi_registers.buf_texadd3[18] ;
 wire \rbzero.spi_registers.buf_texadd3[19] ;
 wire \rbzero.spi_registers.buf_texadd3[1] ;
 wire \rbzero.spi_registers.buf_texadd3[20] ;
 wire \rbzero.spi_registers.buf_texadd3[21] ;
 wire \rbzero.spi_registers.buf_texadd3[22] ;
 wire \rbzero.spi_registers.buf_texadd3[23] ;
 wire \rbzero.spi_registers.buf_texadd3[2] ;
 wire \rbzero.spi_registers.buf_texadd3[3] ;
 wire \rbzero.spi_registers.buf_texadd3[4] ;
 wire \rbzero.spi_registers.buf_texadd3[5] ;
 wire \rbzero.spi_registers.buf_texadd3[6] ;
 wire \rbzero.spi_registers.buf_texadd3[7] ;
 wire \rbzero.spi_registers.buf_texadd3[8] ;
 wire \rbzero.spi_registers.buf_texadd3[9] ;
 wire \rbzero.spi_registers.buf_vinf ;
 wire \rbzero.spi_registers.buf_vshift[0] ;
 wire \rbzero.spi_registers.buf_vshift[1] ;
 wire \rbzero.spi_registers.buf_vshift[2] ;
 wire \rbzero.spi_registers.buf_vshift[3] ;
 wire \rbzero.spi_registers.buf_vshift[4] ;
 wire \rbzero.spi_registers.buf_vshift[5] ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.vsync_n ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_done ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-10] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-11] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-1] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-2] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-3] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-4] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-5] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-6] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-7] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-8] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[-9] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[0] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[10] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[1] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[2] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[3] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[4] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[5] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[6] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[7] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[8] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_data[9] ;
 wire \rbzero.wall_tracer.rcp_fsm.i_start ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-10] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-11] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-1] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-2] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-3] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-4] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-5] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-6] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-7] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-8] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[-9] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[0] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[10] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[1] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[2] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[3] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[4] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[5] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[6] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[7] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[8] ;
 wire \rbzero.wall_tracer.rcp_fsm.o_data[9] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-10] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-11] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-1] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-2] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-3] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-4] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-5] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-6] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-7] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-8] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[-9] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[0] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[10] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[1] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[2] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[3] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[4] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[5] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[6] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[7] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[8] ;
 wire \rbzero.wall_tracer.rcp_fsm.operand[9] ;
 wire \rbzero.wall_tracer.rcp_fsm.state[0] ;
 wire \rbzero.wall_tracer.rcp_fsm.state[1] ;
 wire \rbzero.wall_tracer.rcp_fsm.state[2] ;
 wire \rbzero.wall_tracer.rcp_fsm.state[3] ;
 wire \rbzero.wall_tracer.rcp_fsm.state[4] ;
 wire \rbzero.wall_tracer.side ;
 wire \rbzero.wall_tracer.size[0] ;
 wire \rbzero.wall_tracer.size[10] ;
 wire \rbzero.wall_tracer.size[1] ;
 wire \rbzero.wall_tracer.size[2] ;
 wire \rbzero.wall_tracer.size[3] ;
 wire \rbzero.wall_tracer.size[4] ;
 wire \rbzero.wall_tracer.size[5] ;
 wire \rbzero.wall_tracer.size[6] ;
 wire \rbzero.wall_tracer.size[7] ;
 wire \rbzero.wall_tracer.size[8] ;
 wire \rbzero.wall_tracer.size[9] ;
 wire \rbzero.wall_tracer.size_full[-10] ;
 wire \rbzero.wall_tracer.size_full[-11] ;
 wire \rbzero.wall_tracer.size_full[-9] ;
 wire \rbzero.wall_tracer.size_full[10] ;
 wire \rbzero.wall_tracer.size_full[3] ;
 wire \rbzero.wall_tracer.size_full[4] ;
 wire \rbzero.wall_tracer.size_full[5] ;
 wire \rbzero.wall_tracer.size_full[6] ;
 wire \rbzero.wall_tracer.size_full[7] ;
 wire \rbzero.wall_tracer.size_full[8] ;
 wire \rbzero.wall_tracer.size_full[9] ;
 wire \rbzero.wall_tracer.state[0] ;
 wire \rbzero.wall_tracer.state[1] ;
 wire \rbzero.wall_tracer.state[2] ;
 wire \rbzero.wall_tracer.state[3] ;
 wire \rbzero.wall_tracer.state[4] ;
 wire \rbzero.wall_tracer.state[5] ;
 wire \rbzero.wall_tracer.state[6] ;
 wire \rbzero.wall_tracer.state[7] ;
 wire \rbzero.wall_tracer.state[8] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.texu[0] ;
 wire \rbzero.wall_tracer.texu[1] ;
 wire \rbzero.wall_tracer.texu[2] ;
 wire \rbzero.wall_tracer.texu[3] ;
 wire \rbzero.wall_tracer.texu[4] ;
 wire \rbzero.wall_tracer.texu[5] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \rbzero.wall_tracer.w[0] ;
 wire \rbzero.wall_tracer.w[1] ;
 wire \rbzero.wall_tracer.w[2] ;
 wire \rbzero.wall_tracer.wall[0] ;
 wire \rbzero.wall_tracer.wall[1] ;
 wire \registered_vga_output[0] ;
 wire \registered_vga_output[1] ;
 wire \registered_vga_output[2] ;
 wire \registered_vga_output[3] ;
 wire \registered_vga_output[4] ;
 wire \registered_vga_output[5] ;
 wire \registered_vga_output[6] ;
 wire \registered_vga_output[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_2 _14998_ (.A(rst_n),
    .X(_08409_));
 sg13g2_nand2b_1 _14999_ (.Y(_08410_),
    .B(_08409_),
    .A_N(\rbzero.vga_sync.vsync ));
 sg13g2_buf_1 _15000_ (.A(_08410_),
    .X(_08411_));
 sg13g2_buf_1 _15001_ (.A(_08411_),
    .X(_08412_));
 sg13g2_buf_1 _15002_ (.A(net729),
    .X(_08413_));
 sg13g2_buf_1 _15003_ (.A(\rbzero.wall_tracer.state[5] ),
    .X(_08414_));
 sg13g2_buf_1 _15004_ (.A(\rbzero.wall_tracer.w[0] ),
    .X(_08415_));
 sg13g2_nor2_1 _15005_ (.A(\rbzero.wall_tracer.w[1] ),
    .B(_08415_),
    .Y(_08416_));
 sg13g2_nand2_1 _15006_ (.Y(_08417_),
    .A(_00015_),
    .B(_08416_));
 sg13g2_buf_1 _15007_ (.A(\rbzero.wall_tracer.state[2] ),
    .X(_08418_));
 sg13g2_buf_1 _15008_ (.A(_08418_),
    .X(_08419_));
 sg13g2_buf_1 _15009_ (.A(net800),
    .X(_08420_));
 sg13g2_buf_1 _15010_ (.A(net728),
    .X(_08421_));
 sg13g2_buf_1 _15011_ (.A(_00016_),
    .X(_08422_));
 sg13g2_buf_1 _15012_ (.A(\rbzero.wall_tracer.rcp_done ),
    .X(_08423_));
 sg13g2_and2_1 _15013_ (.A(_08422_),
    .B(_08423_),
    .X(_08424_));
 sg13g2_buf_1 _15014_ (.A(_08424_),
    .X(_08425_));
 sg13g2_and2_1 _15015_ (.A(net685),
    .B(_08425_),
    .X(_08426_));
 sg13g2_buf_1 _15016_ (.A(_08426_),
    .X(_08427_));
 sg13g2_buf_1 _15017_ (.A(_08427_),
    .X(_08428_));
 sg13g2_buf_1 _15018_ (.A(net512),
    .X(_08429_));
 sg13g2_a21oi_1 _15019_ (.A1(_08414_),
    .A2(_08417_),
    .Y(_08430_),
    .B1(net492));
 sg13g2_nor2_1 _15020_ (.A(net686),
    .B(_08430_),
    .Y(_00010_));
 sg13g2_buf_1 _15021_ (.A(\rbzero.wall_tracer.state[6] ),
    .X(_08431_));
 sg13g2_buf_1 _15022_ (.A(_08431_),
    .X(_08432_));
 sg13g2_buf_1 _15023_ (.A(net799),
    .X(_08433_));
 sg13g2_inv_1 _15024_ (.Y(_08434_),
    .A(_08423_));
 sg13g2_buf_1 _15025_ (.A(\rbzero.wall_tracer.rcp_fsm.i_start ),
    .X(_08435_));
 sg13g2_a21o_1 _15026_ (.A2(_08434_),
    .A1(_08422_),
    .B1(net832),
    .X(_08436_));
 sg13g2_buf_1 _15027_ (.A(_08436_),
    .X(_08437_));
 sg13g2_a21oi_1 _15028_ (.A1(_08433_),
    .A2(_08437_),
    .Y(_08438_),
    .B1(\rbzero.wall_tracer.state[0] ));
 sg13g2_nor2_1 _15029_ (.A(net686),
    .B(_08438_),
    .Y(_00011_));
 sg13g2_buf_1 _15030_ (.A(\rbzero.wall_tracer.state[7] ),
    .X(_08439_));
 sg13g2_buf_1 _15031_ (.A(_08439_),
    .X(_08440_));
 sg13g2_buf_1 _15032_ (.A(net798),
    .X(_08441_));
 sg13g2_buf_1 _15033_ (.A(_08441_),
    .X(_08442_));
 sg13g2_buf_1 _15034_ (.A(\rbzero.wall_tracer.state[3] ),
    .X(_08443_));
 sg13g2_buf_1 _15035_ (.A(_08443_),
    .X(_08444_));
 sg13g2_buf_1 _15036_ (.A(net797),
    .X(_08445_));
 sg13g2_buf_1 _15037_ (.A(net725),
    .X(_08446_));
 sg13g2_buf_1 _15038_ (.A(net683),
    .X(_08447_));
 sg13g2_and2_1 _15039_ (.A(net611),
    .B(_08425_),
    .X(_08448_));
 sg13g2_buf_1 _15040_ (.A(_08448_),
    .X(_08449_));
 sg13g2_buf_1 _15041_ (.A(_08449_),
    .X(_08450_));
 sg13g2_a21oi_1 _15042_ (.A1(net684),
    .A2(_08417_),
    .Y(_08451_),
    .B1(net491));
 sg13g2_nor2_1 _15043_ (.A(net686),
    .B(_08451_),
    .Y(_00012_));
 sg13g2_buf_1 _15044_ (.A(\hpos[8] ),
    .X(_08452_));
 sg13g2_buf_1 _15045_ (.A(\hpos[4] ),
    .X(_08453_));
 sg13g2_buf_1 _15046_ (.A(_08453_),
    .X(_08454_));
 sg13g2_buf_1 _15047_ (.A(\hpos[3] ),
    .X(_08455_));
 sg13g2_inv_1 _15048_ (.Y(_08456_),
    .A(net830));
 sg13g2_buf_1 _15049_ (.A(\hpos[2] ),
    .X(_08457_));
 sg13g2_buf_1 _15050_ (.A(\hpos[1] ),
    .X(_08458_));
 sg13g2_buf_1 _15051_ (.A(\hpos[0] ),
    .X(_08459_));
 sg13g2_nand3_1 _15052_ (.B(_08458_),
    .C(net828),
    .A(net829),
    .Y(_08460_));
 sg13g2_buf_1 _15053_ (.A(_08460_),
    .X(_08461_));
 sg13g2_nor2_1 _15054_ (.A(_08456_),
    .B(_08461_),
    .Y(_08462_));
 sg13g2_and2_1 _15055_ (.A(net796),
    .B(_08462_),
    .X(_08463_));
 sg13g2_buf_1 _15056_ (.A(_08463_),
    .X(_08464_));
 sg13g2_buf_2 _15057_ (.A(\hpos[6] ),
    .X(_08465_));
 sg13g2_buf_2 _15058_ (.A(\hpos[7] ),
    .X(_08466_));
 sg13g2_nor2_1 _15059_ (.A(_08465_),
    .B(_08466_),
    .Y(_08467_));
 sg13g2_buf_2 _15060_ (.A(\hpos[5] ),
    .X(_08468_));
 sg13g2_buf_1 _15061_ (.A(\hpos[9] ),
    .X(_08469_));
 sg13g2_inv_2 _15062_ (.Y(_08470_),
    .A(_08469_));
 sg13g2_nor2_1 _15063_ (.A(_08468_),
    .B(_08470_),
    .Y(_08471_));
 sg13g2_nand4_1 _15064_ (.B(_08464_),
    .C(_08467_),
    .A(net831),
    .Y(_08472_),
    .D(_08471_));
 sg13g2_buf_2 _15065_ (.A(_08472_),
    .X(_08473_));
 sg13g2_and2_1 _15066_ (.A(_00015_),
    .B(_08416_),
    .X(_08474_));
 sg13g2_buf_1 _15067_ (.A(_08474_),
    .X(_08475_));
 sg13g2_and2_1 _15068_ (.A(_08414_),
    .B(_08475_),
    .X(_08476_));
 sg13g2_buf_1 _15069_ (.A(_08476_),
    .X(_08477_));
 sg13g2_a21oi_1 _15070_ (.A1(\rbzero.wall_tracer.state[8] ),
    .A2(_08473_),
    .Y(_08478_),
    .B1(_08477_));
 sg13g2_nor2_1 _15071_ (.A(net686),
    .B(_08478_),
    .Y(_00013_));
 sg13g2_buf_1 _15072_ (.A(\rbzero.wall_tracer.state[1] ),
    .X(_08479_));
 sg13g2_buf_1 _15073_ (.A(_08479_),
    .X(_08480_));
 sg13g2_buf_2 _15074_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_08481_));
 sg13g2_buf_2 _15075_ (.A(\rbzero.map_rom.i_col[3] ),
    .X(_08482_));
 sg13g2_buf_2 _15076_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .X(_08483_));
 sg13g2_xnor2_1 _15077_ (.Y(_08484_),
    .A(_08482_),
    .B(_08483_));
 sg13g2_buf_1 _15078_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .X(_08485_));
 sg13g2_buf_2 _15079_ (.A(\rbzero.map_rom.i_row[0] ),
    .X(_08486_));
 sg13g2_xnor2_1 _15080_ (.Y(_08487_),
    .A(_08485_),
    .B(_08486_));
 sg13g2_buf_2 _15081_ (.A(\rbzero.map_rom.i_row[3] ),
    .X(_08488_));
 sg13g2_buf_2 _15082_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .X(_08489_));
 sg13g2_xnor2_1 _15083_ (.Y(_08490_),
    .A(_08488_),
    .B(_08489_));
 sg13g2_buf_2 _15084_ (.A(\rbzero.map_rom.i_row[4] ),
    .X(_08491_));
 sg13g2_buf_2 _15085_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .X(_08492_));
 sg13g2_xor2_1 _15086_ (.B(_08492_),
    .A(_08491_),
    .X(_08493_));
 sg13g2_buf_2 _15087_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .X(_08494_));
 sg13g2_buf_1 _15088_ (.A(\rbzero.map_rom.i_col[0] ),
    .X(_08495_));
 sg13g2_xor2_1 _15089_ (.B(net827),
    .A(_08494_),
    .X(_08496_));
 sg13g2_buf_1 _15090_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .X(_08497_));
 sg13g2_buf_1 _15091_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .X(_08498_));
 sg13g2_xor2_1 _15092_ (.B(_08498_),
    .A(_08497_),
    .X(_08499_));
 sg13g2_buf_1 _15093_ (.A(\rbzero.map_rom.i_col[2] ),
    .X(_08500_));
 sg13g2_buf_1 _15094_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .X(_08501_));
 sg13g2_xor2_1 _15095_ (.B(_08501_),
    .A(_08500_),
    .X(_08502_));
 sg13g2_nor4_1 _15096_ (.A(_08493_),
    .B(_08496_),
    .C(_08499_),
    .D(_08502_),
    .Y(_08503_));
 sg13g2_nand4_1 _15097_ (.B(_08487_),
    .C(_08490_),
    .A(_08484_),
    .Y(_08504_),
    .D(_08503_));
 sg13g2_buf_2 _15098_ (.A(\rbzero.map_rom.i_row[1] ),
    .X(_08505_));
 sg13g2_buf_1 _15099_ (.A(_08505_),
    .X(_08506_));
 sg13g2_buf_1 _15100_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .X(_08507_));
 sg13g2_xnor2_1 _15101_ (.Y(_08508_),
    .A(net794),
    .B(_08507_));
 sg13g2_buf_1 _15102_ (.A(\rbzero.map_rom.i_col[1] ),
    .X(_08509_));
 sg13g2_buf_1 _15103_ (.A(_08509_),
    .X(_08510_));
 sg13g2_buf_2 _15104_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .X(_08511_));
 sg13g2_xnor2_1 _15105_ (.Y(_08512_),
    .A(net793),
    .B(_08511_));
 sg13g2_buf_2 _15106_ (.A(\rbzero.map_rom.i_col[4] ),
    .X(_08513_));
 sg13g2_buf_1 _15107_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .X(_08514_));
 sg13g2_xnor2_1 _15108_ (.Y(_08515_),
    .A(_08513_),
    .B(_08514_));
 sg13g2_buf_1 _15109_ (.A(\rbzero.map_rom.i_row[2] ),
    .X(_08516_));
 sg13g2_buf_1 _15110_ (.A(_08516_),
    .X(_08517_));
 sg13g2_buf_1 _15111_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .X(_08518_));
 sg13g2_xnor2_1 _15112_ (.Y(_08519_),
    .A(net792),
    .B(_08518_));
 sg13g2_nand4_1 _15113_ (.B(_08512_),
    .C(_08515_),
    .A(_08508_),
    .Y(_08520_),
    .D(_08519_));
 sg13g2_buf_2 _15114_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .X(_08521_));
 sg13g2_buf_1 _15115_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .X(_08522_));
 sg13g2_xnor2_1 _15116_ (.Y(_08523_),
    .A(_08521_),
    .B(_08522_));
 sg13g2_buf_1 _15117_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .X(_08524_));
 sg13g2_buf_1 _15118_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .X(_08525_));
 sg13g2_buf_1 _15119_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .X(_08526_));
 sg13g2_nor4_1 _15120_ (.A(_08524_),
    .B(\rbzero.wall_tracer.mapY[6] ),
    .C(_08525_),
    .D(_08526_),
    .Y(_08527_));
 sg13g2_nor2_1 _15121_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(\rbzero.wall_tracer.mapY[10] ),
    .Y(_08528_));
 sg13g2_nor4_1 _15122_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(\rbzero.wall_tracer.mapX[6] ),
    .C(\rbzero.wall_tracer.mapX[9] ),
    .D(\rbzero.wall_tracer.mapX[8] ),
    .Y(_08529_));
 sg13g2_nand4_1 _15123_ (.B(_08527_),
    .C(_08528_),
    .A(_08523_),
    .Y(_08530_),
    .D(_08529_));
 sg13g2_nor3_1 _15124_ (.A(_08504_),
    .B(_08520_),
    .C(_08530_),
    .Y(_08531_));
 sg13g2_buf_1 _15125_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_08532_));
 sg13g2_buf_1 _15126_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_08533_));
 sg13g2_nor2_1 _15127_ (.A(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sg13g2_buf_2 _15128_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_08535_));
 sg13g2_buf_2 _15129_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_08536_));
 sg13g2_buf_2 _15130_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_08537_));
 sg13g2_buf_2 _15131_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_08538_));
 sg13g2_nor4_1 _15132_ (.A(_08535_),
    .B(_08536_),
    .C(_08537_),
    .D(_08538_),
    .Y(_08539_));
 sg13g2_buf_1 _15133_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_08540_));
 sg13g2_buf_1 _15134_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_08541_));
 sg13g2_buf_2 _15135_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_08542_));
 sg13g2_buf_2 _15136_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_08543_));
 sg13g2_nor4_1 _15137_ (.A(_08540_),
    .B(_08541_),
    .C(_08542_),
    .D(_08543_),
    .Y(_08544_));
 sg13g2_buf_2 _15138_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_08545_));
 sg13g2_buf_2 _15139_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_08546_));
 sg13g2_buf_2 _15140_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_08547_));
 sg13g2_nor3_1 _15141_ (.A(_08545_),
    .B(_08546_),
    .C(_08547_),
    .Y(_08548_));
 sg13g2_and4_1 _15142_ (.A(_08534_),
    .B(_08539_),
    .C(_08544_),
    .D(_08548_),
    .X(_08549_));
 sg13g2_nor3_2 _15143_ (.A(_08481_),
    .B(_08531_),
    .C(_08549_),
    .Y(_08550_));
 sg13g2_nor3_1 _15144_ (.A(\rbzero.map_rom.i_col[0] ),
    .B(_08509_),
    .C(_08500_),
    .Y(_08551_));
 sg13g2_nor2b_1 _15145_ (.A(_08513_),
    .B_N(_08551_),
    .Y(_08552_));
 sg13g2_nor3_1 _15146_ (.A(_08482_),
    .B(\rbzero.map_overlay.i_mapdx[3] ),
    .C(_08552_),
    .Y(_08553_));
 sg13g2_and2_1 _15147_ (.A(_08482_),
    .B(\rbzero.map_overlay.i_mapdx[3] ),
    .X(_08554_));
 sg13g2_xor2_1 _15148_ (.B(\rbzero.map_overlay.i_mapdx[4] ),
    .A(_08513_),
    .X(_08555_));
 sg13g2_xor2_1 _15149_ (.B(\rbzero.map_overlay.i_mapdx[1] ),
    .A(_08509_),
    .X(_08556_));
 sg13g2_xor2_1 _15150_ (.B(\rbzero.map_overlay.i_mapdx[0] ),
    .A(net827),
    .X(_08557_));
 sg13g2_buf_1 _15151_ (.A(_08500_),
    .X(_08558_));
 sg13g2_xor2_1 _15152_ (.B(\rbzero.map_overlay.i_mapdx[2] ),
    .A(net791),
    .X(_08559_));
 sg13g2_nor4_1 _15153_ (.A(_08555_),
    .B(_08556_),
    .C(_08557_),
    .D(_08559_),
    .Y(_08560_));
 sg13g2_o21ai_1 _15154_ (.B1(_08560_),
    .Y(_08561_),
    .A1(_08553_),
    .A2(_08554_));
 sg13g2_buf_1 _15155_ (.A(_08561_),
    .X(_08562_));
 sg13g2_nor4_1 _15156_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .C(\rbzero.map_overlay.i_mapdy[2] ),
    .D(\rbzero.map_overlay.i_mapdy[3] ),
    .Y(_08563_));
 sg13g2_nor3_1 _15157_ (.A(_08491_),
    .B(\rbzero.map_overlay.i_mapdy[4] ),
    .C(_08563_),
    .Y(_08564_));
 sg13g2_and2_1 _15158_ (.A(_08491_),
    .B(\rbzero.map_overlay.i_mapdy[4] ),
    .X(_08565_));
 sg13g2_xor2_1 _15159_ (.B(\rbzero.map_overlay.i_mapdy[3] ),
    .A(_08488_),
    .X(_08566_));
 sg13g2_xor2_1 _15160_ (.B(\rbzero.map_overlay.i_mapdy[2] ),
    .A(_08516_),
    .X(_08567_));
 sg13g2_xor2_1 _15161_ (.B(\rbzero.map_overlay.i_mapdy[1] ),
    .A(_08505_),
    .X(_08568_));
 sg13g2_xor2_1 _15162_ (.B(\rbzero.map_overlay.i_mapdy[0] ),
    .A(_08486_),
    .X(_08569_));
 sg13g2_nor4_1 _15163_ (.A(_08566_),
    .B(_08567_),
    .C(_08568_),
    .D(_08569_),
    .Y(_08570_));
 sg13g2_o21ai_1 _15164_ (.B1(_08570_),
    .Y(_08571_),
    .A1(_08564_),
    .A2(_08565_));
 sg13g2_buf_1 _15165_ (.A(_08571_),
    .X(_08572_));
 sg13g2_xnor2_1 _15166_ (.Y(_08573_),
    .A(_08488_),
    .B(\rbzero.map_overlay.i_othery[3] ));
 sg13g2_xnor2_1 _15167_ (.Y(_08574_),
    .A(net791),
    .B(\rbzero.map_overlay.i_otherx[2] ));
 sg13g2_xor2_1 _15168_ (.B(\rbzero.map_overlay.i_othery[4] ),
    .A(_08491_),
    .X(_08575_));
 sg13g2_xor2_1 _15169_ (.B(\rbzero.map_overlay.i_otherx[1] ),
    .A(_08509_),
    .X(_08576_));
 sg13g2_xor2_1 _15170_ (.B(\rbzero.map_overlay.i_othery[2] ),
    .A(_08517_),
    .X(_08577_));
 sg13g2_xor2_1 _15171_ (.B(\rbzero.map_overlay.i_othery[0] ),
    .A(_08486_),
    .X(_08578_));
 sg13g2_nor4_1 _15172_ (.A(_08575_),
    .B(_08576_),
    .C(_08577_),
    .D(_08578_),
    .Y(_08579_));
 sg13g2_xor2_1 _15173_ (.B(\rbzero.map_overlay.i_othery[1] ),
    .A(_08505_),
    .X(_08580_));
 sg13g2_xor2_1 _15174_ (.B(\rbzero.map_overlay.i_otherx[0] ),
    .A(net827),
    .X(_08581_));
 sg13g2_xor2_1 _15175_ (.B(\rbzero.map_overlay.i_otherx[4] ),
    .A(_08513_),
    .X(_08582_));
 sg13g2_xor2_1 _15176_ (.B(\rbzero.map_overlay.i_otherx[3] ),
    .A(_08482_),
    .X(_08583_));
 sg13g2_nor4_1 _15177_ (.A(_08580_),
    .B(_08581_),
    .C(_08582_),
    .D(_08583_),
    .Y(_08584_));
 sg13g2_nand4_1 _15178_ (.B(_08574_),
    .C(_08579_),
    .A(_08573_),
    .Y(_08585_),
    .D(_08584_));
 sg13g2_nand3_1 _15179_ (.B(_08572_),
    .C(_08585_),
    .A(_08562_),
    .Y(_08586_));
 sg13g2_and2_1 _15180_ (.A(_08550_),
    .B(_08586_),
    .X(_08587_));
 sg13g2_buf_1 _15181_ (.A(_08587_),
    .X(_08588_));
 sg13g2_inv_1 _15182_ (.Y(_08589_),
    .A(_08482_));
 sg13g2_buf_1 _15183_ (.A(_08486_),
    .X(_08590_));
 sg13g2_buf_1 _15184_ (.A(_08488_),
    .X(_08591_));
 sg13g2_inv_1 _15185_ (.Y(_08592_),
    .A(_08491_));
 sg13g2_buf_1 _15186_ (.A(_00019_),
    .X(_08593_));
 sg13g2_nand4_1 _15187_ (.B(net789),
    .C(_08592_),
    .A(net794),
    .Y(_08594_),
    .D(_08593_));
 sg13g2_nor4_1 _15188_ (.A(_08589_),
    .B(net790),
    .C(net792),
    .D(_08594_),
    .Y(_08595_));
 sg13g2_xnor2_1 _15189_ (.Y(_08596_),
    .A(_08482_),
    .B(net794));
 sg13g2_xnor2_1 _15190_ (.Y(_08597_),
    .A(net793),
    .B(net790));
 sg13g2_xnor2_1 _15191_ (.Y(_08598_),
    .A(net791),
    .B(net789));
 sg13g2_xnor2_1 _15192_ (.Y(_08599_),
    .A(net827),
    .B(net792));
 sg13g2_nor4_1 _15193_ (.A(_08596_),
    .B(_08597_),
    .C(_08598_),
    .D(_08599_),
    .Y(_08600_));
 sg13g2_a21oi_1 _15194_ (.A1(_08551_),
    .A2(_08595_),
    .Y(_08601_),
    .B1(_08600_));
 sg13g2_xor2_1 _15195_ (.B(_08516_),
    .A(_08558_),
    .X(_08602_));
 sg13g2_inv_1 _15196_ (.Y(_08603_),
    .A(_08488_));
 sg13g2_buf_2 _15197_ (.A(_00021_),
    .X(_08604_));
 sg13g2_xor2_1 _15198_ (.B(_08505_),
    .A(net793),
    .X(_08605_));
 sg13g2_nand4_1 _15199_ (.B(_08604_),
    .C(_08605_),
    .A(_08603_),
    .Y(_08606_),
    .D(_08602_));
 sg13g2_mux2_1 _15200_ (.A0(_08602_),
    .A1(_08606_),
    .S(net790),
    .X(_08607_));
 sg13g2_nor2_1 _15201_ (.A(net827),
    .B(_08607_),
    .Y(_08608_));
 sg13g2_inv_1 _15202_ (.Y(_08609_),
    .A(net827));
 sg13g2_nor3_1 _15203_ (.A(_08609_),
    .B(net790),
    .C(_08606_),
    .Y(_08610_));
 sg13g2_xnor2_1 _15204_ (.Y(_08611_),
    .A(net790),
    .B(net794));
 sg13g2_nand3_1 _15205_ (.B(net792),
    .C(_08611_),
    .A(net791),
    .Y(_08612_));
 sg13g2_or3_1 _15206_ (.A(net791),
    .B(net792),
    .C(_08611_),
    .X(_08613_));
 sg13g2_buf_1 _15207_ (.A(_00022_),
    .X(_08614_));
 sg13g2_nand2b_1 _15208_ (.Y(_08615_),
    .B(net793),
    .A_N(_08614_));
 sg13g2_a21oi_1 _15209_ (.A1(_08612_),
    .A2(_08613_),
    .Y(_08616_),
    .B1(_08615_));
 sg13g2_and4_1 _15210_ (.A(net790),
    .B(_08506_),
    .C(_08488_),
    .D(_08491_),
    .X(_08617_));
 sg13g2_nor4_1 _15211_ (.A(_08590_),
    .B(_08506_),
    .C(net792),
    .D(net789),
    .Y(_08618_));
 sg13g2_buf_2 _15212_ (.A(_00020_),
    .X(_08619_));
 sg13g2_a22oi_1 _15213_ (.Y(_08620_),
    .B1(_08618_),
    .B2(_08619_),
    .A2(_08617_),
    .A1(net792));
 sg13g2_nand2_1 _15214_ (.Y(_08621_),
    .A(_08589_),
    .B(_08552_));
 sg13g2_nand2_1 _15215_ (.Y(_08622_),
    .A(net793),
    .B(net791));
 sg13g2_nor2_1 _15216_ (.A(_08609_),
    .B(_08622_),
    .Y(_08623_));
 sg13g2_nand3_1 _15217_ (.B(_08513_),
    .C(_08623_),
    .A(_08482_),
    .Y(_08624_));
 sg13g2_nand3_1 _15218_ (.B(_08621_),
    .C(_08624_),
    .A(_08620_),
    .Y(_08625_));
 sg13g2_nor4_1 _15219_ (.A(_08608_),
    .B(_08610_),
    .C(_08616_),
    .D(_08625_),
    .Y(_08626_));
 sg13g2_nand2_1 _15220_ (.Y(_08627_),
    .A(_08601_),
    .B(_08626_));
 sg13g2_nand3b_1 _15221_ (.B(_08627_),
    .C(_08550_),
    .Y(_08628_),
    .A_N(_08588_));
 sg13g2_buf_1 _15222_ (.A(_08628_),
    .X(_08629_));
 sg13g2_nand2b_1 _15223_ (.Y(_08630_),
    .B(_08629_),
    .A_N(_08588_));
 sg13g2_buf_1 _15224_ (.A(_08630_),
    .X(_08631_));
 sg13g2_nand2_2 _15225_ (.Y(_08632_),
    .A(_08480_),
    .B(_08631_));
 sg13g2_nor2_1 _15226_ (.A(net686),
    .B(_08632_),
    .Y(_00009_));
 sg13g2_and2_1 _15227_ (.A(_08432_),
    .B(_08425_),
    .X(_08633_));
 sg13g2_buf_1 _15228_ (.A(_08633_),
    .X(_08634_));
 sg13g2_buf_1 _15229_ (.A(_08634_),
    .X(_08635_));
 sg13g2_a21oi_1 _15230_ (.A1(net611),
    .A2(_08437_),
    .Y(_08636_),
    .B1(net546));
 sg13g2_nor2_1 _15231_ (.A(net686),
    .B(_08636_),
    .Y(_00008_));
 sg13g2_inv_1 _15232_ (.Y(_08637_),
    .A(_08409_));
 sg13g2_buf_1 _15233_ (.A(_08637_),
    .X(_08638_));
 sg13g2_nor2_1 _15234_ (.A(_08638_),
    .B(\rbzero.vga_sync.vsync ),
    .Y(_08639_));
 sg13g2_buf_1 _15235_ (.A(_08639_),
    .X(_08640_));
 sg13g2_buf_1 _15236_ (.A(_08640_),
    .X(_08641_));
 sg13g2_buf_1 _15237_ (.A(net610),
    .X(_08642_));
 sg13g2_buf_1 _15238_ (.A(\rbzero.wall_tracer.rcp_fsm.state[0] ),
    .X(_08643_));
 sg13g2_buf_1 _15239_ (.A(\rbzero.wall_tracer.rcp_fsm.state[1] ),
    .X(_08644_));
 sg13g2_buf_1 _15240_ (.A(_08644_),
    .X(_08645_));
 sg13g2_buf_1 _15241_ (.A(net788),
    .X(_08646_));
 sg13g2_a21oi_1 _15242_ (.A1(_08422_),
    .A2(_08643_),
    .Y(_08647_),
    .B1(net724));
 sg13g2_nand2_1 _15243_ (.Y(_00004_),
    .A(_08642_),
    .B(_08647_));
 sg13g2_buf_1 _15244_ (.A(_08466_),
    .X(_08648_));
 sg13g2_buf_2 _15245_ (.A(_00024_),
    .X(_08649_));
 sg13g2_xnor2_1 _15246_ (.Y(_08650_),
    .A(net831),
    .B(_08649_));
 sg13g2_buf_1 _15247_ (.A(_08468_),
    .X(_08651_));
 sg13g2_and2_1 _15248_ (.A(net830),
    .B(net796),
    .X(_08652_));
 sg13g2_buf_1 _15249_ (.A(_08652_),
    .X(_08653_));
 sg13g2_o21ai_1 _15250_ (.B1(_08465_),
    .Y(_08654_),
    .A1(_08651_),
    .A2(_08653_));
 sg13g2_inv_1 _15251_ (.Y(_08655_),
    .A(net831));
 sg13g2_inv_1 _15252_ (.Y(_08656_),
    .A(_08649_));
 sg13g2_nor2_1 _15253_ (.A(_08655_),
    .B(_08656_),
    .Y(_08657_));
 sg13g2_nor3_1 _15254_ (.A(net787),
    .B(net831),
    .C(_08654_),
    .Y(_08658_));
 sg13g2_a221oi_1 _15255_ (.B2(_08657_),
    .C1(_08658_),
    .B1(_08654_),
    .A1(net787),
    .Y(_08659_),
    .A2(_08650_));
 sg13g2_nor3_1 _15256_ (.A(net787),
    .B(_08452_),
    .C(_08649_),
    .Y(_08660_));
 sg13g2_nand3_1 _15257_ (.B(_08654_),
    .C(_08660_),
    .A(_08470_),
    .Y(_08661_));
 sg13g2_o21ai_1 _15258_ (.B1(_08661_),
    .Y(_08662_),
    .A1(_08470_),
    .A2(_08659_));
 sg13g2_buf_1 _15259_ (.A(_08465_),
    .X(_08663_));
 sg13g2_buf_2 _15260_ (.A(_00025_),
    .X(_08664_));
 sg13g2_nor2_1 _15261_ (.A(net785),
    .B(_08664_),
    .Y(_08665_));
 sg13g2_a21oi_1 _15262_ (.A1(net785),
    .A2(_08653_),
    .Y(_08666_),
    .B1(net786));
 sg13g2_o21ai_1 _15263_ (.B1(_08649_),
    .Y(_08667_),
    .A1(_08665_),
    .A2(_08666_));
 sg13g2_nand4_1 _15264_ (.B(net785),
    .C(_08656_),
    .A(net786),
    .Y(_08668_),
    .D(_08664_));
 sg13g2_nand3_1 _15265_ (.B(_08667_),
    .C(_08668_),
    .A(_08662_),
    .Y(\rbzero.o_tex_csb ));
 sg13g2_buf_2 _15266_ (.A(\rbzero.wall_tracer.state[4] ),
    .X(_08669_));
 sg13g2_buf_1 _15267_ (.A(_08669_),
    .X(_08670_));
 sg13g2_a21oi_1 _15268_ (.A1(net685),
    .A2(_08437_),
    .Y(_08671_),
    .B1(net784));
 sg13g2_nor2_1 _15269_ (.A(_08413_),
    .B(_08671_),
    .Y(_00007_));
 sg13g2_inv_2 _15270_ (.Y(_08672_),
    .A(_08479_));
 sg13g2_or2_1 _15271_ (.X(_08673_),
    .B(_08631_),
    .A(_08672_));
 sg13g2_nand2_1 _15272_ (.Y(_08674_),
    .A(net684),
    .B(_08475_));
 sg13g2_buf_2 _15273_ (.A(_08411_),
    .X(_08675_));
 sg13g2_buf_1 _15274_ (.A(_08675_),
    .X(_08676_));
 sg13g2_a21oi_1 _15275_ (.A1(_08673_),
    .A2(_08674_),
    .Y(_00006_),
    .B1(net682));
 sg13g2_and4_1 _15276_ (.A(_08452_),
    .B(_08464_),
    .C(_08467_),
    .D(_08471_),
    .X(_08677_));
 sg13g2_buf_1 _15277_ (.A(_08677_),
    .X(_08678_));
 sg13g2_nand2_1 _15278_ (.Y(_08679_),
    .A(\rbzero.wall_tracer.state[8] ),
    .B(net490));
 sg13g2_buf_2 _15279_ (.A(_08679_),
    .X(_08680_));
 sg13g2_buf_1 _15280_ (.A(_08680_),
    .X(_08681_));
 sg13g2_buf_1 _15281_ (.A(net464),
    .X(_08682_));
 sg13g2_nand2_1 _15282_ (.Y(_00005_),
    .A(net545),
    .B(_08682_));
 sg13g2_inv_1 _15283_ (.Y(_08683_),
    .A(net786));
 sg13g2_nand2_1 _15284_ (.Y(_08684_),
    .A(_08656_),
    .B(_08664_));
 sg13g2_nand3b_1 _15285_ (.B(_08649_),
    .C(net785),
    .Y(_08685_),
    .A_N(_08664_));
 sg13g2_o21ai_1 _15286_ (.B1(_08685_),
    .Y(_08686_),
    .A1(net785),
    .A2(_08684_));
 sg13g2_nand2b_1 _15287_ (.Y(_08687_),
    .B(_08686_),
    .A_N(_08653_));
 sg13g2_nand4_1 _15288_ (.B(net785),
    .C(_08649_),
    .A(_08683_),
    .Y(_08688_),
    .D(_08653_));
 sg13g2_o21ai_1 _15289_ (.B1(_08688_),
    .Y(_08689_),
    .A1(_08683_),
    .A2(_08687_));
 sg13g2_and2_1 _15290_ (.A(_08662_),
    .B(_08689_),
    .X(net13));
 sg13g2_nand2_1 _15291_ (.Y(_08690_),
    .A(net832),
    .B(_08643_));
 sg13g2_buf_1 _15292_ (.A(_08690_),
    .X(_08691_));
 sg13g2_buf_1 _15293_ (.A(_08691_),
    .X(_08692_));
 sg13g2_nor2_1 _15294_ (.A(_08413_),
    .B(_08692_),
    .Y(_00002_));
 sg13g2_buf_1 _15295_ (.A(net610),
    .X(_08693_));
 sg13g2_and2_1 _15296_ (.A(\rbzero.wall_tracer.rcp_fsm.state[2] ),
    .B(net544),
    .X(_00003_));
 sg13g2_and2_1 _15297_ (.A(\rbzero.wall_tracer.rcp_fsm.state[3] ),
    .B(net544),
    .X(_00001_));
 sg13g2_and2_1 _15298_ (.A(\rbzero.wall_tracer.rcp_fsm.state[4] ),
    .B(net544),
    .X(_00000_));
 sg13g2_nand2_1 _15299_ (.Y(_08694_),
    .A(net786),
    .B(_08664_));
 sg13g2_xnor2_1 _15300_ (.Y(_08695_),
    .A(_08656_),
    .B(_08694_));
 sg13g2_and2_1 _15301_ (.A(_08662_),
    .B(_08695_),
    .X(_08696_));
 sg13g2_buf_1 _15302_ (.A(_08696_),
    .X(_08697_));
 sg13g2_nand2_1 _15303_ (.Y(_08698_),
    .A(\rbzero.debug_overlay.h[0] ),
    .B(_08697_));
 sg13g2_buf_2 _15304_ (.A(_08698_),
    .X(_08699_));
 sg13g2_buf_1 _15305_ (.A(_08699_),
    .X(_08700_));
 sg13g2_mux2_1 _15306_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(net437),
    .X(_01069_));
 sg13g2_mux2_1 _15307_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(net437),
    .X(_01070_));
 sg13g2_mux2_1 _15308_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(net437),
    .X(_01071_));
 sg13g2_mux2_1 _15309_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_08700_),
    .X(_01072_));
 sg13g2_mux2_1 _15310_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_08700_),
    .X(_01073_));
 sg13g2_mux2_1 _15311_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(net437),
    .X(_01074_));
 sg13g2_mux2_1 _15312_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(net437),
    .X(_01075_));
 sg13g2_mux2_1 _15313_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(net437),
    .X(_01076_));
 sg13g2_mux2_1 _15314_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(net437),
    .X(_01077_));
 sg13g2_mux2_1 _15315_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(net437),
    .X(_01078_));
 sg13g2_buf_1 _15316_ (.A(_08699_),
    .X(_08701_));
 sg13g2_mux2_1 _15317_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(net436),
    .X(_01079_));
 sg13g2_mux2_1 _15318_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_08701_),
    .X(_01080_));
 sg13g2_mux2_1 _15319_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(net436),
    .X(_01081_));
 sg13g2_mux2_1 _15320_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_08701_),
    .X(_01082_));
 sg13g2_mux2_1 _15321_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(net436),
    .X(_01083_));
 sg13g2_mux2_1 _15322_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(net436),
    .X(_01084_));
 sg13g2_mux2_1 _15323_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(net436),
    .X(_01085_));
 sg13g2_mux2_1 _15324_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(net436),
    .X(_01086_));
 sg13g2_mux2_1 _15325_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(net436),
    .X(_01087_));
 sg13g2_mux2_1 _15326_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(net436),
    .X(_01088_));
 sg13g2_buf_1 _15327_ (.A(_08699_),
    .X(_08702_));
 sg13g2_mux2_1 _15328_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(net435),
    .X(_01089_));
 sg13g2_mux2_1 _15329_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(net435),
    .X(_01090_));
 sg13g2_mux2_1 _15330_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(net435),
    .X(_01091_));
 sg13g2_mux2_1 _15331_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(net435),
    .X(_01092_));
 sg13g2_mux2_1 _15332_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(net435),
    .X(_01093_));
 sg13g2_mux2_1 _15333_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(net435),
    .X(_01094_));
 sg13g2_mux2_1 _15334_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(net435),
    .X(_01095_));
 sg13g2_mux2_1 _15335_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(net435),
    .X(_01096_));
 sg13g2_mux2_1 _15336_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_08702_),
    .X(_01097_));
 sg13g2_mux2_1 _15337_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_08702_),
    .X(_01098_));
 sg13g2_buf_1 _15338_ (.A(_08699_),
    .X(_08703_));
 sg13g2_mux2_1 _15339_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(net434),
    .X(_01099_));
 sg13g2_mux2_1 _15340_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(net434),
    .X(_01100_));
 sg13g2_mux2_1 _15341_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(net434),
    .X(_01101_));
 sg13g2_mux2_1 _15342_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(net434),
    .X(_01102_));
 sg13g2_mux2_1 _15343_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(net434),
    .X(_01103_));
 sg13g2_mux2_1 _15344_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(net434),
    .X(_01104_));
 sg13g2_mux2_1 _15345_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(net434),
    .X(_01105_));
 sg13g2_mux2_1 _15346_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_08703_),
    .X(_01106_));
 sg13g2_mux2_1 _15347_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(net434),
    .X(_01107_));
 sg13g2_mux2_1 _15348_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_08703_),
    .X(_01108_));
 sg13g2_buf_1 _15349_ (.A(_08699_),
    .X(_08704_));
 sg13g2_mux2_1 _15350_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(net433),
    .X(_01109_));
 sg13g2_mux2_1 _15351_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(net433),
    .X(_01110_));
 sg13g2_mux2_1 _15352_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(net433),
    .X(_01111_));
 sg13g2_mux2_1 _15353_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(net433),
    .X(_01112_));
 sg13g2_mux2_1 _15354_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_08704_),
    .X(_01113_));
 sg13g2_mux2_1 _15355_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(net433),
    .X(_01114_));
 sg13g2_mux2_1 _15356_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(net433),
    .X(_01115_));
 sg13g2_mux2_1 _15357_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(net433),
    .X(_01116_));
 sg13g2_mux2_1 _15358_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(net433),
    .X(_01117_));
 sg13g2_mux2_1 _15359_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_08704_),
    .X(_01118_));
 sg13g2_buf_1 _15360_ (.A(_08699_),
    .X(_08705_));
 sg13g2_mux2_1 _15361_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(net432),
    .X(_01119_));
 sg13g2_mux2_1 _15362_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(net432),
    .X(_01120_));
 sg13g2_mux2_1 _15363_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(net432),
    .X(_01121_));
 sg13g2_mux2_1 _15364_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(net432),
    .X(_01122_));
 sg13g2_mux2_1 _15365_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(net432),
    .X(_01123_));
 sg13g2_mux2_1 _15366_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(net432),
    .X(_01124_));
 sg13g2_mux2_1 _15367_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_08705_),
    .X(_01125_));
 sg13g2_mux2_1 _15368_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_08705_),
    .X(_01126_));
 sg13g2_mux2_1 _15369_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(net432),
    .X(_01127_));
 sg13g2_mux2_1 _15370_ (.A0(net12),
    .A1(\rbzero.tex_b0[63] ),
    .S(net432),
    .X(_01128_));
 sg13g2_buf_1 _15371_ (.A(_08698_),
    .X(_08706_));
 sg13g2_buf_1 _15372_ (.A(_08706_),
    .X(_08707_));
 sg13g2_buf_1 _15373_ (.A(_08707_),
    .X(_08708_));
 sg13g2_mux2_1 _15374_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(net402),
    .X(_01129_));
 sg13g2_mux2_1 _15375_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(net402),
    .X(_01130_));
 sg13g2_mux2_1 _15376_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(net402),
    .X(_01131_));
 sg13g2_mux2_1 _15377_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(net402),
    .X(_01132_));
 sg13g2_buf_1 _15378_ (.A(net828),
    .X(_08709_));
 sg13g2_buf_1 _15379_ (.A(net783),
    .X(_08710_));
 sg13g2_nand2_1 _15380_ (.Y(_08711_),
    .A(_08710_),
    .B(_08697_));
 sg13g2_buf_2 _15381_ (.A(_08711_),
    .X(_08712_));
 sg13g2_buf_1 _15382_ (.A(_08712_),
    .X(_08713_));
 sg13g2_mux2_1 _15383_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(net431),
    .X(_01133_));
 sg13g2_mux2_1 _15384_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(net431),
    .X(_01134_));
 sg13g2_mux2_1 _15385_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(net431),
    .X(_01135_));
 sg13g2_mux2_1 _15386_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_08713_),
    .X(_01136_));
 sg13g2_mux2_1 _15387_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(net431),
    .X(_01137_));
 sg13g2_mux2_1 _15388_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(net431),
    .X(_01138_));
 sg13g2_mux2_1 _15389_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_08713_),
    .X(_01139_));
 sg13g2_mux2_1 _15390_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(net431),
    .X(_01140_));
 sg13g2_mux2_1 _15391_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(net431),
    .X(_01141_));
 sg13g2_mux2_1 _15392_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(net431),
    .X(_01142_));
 sg13g2_buf_1 _15393_ (.A(_08712_),
    .X(_08714_));
 sg13g2_mux2_1 _15394_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(net430),
    .X(_01143_));
 sg13g2_mux2_1 _15395_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_08714_),
    .X(_01144_));
 sg13g2_mux2_1 _15396_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(net430),
    .X(_01145_));
 sg13g2_mux2_1 _15397_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(net430),
    .X(_01146_));
 sg13g2_mux2_1 _15398_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(net430),
    .X(_01147_));
 sg13g2_mux2_1 _15399_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_08714_),
    .X(_01148_));
 sg13g2_mux2_1 _15400_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(net430),
    .X(_01149_));
 sg13g2_mux2_1 _15401_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(net430),
    .X(_01150_));
 sg13g2_mux2_1 _15402_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(net430),
    .X(_01151_));
 sg13g2_mux2_1 _15403_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(net430),
    .X(_01152_));
 sg13g2_buf_1 _15404_ (.A(_08712_),
    .X(_08715_));
 sg13g2_mux2_1 _15405_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(net429),
    .X(_01153_));
 sg13g2_mux2_1 _15406_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_08715_),
    .X(_01154_));
 sg13g2_mux2_1 _15407_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(net429),
    .X(_01155_));
 sg13g2_mux2_1 _15408_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_08715_),
    .X(_01156_));
 sg13g2_mux2_1 _15409_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(net429),
    .X(_01157_));
 sg13g2_mux2_1 _15410_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(net429),
    .X(_01158_));
 sg13g2_mux2_1 _15411_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(net429),
    .X(_01159_));
 sg13g2_mux2_1 _15412_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(net429),
    .X(_01160_));
 sg13g2_mux2_1 _15413_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(net429),
    .X(_01161_));
 sg13g2_mux2_1 _15414_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(net429),
    .X(_01162_));
 sg13g2_buf_1 _15415_ (.A(_08712_),
    .X(_08716_));
 sg13g2_mux2_1 _15416_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(net428),
    .X(_01163_));
 sg13g2_mux2_1 _15417_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_08716_),
    .X(_01164_));
 sg13g2_mux2_1 _15418_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(net428),
    .X(_01165_));
 sg13g2_mux2_1 _15419_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_08716_),
    .X(_01166_));
 sg13g2_mux2_1 _15420_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(net428),
    .X(_01167_));
 sg13g2_mux2_1 _15421_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(net428),
    .X(_01168_));
 sg13g2_mux2_1 _15422_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(net428),
    .X(_01169_));
 sg13g2_mux2_1 _15423_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(net428),
    .X(_01170_));
 sg13g2_mux2_1 _15424_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(net428),
    .X(_01171_));
 sg13g2_mux2_1 _15425_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(net428),
    .X(_01172_));
 sg13g2_buf_1 _15426_ (.A(_08712_),
    .X(_08717_));
 sg13g2_mux2_1 _15427_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(net427),
    .X(_01173_));
 sg13g2_mux2_1 _15428_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(net427),
    .X(_01174_));
 sg13g2_mux2_1 _15429_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(net427),
    .X(_01175_));
 sg13g2_mux2_1 _15430_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(net427),
    .X(_01176_));
 sg13g2_mux2_1 _15431_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_08717_),
    .X(_01177_));
 sg13g2_mux2_1 _15432_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_08717_),
    .X(_01178_));
 sg13g2_mux2_1 _15433_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(net427),
    .X(_01179_));
 sg13g2_mux2_1 _15434_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(net427),
    .X(_01180_));
 sg13g2_mux2_1 _15435_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(net427),
    .X(_01181_));
 sg13g2_mux2_1 _15436_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(net427),
    .X(_01182_));
 sg13g2_buf_1 _15437_ (.A(_08712_),
    .X(_08718_));
 sg13g2_mux2_1 _15438_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(net426),
    .X(_01183_));
 sg13g2_mux2_1 _15439_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(net426),
    .X(_01184_));
 sg13g2_mux2_1 _15440_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(net426),
    .X(_01185_));
 sg13g2_mux2_1 _15441_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(net426),
    .X(_01186_));
 sg13g2_mux2_1 _15442_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(net426),
    .X(_01187_));
 sg13g2_mux2_1 _15443_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_08718_),
    .X(_01188_));
 sg13g2_mux2_1 _15444_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_08718_),
    .X(_01189_));
 sg13g2_mux2_1 _15445_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(net426),
    .X(_01190_));
 sg13g2_mux2_1 _15446_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(net426),
    .X(_01191_));
 sg13g2_mux2_1 _15447_ (.A0(net12),
    .A1(\rbzero.tex_b1[63] ),
    .S(net426),
    .X(_01192_));
 sg13g2_buf_1 _15448_ (.A(_08711_),
    .X(_08719_));
 sg13g2_buf_1 _15449_ (.A(_08719_),
    .X(_08720_));
 sg13g2_buf_1 _15450_ (.A(_08720_),
    .X(_08721_));
 sg13g2_mux2_1 _15451_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(net401),
    .X(_01193_));
 sg13g2_mux2_1 _15452_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(net401),
    .X(_01194_));
 sg13g2_mux2_1 _15453_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_08721_),
    .X(_01195_));
 sg13g2_mux2_1 _15454_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_08721_),
    .X(_01196_));
 sg13g2_mux2_1 _15455_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(net402),
    .X(_01197_));
 sg13g2_mux2_1 _15456_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_08708_),
    .X(_01198_));
 sg13g2_mux2_1 _15457_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_08708_),
    .X(_01199_));
 sg13g2_mux2_1 _15458_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(net402),
    .X(_01200_));
 sg13g2_mux2_1 _15459_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(net402),
    .X(_01201_));
 sg13g2_mux2_1 _15460_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(net402),
    .X(_01202_));
 sg13g2_buf_1 _15461_ (.A(_08707_),
    .X(_08722_));
 sg13g2_mux2_1 _15462_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(net400),
    .X(_01203_));
 sg13g2_mux2_1 _15463_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_08722_),
    .X(_01204_));
 sg13g2_mux2_1 _15464_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(net400),
    .X(_01205_));
 sg13g2_mux2_1 _15465_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(net400),
    .X(_01206_));
 sg13g2_mux2_1 _15466_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(net400),
    .X(_01207_));
 sg13g2_mux2_1 _15467_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_08722_),
    .X(_01208_));
 sg13g2_mux2_1 _15468_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(net400),
    .X(_01209_));
 sg13g2_mux2_1 _15469_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(net400),
    .X(_01210_));
 sg13g2_mux2_1 _15470_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(net400),
    .X(_01211_));
 sg13g2_mux2_1 _15471_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(net400),
    .X(_01212_));
 sg13g2_buf_1 _15472_ (.A(_08707_),
    .X(_08723_));
 sg13g2_mux2_1 _15473_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(net399),
    .X(_01213_));
 sg13g2_mux2_1 _15474_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(net399),
    .X(_01214_));
 sg13g2_mux2_1 _15475_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(net399),
    .X(_01215_));
 sg13g2_mux2_1 _15476_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(net399),
    .X(_01216_));
 sg13g2_mux2_1 _15477_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(net399),
    .X(_01217_));
 sg13g2_mux2_1 _15478_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(net399),
    .X(_01218_));
 sg13g2_mux2_1 _15479_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_08723_),
    .X(_01219_));
 sg13g2_mux2_1 _15480_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(net399),
    .X(_01220_));
 sg13g2_mux2_1 _15481_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(net399),
    .X(_01221_));
 sg13g2_mux2_1 _15482_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_08723_),
    .X(_01222_));
 sg13g2_buf_1 _15483_ (.A(_08707_),
    .X(_08724_));
 sg13g2_mux2_1 _15484_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(net398),
    .X(_01223_));
 sg13g2_mux2_1 _15485_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(net398),
    .X(_01224_));
 sg13g2_mux2_1 _15486_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(net398),
    .X(_01225_));
 sg13g2_mux2_1 _15487_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(net398),
    .X(_01226_));
 sg13g2_mux2_1 _15488_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(net398),
    .X(_01227_));
 sg13g2_mux2_1 _15489_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(net398),
    .X(_01228_));
 sg13g2_mux2_1 _15490_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(net398),
    .X(_01229_));
 sg13g2_mux2_1 _15491_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(net398),
    .X(_01230_));
 sg13g2_mux2_1 _15492_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_08724_),
    .X(_01231_));
 sg13g2_mux2_1 _15493_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_08724_),
    .X(_01232_));
 sg13g2_buf_1 _15494_ (.A(_08707_),
    .X(_08725_));
 sg13g2_mux2_1 _15495_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(net397),
    .X(_01233_));
 sg13g2_mux2_1 _15496_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(net397),
    .X(_01234_));
 sg13g2_mux2_1 _15497_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(net397),
    .X(_01235_));
 sg13g2_mux2_1 _15498_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(net397),
    .X(_01236_));
 sg13g2_mux2_1 _15499_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(net397),
    .X(_01237_));
 sg13g2_mux2_1 _15500_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(net397),
    .X(_01238_));
 sg13g2_mux2_1 _15501_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_08725_),
    .X(_01239_));
 sg13g2_mux2_1 _15502_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(net397),
    .X(_01240_));
 sg13g2_mux2_1 _15503_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(net397),
    .X(_01241_));
 sg13g2_mux2_1 _15504_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_08725_),
    .X(_01242_));
 sg13g2_buf_1 _15505_ (.A(_08707_),
    .X(_08726_));
 sg13g2_mux2_1 _15506_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(net396),
    .X(_01243_));
 sg13g2_mux2_1 _15507_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(net396),
    .X(_01244_));
 sg13g2_mux2_1 _15508_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(net396),
    .X(_01245_));
 sg13g2_mux2_1 _15509_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(net396),
    .X(_01246_));
 sg13g2_mux2_1 _15510_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(net396),
    .X(_01247_));
 sg13g2_mux2_1 _15511_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(net396),
    .X(_01248_));
 sg13g2_mux2_1 _15512_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(net396),
    .X(_01249_));
 sg13g2_mux2_1 _15513_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_08726_),
    .X(_01250_));
 sg13g2_mux2_1 _15514_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_08726_),
    .X(_01251_));
 sg13g2_mux2_1 _15515_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(net396),
    .X(_01252_));
 sg13g2_buf_1 _15516_ (.A(_08707_),
    .X(_08727_));
 sg13g2_mux2_1 _15517_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(net395),
    .X(_01253_));
 sg13g2_mux2_1 _15518_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(net395),
    .X(_01254_));
 sg13g2_mux2_1 _15519_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(net395),
    .X(_01255_));
 sg13g2_mux2_1 _15520_ (.A0(net11),
    .A1(\rbzero.tex_g0[63] ),
    .S(net395),
    .X(_01256_));
 sg13g2_mux2_1 _15521_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(net395),
    .X(_01257_));
 sg13g2_mux2_1 _15522_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(net395),
    .X(_01258_));
 sg13g2_mux2_1 _15523_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(net395),
    .X(_01259_));
 sg13g2_mux2_1 _15524_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(net395),
    .X(_01260_));
 sg13g2_mux2_1 _15525_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[0] ),
    .S(net401),
    .X(_01261_));
 sg13g2_mux2_1 _15526_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(net401),
    .X(_01262_));
 sg13g2_mux2_1 _15527_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(net401),
    .X(_01263_));
 sg13g2_mux2_1 _15528_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(net401),
    .X(_01264_));
 sg13g2_mux2_1 _15529_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(net401),
    .X(_01265_));
 sg13g2_mux2_1 _15530_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(net401),
    .X(_01266_));
 sg13g2_buf_1 _15531_ (.A(_08720_),
    .X(_08728_));
 sg13g2_mux2_1 _15532_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(net394),
    .X(_01267_));
 sg13g2_mux2_1 _15533_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_08728_),
    .X(_01268_));
 sg13g2_mux2_1 _15534_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(net394),
    .X(_01269_));
 sg13g2_mux2_1 _15535_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(net394),
    .X(_01270_));
 sg13g2_mux2_1 _15536_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(net394),
    .X(_01271_));
 sg13g2_mux2_1 _15537_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_08728_),
    .X(_01272_));
 sg13g2_mux2_1 _15538_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(net394),
    .X(_01273_));
 sg13g2_mux2_1 _15539_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(net394),
    .X(_01274_));
 sg13g2_mux2_1 _15540_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(net394),
    .X(_01275_));
 sg13g2_mux2_1 _15541_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(net394),
    .X(_01276_));
 sg13g2_buf_1 _15542_ (.A(_08720_),
    .X(_08729_));
 sg13g2_mux2_1 _15543_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(net393),
    .X(_01277_));
 sg13g2_mux2_1 _15544_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(net393),
    .X(_01278_));
 sg13g2_mux2_1 _15545_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(net393),
    .X(_01279_));
 sg13g2_mux2_1 _15546_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(net393),
    .X(_01280_));
 sg13g2_mux2_1 _15547_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(net393),
    .X(_01281_));
 sg13g2_mux2_1 _15548_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(net393),
    .X(_01282_));
 sg13g2_mux2_1 _15549_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_08729_),
    .X(_01283_));
 sg13g2_mux2_1 _15550_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(net393),
    .X(_01284_));
 sg13g2_mux2_1 _15551_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(net393),
    .X(_01285_));
 sg13g2_mux2_1 _15552_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_08729_),
    .X(_01286_));
 sg13g2_buf_1 _15553_ (.A(_08720_),
    .X(_08730_));
 sg13g2_mux2_1 _15554_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(net392),
    .X(_01287_));
 sg13g2_mux2_1 _15555_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(net392),
    .X(_01288_));
 sg13g2_mux2_1 _15556_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(net392),
    .X(_01289_));
 sg13g2_mux2_1 _15557_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(net392),
    .X(_01290_));
 sg13g2_mux2_1 _15558_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(net392),
    .X(_01291_));
 sg13g2_mux2_1 _15559_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(net392),
    .X(_01292_));
 sg13g2_mux2_1 _15560_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(net392),
    .X(_01293_));
 sg13g2_mux2_1 _15561_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(net392),
    .X(_01294_));
 sg13g2_mux2_1 _15562_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_08730_),
    .X(_01295_));
 sg13g2_mux2_1 _15563_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_08730_),
    .X(_01296_));
 sg13g2_buf_1 _15564_ (.A(_08720_),
    .X(_08731_));
 sg13g2_mux2_1 _15565_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(net391),
    .X(_01297_));
 sg13g2_mux2_1 _15566_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(net391),
    .X(_01298_));
 sg13g2_mux2_1 _15567_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(net391),
    .X(_01299_));
 sg13g2_mux2_1 _15568_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(net391),
    .X(_01300_));
 sg13g2_mux2_1 _15569_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(net391),
    .X(_01301_));
 sg13g2_mux2_1 _15570_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(net391),
    .X(_01302_));
 sg13g2_mux2_1 _15571_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(net391),
    .X(_01303_));
 sg13g2_mux2_1 _15572_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_08731_),
    .X(_01304_));
 sg13g2_mux2_1 _15573_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_08731_),
    .X(_01305_));
 sg13g2_mux2_1 _15574_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(net391),
    .X(_01306_));
 sg13g2_buf_1 _15575_ (.A(_08720_),
    .X(_08732_));
 sg13g2_mux2_1 _15576_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(net390),
    .X(_01307_));
 sg13g2_mux2_1 _15577_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(net390),
    .X(_01308_));
 sg13g2_mux2_1 _15578_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(net390),
    .X(_01309_));
 sg13g2_mux2_1 _15579_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(net390),
    .X(_01310_));
 sg13g2_mux2_1 _15580_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(net390),
    .X(_01311_));
 sg13g2_mux2_1 _15581_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(net390),
    .X(_01312_));
 sg13g2_mux2_1 _15582_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(net390),
    .X(_01313_));
 sg13g2_mux2_1 _15583_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_08732_),
    .X(_01314_));
 sg13g2_mux2_1 _15584_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_08732_),
    .X(_01315_));
 sg13g2_mux2_1 _15585_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(net390),
    .X(_01316_));
 sg13g2_buf_1 _15586_ (.A(_08720_),
    .X(_08733_));
 sg13g2_mux2_1 _15587_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(net389),
    .X(_01317_));
 sg13g2_mux2_1 _15588_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(net389),
    .X(_01318_));
 sg13g2_mux2_1 _15589_ (.A0(\rbzero.tex_g1[63] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(net389),
    .X(_01319_));
 sg13g2_mux2_1 _15590_ (.A0(net11),
    .A1(\rbzero.tex_g1[63] ),
    .S(net389),
    .X(_01320_));
 sg13g2_mux2_1 _15591_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(net389),
    .X(_01321_));
 sg13g2_mux2_1 _15592_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(net389),
    .X(_01322_));
 sg13g2_mux2_1 _15593_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(net389),
    .X(_01323_));
 sg13g2_mux2_1 _15594_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(net389),
    .X(_01324_));
 sg13g2_mux2_1 _15595_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_08727_),
    .X(_01325_));
 sg13g2_mux2_1 _15596_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_08727_),
    .X(_01326_));
 sg13g2_buf_1 _15597_ (.A(_08706_),
    .X(_08734_));
 sg13g2_mux2_1 _15598_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(net425),
    .X(_01327_));
 sg13g2_mux2_1 _15599_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(net425),
    .X(_01328_));
 sg13g2_mux2_1 _15600_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(net425),
    .X(_01329_));
 sg13g2_mux2_1 _15601_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(net425),
    .X(_01330_));
 sg13g2_mux2_1 _15602_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(net425),
    .X(_01331_));
 sg13g2_mux2_1 _15603_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(net425),
    .X(_01332_));
 sg13g2_mux2_1 _15604_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(net425),
    .X(_01333_));
 sg13g2_mux2_1 _15605_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_08734_),
    .X(_01334_));
 sg13g2_mux2_1 _15606_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(net425),
    .X(_01335_));
 sg13g2_mux2_1 _15607_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_08734_),
    .X(_01336_));
 sg13g2_buf_1 _15608_ (.A(_08706_),
    .X(_08735_));
 sg13g2_mux2_1 _15609_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(net424),
    .X(_01337_));
 sg13g2_mux2_1 _15610_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(net424),
    .X(_01338_));
 sg13g2_mux2_1 _15611_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(net424),
    .X(_01339_));
 sg13g2_mux2_1 _15612_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(net424),
    .X(_01340_));
 sg13g2_mux2_1 _15613_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(net424),
    .X(_01341_));
 sg13g2_mux2_1 _15614_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(net424),
    .X(_01342_));
 sg13g2_mux2_1 _15615_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_08735_),
    .X(_01343_));
 sg13g2_mux2_1 _15616_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_08735_),
    .X(_01344_));
 sg13g2_mux2_1 _15617_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(net424),
    .X(_01345_));
 sg13g2_mux2_1 _15618_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(net424),
    .X(_01346_));
 sg13g2_buf_1 _15619_ (.A(_08706_),
    .X(_08736_));
 sg13g2_mux2_1 _15620_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(net423),
    .X(_01347_));
 sg13g2_mux2_1 _15621_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_08736_),
    .X(_01348_));
 sg13g2_mux2_1 _15622_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(net423),
    .X(_01349_));
 sg13g2_mux2_1 _15623_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(net423),
    .X(_01350_));
 sg13g2_mux2_1 _15624_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_08736_),
    .X(_01351_));
 sg13g2_mux2_1 _15625_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(net423),
    .X(_01352_));
 sg13g2_mux2_1 _15626_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(net423),
    .X(_01353_));
 sg13g2_mux2_1 _15627_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(net423),
    .X(_01354_));
 sg13g2_mux2_1 _15628_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(net423),
    .X(_01355_));
 sg13g2_mux2_1 _15629_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(net423),
    .X(_01356_));
 sg13g2_buf_1 _15630_ (.A(_08706_),
    .X(_08737_));
 sg13g2_mux2_1 _15631_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(net422),
    .X(_01357_));
 sg13g2_mux2_1 _15632_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(net422),
    .X(_01358_));
 sg13g2_mux2_1 _15633_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(net422),
    .X(_01359_));
 sg13g2_mux2_1 _15634_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(net422),
    .X(_01360_));
 sg13g2_mux2_1 _15635_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(net422),
    .X(_01361_));
 sg13g2_mux2_1 _15636_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(net422),
    .X(_01362_));
 sg13g2_mux2_1 _15637_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(net422),
    .X(_01363_));
 sg13g2_mux2_1 _15638_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_08737_),
    .X(_01364_));
 sg13g2_mux2_1 _15639_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_08737_),
    .X(_01365_));
 sg13g2_mux2_1 _15640_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(net422),
    .X(_01366_));
 sg13g2_buf_1 _15641_ (.A(_08706_),
    .X(_08738_));
 sg13g2_mux2_1 _15642_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(net421),
    .X(_01367_));
 sg13g2_mux2_1 _15643_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(net421),
    .X(_01368_));
 sg13g2_mux2_1 _15644_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_08738_),
    .X(_01369_));
 sg13g2_mux2_1 _15645_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(net421),
    .X(_01370_));
 sg13g2_mux2_1 _15646_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_08738_),
    .X(_01371_));
 sg13g2_mux2_1 _15647_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(net421),
    .X(_01372_));
 sg13g2_mux2_1 _15648_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(net421),
    .X(_01373_));
 sg13g2_mux2_1 _15649_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(net421),
    .X(_01374_));
 sg13g2_mux2_1 _15650_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(net421),
    .X(_01375_));
 sg13g2_mux2_1 _15651_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(net421),
    .X(_01376_));
 sg13g2_buf_1 _15652_ (.A(_08706_),
    .X(_08739_));
 sg13g2_mux2_1 _15653_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(net420),
    .X(_01377_));
 sg13g2_mux2_1 _15654_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(net420),
    .X(_01378_));
 sg13g2_mux2_1 _15655_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(net420),
    .X(_01379_));
 sg13g2_mux2_1 _15656_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(net420),
    .X(_01380_));
 sg13g2_mux2_1 _15657_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(net420),
    .X(_01381_));
 sg13g2_mux2_1 _15658_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_08739_),
    .X(_01382_));
 sg13g2_mux2_1 _15659_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_08739_),
    .X(_01383_));
 sg13g2_mux2_1 _15660_ (.A0(net10),
    .A1(\rbzero.tex_r0[63] ),
    .S(net420),
    .X(_01384_));
 sg13g2_mux2_1 _15661_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(net420),
    .X(_01385_));
 sg13g2_mux2_1 _15662_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(net420),
    .X(_01386_));
 sg13g2_mux2_1 _15663_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_08699_),
    .X(_01387_));
 sg13g2_mux2_1 _15664_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_08699_),
    .X(_01388_));
 sg13g2_mux2_1 _15665_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[0] ),
    .S(_08733_),
    .X(_01389_));
 sg13g2_mux2_1 _15666_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_08733_),
    .X(_01390_));
 sg13g2_buf_1 _15667_ (.A(_08719_),
    .X(_08740_));
 sg13g2_mux2_1 _15668_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(net419),
    .X(_01391_));
 sg13g2_mux2_1 _15669_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(net419),
    .X(_01392_));
 sg13g2_mux2_1 _15670_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_08740_),
    .X(_01393_));
 sg13g2_mux2_1 _15671_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_08740_),
    .X(_01394_));
 sg13g2_mux2_1 _15672_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(net419),
    .X(_01395_));
 sg13g2_mux2_1 _15673_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(net419),
    .X(_01396_));
 sg13g2_mux2_1 _15674_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(net419),
    .X(_01397_));
 sg13g2_mux2_1 _15675_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(net419),
    .X(_01398_));
 sg13g2_mux2_1 _15676_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(net419),
    .X(_01399_));
 sg13g2_mux2_1 _15677_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(net419),
    .X(_01400_));
 sg13g2_buf_1 _15678_ (.A(_08719_),
    .X(_08741_));
 sg13g2_mux2_1 _15679_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_08741_),
    .X(_01401_));
 sg13g2_mux2_1 _15680_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(net418),
    .X(_01402_));
 sg13g2_mux2_1 _15681_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(net418),
    .X(_01403_));
 sg13g2_mux2_1 _15682_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(net418),
    .X(_01404_));
 sg13g2_mux2_1 _15683_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(net418),
    .X(_01405_));
 sg13g2_mux2_1 _15684_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(net418),
    .X(_01406_));
 sg13g2_mux2_1 _15685_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_08741_),
    .X(_01407_));
 sg13g2_mux2_1 _15686_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(net418),
    .X(_01408_));
 sg13g2_mux2_1 _15687_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(net418),
    .X(_01409_));
 sg13g2_mux2_1 _15688_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(net418),
    .X(_01410_));
 sg13g2_buf_1 _15689_ (.A(_08719_),
    .X(_08742_));
 sg13g2_mux2_1 _15690_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(net417),
    .X(_01411_));
 sg13g2_mux2_1 _15691_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(net417),
    .X(_01412_));
 sg13g2_mux2_1 _15692_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(net417),
    .X(_01413_));
 sg13g2_mux2_1 _15693_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(net417),
    .X(_01414_));
 sg13g2_mux2_1 _15694_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(net417),
    .X(_01415_));
 sg13g2_mux2_1 _15695_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(net417),
    .X(_01416_));
 sg13g2_mux2_1 _15696_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(net417),
    .X(_01417_));
 sg13g2_mux2_1 _15697_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(net417),
    .X(_01418_));
 sg13g2_mux2_1 _15698_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_08742_),
    .X(_01419_));
 sg13g2_mux2_1 _15699_ (.A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_08742_),
    .X(_01420_));
 sg13g2_buf_1 _15700_ (.A(_08719_),
    .X(_08743_));
 sg13g2_mux2_1 _15701_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(net416),
    .X(_01421_));
 sg13g2_mux2_1 _15702_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_08743_),
    .X(_01422_));
 sg13g2_mux2_1 _15703_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(net416),
    .X(_01423_));
 sg13g2_mux2_1 _15704_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(net416),
    .X(_01424_));
 sg13g2_mux2_1 _15705_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(net416),
    .X(_01425_));
 sg13g2_mux2_1 _15706_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(net416),
    .X(_01426_));
 sg13g2_mux2_1 _15707_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(net416),
    .X(_01427_));
 sg13g2_mux2_1 _15708_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(net416),
    .X(_01428_));
 sg13g2_mux2_1 _15709_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_08743_),
    .X(_01429_));
 sg13g2_mux2_1 _15710_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(net416),
    .X(_01430_));
 sg13g2_buf_1 _15711_ (.A(_08719_),
    .X(_08744_));
 sg13g2_mux2_1 _15712_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(net415),
    .X(_01431_));
 sg13g2_mux2_1 _15713_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(net415),
    .X(_01432_));
 sg13g2_mux2_1 _15714_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(net415),
    .X(_01433_));
 sg13g2_mux2_1 _15715_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_08744_),
    .X(_01434_));
 sg13g2_mux2_1 _15716_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_08744_),
    .X(_01435_));
 sg13g2_mux2_1 _15717_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(net415),
    .X(_01436_));
 sg13g2_mux2_1 _15718_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(net415),
    .X(_01437_));
 sg13g2_mux2_1 _15719_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(net415),
    .X(_01438_));
 sg13g2_mux2_1 _15720_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(net415),
    .X(_01439_));
 sg13g2_mux2_1 _15721_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(net415),
    .X(_01440_));
 sg13g2_buf_1 _15722_ (.A(_08719_),
    .X(_08745_));
 sg13g2_mux2_1 _15723_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(net414),
    .X(_01441_));
 sg13g2_mux2_1 _15724_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_08745_),
    .X(_01442_));
 sg13g2_mux2_1 _15725_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_08745_),
    .X(_01443_));
 sg13g2_mux2_1 _15726_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(net414),
    .X(_01444_));
 sg13g2_mux2_1 _15727_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(net414),
    .X(_01445_));
 sg13g2_mux2_1 _15728_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(net414),
    .X(_01446_));
 sg13g2_mux2_1 _15729_ (.A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(net414),
    .X(_01447_));
 sg13g2_mux2_1 _15730_ (.A0(net10),
    .A1(\rbzero.tex_r1[63] ),
    .S(net414),
    .X(_01448_));
 sg13g2_mux2_1 _15731_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(net414),
    .X(_01449_));
 sg13g2_mux2_1 _15732_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(net414),
    .X(_01450_));
 sg13g2_mux2_1 _15733_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_08712_),
    .X(_01451_));
 sg13g2_mux2_1 _15734_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_08712_),
    .X(_01452_));
 sg13g2_buf_1 _15735_ (.A(_08411_),
    .X(_08746_));
 sg13g2_buf_1 _15736_ (.A(_08746_),
    .X(_08747_));
 sg13g2_buf_2 _15737_ (.A(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_08748_));
 sg13g2_buf_1 _15738_ (.A(_08680_),
    .X(_08749_));
 sg13g2_buf_2 _15739_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_08750_));
 sg13g2_inv_2 _15740_ (.Y(_08751_),
    .A(_08750_));
 sg13g2_buf_1 _15741_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_08752_));
 sg13g2_buf_1 _15742_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_08753_));
 sg13g2_inv_1 _15743_ (.Y(_08754_),
    .A(_08753_));
 sg13g2_inv_1 _15744_ (.Y(_08755_),
    .A(\rbzero.wall_tracer.rayAddendX[-5] ));
 sg13g2_buf_1 _15745_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_08756_));
 sg13g2_inv_1 _15746_ (.Y(_08757_),
    .A(_08756_));
 sg13g2_buf_1 _15747_ (.A(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_08758_));
 sg13g2_buf_1 _15748_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_08759_));
 sg13g2_a21oi_1 _15749_ (.A1(_08758_),
    .A2(net826),
    .Y(_08760_),
    .B1(\rbzero.wall_tracer.rayAddendX[-8] ));
 sg13g2_nand3_1 _15750_ (.B(_08758_),
    .C(net826),
    .A(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_08761_));
 sg13g2_o21ai_1 _15751_ (.B1(_08761_),
    .Y(_08762_),
    .A1(_08757_),
    .A2(_08760_));
 sg13g2_buf_1 _15752_ (.A(_08762_),
    .X(_08763_));
 sg13g2_nor2_1 _15753_ (.A(\rbzero.wall_tracer.rayAddendX[-7] ),
    .B(_08763_),
    .Y(_08764_));
 sg13g2_buf_1 _15754_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_08765_));
 sg13g2_a21oi_1 _15755_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_08763_),
    .Y(_08766_),
    .B1(_08765_));
 sg13g2_nor2_1 _15756_ (.A(_08764_),
    .B(_08766_),
    .Y(_08767_));
 sg13g2_buf_2 _15757_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_08768_));
 sg13g2_a21o_1 _15758_ (.A2(_08767_),
    .A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_08768_),
    .X(_08769_));
 sg13g2_o21ai_1 _15759_ (.B1(_08769_),
    .Y(_08770_),
    .A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_08767_));
 sg13g2_buf_1 _15760_ (.A(_08770_),
    .X(_08771_));
 sg13g2_inv_1 _15761_ (.Y(_08772_),
    .A(_08771_));
 sg13g2_buf_1 _15762_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_08773_));
 sg13g2_a21oi_1 _15763_ (.A1(\rbzero.wall_tracer.rayAddendX[-5] ),
    .A2(_08772_),
    .Y(_08774_),
    .B1(_08773_));
 sg13g2_a21oi_1 _15764_ (.A1(_08755_),
    .A2(_08771_),
    .Y(_08775_),
    .B1(_08774_));
 sg13g2_buf_2 _15765_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_08776_));
 sg13g2_a21o_1 _15766_ (.A2(_08775_),
    .A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B1(_08776_),
    .X(_08777_));
 sg13g2_o21ai_1 _15767_ (.B1(_08777_),
    .Y(_08778_),
    .A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_08775_));
 sg13g2_buf_1 _15768_ (.A(_08778_),
    .X(_08779_));
 sg13g2_inv_1 _15769_ (.Y(_08780_),
    .A(_08779_));
 sg13g2_buf_1 _15770_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_08781_));
 sg13g2_a21oi_1 _15771_ (.A1(_08753_),
    .A2(_08780_),
    .Y(_08782_),
    .B1(_08781_));
 sg13g2_a21oi_1 _15772_ (.A1(_08754_),
    .A2(_08779_),
    .Y(_08783_),
    .B1(_08782_));
 sg13g2_buf_1 _15773_ (.A(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_08784_));
 sg13g2_a21o_1 _15774_ (.A2(_08783_),
    .A1(_08752_),
    .B1(_08784_),
    .X(_08785_));
 sg13g2_o21ai_1 _15775_ (.B1(_08785_),
    .Y(_08786_),
    .A1(_08752_),
    .A2(_08783_));
 sg13g2_buf_1 _15776_ (.A(_08786_),
    .X(_08787_));
 sg13g2_xnor2_1 _15777_ (.Y(_08788_),
    .A(_08751_),
    .B(_08787_));
 sg13g2_nor2_1 _15778_ (.A(_08749_),
    .B(_08788_),
    .Y(_08789_));
 sg13g2_xnor2_1 _15779_ (.Y(_08790_),
    .A(_08748_),
    .B(_08789_));
 sg13g2_buf_1 _15780_ (.A(_08746_),
    .X(_08791_));
 sg13g2_buf_1 _15781_ (.A(_08773_),
    .X(_08792_));
 sg13g2_buf_1 _15782_ (.A(net782),
    .X(_08793_));
 sg13g2_buf_1 _15783_ (.A(_08756_),
    .X(_08794_));
 sg13g2_buf_1 _15784_ (.A(_08765_),
    .X(_08795_));
 sg13g2_nor3_1 _15785_ (.A(net781),
    .B(net780),
    .C(_08768_),
    .Y(_08796_));
 sg13g2_nor2_1 _15786_ (.A(net826),
    .B(_08796_),
    .Y(_08797_));
 sg13g2_xor2_1 _15787_ (.B(_08797_),
    .A(net722),
    .X(_08798_));
 sg13g2_nand2_1 _15788_ (.Y(_08799_),
    .A(net679),
    .B(_08798_));
 sg13g2_o21ai_1 _15789_ (.B1(_08799_),
    .Y(_01558_),
    .A1(net680),
    .A2(_08790_));
 sg13g2_buf_2 _15790_ (.A(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_08800_));
 sg13g2_buf_1 _15791_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_08801_));
 sg13g2_inv_1 _15792_ (.Y(_08802_),
    .A(_08787_));
 sg13g2_a21oi_1 _15793_ (.A1(_08750_),
    .A2(_08802_),
    .Y(_08803_),
    .B1(_08748_));
 sg13g2_a21oi_1 _15794_ (.A1(_08751_),
    .A2(_08787_),
    .Y(_08804_),
    .B1(_08803_));
 sg13g2_and2_1 _15795_ (.A(_08801_),
    .B(_08804_),
    .X(_08805_));
 sg13g2_and2_1 _15796_ (.A(\rbzero.wall_tracer.state[8] ),
    .B(net490),
    .X(_08806_));
 sg13g2_buf_1 _15797_ (.A(_08806_),
    .X(_08807_));
 sg13g2_buf_1 _15798_ (.A(_08807_),
    .X(_08808_));
 sg13g2_or2_1 _15799_ (.X(_08809_),
    .B(_08804_),
    .A(_08801_));
 sg13g2_nand3b_1 _15800_ (.B(net462),
    .C(_08809_),
    .Y(_08810_),
    .A_N(_08805_));
 sg13g2_xor2_1 _15801_ (.B(_08810_),
    .A(_08800_),
    .X(_08811_));
 sg13g2_buf_1 _15802_ (.A(_08776_),
    .X(_08812_));
 sg13g2_inv_1 _15803_ (.Y(_08813_),
    .A(net780));
 sg13g2_buf_1 _15804_ (.A(_08768_),
    .X(_08814_));
 sg13g2_buf_1 _15805_ (.A(net826),
    .X(_08815_));
 sg13g2_o21ai_1 _15806_ (.B1(_08757_),
    .Y(_08816_),
    .A1(net778),
    .A2(net777));
 sg13g2_buf_1 _15807_ (.A(_00060_),
    .X(_08817_));
 sg13g2_nand2_1 _15808_ (.Y(_08818_),
    .A(_08817_),
    .B(net778));
 sg13g2_a22oi_1 _15809_ (.Y(_08819_),
    .B1(_08818_),
    .B2(net781),
    .A2(_08816_),
    .A1(_08813_));
 sg13g2_nor2b_1 _15810_ (.A(net781),
    .B_N(net777),
    .Y(_08820_));
 sg13g2_nor2_1 _15811_ (.A(_08757_),
    .B(net777),
    .Y(_08821_));
 sg13g2_a21oi_1 _15812_ (.A1(net722),
    .A2(_08820_),
    .Y(_08822_),
    .B1(_08821_));
 sg13g2_o21ai_1 _15813_ (.B1(_08822_),
    .Y(_08823_),
    .A1(net722),
    .A2(_08819_));
 sg13g2_xnor2_1 _15814_ (.Y(_08824_),
    .A(net779),
    .B(_08823_));
 sg13g2_nor2_1 _15815_ (.A(net544),
    .B(_08824_),
    .Y(_08825_));
 sg13g2_a21oi_1 _15816_ (.A1(net545),
    .A2(_08811_),
    .Y(_01559_),
    .B1(_08825_));
 sg13g2_buf_2 _15817_ (.A(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_08826_));
 sg13g2_a21oi_2 _15818_ (.B1(_08805_),
    .Y(_08827_),
    .A2(_08809_),
    .A1(_08800_));
 sg13g2_nor2_1 _15819_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(_08827_),
    .Y(_08828_));
 sg13g2_inv_1 _15820_ (.Y(_08829_),
    .A(_08828_));
 sg13g2_buf_1 _15821_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_08830_));
 sg13g2_buf_1 _15822_ (.A(net825),
    .X(_08831_));
 sg13g2_nand2_1 _15823_ (.Y(_08832_),
    .A(net776),
    .B(_08827_));
 sg13g2_a21oi_1 _15824_ (.A1(_08829_),
    .A2(_08832_),
    .Y(_08833_),
    .B1(_08749_));
 sg13g2_xnor2_1 _15825_ (.Y(_08834_),
    .A(_08826_),
    .B(_08833_));
 sg13g2_nand2_1 _15826_ (.Y(_08835_),
    .A(net781),
    .B(_08776_));
 sg13g2_nor2_1 _15827_ (.A(_08756_),
    .B(_08776_),
    .Y(_08836_));
 sg13g2_buf_2 _15828_ (.A(_08836_),
    .X(_08837_));
 sg13g2_o21ai_1 _15829_ (.B1(net826),
    .Y(_08838_),
    .A1(net782),
    .A2(_08837_));
 sg13g2_nor3_1 _15830_ (.A(_08765_),
    .B(_08768_),
    .C(_08773_),
    .Y(_08839_));
 sg13g2_nand2b_1 _15831_ (.Y(_08840_),
    .B(_08837_),
    .A_N(_08839_));
 sg13g2_nand3_1 _15832_ (.B(_08838_),
    .C(_08840_),
    .A(_08835_),
    .Y(_08841_));
 sg13g2_xnor2_1 _15833_ (.Y(_08842_),
    .A(_08765_),
    .B(_08753_));
 sg13g2_xnor2_1 _15834_ (.Y(_08843_),
    .A(_08837_),
    .B(_08842_));
 sg13g2_xnor2_1 _15835_ (.Y(_08844_),
    .A(_08841_),
    .B(_08843_));
 sg13g2_nor2_1 _15836_ (.A(net544),
    .B(_08844_),
    .Y(_08845_));
 sg13g2_a21oi_1 _15837_ (.A1(net545),
    .A2(_08834_),
    .Y(_01560_),
    .B1(_08845_));
 sg13g2_buf_2 _15838_ (.A(\rbzero.wall_tracer.rayAddendX[2] ),
    .X(_08846_));
 sg13g2_nor2_1 _15839_ (.A(_08826_),
    .B(_08832_),
    .Y(_08847_));
 sg13g2_a21oi_1 _15840_ (.A1(_08826_),
    .A2(_08828_),
    .Y(_08848_),
    .B1(_08847_));
 sg13g2_nor2_1 _15841_ (.A(net463),
    .B(_08848_),
    .Y(_08849_));
 sg13g2_xnor2_1 _15842_ (.Y(_08850_),
    .A(_08846_),
    .B(_08849_));
 sg13g2_o21ai_1 _15843_ (.B1(_08776_),
    .Y(_08851_),
    .A1(net782),
    .A2(net826));
 sg13g2_nor3_1 _15844_ (.A(net782),
    .B(_08776_),
    .C(net826),
    .Y(_08852_));
 sg13g2_a21oi_1 _15845_ (.A1(_08757_),
    .A2(_08851_),
    .Y(_08853_),
    .B1(_08852_));
 sg13g2_nor2_1 _15846_ (.A(_08842_),
    .B(_08853_),
    .Y(_08854_));
 sg13g2_nor2_1 _15847_ (.A(_08792_),
    .B(net826),
    .Y(_08855_));
 sg13g2_nand2_1 _15848_ (.Y(_08856_),
    .A(_08817_),
    .B(_08796_));
 sg13g2_and2_1 _15849_ (.A(net781),
    .B(_08776_),
    .X(_08857_));
 sg13g2_and2_1 _15850_ (.A(net782),
    .B(_08759_),
    .X(_08858_));
 sg13g2_nor4_1 _15851_ (.A(_08858_),
    .B(_08857_),
    .C(_08837_),
    .D(_08855_),
    .Y(_08859_));
 sg13g2_a21oi_1 _15852_ (.A1(_08857_),
    .A2(_08855_),
    .Y(_08860_),
    .B1(_08859_));
 sg13g2_nand2_1 _15853_ (.Y(_08861_),
    .A(_08837_),
    .B(_08855_));
 sg13g2_mux2_1 _15854_ (.A0(_08860_),
    .A1(_08861_),
    .S(_08842_),
    .X(_08862_));
 sg13g2_a21oi_1 _15855_ (.A1(_08855_),
    .A2(_08856_),
    .Y(_08863_),
    .B1(_08862_));
 sg13g2_nor2_1 _15856_ (.A(_08854_),
    .B(_08863_),
    .Y(_08864_));
 sg13g2_buf_1 _15857_ (.A(_08753_),
    .X(_08865_));
 sg13g2_nor2_1 _15858_ (.A(net780),
    .B(net775),
    .Y(_08866_));
 sg13g2_buf_1 _15859_ (.A(_08866_),
    .X(_08867_));
 sg13g2_xnor2_1 _15860_ (.Y(_08868_),
    .A(_08768_),
    .B(_08752_));
 sg13g2_xnor2_1 _15861_ (.Y(_08869_),
    .A(_08867_),
    .B(_08868_));
 sg13g2_xnor2_1 _15862_ (.Y(_08870_),
    .A(_08864_),
    .B(_08869_));
 sg13g2_nand2_1 _15863_ (.Y(_08871_),
    .A(net679),
    .B(_08870_));
 sg13g2_o21ai_1 _15864_ (.B1(_08871_),
    .Y(_01561_),
    .A1(net680),
    .A2(_08850_));
 sg13g2_buf_2 _15865_ (.A(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_08872_));
 sg13g2_inv_1 _15866_ (.Y(_08873_),
    .A(_08846_));
 sg13g2_inv_1 _15867_ (.Y(_08874_),
    .A(net825));
 sg13g2_o21ai_1 _15868_ (.B1(net774),
    .Y(_08875_),
    .A1(_08873_),
    .A2(_08827_));
 sg13g2_a21oi_1 _15869_ (.A1(_08873_),
    .A2(_08827_),
    .Y(_08876_),
    .B1(net774));
 sg13g2_a21o_1 _15870_ (.A2(_08875_),
    .A1(_08826_),
    .B1(_08876_),
    .X(_08877_));
 sg13g2_buf_1 _15871_ (.A(_08877_),
    .X(_08878_));
 sg13g2_xnor2_1 _15872_ (.Y(_08879_),
    .A(net776),
    .B(_08878_));
 sg13g2_nor2_1 _15873_ (.A(net463),
    .B(_08879_),
    .Y(_08880_));
 sg13g2_xnor2_1 _15874_ (.Y(_08881_),
    .A(_08872_),
    .B(_08880_));
 sg13g2_inv_1 _15875_ (.Y(_08882_),
    .A(_08868_));
 sg13g2_a21oi_1 _15876_ (.A1(_08835_),
    .A2(_08838_),
    .Y(_08883_),
    .B1(_08837_));
 sg13g2_nand4_1 _15877_ (.B(_08837_),
    .C(_08838_),
    .A(_08835_),
    .Y(_08884_),
    .D(_08840_));
 sg13g2_o21ai_1 _15878_ (.B1(_08884_),
    .Y(_08885_),
    .A1(net775),
    .A2(_08883_));
 sg13g2_a21o_1 _15879_ (.A2(_08884_),
    .A1(_08868_),
    .B1(net775),
    .X(_08886_));
 sg13g2_o21ai_1 _15880_ (.B1(_08886_),
    .Y(_08887_),
    .A1(_08868_),
    .A2(_08883_));
 sg13g2_a22oi_1 _15881_ (.Y(_08888_),
    .B1(_08887_),
    .B2(_08813_),
    .A2(_08885_),
    .A1(_08882_));
 sg13g2_buf_1 _15882_ (.A(_08888_),
    .X(_08889_));
 sg13g2_buf_1 _15883_ (.A(_08752_),
    .X(_08890_));
 sg13g2_nor2_1 _15884_ (.A(_08768_),
    .B(net773),
    .Y(_08891_));
 sg13g2_nand2_1 _15885_ (.Y(_08892_),
    .A(net782),
    .B(_08751_));
 sg13g2_nand2b_1 _15886_ (.Y(_08893_),
    .B(_08750_),
    .A_N(net782));
 sg13g2_nand2_2 _15887_ (.Y(_08894_),
    .A(_08892_),
    .B(_08893_));
 sg13g2_xor2_1 _15888_ (.B(_08894_),
    .A(_08891_),
    .X(_08895_));
 sg13g2_xnor2_1 _15889_ (.Y(_08896_),
    .A(_08889_),
    .B(_08895_));
 sg13g2_nand2_1 _15890_ (.Y(_08897_),
    .A(net679),
    .B(_08896_));
 sg13g2_o21ai_1 _15891_ (.B1(_08897_),
    .Y(_01562_),
    .A1(net680),
    .A2(_08881_));
 sg13g2_buf_1 _15892_ (.A(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_08898_));
 sg13g2_inv_1 _15893_ (.Y(_08899_),
    .A(_08898_));
 sg13g2_nand2_1 _15894_ (.Y(_08900_),
    .A(_08873_),
    .B(net825));
 sg13g2_nor2_1 _15895_ (.A(_08872_),
    .B(_08900_),
    .Y(_08901_));
 sg13g2_inv_1 _15896_ (.Y(_08902_),
    .A(_08872_));
 sg13g2_nor2_1 _15897_ (.A(_08902_),
    .B(net776),
    .Y(_08903_));
 sg13g2_o21ai_1 _15898_ (.B1(_08900_),
    .Y(_08904_),
    .A1(_08873_),
    .A2(_08829_));
 sg13g2_nand2_1 _15899_ (.Y(_08905_),
    .A(_08826_),
    .B(_08904_));
 sg13g2_o21ai_1 _15900_ (.B1(_08905_),
    .Y(_08906_),
    .A1(_08827_),
    .A2(_08900_));
 sg13g2_mux2_1 _15901_ (.A0(_08901_),
    .A1(_08903_),
    .S(_08906_),
    .X(_08907_));
 sg13g2_nand2_1 _15902_ (.Y(_08908_),
    .A(net462),
    .B(_08907_));
 sg13g2_xnor2_1 _15903_ (.Y(_08909_),
    .A(_08899_),
    .B(_08908_));
 sg13g2_and2_1 _15904_ (.A(_08867_),
    .B(_08891_),
    .X(_08910_));
 sg13g2_buf_1 _15905_ (.A(_08750_),
    .X(_08911_));
 sg13g2_nor2_1 _15906_ (.A(_08792_),
    .B(_08750_),
    .Y(_08912_));
 sg13g2_buf_1 _15907_ (.A(_08912_),
    .X(_08913_));
 sg13g2_nor2b_1 _15908_ (.A(_08797_),
    .B_N(_08913_),
    .Y(_08914_));
 sg13g2_a21o_1 _15909_ (.A2(net772),
    .A1(net722),
    .B1(_08914_),
    .X(_08915_));
 sg13g2_o21ai_1 _15910_ (.B1(_08892_),
    .Y(_08916_),
    .A1(_08797_),
    .A2(_08893_));
 sg13g2_o21ai_1 _15911_ (.B1(net773),
    .Y(_08917_),
    .A1(net780),
    .A2(net775));
 sg13g2_inv_1 _15912_ (.Y(_08918_),
    .A(net773));
 sg13g2_nand2_1 _15913_ (.Y(_08919_),
    .A(_08918_),
    .B(_08867_));
 sg13g2_nand3_1 _15914_ (.B(_08917_),
    .C(_08919_),
    .A(net778),
    .Y(_08920_));
 sg13g2_o21ai_1 _15915_ (.B1(_08920_),
    .Y(_08921_),
    .A1(net778),
    .A2(_08917_));
 sg13g2_a22oi_1 _15916_ (.Y(_08922_),
    .B1(_08916_),
    .B2(_08921_),
    .A2(_08915_),
    .A1(_08910_));
 sg13g2_nor2_1 _15917_ (.A(_08854_),
    .B(_08867_),
    .Y(_08923_));
 sg13g2_a21oi_1 _15918_ (.A1(net773),
    .A2(_08923_),
    .Y(_08924_),
    .B1(net778));
 sg13g2_nor2_1 _15919_ (.A(net773),
    .B(_08923_),
    .Y(_08925_));
 sg13g2_o21ai_1 _15920_ (.B1(_08894_),
    .Y(_08926_),
    .A1(_08924_),
    .A2(_08925_));
 sg13g2_o21ai_1 _15921_ (.B1(_08926_),
    .Y(_08927_),
    .A1(_08862_),
    .A2(_08922_));
 sg13g2_buf_1 _15922_ (.A(_08801_),
    .X(_08928_));
 sg13g2_xor2_1 _15923_ (.B(net771),
    .A(_08776_),
    .X(_08929_));
 sg13g2_xnor2_1 _15924_ (.Y(_08930_),
    .A(_08913_),
    .B(_08929_));
 sg13g2_xnor2_1 _15925_ (.Y(_08931_),
    .A(_08927_),
    .B(_08930_));
 sg13g2_nand2_1 _15926_ (.Y(_08932_),
    .A(net679),
    .B(_08931_));
 sg13g2_o21ai_1 _15927_ (.B1(_08932_),
    .Y(_01563_),
    .A1(net680),
    .A2(_08909_));
 sg13g2_buf_2 _15928_ (.A(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_08933_));
 sg13g2_nand3_1 _15929_ (.B(_08878_),
    .C(_08903_),
    .A(net824),
    .Y(_08934_));
 sg13g2_or4_1 _15930_ (.A(_08872_),
    .B(net824),
    .C(net774),
    .D(_08878_),
    .X(_08935_));
 sg13g2_a21oi_1 _15931_ (.A1(_08934_),
    .A2(_08935_),
    .Y(_08936_),
    .B1(_08680_));
 sg13g2_xnor2_1 _15932_ (.Y(_08937_),
    .A(_08933_),
    .B(_08936_));
 sg13g2_or2_1 _15933_ (.X(_08938_),
    .B(_08889_),
    .A(net772));
 sg13g2_a21o_1 _15934_ (.A2(_08889_),
    .A1(net772),
    .B1(net722),
    .X(_08939_));
 sg13g2_inv_1 _15935_ (.Y(_08940_),
    .A(_08929_));
 sg13g2_a21oi_1 _15936_ (.A1(_08938_),
    .A2(_08939_),
    .Y(_08941_),
    .B1(_08940_));
 sg13g2_a21oi_1 _15937_ (.A1(_08940_),
    .A2(_08938_),
    .Y(_08942_),
    .B1(_08793_));
 sg13g2_a21oi_1 _15938_ (.A1(net772),
    .A2(_08889_),
    .Y(_08943_),
    .B1(_08940_));
 sg13g2_o21ai_1 _15939_ (.B1(_08891_),
    .Y(_08944_),
    .A1(_08942_),
    .A2(_08943_));
 sg13g2_nand2b_1 _15940_ (.Y(_08945_),
    .B(_08944_),
    .A_N(_08941_));
 sg13g2_buf_1 _15941_ (.A(_08945_),
    .X(_08946_));
 sg13g2_nor2_2 _15942_ (.A(net779),
    .B(net771),
    .Y(_08947_));
 sg13g2_xor2_1 _15943_ (.B(net825),
    .A(net775),
    .X(_08948_));
 sg13g2_buf_1 _15944_ (.A(_08948_),
    .X(_08949_));
 sg13g2_xnor2_1 _15945_ (.Y(_08950_),
    .A(_08947_),
    .B(_08949_));
 sg13g2_xnor2_1 _15946_ (.Y(_08951_),
    .A(_08946_),
    .B(_08950_));
 sg13g2_nand2_1 _15947_ (.Y(_08952_),
    .A(_08791_),
    .B(_08951_));
 sg13g2_o21ai_1 _15948_ (.B1(_08952_),
    .Y(_01564_),
    .A1(net680),
    .A2(_08937_));
 sg13g2_buf_2 _15949_ (.A(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_08953_));
 sg13g2_nor4_1 _15950_ (.A(_08846_),
    .B(net824),
    .C(_08933_),
    .D(_08906_),
    .Y(_08954_));
 sg13g2_nand2b_1 _15951_ (.Y(_08955_),
    .B(_08830_),
    .A_N(_08954_));
 sg13g2_nand3_1 _15952_ (.B(_08933_),
    .C(_08906_),
    .A(net824),
    .Y(_08956_));
 sg13g2_a22oi_1 _15953_ (.Y(_08957_),
    .B1(_08956_),
    .B2(_08874_),
    .A2(_08955_),
    .A1(_08902_));
 sg13g2_xnor2_1 _15954_ (.Y(_08958_),
    .A(net776),
    .B(_08957_));
 sg13g2_nor2_1 _15955_ (.A(net463),
    .B(_08958_),
    .Y(_08959_));
 sg13g2_xnor2_1 _15956_ (.Y(_08960_),
    .A(_08953_),
    .B(_08959_));
 sg13g2_inv_1 _15957_ (.Y(_08961_),
    .A(net771));
 sg13g2_nand2b_1 _15958_ (.Y(_08962_),
    .B(_08864_),
    .A_N(_08867_));
 sg13g2_nor2b_1 _15959_ (.A(_08864_),
    .B_N(_08867_),
    .Y(_08963_));
 sg13g2_or2_1 _15960_ (.X(_08964_),
    .B(_08963_),
    .A(_08894_));
 sg13g2_a22oi_1 _15961_ (.Y(_08965_),
    .B1(_08964_),
    .B2(_08918_),
    .A2(_08962_),
    .A1(_08894_));
 sg13g2_and2_1 _15962_ (.A(_08918_),
    .B(_08962_),
    .X(_08966_));
 sg13g2_o21ai_1 _15963_ (.B1(_08894_),
    .Y(_08967_),
    .A1(_08963_),
    .A2(_08966_));
 sg13g2_o21ai_1 _15964_ (.B1(_08967_),
    .Y(_08968_),
    .A1(_08814_),
    .A2(_08965_));
 sg13g2_or2_1 _15965_ (.X(_08969_),
    .B(_08968_),
    .A(_08913_));
 sg13g2_and2_1 _15966_ (.A(_08913_),
    .B(_08968_),
    .X(_08970_));
 sg13g2_a21o_1 _15967_ (.A2(_08969_),
    .A1(_08961_),
    .B1(_08970_),
    .X(_08971_));
 sg13g2_o21ai_1 _15968_ (.B1(_08961_),
    .Y(_08972_),
    .A1(_08949_),
    .A2(_08970_));
 sg13g2_nand2_1 _15969_ (.Y(_08973_),
    .A(_08949_),
    .B(_08969_));
 sg13g2_a21oi_1 _15970_ (.A1(_08972_),
    .A2(_08973_),
    .Y(_08974_),
    .B1(net779));
 sg13g2_a21oi_1 _15971_ (.A1(_08949_),
    .A2(_08971_),
    .Y(_08975_),
    .B1(_08974_));
 sg13g2_nor2_1 _15972_ (.A(_08754_),
    .B(net776),
    .Y(_08976_));
 sg13g2_xnor2_1 _15973_ (.Y(_08977_),
    .A(net773),
    .B(_08976_));
 sg13g2_xnor2_1 _15974_ (.Y(_08978_),
    .A(_08975_),
    .B(_08977_));
 sg13g2_nand2_1 _15975_ (.Y(_08979_),
    .A(_08791_),
    .B(_08978_));
 sg13g2_o21ai_1 _15976_ (.B1(_08979_),
    .Y(_01565_),
    .A1(net680),
    .A2(_08960_));
 sg13g2_buf_2 _15977_ (.A(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_08980_));
 sg13g2_buf_1 _15978_ (.A(_08680_),
    .X(_08981_));
 sg13g2_nand4_1 _15979_ (.B(_08933_),
    .C(_08953_),
    .A(net824),
    .Y(_08982_),
    .D(_08878_));
 sg13g2_or4_1 _15980_ (.A(net824),
    .B(_08933_),
    .C(_08953_),
    .D(_08878_),
    .X(_08983_));
 sg13g2_a21oi_1 _15981_ (.A1(_08830_),
    .A2(_08983_),
    .Y(_08984_),
    .B1(_08872_));
 sg13g2_a21oi_2 _15982_ (.B1(_08984_),
    .Y(_08985_),
    .A2(_08982_),
    .A1(net774));
 sg13g2_xnor2_1 _15983_ (.Y(_08986_),
    .A(net776),
    .B(_08985_));
 sg13g2_nor2_1 _15984_ (.A(_08981_),
    .B(_08986_),
    .Y(_08987_));
 sg13g2_xnor2_1 _15985_ (.Y(_08988_),
    .A(_08980_),
    .B(_08987_));
 sg13g2_nor2_1 _15986_ (.A(net775),
    .B(_08890_),
    .Y(_08989_));
 sg13g2_inv_1 _15987_ (.Y(_08990_),
    .A(_08946_));
 sg13g2_o21ai_1 _15988_ (.B1(_08947_),
    .Y(_08991_),
    .A1(net825),
    .A2(_08946_));
 sg13g2_o21ai_1 _15989_ (.B1(_08991_),
    .Y(_08992_),
    .A1(net774),
    .A2(_08990_));
 sg13g2_nor4_1 _15990_ (.A(_08754_),
    .B(_08918_),
    .C(net825),
    .D(_08947_),
    .Y(_08993_));
 sg13g2_a22oi_1 _15991_ (.Y(_08994_),
    .B1(_08993_),
    .B2(_08990_),
    .A2(_08992_),
    .A1(_08989_));
 sg13g2_xnor2_1 _15992_ (.Y(_08995_),
    .A(_08751_),
    .B(_08994_));
 sg13g2_nor2_1 _15993_ (.A(_08693_),
    .B(_08995_),
    .Y(_08996_));
 sg13g2_a21oi_1 _15994_ (.A1(net545),
    .A2(_08988_),
    .Y(_01566_),
    .B1(_08996_));
 sg13g2_buf_1 _15995_ (.A(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_08997_));
 sg13g2_nor2b_1 _15996_ (.A(net776),
    .B_N(_08980_),
    .Y(_08998_));
 sg13g2_nand3_1 _15997_ (.B(_08957_),
    .C(_08998_),
    .A(_08953_),
    .Y(_08999_));
 sg13g2_nand2b_1 _15998_ (.Y(_09000_),
    .B(net825),
    .A_N(_08980_));
 sg13g2_or3_1 _15999_ (.A(_08953_),
    .B(_08957_),
    .C(_09000_),
    .X(_09001_));
 sg13g2_a21oi_1 _16000_ (.A1(_08999_),
    .A2(_09001_),
    .Y(_09002_),
    .B1(net463));
 sg13g2_xnor2_1 _16001_ (.Y(_09003_),
    .A(net823),
    .B(_09002_));
 sg13g2_nand2_1 _16002_ (.Y(_09004_),
    .A(_08961_),
    .B(_08913_));
 sg13g2_o21ai_1 _16003_ (.B1(net771),
    .Y(_09005_),
    .A1(net782),
    .A2(_08750_));
 sg13g2_nand2b_1 _16004_ (.Y(_09006_),
    .B(_09005_),
    .A_N(net779));
 sg13g2_and2_1 _16005_ (.A(_09004_),
    .B(_09006_),
    .X(_09007_));
 sg13g2_nand2_1 _16006_ (.Y(_09008_),
    .A(_08913_),
    .B(_08947_));
 sg13g2_nand3_1 _16007_ (.B(_09004_),
    .C(_09005_),
    .A(net779),
    .Y(_09009_));
 sg13g2_o21ai_1 _16008_ (.B1(_09009_),
    .Y(_09010_),
    .A1(net779),
    .A2(_09005_));
 sg13g2_nand2_1 _16009_ (.Y(_09011_),
    .A(_08949_),
    .B(_09010_));
 sg13g2_o21ai_1 _16010_ (.B1(_09011_),
    .Y(_09012_),
    .A1(_08949_),
    .A2(_09008_));
 sg13g2_nand3_1 _16011_ (.B(net780),
    .C(net778),
    .A(net781),
    .Y(_09013_));
 sg13g2_nand2b_1 _16012_ (.Y(_09014_),
    .B(_09013_),
    .A_N(_08793_));
 sg13g2_nand4_1 _16013_ (.B(net777),
    .C(_08926_),
    .A(_08817_),
    .Y(_09015_),
    .D(_09014_));
 sg13g2_nand3_1 _16014_ (.B(_09012_),
    .C(_09015_),
    .A(_08927_),
    .Y(_09016_));
 sg13g2_o21ai_1 _16015_ (.B1(_09016_),
    .Y(_09017_),
    .A1(net774),
    .A2(_09007_));
 sg13g2_nand2_1 _16016_ (.Y(_09018_),
    .A(_08989_),
    .B(_09017_));
 sg13g2_nand3_1 _16017_ (.B(_08993_),
    .C(_09016_),
    .A(net772),
    .Y(_09019_));
 sg13g2_o21ai_1 _16018_ (.B1(_09019_),
    .Y(_09020_),
    .A1(net772),
    .A2(_09018_));
 sg13g2_xnor2_1 _16019_ (.Y(_09021_),
    .A(net771),
    .B(_09020_));
 sg13g2_nor2_1 _16020_ (.A(_08693_),
    .B(_09021_),
    .Y(_09022_));
 sg13g2_a21oi_1 _16021_ (.A1(net545),
    .A2(_09003_),
    .Y(_01567_),
    .B1(_09022_));
 sg13g2_buf_2 _16022_ (.A(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_09023_));
 sg13g2_or2_1 _16023_ (.X(_09024_),
    .B(_09000_),
    .A(net823));
 sg13g2_or2_1 _16024_ (.X(_09025_),
    .B(_09024_),
    .A(_08985_));
 sg13g2_nand3_1 _16025_ (.B(_08985_),
    .C(_08998_),
    .A(net823),
    .Y(_09026_));
 sg13g2_a21oi_1 _16026_ (.A1(_09025_),
    .A2(_09026_),
    .Y(_09027_),
    .B1(_08680_));
 sg13g2_xnor2_1 _16027_ (.Y(_09028_),
    .A(_09023_),
    .B(_09027_));
 sg13g2_nand4_1 _16028_ (.B(_08911_),
    .C(net771),
    .A(_08865_),
    .Y(_09029_),
    .D(_08990_));
 sg13g2_a21o_1 _16029_ (.A2(_09029_),
    .A1(net774),
    .B1(_08918_),
    .X(_09030_));
 sg13g2_nor3_1 _16030_ (.A(_08865_),
    .B(_08911_),
    .C(_08928_),
    .Y(_09031_));
 sg13g2_o21ai_1 _16031_ (.B1(_09031_),
    .Y(_09032_),
    .A1(_08946_),
    .A2(_08947_));
 sg13g2_nand3_1 _16032_ (.B(_08961_),
    .C(_08989_),
    .A(_08751_),
    .Y(_09033_));
 sg13g2_nor4_1 _16033_ (.A(_08812_),
    .B(_08928_),
    .C(_08831_),
    .D(_09033_),
    .Y(_09034_));
 sg13g2_a22oi_1 _16034_ (.Y(_09035_),
    .B1(_09034_),
    .B2(_08946_),
    .A2(_09032_),
    .A1(net776));
 sg13g2_nand3_1 _16035_ (.B(_09030_),
    .C(_09035_),
    .A(net729),
    .Y(_09036_));
 sg13g2_o21ai_1 _16036_ (.B1(_09036_),
    .Y(_01568_),
    .A1(net680),
    .A2(_09028_));
 sg13g2_buf_2 _16037_ (.A(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(_09037_));
 sg13g2_or3_1 _16038_ (.A(_09023_),
    .B(_08985_),
    .C(_09024_),
    .X(_09038_));
 sg13g2_nand4_1 _16039_ (.B(_09023_),
    .C(_08985_),
    .A(net823),
    .Y(_09039_),
    .D(_08998_));
 sg13g2_a21oi_1 _16040_ (.A1(_09038_),
    .A2(_09039_),
    .Y(_09040_),
    .B1(net463));
 sg13g2_xnor2_1 _16041_ (.Y(_09041_),
    .A(_09037_),
    .B(_09040_));
 sg13g2_or2_1 _16042_ (.X(_09042_),
    .B(_09033_),
    .A(_08975_));
 sg13g2_buf_1 _16043_ (.A(_08640_),
    .X(_09043_));
 sg13g2_a21oi_1 _16044_ (.A1(net774),
    .A2(_09042_),
    .Y(_09044_),
    .B1(net609));
 sg13g2_a21oi_1 _16045_ (.A1(_08642_),
    .A2(_09041_),
    .Y(_01569_),
    .B1(_09044_));
 sg13g2_nand2_1 _16046_ (.Y(_09045_),
    .A(net777),
    .B(net462));
 sg13g2_xor2_1 _16047_ (.B(_09045_),
    .A(_08758_),
    .X(_09046_));
 sg13g2_nor2_1 _16048_ (.A(net686),
    .B(_09046_),
    .Y(_01570_));
 sg13g2_nand2_1 _16049_ (.Y(_09047_),
    .A(_08758_),
    .B(net777));
 sg13g2_xnor2_1 _16050_ (.Y(_09048_),
    .A(_08757_),
    .B(_09047_));
 sg13g2_nor2_1 _16051_ (.A(net461),
    .B(_09048_),
    .Y(_09049_));
 sg13g2_xnor2_1 _16052_ (.Y(_09050_),
    .A(\rbzero.wall_tracer.rayAddendX[-8] ),
    .B(_09049_));
 sg13g2_nor2_1 _16053_ (.A(net686),
    .B(_09050_),
    .Y(_01571_));
 sg13g2_buf_1 _16054_ (.A(net729),
    .X(_09051_));
 sg13g2_xnor2_1 _16055_ (.Y(_09052_),
    .A(net780),
    .B(_08763_));
 sg13g2_nor2_1 _16056_ (.A(net461),
    .B(_09052_),
    .Y(_09053_));
 sg13g2_xnor2_1 _16057_ (.Y(_09054_),
    .A(\rbzero.wall_tracer.rayAddendX[-7] ),
    .B(_09053_));
 sg13g2_nor2_1 _16058_ (.A(net678),
    .B(_09054_),
    .Y(_01572_));
 sg13g2_xnor2_1 _16059_ (.Y(_09055_),
    .A(net778),
    .B(_08767_));
 sg13g2_nor2_1 _16060_ (.A(net461),
    .B(_09055_),
    .Y(_09056_));
 sg13g2_xnor2_1 _16061_ (.Y(_09057_),
    .A(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B(_09056_));
 sg13g2_nor2_1 _16062_ (.A(net678),
    .B(_09057_),
    .Y(_01573_));
 sg13g2_buf_1 _16063_ (.A(_08746_),
    .X(_09058_));
 sg13g2_xor2_1 _16064_ (.B(_08771_),
    .A(net722),
    .X(_09059_));
 sg13g2_nor2_1 _16065_ (.A(net463),
    .B(_09059_),
    .Y(_09060_));
 sg13g2_xnor2_1 _16066_ (.Y(_09061_),
    .A(\rbzero.wall_tracer.rayAddendX[-5] ),
    .B(_09060_));
 sg13g2_nand2_1 _16067_ (.Y(_09062_),
    .A(net777),
    .B(net729));
 sg13g2_o21ai_1 _16068_ (.B1(_09062_),
    .Y(_01574_),
    .A1(net677),
    .A2(_09061_));
 sg13g2_buf_1 _16069_ (.A(_08680_),
    .X(_09063_));
 sg13g2_xnor2_1 _16070_ (.Y(_09064_),
    .A(_08812_),
    .B(_08775_));
 sg13g2_nor2_1 _16071_ (.A(net460),
    .B(_09064_),
    .Y(_09065_));
 sg13g2_xnor2_1 _16072_ (.Y(_09066_),
    .A(\rbzero.wall_tracer.rayAddendX[-4] ),
    .B(_09065_));
 sg13g2_o21ai_1 _16073_ (.B1(net729),
    .Y(_09067_),
    .A1(_08820_),
    .A2(_08821_));
 sg13g2_o21ai_1 _16074_ (.B1(_09067_),
    .Y(_01575_),
    .A1(net677),
    .A2(_09066_));
 sg13g2_xnor2_1 _16075_ (.Y(_09068_),
    .A(_08754_),
    .B(_08779_));
 sg13g2_nor2_1 _16076_ (.A(net460),
    .B(_09068_),
    .Y(_09069_));
 sg13g2_xnor2_1 _16077_ (.Y(_09070_),
    .A(_08781_),
    .B(_09069_));
 sg13g2_buf_1 _16078_ (.A(_08746_),
    .X(_09071_));
 sg13g2_nor2_1 _16079_ (.A(_08794_),
    .B(net777),
    .Y(_09072_));
 sg13g2_xnor2_1 _16080_ (.Y(_09073_),
    .A(_08795_),
    .B(_09072_));
 sg13g2_nand2_1 _16081_ (.Y(_09074_),
    .A(net676),
    .B(_09073_));
 sg13g2_o21ai_1 _16082_ (.B1(_09074_),
    .Y(_01576_),
    .A1(net677),
    .A2(_09070_));
 sg13g2_xnor2_1 _16083_ (.Y(_09075_),
    .A(_08890_),
    .B(_08783_));
 sg13g2_nor2_1 _16084_ (.A(net461),
    .B(_09075_),
    .Y(_09076_));
 sg13g2_xnor2_1 _16085_ (.Y(_09077_),
    .A(_08784_),
    .B(_09076_));
 sg13g2_buf_1 _16086_ (.A(_08640_),
    .X(_09078_));
 sg13g2_inv_1 _16087_ (.Y(_09079_),
    .A(_08817_));
 sg13g2_nor4_1 _16088_ (.A(_09079_),
    .B(_08794_),
    .C(_08795_),
    .D(_08815_),
    .Y(_09080_));
 sg13g2_xnor2_1 _16089_ (.Y(_09081_),
    .A(_08814_),
    .B(_09080_));
 sg13g2_nor2_1 _16090_ (.A(net608),
    .B(_09081_),
    .Y(_09082_));
 sg13g2_a21oi_1 _16091_ (.A1(net545),
    .A2(_09077_),
    .Y(_01577_),
    .B1(_09082_));
 sg13g2_buf_1 _16092_ (.A(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_09083_));
 sg13g2_buf_1 _16093_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_09084_));
 sg13g2_inv_1 _16094_ (.Y(_09085_),
    .A(_09084_));
 sg13g2_buf_1 _16095_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_09086_));
 sg13g2_buf_1 _16096_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_09087_));
 sg13g2_inv_2 _16097_ (.Y(_09088_),
    .A(_09087_));
 sg13g2_inv_1 _16098_ (.Y(_09089_),
    .A(\rbzero.wall_tracer.rayAddendY[-5] ));
 sg13g2_buf_1 _16099_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_09090_));
 sg13g2_inv_1 _16100_ (.Y(_09091_),
    .A(_09090_));
 sg13g2_buf_1 _16101_ (.A(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_09092_));
 sg13g2_buf_1 _16102_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_09093_));
 sg13g2_a21oi_1 _16103_ (.A1(_09092_),
    .A2(_09093_),
    .Y(_09094_),
    .B1(\rbzero.wall_tracer.rayAddendY[-8] ));
 sg13g2_nand3_1 _16104_ (.B(_09092_),
    .C(_09093_),
    .A(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_09095_));
 sg13g2_o21ai_1 _16105_ (.B1(_09095_),
    .Y(_09096_),
    .A1(_09091_),
    .A2(_09094_));
 sg13g2_buf_1 _16106_ (.A(_09096_),
    .X(_09097_));
 sg13g2_nor2_1 _16107_ (.A(\rbzero.wall_tracer.rayAddendY[-7] ),
    .B(_09097_),
    .Y(_09098_));
 sg13g2_buf_1 _16108_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_09099_));
 sg13g2_a21oi_1 _16109_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_09097_),
    .Y(_09100_),
    .B1(_09099_));
 sg13g2_nor2_1 _16110_ (.A(_09098_),
    .B(_09100_),
    .Y(_09101_));
 sg13g2_buf_1 _16111_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_09102_));
 sg13g2_a21o_1 _16112_ (.A2(_09101_),
    .A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_09102_),
    .X(_09103_));
 sg13g2_o21ai_1 _16113_ (.B1(_09103_),
    .Y(_09104_),
    .A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_09101_));
 sg13g2_buf_1 _16114_ (.A(_09104_),
    .X(_09105_));
 sg13g2_inv_1 _16115_ (.Y(_09106_),
    .A(_09105_));
 sg13g2_buf_2 _16116_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_09107_));
 sg13g2_a21oi_1 _16117_ (.A1(\rbzero.wall_tracer.rayAddendY[-5] ),
    .A2(_09106_),
    .Y(_09108_),
    .B1(_09107_));
 sg13g2_a21oi_1 _16118_ (.A1(_09089_),
    .A2(_09105_),
    .Y(_09109_),
    .B1(_09108_));
 sg13g2_buf_1 _16119_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_09110_));
 sg13g2_a21o_1 _16120_ (.A2(_09109_),
    .A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B1(_09110_),
    .X(_09111_));
 sg13g2_o21ai_1 _16121_ (.B1(_09111_),
    .Y(_09112_),
    .A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_09109_));
 sg13g2_buf_1 _16122_ (.A(_09112_),
    .X(_09113_));
 sg13g2_inv_1 _16123_ (.Y(_09114_),
    .A(_09113_));
 sg13g2_buf_1 _16124_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_09115_));
 sg13g2_a21oi_1 _16125_ (.A1(_09087_),
    .A2(_09114_),
    .Y(_09116_),
    .B1(_09115_));
 sg13g2_a21oi_1 _16126_ (.A1(_09088_),
    .A2(_09113_),
    .Y(_09117_),
    .B1(_09116_));
 sg13g2_buf_1 _16127_ (.A(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_09118_));
 sg13g2_a21o_1 _16128_ (.A2(_09117_),
    .A1(net822),
    .B1(_09118_),
    .X(_09119_));
 sg13g2_o21ai_1 _16129_ (.B1(_09119_),
    .Y(_09120_),
    .A1(net822),
    .A2(_09117_));
 sg13g2_buf_1 _16130_ (.A(_09120_),
    .X(_09121_));
 sg13g2_xnor2_1 _16131_ (.Y(_09122_),
    .A(_09085_),
    .B(_09121_));
 sg13g2_nor2_1 _16132_ (.A(net461),
    .B(_09122_),
    .Y(_09123_));
 sg13g2_xnor2_1 _16133_ (.Y(_09124_),
    .A(_09083_),
    .B(_09123_));
 sg13g2_buf_1 _16134_ (.A(_09107_),
    .X(_09125_));
 sg13g2_buf_1 _16135_ (.A(_09093_),
    .X(_09126_));
 sg13g2_buf_1 _16136_ (.A(_09090_),
    .X(_09127_));
 sg13g2_nor3_1 _16137_ (.A(net768),
    .B(_09099_),
    .C(_09102_),
    .Y(_09128_));
 sg13g2_nor2_1 _16138_ (.A(net769),
    .B(_09128_),
    .Y(_09129_));
 sg13g2_xor2_1 _16139_ (.B(_09129_),
    .A(net770),
    .X(_09130_));
 sg13g2_nor2_1 _16140_ (.A(net608),
    .B(_09130_),
    .Y(_09131_));
 sg13g2_a21oi_1 _16141_ (.A1(net545),
    .A2(_09124_),
    .Y(_01578_),
    .B1(_09131_));
 sg13g2_buf_2 _16142_ (.A(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_09132_));
 sg13g2_buf_1 _16143_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_09133_));
 sg13g2_inv_1 _16144_ (.Y(_09134_),
    .A(_09121_));
 sg13g2_a21oi_1 _16145_ (.A1(_09084_),
    .A2(_09134_),
    .Y(_09135_),
    .B1(_09083_));
 sg13g2_a21oi_1 _16146_ (.A1(_09085_),
    .A2(_09121_),
    .Y(_09136_),
    .B1(_09135_));
 sg13g2_and2_1 _16147_ (.A(net821),
    .B(_09136_),
    .X(_09137_));
 sg13g2_or2_1 _16148_ (.X(_09138_),
    .B(_09136_),
    .A(\rbzero.debug_overlay.vplaneY[0] ));
 sg13g2_nand3b_1 _16149_ (.B(_08807_),
    .C(_09138_),
    .Y(_09139_),
    .A_N(_09137_));
 sg13g2_xor2_1 _16150_ (.B(_09139_),
    .A(_09132_),
    .X(_09140_));
 sg13g2_buf_1 _16151_ (.A(_09110_),
    .X(_09141_));
 sg13g2_buf_1 _16152_ (.A(_09099_),
    .X(_09142_));
 sg13g2_inv_1 _16153_ (.Y(_09143_),
    .A(net766));
 sg13g2_buf_1 _16154_ (.A(_09102_),
    .X(_09144_));
 sg13g2_o21ai_1 _16155_ (.B1(_09091_),
    .Y(_09145_),
    .A1(net765),
    .A2(net769));
 sg13g2_buf_2 _16156_ (.A(_00061_),
    .X(_09146_));
 sg13g2_nand2_1 _16157_ (.Y(_09147_),
    .A(_09146_),
    .B(net765));
 sg13g2_a22oi_1 _16158_ (.Y(_09148_),
    .B1(_09147_),
    .B2(net768),
    .A2(_09145_),
    .A1(_09143_));
 sg13g2_and2_1 _16159_ (.A(_09107_),
    .B(_09093_),
    .X(_09149_));
 sg13g2_buf_1 _16160_ (.A(_09149_),
    .X(_09150_));
 sg13g2_nand2_1 _16161_ (.Y(_09151_),
    .A(net768),
    .B(net769));
 sg13g2_o21ai_1 _16162_ (.B1(_09151_),
    .Y(_09152_),
    .A1(net768),
    .A2(_09150_));
 sg13g2_o21ai_1 _16163_ (.B1(_09152_),
    .Y(_09153_),
    .A1(net770),
    .A2(_09148_));
 sg13g2_xnor2_1 _16164_ (.Y(_09154_),
    .A(net767),
    .B(_09153_));
 sg13g2_nor2_1 _16165_ (.A(net608),
    .B(_09154_),
    .Y(_09155_));
 sg13g2_a21oi_1 _16166_ (.A1(net545),
    .A2(_09140_),
    .Y(_01579_),
    .B1(_09155_));
 sg13g2_buf_2 _16167_ (.A(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_09156_));
 sg13g2_buf_1 _16168_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_09157_));
 sg13g2_buf_1 _16169_ (.A(net820),
    .X(_09158_));
 sg13g2_a21o_1 _16170_ (.A2(_09138_),
    .A1(_09132_),
    .B1(_09137_),
    .X(_09159_));
 sg13g2_buf_2 _16171_ (.A(_09159_),
    .X(_09160_));
 sg13g2_xnor2_1 _16172_ (.Y(_09161_),
    .A(net764),
    .B(_09160_));
 sg13g2_nor2_1 _16173_ (.A(net460),
    .B(_09161_),
    .Y(_09162_));
 sg13g2_xnor2_1 _16174_ (.Y(_09163_),
    .A(_09156_),
    .B(_09162_));
 sg13g2_buf_1 _16175_ (.A(_09087_),
    .X(_09164_));
 sg13g2_xor2_1 _16176_ (.B(net763),
    .A(net766),
    .X(_09165_));
 sg13g2_nor3_1 _16177_ (.A(_09107_),
    .B(_09110_),
    .C(_09093_),
    .Y(_09166_));
 sg13g2_nand2_1 _16178_ (.Y(_09167_),
    .A(_09128_),
    .B(_09166_));
 sg13g2_a21o_1 _16179_ (.A2(_09150_),
    .A1(_09110_),
    .B1(_09090_),
    .X(_09168_));
 sg13g2_o21ai_1 _16180_ (.B1(_09168_),
    .Y(_09169_),
    .A1(_09110_),
    .A2(_09150_));
 sg13g2_buf_1 _16181_ (.A(_09169_),
    .X(_09170_));
 sg13g2_nand2_1 _16182_ (.Y(_09171_),
    .A(_09167_),
    .B(_09170_));
 sg13g2_xnor2_1 _16183_ (.Y(_09172_),
    .A(_09165_),
    .B(_09171_));
 sg13g2_nand2_1 _16184_ (.Y(_09173_),
    .A(net676),
    .B(_09172_));
 sg13g2_o21ai_1 _16185_ (.B1(_09173_),
    .Y(_01580_),
    .A1(_09058_),
    .A2(_09163_));
 sg13g2_buf_1 _16186_ (.A(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_09174_));
 sg13g2_inv_1 _16187_ (.Y(_09175_),
    .A(net820));
 sg13g2_and2_1 _16188_ (.A(_09175_),
    .B(_09160_),
    .X(_09176_));
 sg13g2_buf_1 _16189_ (.A(_09175_),
    .X(_09177_));
 sg13g2_nor3_1 _16190_ (.A(_09156_),
    .B(net721),
    .C(_09160_),
    .Y(_09178_));
 sg13g2_a21oi_1 _16191_ (.A1(_09156_),
    .A2(_09176_),
    .Y(_09179_),
    .B1(_09178_));
 sg13g2_nor2_1 _16192_ (.A(net460),
    .B(_09179_),
    .Y(_09180_));
 sg13g2_xnor2_1 _16193_ (.Y(_09181_),
    .A(net819),
    .B(_09180_));
 sg13g2_xor2_1 _16194_ (.B(net822),
    .A(_09102_),
    .X(_09182_));
 sg13g2_nor2_2 _16195_ (.A(_09087_),
    .B(_09167_),
    .Y(_09183_));
 sg13g2_inv_1 _16196_ (.Y(_09184_),
    .A(_09170_));
 sg13g2_a21oi_1 _16197_ (.A1(_09087_),
    .A2(_09184_),
    .Y(_09185_),
    .B1(_09099_));
 sg13g2_a21oi_1 _16198_ (.A1(_09088_),
    .A2(_09170_),
    .Y(_09186_),
    .B1(_09185_));
 sg13g2_a21oi_1 _16199_ (.A1(_09146_),
    .A2(_09183_),
    .Y(_09187_),
    .B1(_09186_));
 sg13g2_xor2_1 _16200_ (.B(_09187_),
    .A(_09182_),
    .X(_09188_));
 sg13g2_nand2_1 _16201_ (.Y(_09189_),
    .A(net676),
    .B(_09188_));
 sg13g2_o21ai_1 _16202_ (.B1(_09189_),
    .Y(_01581_),
    .A1(net677),
    .A2(_09181_));
 sg13g2_buf_1 _16203_ (.A(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_09190_));
 sg13g2_inv_1 _16204_ (.Y(_09191_),
    .A(_09156_));
 sg13g2_a21oi_1 _16205_ (.A1(net819),
    .A2(_09160_),
    .Y(_09192_),
    .B1(net820));
 sg13g2_o21ai_1 _16206_ (.B1(net764),
    .Y(_09193_),
    .A1(net819),
    .A2(_09160_));
 sg13g2_o21ai_1 _16207_ (.B1(_09193_),
    .Y(_09194_),
    .A1(_09191_),
    .A2(_09192_));
 sg13g2_xnor2_1 _16208_ (.Y(_09195_),
    .A(net764),
    .B(_09194_));
 sg13g2_nor2_1 _16209_ (.A(net460),
    .B(_09195_),
    .Y(_09196_));
 sg13g2_xnor2_1 _16210_ (.Y(_09197_),
    .A(net818),
    .B(_09196_));
 sg13g2_inv_1 _16211_ (.Y(_09198_),
    .A(_09186_));
 sg13g2_a21o_1 _16212_ (.A2(_09198_),
    .A1(_09182_),
    .B1(_09183_),
    .X(_09199_));
 sg13g2_buf_1 _16213_ (.A(_09199_),
    .X(_09200_));
 sg13g2_xnor2_1 _16214_ (.Y(_09201_),
    .A(_09107_),
    .B(_09084_));
 sg13g2_buf_1 _16215_ (.A(_09201_),
    .X(_09202_));
 sg13g2_nor2_1 _16216_ (.A(net765),
    .B(net822),
    .Y(_09203_));
 sg13g2_xor2_1 _16217_ (.B(_09203_),
    .A(_09202_),
    .X(_09204_));
 sg13g2_xnor2_1 _16218_ (.Y(_09205_),
    .A(_09200_),
    .B(_09204_));
 sg13g2_nand2_1 _16219_ (.Y(_09206_),
    .A(net676),
    .B(_09205_));
 sg13g2_o21ai_1 _16220_ (.B1(_09206_),
    .Y(_01582_),
    .A1(_09058_),
    .A2(_09197_));
 sg13g2_buf_1 _16221_ (.A(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_09207_));
 sg13g2_inv_1 _16222_ (.Y(_09208_),
    .A(net817));
 sg13g2_nor2_1 _16223_ (.A(net819),
    .B(_09175_),
    .Y(_09209_));
 sg13g2_a21oi_1 _16224_ (.A1(net819),
    .A2(_09176_),
    .Y(_09210_),
    .B1(_09209_));
 sg13g2_nand2_1 _16225_ (.Y(_09211_),
    .A(_09160_),
    .B(_09209_));
 sg13g2_o21ai_1 _16226_ (.B1(_09211_),
    .Y(_09212_),
    .A1(_09191_),
    .A2(_09210_));
 sg13g2_buf_1 _16227_ (.A(_09212_),
    .X(_09213_));
 sg13g2_nor4_1 _16228_ (.A(net819),
    .B(_09190_),
    .C(net721),
    .D(_09213_),
    .Y(_09214_));
 sg13g2_and3_1 _16229_ (.X(_09215_),
    .A(net818),
    .B(net721),
    .C(_09213_));
 sg13g2_o21ai_1 _16230_ (.B1(net462),
    .Y(_09216_),
    .A1(_09214_),
    .A2(_09215_));
 sg13g2_xnor2_1 _16231_ (.Y(_09217_),
    .A(_09208_),
    .B(_09216_));
 sg13g2_inv_1 _16232_ (.Y(_09218_),
    .A(net822));
 sg13g2_nor2_1 _16233_ (.A(_09099_),
    .B(net763),
    .Y(_09219_));
 sg13g2_buf_1 _16234_ (.A(_09219_),
    .X(_09220_));
 sg13g2_nor2_1 _16235_ (.A(_09220_),
    .B(_09202_),
    .Y(_09221_));
 sg13g2_a21oi_1 _16236_ (.A1(_09218_),
    .A2(_09220_),
    .Y(_09222_),
    .B1(_09221_));
 sg13g2_nand3_1 _16237_ (.B(_09086_),
    .C(_09220_),
    .A(_09102_),
    .Y(_09223_));
 sg13g2_o21ai_1 _16238_ (.B1(_09223_),
    .Y(_09224_),
    .A1(_09086_),
    .A2(_09220_));
 sg13g2_nand2b_1 _16239_ (.Y(_09225_),
    .B(_09224_),
    .A_N(_09202_));
 sg13g2_o21ai_1 _16240_ (.B1(_09225_),
    .Y(_09226_),
    .A1(net765),
    .A2(_09222_));
 sg13g2_nor2_1 _16241_ (.A(_09107_),
    .B(_09093_),
    .Y(_09227_));
 sg13g2_xnor2_1 _16242_ (.Y(_09228_),
    .A(net768),
    .B(net767));
 sg13g2_nor3_1 _16243_ (.A(_09150_),
    .B(_09227_),
    .C(_09228_),
    .Y(_09229_));
 sg13g2_a21oi_1 _16244_ (.A1(net763),
    .A2(_09229_),
    .Y(_09230_),
    .B1(_09183_));
 sg13g2_nand3_1 _16245_ (.B(_09088_),
    .C(_09229_),
    .A(net766),
    .Y(_09231_));
 sg13g2_o21ai_1 _16246_ (.B1(_09231_),
    .Y(_09232_),
    .A1(net766),
    .A2(_09230_));
 sg13g2_o21ai_1 _16247_ (.B1(net767),
    .Y(_09233_),
    .A1(_09107_),
    .A2(_09093_));
 sg13g2_a21oi_1 _16248_ (.A1(_09091_),
    .A2(_09233_),
    .Y(_09234_),
    .B1(_09166_));
 sg13g2_a21oi_1 _16249_ (.A1(net766),
    .A2(net763),
    .Y(_09235_),
    .B1(_09234_));
 sg13g2_nor3_1 _16250_ (.A(_09218_),
    .B(_09220_),
    .C(_09235_),
    .Y(_09236_));
 sg13g2_or2_1 _16251_ (.X(_09237_),
    .B(_09236_),
    .A(_09102_));
 sg13g2_o21ai_1 _16252_ (.B1(_09218_),
    .Y(_09238_),
    .A1(_09220_),
    .A2(_09235_));
 sg13g2_a21oi_1 _16253_ (.A1(_09237_),
    .A2(_09238_),
    .Y(_09239_),
    .B1(_09202_));
 sg13g2_a21oi_1 _16254_ (.A1(_09226_),
    .A2(_09232_),
    .Y(_09240_),
    .B1(_09239_));
 sg13g2_xor2_1 _16255_ (.B(_09133_),
    .A(_09141_),
    .X(_09241_));
 sg13g2_buf_1 _16256_ (.A(_09084_),
    .X(_09242_));
 sg13g2_nor2_2 _16257_ (.A(net770),
    .B(net762),
    .Y(_09243_));
 sg13g2_xor2_1 _16258_ (.B(_09243_),
    .A(_09241_),
    .X(_09244_));
 sg13g2_xnor2_1 _16259_ (.Y(_09245_),
    .A(_09240_),
    .B(_09244_));
 sg13g2_nand2_1 _16260_ (.Y(_09246_),
    .A(net676),
    .B(_09245_));
 sg13g2_o21ai_1 _16261_ (.B1(_09246_),
    .Y(_01583_),
    .A1(net677),
    .A2(_09217_));
 sg13g2_buf_1 _16262_ (.A(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_09247_));
 sg13g2_buf_1 _16263_ (.A(_09247_),
    .X(_09248_));
 sg13g2_and2_1 _16264_ (.A(net818),
    .B(net817),
    .X(_09249_));
 sg13g2_nand3_1 _16265_ (.B(_09160_),
    .C(_09249_),
    .A(net819),
    .Y(_09250_));
 sg13g2_or4_1 _16266_ (.A(_09174_),
    .B(net818),
    .C(net817),
    .D(_09160_),
    .X(_09251_));
 sg13g2_a21oi_1 _16267_ (.A1(net820),
    .A2(_09251_),
    .Y(_09252_),
    .B1(_09156_));
 sg13g2_a21oi_1 _16268_ (.A1(net721),
    .A2(_09250_),
    .Y(_09253_),
    .B1(_09252_));
 sg13g2_xnor2_1 _16269_ (.Y(_09254_),
    .A(net764),
    .B(_09253_));
 sg13g2_nor2_1 _16270_ (.A(_09063_),
    .B(_09254_),
    .Y(_09255_));
 sg13g2_xnor2_1 _16271_ (.Y(_09256_),
    .A(net761),
    .B(_09255_));
 sg13g2_inv_1 _16272_ (.Y(_09257_),
    .A(_09200_));
 sg13g2_a21oi_1 _16273_ (.A1(_09084_),
    .A2(_09257_),
    .Y(_09258_),
    .B1(net770));
 sg13g2_a21o_1 _16274_ (.A2(_09200_),
    .A1(_09085_),
    .B1(_09258_),
    .X(_09259_));
 sg13g2_a21oi_1 _16275_ (.A1(_09085_),
    .A2(_09200_),
    .Y(_09260_),
    .B1(_09241_));
 sg13g2_o21ai_1 _16276_ (.B1(_09241_),
    .Y(_09261_),
    .A1(_09085_),
    .A2(_09200_));
 sg13g2_o21ai_1 _16277_ (.B1(_09261_),
    .Y(_09262_),
    .A1(net770),
    .A2(_09260_));
 sg13g2_a22oi_1 _16278_ (.Y(_09263_),
    .B1(_09262_),
    .B2(_09203_),
    .A2(_09259_),
    .A1(_09241_));
 sg13g2_buf_1 _16279_ (.A(_09263_),
    .X(_09264_));
 sg13g2_xor2_1 _16280_ (.B(_09157_),
    .A(_09164_),
    .X(_09265_));
 sg13g2_buf_2 _16281_ (.A(_09265_),
    .X(_09266_));
 sg13g2_nor2_1 _16282_ (.A(net767),
    .B(net821),
    .Y(_09267_));
 sg13g2_xor2_1 _16283_ (.B(_09267_),
    .A(_09266_),
    .X(_09268_));
 sg13g2_xnor2_1 _16284_ (.Y(_09269_),
    .A(_09264_),
    .B(_09268_));
 sg13g2_nand2_1 _16285_ (.Y(_09270_),
    .A(_09071_),
    .B(_09269_));
 sg13g2_o21ai_1 _16286_ (.B1(_09270_),
    .Y(_01584_),
    .A1(net677),
    .A2(_09256_));
 sg13g2_buf_2 _16287_ (.A(\rbzero.wall_tracer.rayAddendY[6] ),
    .X(_09271_));
 sg13g2_nand3_1 _16288_ (.B(net761),
    .C(_09213_),
    .A(net817),
    .Y(_09272_));
 sg13g2_or4_1 _16289_ (.A(_09174_),
    .B(net817),
    .C(net761),
    .D(_09213_),
    .X(_09273_));
 sg13g2_a21oi_1 _16290_ (.A1(net820),
    .A2(_09273_),
    .Y(_09274_),
    .B1(net818));
 sg13g2_a21oi_2 _16291_ (.B1(_09274_),
    .Y(_09275_),
    .A2(_09272_),
    .A1(net721));
 sg13g2_xnor2_1 _16292_ (.Y(_09276_),
    .A(net764),
    .B(_09275_));
 sg13g2_nor2_1 _16293_ (.A(_09063_),
    .B(_09276_),
    .Y(_09277_));
 sg13g2_xnor2_1 _16294_ (.Y(_09278_),
    .A(_09271_),
    .B(_09277_));
 sg13g2_nand3_1 _16295_ (.B(_09183_),
    .C(_09203_),
    .A(_09146_),
    .Y(_09279_));
 sg13g2_nor3_1 _16296_ (.A(net770),
    .B(net762),
    .C(_09279_),
    .Y(_09280_));
 sg13g2_a21oi_1 _16297_ (.A1(net822),
    .A2(_09186_),
    .Y(_09281_),
    .B1(net765));
 sg13g2_a221oi_1 _16298_ (.B2(_09146_),
    .C1(_09281_),
    .B1(_09183_),
    .A1(_09218_),
    .Y(_09282_),
    .A2(_09198_));
 sg13g2_o21ai_1 _16299_ (.B1(_09279_),
    .Y(_09283_),
    .A1(_09202_),
    .A2(_09282_));
 sg13g2_inv_1 _16300_ (.Y(_09284_),
    .A(net821));
 sg13g2_o21ai_1 _16301_ (.B1(_09284_),
    .Y(_09285_),
    .A1(_09243_),
    .A2(_09283_));
 sg13g2_nand2b_1 _16302_ (.Y(_09286_),
    .B(_09285_),
    .A_N(_09280_));
 sg13g2_and2_1 _16303_ (.A(_09266_),
    .B(_09286_),
    .X(_09287_));
 sg13g2_o21ai_1 _16304_ (.B1(_09284_),
    .Y(_09288_),
    .A1(_09266_),
    .A2(_09280_));
 sg13g2_o21ai_1 _16305_ (.B1(_09266_),
    .Y(_09289_),
    .A1(_09243_),
    .A2(_09283_));
 sg13g2_a21oi_1 _16306_ (.A1(_09288_),
    .A2(_09289_),
    .Y(_09290_),
    .B1(net767));
 sg13g2_nor2_1 _16307_ (.A(_09287_),
    .B(_09290_),
    .Y(_09291_));
 sg13g2_buf_1 _16308_ (.A(net822),
    .X(_09292_));
 sg13g2_nor2_1 _16309_ (.A(_09088_),
    .B(_09158_),
    .Y(_09293_));
 sg13g2_xnor2_1 _16310_ (.Y(_09294_),
    .A(net760),
    .B(_09293_));
 sg13g2_xnor2_1 _16311_ (.Y(_09295_),
    .A(_09291_),
    .B(_09294_));
 sg13g2_nand2_1 _16312_ (.Y(_09296_),
    .A(_09071_),
    .B(_09295_));
 sg13g2_o21ai_1 _16313_ (.B1(_09296_),
    .Y(_01585_),
    .A1(net677),
    .A2(_09278_));
 sg13g2_buf_1 _16314_ (.A(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_09297_));
 sg13g2_nor2b_1 _16315_ (.A(net820),
    .B_N(_09271_),
    .Y(_09298_));
 sg13g2_nand4_1 _16316_ (.B(_09194_),
    .C(_09249_),
    .A(net761),
    .Y(_09299_),
    .D(_09298_));
 sg13g2_nand2b_1 _16317_ (.Y(_09300_),
    .B(net820),
    .A_N(_09271_));
 sg13g2_nor4_1 _16318_ (.A(net818),
    .B(net817),
    .C(net761),
    .D(_09300_),
    .Y(_09301_));
 sg13g2_nand2b_1 _16319_ (.Y(_09302_),
    .B(_09301_),
    .A_N(_09194_));
 sg13g2_a21oi_1 _16320_ (.A1(_09299_),
    .A2(_09302_),
    .Y(_09303_),
    .B1(net463));
 sg13g2_xnor2_1 _16321_ (.Y(_09304_),
    .A(_09297_),
    .B(_09303_));
 sg13g2_nor2_1 _16322_ (.A(net721),
    .B(_09264_),
    .Y(_09305_));
 sg13g2_a21oi_1 _16323_ (.A1(net721),
    .A2(_09264_),
    .Y(_09306_),
    .B1(net763));
 sg13g2_o21ai_1 _16324_ (.B1(_09267_),
    .Y(_09307_),
    .A1(_09305_),
    .A2(_09306_));
 sg13g2_nand2_1 _16325_ (.Y(_09308_),
    .A(_09088_),
    .B(_09305_));
 sg13g2_nand2_1 _16326_ (.Y(_09309_),
    .A(_09307_),
    .B(_09308_));
 sg13g2_nand2_1 _16327_ (.Y(_09310_),
    .A(net763),
    .B(_09264_));
 sg13g2_o21ai_1 _16328_ (.B1(net721),
    .Y(_09311_),
    .A1(_09267_),
    .A2(_09310_));
 sg13g2_nand2_1 _16329_ (.Y(_09312_),
    .A(net760),
    .B(_09311_));
 sg13g2_o21ai_1 _16330_ (.B1(_09312_),
    .Y(_09313_),
    .A1(net760),
    .A2(_09309_));
 sg13g2_buf_1 _16331_ (.A(_09313_),
    .X(_09314_));
 sg13g2_nor2_1 _16332_ (.A(_09218_),
    .B(net764),
    .Y(_09315_));
 sg13g2_xnor2_1 _16333_ (.Y(_09316_),
    .A(net762),
    .B(_09315_));
 sg13g2_xnor2_1 _16334_ (.Y(_09317_),
    .A(_09314_),
    .B(_09316_));
 sg13g2_nor2_1 _16335_ (.A(net608),
    .B(_09317_),
    .Y(_09318_));
 sg13g2_a21oi_1 _16336_ (.A1(net544),
    .A2(_09304_),
    .Y(_01586_),
    .B1(_09318_));
 sg13g2_buf_2 _16337_ (.A(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_09319_));
 sg13g2_inv_1 _16338_ (.Y(_09320_),
    .A(_09297_));
 sg13g2_nand2b_1 _16339_ (.Y(_09321_),
    .B(_09320_),
    .A_N(_09300_));
 sg13g2_nand2_1 _16340_ (.Y(_09322_),
    .A(_09297_),
    .B(_09298_));
 sg13g2_mux2_1 _16341_ (.A0(_09321_),
    .A1(_09322_),
    .S(_09275_),
    .X(_09323_));
 sg13g2_nor2_1 _16342_ (.A(net463),
    .B(_09323_),
    .Y(_09324_));
 sg13g2_xnor2_1 _16343_ (.Y(_09325_),
    .A(_09319_),
    .B(_09324_));
 sg13g2_nand3_1 _16344_ (.B(net762),
    .C(_09293_),
    .A(net760),
    .Y(_09326_));
 sg13g2_or3_1 _16345_ (.A(_09292_),
    .B(net762),
    .C(_09293_),
    .X(_09327_));
 sg13g2_nand2_1 _16346_ (.Y(_09328_),
    .A(_09146_),
    .B(_09126_));
 sg13g2_nand3_1 _16347_ (.B(_09142_),
    .C(_09144_),
    .A(_09127_),
    .Y(_09329_));
 sg13g2_nor2b_1 _16348_ (.A(_09125_),
    .B_N(_09329_),
    .Y(_09330_));
 sg13g2_nor3_1 _16349_ (.A(_09239_),
    .B(_09328_),
    .C(_09330_),
    .Y(_09331_));
 sg13g2_nor2_1 _16350_ (.A(_09240_),
    .B(_09331_),
    .Y(_09332_));
 sg13g2_or2_1 _16351_ (.X(_09333_),
    .B(_09332_),
    .A(_09243_));
 sg13g2_and2_1 _16352_ (.A(_09243_),
    .B(_09332_),
    .X(_09334_));
 sg13g2_or2_1 _16353_ (.X(_09335_),
    .B(_09334_),
    .A(_09266_));
 sg13g2_a22oi_1 _16354_ (.Y(_09336_),
    .B1(_09335_),
    .B2(_09284_),
    .A2(_09333_),
    .A1(_09266_));
 sg13g2_and2_1 _16355_ (.A(_09284_),
    .B(_09333_),
    .X(_09337_));
 sg13g2_o21ai_1 _16356_ (.B1(_09266_),
    .Y(_09338_),
    .A1(_09334_),
    .A2(_09337_));
 sg13g2_o21ai_1 _16357_ (.B1(_09338_),
    .Y(_09339_),
    .A1(net767),
    .A2(_09336_));
 sg13g2_mux2_1 _16358_ (.A0(_09326_),
    .A1(_09327_),
    .S(_09339_),
    .X(_09340_));
 sg13g2_xnor2_1 _16359_ (.Y(_09341_),
    .A(_09284_),
    .B(_09340_));
 sg13g2_nor2_1 _16360_ (.A(net608),
    .B(_09341_),
    .Y(_09342_));
 sg13g2_a21oi_1 _16361_ (.A1(net544),
    .A2(_09325_),
    .Y(_01587_),
    .B1(_09342_));
 sg13g2_buf_2 _16362_ (.A(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_09343_));
 sg13g2_inv_1 _16363_ (.Y(_09344_),
    .A(_09319_));
 sg13g2_nor2_1 _16364_ (.A(_09344_),
    .B(_09322_),
    .Y(_09345_));
 sg13g2_and3_1 _16365_ (.X(_09346_),
    .A(net761),
    .B(_09253_),
    .C(_09345_));
 sg13g2_nor4_1 _16366_ (.A(net761),
    .B(_09319_),
    .C(_09253_),
    .D(_09321_),
    .Y(_09347_));
 sg13g2_o21ai_1 _16367_ (.B1(net462),
    .Y(_09348_),
    .A1(_09346_),
    .A2(_09347_));
 sg13g2_xor2_1 _16368_ (.B(_09348_),
    .A(_09343_),
    .X(_09349_));
 sg13g2_o21ai_1 _16369_ (.B1(_09158_),
    .Y(_09350_),
    .A1(net821),
    .A2(_09314_));
 sg13g2_nand2_1 _16370_ (.Y(_09351_),
    .A(net760),
    .B(net821));
 sg13g2_o21ai_1 _16371_ (.B1(_09177_),
    .Y(_09352_),
    .A1(_09310_),
    .A2(_09351_));
 sg13g2_nor2_1 _16372_ (.A(_09133_),
    .B(_09314_),
    .Y(_09353_));
 sg13g2_nor3_1 _16373_ (.A(net760),
    .B(net762),
    .C(net764),
    .Y(_09354_));
 sg13g2_a22oi_1 _16374_ (.Y(_09355_),
    .B1(_09353_),
    .B2(_09354_),
    .A2(_09352_),
    .A1(_09242_));
 sg13g2_a21oi_1 _16375_ (.A1(_09350_),
    .A2(_09355_),
    .Y(_09356_),
    .B1(net609));
 sg13g2_a21oi_1 _16376_ (.A1(net544),
    .A2(_09349_),
    .Y(_01588_),
    .B1(_09356_));
 sg13g2_buf_2 _16377_ (.A(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_09357_));
 sg13g2_and3_1 _16378_ (.X(_09358_),
    .A(_09343_),
    .B(_09275_),
    .C(_09345_));
 sg13g2_nor4_1 _16379_ (.A(_09319_),
    .B(_09343_),
    .C(_09275_),
    .D(_09321_),
    .Y(_09359_));
 sg13g2_o21ai_1 _16380_ (.B1(net462),
    .Y(_09360_),
    .A1(_09358_),
    .A2(_09359_));
 sg13g2_xor2_1 _16381_ (.B(_09360_),
    .A(_09357_),
    .X(_09361_));
 sg13g2_nor4_1 _16382_ (.A(_09164_),
    .B(net760),
    .C(_09242_),
    .D(net821),
    .Y(_09362_));
 sg13g2_o21ai_1 _16383_ (.B1(_09362_),
    .Y(_09363_),
    .A1(_09287_),
    .A2(_09290_));
 sg13g2_nand3_1 _16384_ (.B(_08412_),
    .C(_09363_),
    .A(_09177_),
    .Y(_09364_));
 sg13g2_o21ai_1 _16385_ (.B1(_09364_),
    .Y(_01589_),
    .A1(net677),
    .A2(_09361_));
 sg13g2_nand2_1 _16386_ (.Y(_09365_),
    .A(_09126_),
    .B(net462));
 sg13g2_xor2_1 _16387_ (.B(_09365_),
    .A(_09092_),
    .X(_09366_));
 sg13g2_nor2_1 _16388_ (.A(net678),
    .B(_09366_),
    .Y(_01590_));
 sg13g2_nand2_1 _16389_ (.Y(_09367_),
    .A(_09092_),
    .B(net769));
 sg13g2_xnor2_1 _16390_ (.Y(_09368_),
    .A(_09091_),
    .B(_09367_));
 sg13g2_nor2_1 _16391_ (.A(net461),
    .B(_09368_),
    .Y(_09369_));
 sg13g2_xnor2_1 _16392_ (.Y(_09370_),
    .A(\rbzero.wall_tracer.rayAddendY[-8] ),
    .B(_09369_));
 sg13g2_nor2_1 _16393_ (.A(net678),
    .B(_09370_),
    .Y(_01591_));
 sg13g2_xnor2_1 _16394_ (.Y(_09371_),
    .A(_09142_),
    .B(_09097_));
 sg13g2_nor2_1 _16395_ (.A(net461),
    .B(_09371_),
    .Y(_09372_));
 sg13g2_xnor2_1 _16396_ (.Y(_09373_),
    .A(\rbzero.wall_tracer.rayAddendY[-7] ),
    .B(_09372_));
 sg13g2_nor2_1 _16397_ (.A(net678),
    .B(_09373_),
    .Y(_01592_));
 sg13g2_xnor2_1 _16398_ (.Y(_09374_),
    .A(_09144_),
    .B(_09101_));
 sg13g2_nor2_1 _16399_ (.A(net461),
    .B(_09374_),
    .Y(_09375_));
 sg13g2_xnor2_1 _16400_ (.Y(_09376_),
    .A(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B(_09375_));
 sg13g2_nor2_1 _16401_ (.A(net678),
    .B(_09376_),
    .Y(_01593_));
 sg13g2_xor2_1 _16402_ (.B(_09105_),
    .A(_09125_),
    .X(_09377_));
 sg13g2_nor2_1 _16403_ (.A(net460),
    .B(_09377_),
    .Y(_09378_));
 sg13g2_xnor2_1 _16404_ (.Y(_09379_),
    .A(\rbzero.wall_tracer.rayAddendY[-5] ),
    .B(_09378_));
 sg13g2_nand2_1 _16405_ (.Y(_09380_),
    .A(net769),
    .B(_08412_));
 sg13g2_o21ai_1 _16406_ (.B1(_09380_),
    .Y(_01594_),
    .A1(net679),
    .A2(_09379_));
 sg13g2_xnor2_1 _16407_ (.Y(_09381_),
    .A(_09141_),
    .B(_09109_));
 sg13g2_nor2_1 _16408_ (.A(net460),
    .B(_09381_),
    .Y(_09382_));
 sg13g2_xnor2_1 _16409_ (.Y(_09383_),
    .A(\rbzero.wall_tracer.rayAddendY[-4] ),
    .B(_09382_));
 sg13g2_xor2_1 _16410_ (.B(net769),
    .A(_09127_),
    .X(_09384_));
 sg13g2_nand2_1 _16411_ (.Y(_09385_),
    .A(net676),
    .B(_09384_));
 sg13g2_o21ai_1 _16412_ (.B1(_09385_),
    .Y(_01595_),
    .A1(net679),
    .A2(_09383_));
 sg13g2_xnor2_1 _16413_ (.Y(_09386_),
    .A(_09088_),
    .B(_09113_));
 sg13g2_nor2_1 _16414_ (.A(net460),
    .B(_09386_),
    .Y(_09387_));
 sg13g2_xnor2_1 _16415_ (.Y(_09388_),
    .A(_09115_),
    .B(_09387_));
 sg13g2_nor2_1 _16416_ (.A(net768),
    .B(net769),
    .Y(_09389_));
 sg13g2_xnor2_1 _16417_ (.Y(_09390_),
    .A(net766),
    .B(_09389_));
 sg13g2_nand2_1 _16418_ (.Y(_09391_),
    .A(net676),
    .B(_09390_));
 sg13g2_o21ai_1 _16419_ (.B1(_09391_),
    .Y(_01596_),
    .A1(net679),
    .A2(_09388_));
 sg13g2_xnor2_1 _16420_ (.Y(_09392_),
    .A(net760),
    .B(_09117_));
 sg13g2_nor2_1 _16421_ (.A(_08680_),
    .B(_09392_),
    .Y(_09393_));
 sg13g2_xnor2_1 _16422_ (.Y(_09394_),
    .A(_09118_),
    .B(_09393_));
 sg13g2_nand3_1 _16423_ (.B(_09143_),
    .C(_09389_),
    .A(_09146_),
    .Y(_09395_));
 sg13g2_xor2_1 _16424_ (.B(_09395_),
    .A(net765),
    .X(_09396_));
 sg13g2_nand2_1 _16425_ (.Y(_09397_),
    .A(net676),
    .B(_09396_));
 sg13g2_o21ai_1 _16426_ (.B1(_09397_),
    .Y(_01597_),
    .A1(net679),
    .A2(_09394_));
 sg13g2_buf_2 _16427_ (.A(\rbzero.debug_overlay.vpos[5] ),
    .X(_09398_));
 sg13g2_buf_2 _16428_ (.A(\rbzero.debug_overlay.vpos[9] ),
    .X(_09399_));
 sg13g2_buf_2 _16429_ (.A(\rbzero.debug_overlay.vpos[1] ),
    .X(_09400_));
 sg13g2_buf_1 _16430_ (.A(\rbzero.debug_overlay.vpos[0] ),
    .X(_09401_));
 sg13g2_buf_1 _16431_ (.A(\rbzero.debug_overlay.vpos[4] ),
    .X(_09402_));
 sg13g2_buf_2 _16432_ (.A(\rbzero.debug_overlay.vpos[3] ),
    .X(_09403_));
 sg13g2_inv_2 _16433_ (.Y(_09404_),
    .A(_09403_));
 sg13g2_buf_1 _16434_ (.A(\rbzero.debug_overlay.vpos[2] ),
    .X(_09405_));
 sg13g2_inv_1 _16435_ (.Y(_09406_),
    .A(_09405_));
 sg13g2_nor2_1 _16436_ (.A(_09404_),
    .B(_09406_),
    .Y(_09407_));
 sg13g2_nand4_1 _16437_ (.B(net816),
    .C(_09402_),
    .A(_09400_),
    .Y(_09408_),
    .D(_09407_));
 sg13g2_or2_1 _16438_ (.X(_09409_),
    .B(_09408_),
    .A(_08473_));
 sg13g2_buf_1 _16439_ (.A(_09409_),
    .X(_09410_));
 sg13g2_buf_1 _16440_ (.A(\rbzero.debug_overlay.vpos[7] ),
    .X(_09411_));
 sg13g2_buf_1 _16441_ (.A(\rbzero.debug_overlay.vpos[6] ),
    .X(_09412_));
 sg13g2_nand3_1 _16442_ (.B(_09412_),
    .C(\rbzero.debug_overlay.vpos[8] ),
    .A(_09411_),
    .Y(_09413_));
 sg13g2_buf_1 _16443_ (.A(_09413_),
    .X(_09414_));
 sg13g2_or4_1 _16444_ (.A(_09398_),
    .B(_09399_),
    .C(_09410_),
    .D(_09414_),
    .X(_09415_));
 sg13g2_buf_1 _16445_ (.A(_09415_),
    .X(_09416_));
 sg13g2_nor2_1 _16446_ (.A(net6),
    .B(net5),
    .Y(_09417_));
 sg13g2_nor2_1 _16447_ (.A(_09416_),
    .B(_09417_),
    .Y(_09418_));
 sg13g2_buf_1 _16448_ (.A(_09418_),
    .X(_09419_));
 sg13g2_buf_1 _16449_ (.A(_09419_),
    .X(_09420_));
 sg13g2_buf_1 _16450_ (.A(net359),
    .X(_09421_));
 sg13g2_buf_1 _16451_ (.A(\rbzero.pov.spi_done ),
    .X(_09422_));
 sg13g2_buf_1 _16452_ (.A(_09422_),
    .X(_09423_));
 sg13g2_buf_2 _16453_ (.A(_08409_),
    .X(_09424_));
 sg13g2_buf_1 _16454_ (.A(_09424_),
    .X(_09425_));
 sg13g2_o21ai_1 _16455_ (.B1(net758),
    .Y(_09426_),
    .A1(net759),
    .A2(\rbzero.pov.ready ));
 sg13g2_nor2_1 _16456_ (.A(net340),
    .B(_09426_),
    .Y(_00530_));
 sg13g2_nand2b_1 _16457_ (.Y(_09427_),
    .B(_08409_),
    .A_N(\rbzero.pov.ss_buffer[1] ));
 sg13g2_nor2b_1 _16458_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_09428_));
 sg13g2_buf_1 _16459_ (.A(_09428_),
    .X(_09429_));
 sg13g2_xnor2_1 _16460_ (.Y(_09430_),
    .A(\rbzero.pov.spi_counter[0] ),
    .B(_09429_));
 sg13g2_nor2_1 _16461_ (.A(_09427_),
    .B(_09430_),
    .Y(_00682_));
 sg13g2_buf_1 _16462_ (.A(\rbzero.pov.spi_counter[1] ),
    .X(_09431_));
 sg13g2_inv_1 _16463_ (.Y(_09432_),
    .A(_09431_));
 sg13g2_buf_1 _16464_ (.A(\rbzero.pov.spi_counter[3] ),
    .X(_09433_));
 sg13g2_and2_1 _16465_ (.A(\rbzero.pov.spi_counter[0] ),
    .B(_09429_),
    .X(_09434_));
 sg13g2_buf_1 _16466_ (.A(_09434_),
    .X(_09435_));
 sg13g2_buf_1 _16467_ (.A(\rbzero.pov.spi_counter[2] ),
    .X(_09436_));
 sg13g2_buf_1 _16468_ (.A(\rbzero.pov.spi_counter[4] ),
    .X(_09437_));
 sg13g2_nor4_1 _16469_ (.A(_09436_),
    .B(\rbzero.pov.spi_counter[5] ),
    .C(_09437_),
    .D(_00026_),
    .Y(_09438_));
 sg13g2_nand4_1 _16470_ (.B(_09433_),
    .C(_09435_),
    .A(_09432_),
    .Y(_09439_),
    .D(_09438_));
 sg13g2_nand2b_1 _16471_ (.Y(_09440_),
    .B(_09439_),
    .A_N(_09427_));
 sg13g2_buf_1 _16472_ (.A(_09440_),
    .X(_09441_));
 sg13g2_xnor2_1 _16473_ (.Y(_09442_),
    .A(_09431_),
    .B(_09435_));
 sg13g2_nor2_1 _16474_ (.A(_09441_),
    .B(_09442_),
    .Y(_00683_));
 sg13g2_nand2_1 _16475_ (.Y(_09443_),
    .A(_09431_),
    .B(_09435_));
 sg13g2_xor2_1 _16476_ (.B(_09443_),
    .A(_09436_),
    .X(_09444_));
 sg13g2_nor2_1 _16477_ (.A(_09441_),
    .B(_09444_),
    .Y(_00684_));
 sg13g2_and3_1 _16478_ (.X(_09445_),
    .A(_09431_),
    .B(_09436_),
    .C(_09435_));
 sg13g2_xnor2_1 _16479_ (.Y(_09446_),
    .A(_09433_),
    .B(_09445_));
 sg13g2_nor2_1 _16480_ (.A(_09441_),
    .B(_09446_),
    .Y(_00685_));
 sg13g2_and2_1 _16481_ (.A(_09433_),
    .B(_09445_),
    .X(_09447_));
 sg13g2_xnor2_1 _16482_ (.Y(_09448_),
    .A(_09437_),
    .B(_09447_));
 sg13g2_nor2_1 _16483_ (.A(_09441_),
    .B(_09448_),
    .Y(_00686_));
 sg13g2_nand2_1 _16484_ (.Y(_09449_),
    .A(_09437_),
    .B(_09447_));
 sg13g2_xor2_1 _16485_ (.B(_09449_),
    .A(\rbzero.pov.spi_counter[5] ),
    .X(_09450_));
 sg13g2_nor2_1 _16486_ (.A(_09441_),
    .B(_09450_),
    .Y(_00687_));
 sg13g2_and4_1 _16487_ (.A(_09431_),
    .B(_09436_),
    .C(\rbzero.pov.spi_counter[5] ),
    .D(_09437_),
    .X(_09451_));
 sg13g2_nand3_1 _16488_ (.B(_09433_),
    .C(_09451_),
    .A(\rbzero.pov.spi_counter[0] ),
    .Y(_09452_));
 sg13g2_xor2_1 _16489_ (.B(_09452_),
    .A(_00026_),
    .X(_09453_));
 sg13g2_nor2b_1 _16490_ (.A(_09429_),
    .B_N(\rbzero.pov.spi_counter[6] ),
    .Y(_09454_));
 sg13g2_a21oi_1 _16491_ (.A1(_09429_),
    .A2(_09453_),
    .Y(_09455_),
    .B1(_09454_));
 sg13g2_nor2_1 _16492_ (.A(_09441_),
    .B(_09455_),
    .Y(_00688_));
 sg13g2_buf_1 _16493_ (.A(_09422_),
    .X(_09456_));
 sg13g2_buf_1 _16494_ (.A(_09456_),
    .X(_09457_));
 sg13g2_nor3_1 _16495_ (.A(net720),
    .B(_09427_),
    .C(_09439_),
    .Y(_00689_));
 sg13g2_nand2b_1 _16496_ (.Y(_09458_),
    .B(_08409_),
    .A_N(\rbzero.spi_registers.ss_buffer[1] ));
 sg13g2_buf_1 _16497_ (.A(_09458_),
    .X(_09459_));
 sg13g2_buf_1 _16498_ (.A(_09459_),
    .X(_09460_));
 sg13g2_buf_1 _16499_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_09461_));
 sg13g2_buf_1 _16500_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .X(_09462_));
 sg13g2_buf_2 _16501_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .X(_09463_));
 sg13g2_buf_1 _16502_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .X(_09464_));
 sg13g2_nand3b_1 _16503_ (.B(_09464_),
    .C(_00475_),
    .Y(_09465_),
    .A_N(_09463_));
 sg13g2_buf_1 _16504_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .X(_09466_));
 sg13g2_buf_1 _16505_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .X(_09467_));
 sg13g2_or4_1 _16506_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_09466_),
    .C(_09467_),
    .D(\rbzero.spi_registers.spi_counter[6] ),
    .X(_09468_));
 sg13g2_a21oi_1 _16507_ (.A1(_09462_),
    .A2(_09465_),
    .Y(_09469_),
    .B1(_09468_));
 sg13g2_nor2b_1 _16508_ (.A(\rbzero.spi_registers.sclk_buffer[2] ),
    .B_N(\rbzero.spi_registers.sclk_buffer[1] ),
    .Y(_09470_));
 sg13g2_nand2_1 _16509_ (.Y(_09471_),
    .A(_09469_),
    .B(_09470_));
 sg13g2_buf_2 _16510_ (.A(_09471_),
    .X(_09472_));
 sg13g2_mux2_1 _16511_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(net815),
    .S(_09472_),
    .X(_09473_));
 sg13g2_nor2b_1 _16512_ (.A(net719),
    .B_N(_09473_),
    .Y(_00930_));
 sg13g2_inv_1 _16513_ (.Y(_09474_),
    .A(net815));
 sg13g2_buf_1 _16514_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_09475_));
 sg13g2_buf_1 _16515_ (.A(_09475_),
    .X(_09476_));
 sg13g2_nand2_1 _16516_ (.Y(_09477_),
    .A(net757),
    .B(_09472_));
 sg13g2_o21ai_1 _16517_ (.B1(_09477_),
    .Y(_09478_),
    .A1(_09474_),
    .A2(_09472_));
 sg13g2_nor2b_1 _16518_ (.A(net719),
    .B_N(_09478_),
    .Y(_00931_));
 sg13g2_buf_1 _16519_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_09479_));
 sg13g2_buf_1 _16520_ (.A(_09479_),
    .X(_09480_));
 sg13g2_mux2_1 _16521_ (.A0(net757),
    .A1(net756),
    .S(_09472_),
    .X(_09481_));
 sg13g2_nor2b_1 _16522_ (.A(net719),
    .B_N(_09481_),
    .Y(_00932_));
 sg13g2_buf_2 _16523_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_09482_));
 sg13g2_mux2_1 _16524_ (.A0(net756),
    .A1(_09482_),
    .S(_09472_),
    .X(_09483_));
 sg13g2_nor2b_1 _16525_ (.A(net719),
    .B_N(_09483_),
    .Y(_00933_));
 sg13g2_inv_1 _16526_ (.Y(_09484_),
    .A(\rbzero.spi_registers.spi_counter[3] ));
 sg13g2_o21ai_1 _16527_ (.B1(net756),
    .Y(_09485_),
    .A1(net757),
    .A2(_09482_));
 sg13g2_and2_1 _16528_ (.A(net815),
    .B(net757),
    .X(_09486_));
 sg13g2_inv_1 _16529_ (.Y(_09487_),
    .A(_09482_));
 sg13g2_nor2_1 _16530_ (.A(_09475_),
    .B(net756),
    .Y(_09488_));
 sg13g2_a221oi_1 _16531_ (.B2(_09487_),
    .C1(_09488_),
    .B1(_09486_),
    .A1(_09474_),
    .Y(_09489_),
    .A2(_09485_));
 sg13g2_xnor2_1 _16532_ (.Y(_09490_),
    .A(_09484_),
    .B(_09489_));
 sg13g2_xor2_1 _16533_ (.B(net756),
    .A(net757),
    .X(_09491_));
 sg13g2_nand2_1 _16534_ (.Y(_09492_),
    .A(_09479_),
    .B(_09482_));
 sg13g2_nand2_1 _16535_ (.Y(_09493_),
    .A(_09462_),
    .B(_09492_));
 sg13g2_a21oi_1 _16536_ (.A1(net815),
    .A2(_09491_),
    .Y(_09494_),
    .B1(_09493_));
 sg13g2_nor4_1 _16537_ (.A(_09466_),
    .B(\rbzero.spi_registers.spi_counter[6] ),
    .C(_09469_),
    .D(_09494_),
    .Y(_09495_));
 sg13g2_mux2_1 _16538_ (.A0(_09479_),
    .A1(_09482_),
    .S(_09475_),
    .X(_09496_));
 sg13g2_a22oi_1 _16539_ (.Y(_09497_),
    .B1(_09496_),
    .B2(net815),
    .A2(_09482_),
    .A1(_09480_));
 sg13g2_nor2b_1 _16540_ (.A(_09482_),
    .B_N(_09475_),
    .Y(_09498_));
 sg13g2_nand2_1 _16541_ (.Y(_09499_),
    .A(_09464_),
    .B(_09498_));
 sg13g2_o21ai_1 _16542_ (.B1(_09499_),
    .Y(_09500_),
    .A1(_09464_),
    .A2(_09497_));
 sg13g2_a22oi_1 _16543_ (.Y(_09501_),
    .B1(_09492_),
    .B2(_09474_),
    .A2(_09498_),
    .A1(net756));
 sg13g2_nand2b_1 _16544_ (.Y(_09502_),
    .B(_09501_),
    .A_N(_09488_));
 sg13g2_a22oi_1 _16545_ (.Y(_09503_),
    .B1(_09502_),
    .B2(_09464_),
    .A2(_09500_),
    .A1(_09462_));
 sg13g2_inv_1 _16546_ (.Y(_09504_),
    .A(_09503_));
 sg13g2_nor2_1 _16547_ (.A(_09479_),
    .B(_09482_),
    .Y(_09505_));
 sg13g2_nand2_1 _16548_ (.Y(_09506_),
    .A(_09463_),
    .B(_09505_));
 sg13g2_o21ai_1 _16549_ (.B1(_09506_),
    .Y(_09507_),
    .A1(_09487_),
    .A2(_09463_));
 sg13g2_o21ai_1 _16550_ (.B1(_09475_),
    .Y(_09508_),
    .A1(net815),
    .A2(_09479_));
 sg13g2_nand2_1 _16551_ (.Y(_09509_),
    .A(_09487_),
    .B(_09508_));
 sg13g2_a21oi_1 _16552_ (.A1(_09492_),
    .A2(_09509_),
    .Y(_09510_),
    .B1(_09463_));
 sg13g2_a21oi_1 _16553_ (.A1(_09486_),
    .A2(_09507_),
    .Y(_09511_),
    .B1(_09510_));
 sg13g2_nand2_1 _16554_ (.Y(_09512_),
    .A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_09475_));
 sg13g2_buf_1 _16555_ (.A(_09512_),
    .X(_09513_));
 sg13g2_nor2_1 _16556_ (.A(net756),
    .B(_09487_),
    .Y(_09514_));
 sg13g2_a22oi_1 _16557_ (.Y(_09515_),
    .B1(_09513_),
    .B2(_09514_),
    .A2(_09498_),
    .A1(_09480_));
 sg13g2_nand3b_1 _16558_ (.B(_09467_),
    .C(_09463_),
    .Y(_09516_),
    .A_N(_09515_));
 sg13g2_o21ai_1 _16559_ (.B1(_09516_),
    .Y(_09517_),
    .A1(_09467_),
    .A2(_09511_));
 sg13g2_nand4_1 _16560_ (.B(_09495_),
    .C(_09504_),
    .A(_09490_),
    .Y(_09518_),
    .D(_09517_));
 sg13g2_and2_1 _16561_ (.A(_09470_),
    .B(_09518_),
    .X(_09519_));
 sg13g2_buf_1 _16562_ (.A(_09519_),
    .X(_09520_));
 sg13g2_nand2_1 _16563_ (.Y(_09521_),
    .A(_00475_),
    .B(_09520_));
 sg13g2_nand2b_1 _16564_ (.Y(_09522_),
    .B(_09464_),
    .A_N(_09520_));
 sg13g2_a21oi_1 _16565_ (.A1(_09521_),
    .A2(_09522_),
    .Y(_00934_),
    .B1(_09459_));
 sg13g2_and2_1 _16566_ (.A(_09464_),
    .B(_09520_),
    .X(_09523_));
 sg13g2_buf_1 _16567_ (.A(_09523_),
    .X(_09524_));
 sg13g2_xnor2_1 _16568_ (.Y(_09525_),
    .A(_09463_),
    .B(_09524_));
 sg13g2_nor2_1 _16569_ (.A(net719),
    .B(_09525_),
    .Y(_00935_));
 sg13g2_nand2_1 _16570_ (.Y(_09526_),
    .A(_09463_),
    .B(_09524_));
 sg13g2_xor2_1 _16571_ (.B(_09526_),
    .A(_09462_),
    .X(_09527_));
 sg13g2_nor2_1 _16572_ (.A(net719),
    .B(_09527_),
    .Y(_00936_));
 sg13g2_nand3_1 _16573_ (.B(_09463_),
    .C(_09524_),
    .A(_09462_),
    .Y(_09528_));
 sg13g2_xnor2_1 _16574_ (.Y(_09529_),
    .A(_09484_),
    .B(_09528_));
 sg13g2_nor2_1 _16575_ (.A(_09460_),
    .B(_09529_),
    .Y(_00937_));
 sg13g2_nor2_1 _16576_ (.A(_09484_),
    .B(_09528_),
    .Y(_09530_));
 sg13g2_xnor2_1 _16577_ (.Y(_09531_),
    .A(_09467_),
    .B(_09530_));
 sg13g2_nor2_1 _16578_ (.A(_09460_),
    .B(_09531_),
    .Y(_00938_));
 sg13g2_nand2_1 _16579_ (.Y(_09532_),
    .A(_09467_),
    .B(_09530_));
 sg13g2_xor2_1 _16580_ (.B(_09532_),
    .A(_09466_),
    .X(_09533_));
 sg13g2_nor2_1 _16581_ (.A(net719),
    .B(_09533_),
    .Y(_00939_));
 sg13g2_nand3_1 _16582_ (.B(_09467_),
    .C(_09530_),
    .A(_09466_),
    .Y(_09534_));
 sg13g2_xor2_1 _16583_ (.B(_09534_),
    .A(\rbzero.spi_registers.spi_counter[6] ),
    .X(_09535_));
 sg13g2_nor2_1 _16584_ (.A(net719),
    .B(_09535_),
    .Y(_00940_));
 sg13g2_buf_1 _16585_ (.A(\rbzero.spi_registers.spi_done ),
    .X(_09536_));
 sg13g2_nand2b_1 _16586_ (.Y(_09537_),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .A_N(\rbzero.spi_registers.sclk_buffer[2] ));
 sg13g2_nor4_1 _16587_ (.A(_09536_),
    .B(_09459_),
    .C(_09537_),
    .D(_09518_),
    .Y(_00941_));
 sg13g2_buf_1 _16588_ (.A(_08678_),
    .X(_09538_));
 sg13g2_buf_1 _16589_ (.A(\rbzero.texV[-11] ),
    .X(_09539_));
 sg13g2_buf_1 _16590_ (.A(\rbzero.traced_texa[-11] ),
    .X(_09540_));
 sg13g2_xnor2_1 _16591_ (.Y(_09541_),
    .A(_09539_),
    .B(_09540_));
 sg13g2_nor2_1 _16592_ (.A(_09538_),
    .B(_09541_),
    .Y(_01047_));
 sg13g2_buf_1 _16593_ (.A(\rbzero.traced_texa[-2] ),
    .X(_09542_));
 sg13g2_buf_1 _16594_ (.A(\rbzero.traced_texa[-3] ),
    .X(_09543_));
 sg13g2_inv_1 _16595_ (.Y(_09544_),
    .A(_09543_));
 sg13g2_buf_1 _16596_ (.A(\rbzero.traced_texa[-4] ),
    .X(_09545_));
 sg13g2_buf_1 _16597_ (.A(\rbzero.traced_texa[-5] ),
    .X(_09546_));
 sg13g2_inv_1 _16598_ (.Y(_09547_),
    .A(_09546_));
 sg13g2_buf_1 _16599_ (.A(\rbzero.traced_texa[-6] ),
    .X(_09548_));
 sg13g2_buf_1 _16600_ (.A(\rbzero.traced_texa[-7] ),
    .X(_09549_));
 sg13g2_inv_1 _16601_ (.Y(_09550_),
    .A(_09549_));
 sg13g2_buf_1 _16602_ (.A(\rbzero.traced_texa[-8] ),
    .X(_09551_));
 sg13g2_buf_1 _16603_ (.A(\rbzero.traced_texa[-9] ),
    .X(_09552_));
 sg13g2_inv_1 _16604_ (.Y(_09553_),
    .A(\rbzero.texV[-10] ));
 sg13g2_buf_1 _16605_ (.A(\rbzero.traced_texa[-10] ),
    .X(_09554_));
 sg13g2_a21oi_1 _16606_ (.A1(_09539_),
    .A2(_09540_),
    .Y(_09555_),
    .B1(_09554_));
 sg13g2_nand3_1 _16607_ (.B(_09540_),
    .C(_09554_),
    .A(_09539_),
    .Y(_09556_));
 sg13g2_o21ai_1 _16608_ (.B1(_09556_),
    .Y(_09557_),
    .A1(_09553_),
    .A2(_09555_));
 sg13g2_buf_1 _16609_ (.A(_09557_),
    .X(_09558_));
 sg13g2_nor2_1 _16610_ (.A(_09552_),
    .B(_09558_),
    .Y(_09559_));
 sg13g2_a21oi_1 _16611_ (.A1(_09552_),
    .A2(_09558_),
    .Y(_09560_),
    .B1(\rbzero.texV[-9] ));
 sg13g2_nor2_1 _16612_ (.A(_09559_),
    .B(_09560_),
    .Y(_09561_));
 sg13g2_a21o_1 _16613_ (.A2(_09561_),
    .A1(_09551_),
    .B1(\rbzero.texV[-8] ),
    .X(_09562_));
 sg13g2_o21ai_1 _16614_ (.B1(_09562_),
    .Y(_09563_),
    .A1(_09551_),
    .A2(_09561_));
 sg13g2_buf_1 _16615_ (.A(_09563_),
    .X(_09564_));
 sg13g2_inv_1 _16616_ (.Y(_09565_),
    .A(_09564_));
 sg13g2_a21oi_1 _16617_ (.A1(_09549_),
    .A2(_09565_),
    .Y(_09566_),
    .B1(\rbzero.texV[-7] ));
 sg13g2_a21oi_2 _16618_ (.B1(_09566_),
    .Y(_09567_),
    .A2(_09564_),
    .A1(_09550_));
 sg13g2_a21o_1 _16619_ (.A2(_09567_),
    .A1(_09548_),
    .B1(\rbzero.texV[-6] ),
    .X(_09568_));
 sg13g2_o21ai_1 _16620_ (.B1(_09568_),
    .Y(_09569_),
    .A1(_09548_),
    .A2(_09567_));
 sg13g2_buf_1 _16621_ (.A(_09569_),
    .X(_09570_));
 sg13g2_inv_1 _16622_ (.Y(_09571_),
    .A(_09570_));
 sg13g2_a21oi_1 _16623_ (.A1(_09546_),
    .A2(_09571_),
    .Y(_09572_),
    .B1(\rbzero.texV[-5] ));
 sg13g2_a21oi_2 _16624_ (.B1(_09572_),
    .Y(_09573_),
    .A2(_09570_),
    .A1(_09547_));
 sg13g2_a21o_1 _16625_ (.A2(_09573_),
    .A1(_09545_),
    .B1(\rbzero.texV[-4] ),
    .X(_09574_));
 sg13g2_o21ai_1 _16626_ (.B1(_09574_),
    .Y(_09575_),
    .A1(_09545_),
    .A2(_09573_));
 sg13g2_buf_1 _16627_ (.A(_09575_),
    .X(_09576_));
 sg13g2_inv_1 _16628_ (.Y(_09577_),
    .A(_09576_));
 sg13g2_a21oi_1 _16629_ (.A1(_09543_),
    .A2(_09577_),
    .Y(_09578_),
    .B1(\rbzero.texV[-3] ));
 sg13g2_a21oi_2 _16630_ (.B1(_09578_),
    .Y(_09579_),
    .A2(_09576_),
    .A1(_09544_));
 sg13g2_a21o_1 _16631_ (.A2(_09579_),
    .A1(_09542_),
    .B1(\rbzero.texV[-2] ),
    .X(_09580_));
 sg13g2_o21ai_1 _16632_ (.B1(_09580_),
    .Y(_09581_),
    .A1(_09542_),
    .A2(_09579_));
 sg13g2_buf_1 _16633_ (.A(_09581_),
    .X(_09582_));
 sg13g2_buf_1 _16634_ (.A(\rbzero.traced_texa[-1] ),
    .X(_09583_));
 sg13g2_xnor2_1 _16635_ (.Y(_09584_),
    .A(\rbzero.texV[-1] ),
    .B(_09583_));
 sg13g2_xnor2_1 _16636_ (.Y(_09585_),
    .A(_09582_),
    .B(_09584_));
 sg13g2_nor2_1 _16637_ (.A(net473),
    .B(_09585_),
    .Y(_01048_));
 sg13g2_inv_1 _16638_ (.Y(_09586_),
    .A(_09583_));
 sg13g2_inv_1 _16639_ (.Y(_09587_),
    .A(_09582_));
 sg13g2_a21oi_1 _16640_ (.A1(_09583_),
    .A2(_09587_),
    .Y(_09588_),
    .B1(\rbzero.texV[-1] ));
 sg13g2_a21oi_2 _16641_ (.B1(_09588_),
    .Y(_09589_),
    .A2(_09582_),
    .A1(_09586_));
 sg13g2_buf_1 _16642_ (.A(\rbzero.texV[0] ),
    .X(_09590_));
 sg13g2_buf_1 _16643_ (.A(\rbzero.traced_texa[0] ),
    .X(_09591_));
 sg13g2_xor2_1 _16644_ (.B(_09591_),
    .A(_09590_),
    .X(_09592_));
 sg13g2_xnor2_1 _16645_ (.Y(_09593_),
    .A(_09589_),
    .B(_09592_));
 sg13g2_nor2_1 _16646_ (.A(_09538_),
    .B(_09593_),
    .Y(_01049_));
 sg13g2_buf_1 _16647_ (.A(\rbzero.texV[1] ),
    .X(_09594_));
 sg13g2_buf_1 _16648_ (.A(\rbzero.traced_texa[1] ),
    .X(_09595_));
 sg13g2_xnor2_1 _16649_ (.Y(_09596_),
    .A(_09594_),
    .B(_09595_));
 sg13g2_a21o_1 _16650_ (.A2(_09589_),
    .A1(_09591_),
    .B1(_09590_),
    .X(_09597_));
 sg13g2_o21ai_1 _16651_ (.B1(_09597_),
    .Y(_09598_),
    .A1(_09591_),
    .A2(_09589_));
 sg13g2_xnor2_1 _16652_ (.Y(_09599_),
    .A(_09596_),
    .B(_09598_));
 sg13g2_nor2_1 _16653_ (.A(net473),
    .B(_09599_),
    .Y(_01050_));
 sg13g2_nor2_1 _16654_ (.A(_09594_),
    .B(_09595_),
    .Y(_09600_));
 sg13g2_nand2_1 _16655_ (.Y(_09601_),
    .A(_09594_),
    .B(_09595_));
 sg13g2_o21ai_1 _16656_ (.B1(_09601_),
    .Y(_09602_),
    .A1(_09600_),
    .A2(_09598_));
 sg13g2_buf_1 _16657_ (.A(_09602_),
    .X(_09603_));
 sg13g2_buf_1 _16658_ (.A(\rbzero.texV[2] ),
    .X(_09604_));
 sg13g2_buf_1 _16659_ (.A(\rbzero.traced_texa[2] ),
    .X(_09605_));
 sg13g2_xor2_1 _16660_ (.B(_09605_),
    .A(_09604_),
    .X(_09606_));
 sg13g2_xnor2_1 _16661_ (.Y(_09607_),
    .A(_09603_),
    .B(_09606_));
 sg13g2_nor2_1 _16662_ (.A(net473),
    .B(_09607_),
    .Y(_01051_));
 sg13g2_a21o_1 _16663_ (.A2(_09603_),
    .A1(_09605_),
    .B1(_09604_),
    .X(_09608_));
 sg13g2_o21ai_1 _16664_ (.B1(_09608_),
    .Y(_09609_),
    .A1(_09605_),
    .A2(_09603_));
 sg13g2_buf_1 _16665_ (.A(_09609_),
    .X(_09610_));
 sg13g2_buf_1 _16666_ (.A(\rbzero.texV[3] ),
    .X(_09611_));
 sg13g2_buf_1 _16667_ (.A(\rbzero.traced_texa[3] ),
    .X(_09612_));
 sg13g2_xnor2_1 _16668_ (.Y(_09613_),
    .A(_09611_),
    .B(_09612_));
 sg13g2_xnor2_1 _16669_ (.Y(_09614_),
    .A(_09610_),
    .B(_09613_));
 sg13g2_nor2_1 _16670_ (.A(net473),
    .B(_09614_),
    .Y(_01052_));
 sg13g2_inv_1 _16671_ (.Y(_09615_),
    .A(_09612_));
 sg13g2_inv_1 _16672_ (.Y(_09616_),
    .A(_09610_));
 sg13g2_a21oi_1 _16673_ (.A1(_09612_),
    .A2(_09616_),
    .Y(_09617_),
    .B1(_09611_));
 sg13g2_a21oi_2 _16674_ (.B1(_09617_),
    .Y(_09618_),
    .A2(_09610_),
    .A1(_09615_));
 sg13g2_buf_1 _16675_ (.A(\rbzero.texV[4] ),
    .X(_09619_));
 sg13g2_buf_1 _16676_ (.A(\rbzero.traced_texa[4] ),
    .X(_09620_));
 sg13g2_xor2_1 _16677_ (.B(_09620_),
    .A(_09619_),
    .X(_09621_));
 sg13g2_xnor2_1 _16678_ (.Y(_09622_),
    .A(_09618_),
    .B(_09621_));
 sg13g2_nor2_1 _16679_ (.A(net473),
    .B(_09622_),
    .Y(_01053_));
 sg13g2_a21o_1 _16680_ (.A2(_09618_),
    .A1(_09620_),
    .B1(_09619_),
    .X(_09623_));
 sg13g2_o21ai_1 _16681_ (.B1(_09623_),
    .Y(_09624_),
    .A1(_09620_),
    .A2(_09618_));
 sg13g2_buf_1 _16682_ (.A(_09624_),
    .X(_09625_));
 sg13g2_buf_1 _16683_ (.A(\rbzero.texV[5] ),
    .X(_09626_));
 sg13g2_buf_1 _16684_ (.A(_09626_),
    .X(_09627_));
 sg13g2_buf_1 _16685_ (.A(\rbzero.traced_texa[5] ),
    .X(_09628_));
 sg13g2_xnor2_1 _16686_ (.Y(_09629_),
    .A(net755),
    .B(_09628_));
 sg13g2_xnor2_1 _16687_ (.Y(_09630_),
    .A(_09625_),
    .B(_09629_));
 sg13g2_nor2_1 _16688_ (.A(net473),
    .B(_09630_),
    .Y(_01054_));
 sg13g2_buf_2 _16689_ (.A(\rbzero.texV[6] ),
    .X(_09631_));
 sg13g2_buf_1 _16690_ (.A(\rbzero.traced_texa[6] ),
    .X(_09632_));
 sg13g2_xor2_1 _16691_ (.B(_09632_),
    .A(_09631_),
    .X(_09633_));
 sg13g2_nor2_1 _16692_ (.A(net755),
    .B(_09628_),
    .Y(_09634_));
 sg13g2_nand2_1 _16693_ (.Y(_09635_),
    .A(net755),
    .B(_09628_));
 sg13g2_o21ai_1 _16694_ (.B1(_09635_),
    .Y(_09636_),
    .A1(_09625_),
    .A2(_09634_));
 sg13g2_xnor2_1 _16695_ (.Y(_09637_),
    .A(_09633_),
    .B(_09636_));
 sg13g2_nor2_1 _16696_ (.A(net473),
    .B(_09637_),
    .Y(_01055_));
 sg13g2_inv_1 _16697_ (.Y(_09638_),
    .A(_09631_));
 sg13g2_inv_1 _16698_ (.Y(_09639_),
    .A(_09632_));
 sg13g2_a21oi_1 _16699_ (.A1(_09631_),
    .A2(_09632_),
    .Y(_09640_),
    .B1(_09636_));
 sg13g2_a21oi_1 _16700_ (.A1(_09638_),
    .A2(_09639_),
    .Y(_09641_),
    .B1(_09640_));
 sg13g2_buf_2 _16701_ (.A(\rbzero.texV[7] ),
    .X(_09642_));
 sg13g2_buf_2 _16702_ (.A(\rbzero.traced_texa[7] ),
    .X(_09643_));
 sg13g2_xnor2_1 _16703_ (.Y(_09644_),
    .A(_09642_),
    .B(_09643_));
 sg13g2_xnor2_1 _16704_ (.Y(_09645_),
    .A(_09641_),
    .B(_09644_));
 sg13g2_and2_1 _16705_ (.A(_08473_),
    .B(_09645_),
    .X(_01056_));
 sg13g2_buf_2 _16706_ (.A(\rbzero.texV[8] ),
    .X(_09646_));
 sg13g2_buf_1 _16707_ (.A(\rbzero.traced_texa[8] ),
    .X(_09647_));
 sg13g2_xnor2_1 _16708_ (.Y(_09648_),
    .A(_09646_),
    .B(_09647_));
 sg13g2_o21ai_1 _16709_ (.B1(_09641_),
    .Y(_09649_),
    .A1(_09642_),
    .A2(_09643_));
 sg13g2_inv_1 _16710_ (.Y(_09650_),
    .A(_09649_));
 sg13g2_a21oi_1 _16711_ (.A1(_09642_),
    .A2(_09643_),
    .Y(_09651_),
    .B1(_09650_));
 sg13g2_xnor2_1 _16712_ (.Y(_09652_),
    .A(_09648_),
    .B(_09651_));
 sg13g2_nor2_1 _16713_ (.A(net473),
    .B(_09652_),
    .Y(_01057_));
 sg13g2_buf_1 _16714_ (.A(net490),
    .X(_09653_));
 sg13g2_nand2_1 _16715_ (.Y(_09654_),
    .A(_09539_),
    .B(_09540_));
 sg13g2_xnor2_1 _16716_ (.Y(_09655_),
    .A(\rbzero.texV[-10] ),
    .B(_09554_));
 sg13g2_xnor2_1 _16717_ (.Y(_09656_),
    .A(_09654_),
    .B(_09655_));
 sg13g2_nor2_1 _16718_ (.A(net472),
    .B(_09656_),
    .Y(_01058_));
 sg13g2_nor2_1 _16719_ (.A(_09644_),
    .B(_09648_),
    .Y(_09657_));
 sg13g2_nand3b_1 _16720_ (.B(_09633_),
    .C(_09657_),
    .Y(_09658_),
    .A_N(_09629_));
 sg13g2_a21oi_1 _16721_ (.A1(_09627_),
    .A2(_09628_),
    .Y(_09659_),
    .B1(_09632_));
 sg13g2_nand3_1 _16722_ (.B(_09628_),
    .C(_09632_),
    .A(_09627_),
    .Y(_09660_));
 sg13g2_o21ai_1 _16723_ (.B1(_09660_),
    .Y(_09661_),
    .A1(_09638_),
    .A2(_09659_));
 sg13g2_a21oi_1 _16724_ (.A1(_09643_),
    .A2(_09661_),
    .Y(_09662_),
    .B1(_09642_));
 sg13g2_nor2_1 _16725_ (.A(_09643_),
    .B(_09661_),
    .Y(_09663_));
 sg13g2_nand2_1 _16726_ (.Y(_09664_),
    .A(_09646_),
    .B(_09647_));
 sg13g2_o21ai_1 _16727_ (.B1(_09664_),
    .Y(_09665_),
    .A1(_09662_),
    .A2(_09663_));
 sg13g2_o21ai_1 _16728_ (.B1(_09665_),
    .Y(_09666_),
    .A1(_09646_),
    .A2(_09647_));
 sg13g2_o21ai_1 _16729_ (.B1(_09666_),
    .Y(_09667_),
    .A1(_09625_),
    .A2(_09658_));
 sg13g2_buf_1 _16730_ (.A(\rbzero.texV[9] ),
    .X(_09668_));
 sg13g2_buf_1 _16731_ (.A(\rbzero.traced_texa[9] ),
    .X(_09669_));
 sg13g2_xor2_1 _16732_ (.B(_09669_),
    .A(_09668_),
    .X(_09670_));
 sg13g2_xnor2_1 _16733_ (.Y(_09671_),
    .A(_09667_),
    .B(_09670_));
 sg13g2_nor2_1 _16734_ (.A(net472),
    .B(_09671_),
    .Y(_01059_));
 sg13g2_xor2_1 _16735_ (.B(\rbzero.traced_texa[10] ),
    .A(\rbzero.texV[10] ),
    .X(_09672_));
 sg13g2_nand2_1 _16736_ (.Y(_09673_),
    .A(_09668_),
    .B(_09669_));
 sg13g2_o21ai_1 _16737_ (.B1(_09667_),
    .Y(_09674_),
    .A1(_09668_),
    .A2(_09669_));
 sg13g2_nand2_1 _16738_ (.Y(_09675_),
    .A(_09673_),
    .B(_09674_));
 sg13g2_xnor2_1 _16739_ (.Y(_09676_),
    .A(_09672_),
    .B(_09675_));
 sg13g2_nor2_1 _16740_ (.A(net472),
    .B(_09676_),
    .Y(_01060_));
 sg13g2_xor2_1 _16741_ (.B(_09552_),
    .A(\rbzero.texV[-9] ),
    .X(_09677_));
 sg13g2_xnor2_1 _16742_ (.Y(_09678_),
    .A(_09558_),
    .B(_09677_));
 sg13g2_nor2_1 _16743_ (.A(net472),
    .B(_09678_),
    .Y(_01061_));
 sg13g2_xor2_1 _16744_ (.B(_09551_),
    .A(\rbzero.texV[-8] ),
    .X(_09679_));
 sg13g2_xnor2_1 _16745_ (.Y(_09680_),
    .A(_09561_),
    .B(_09679_));
 sg13g2_nor2_1 _16746_ (.A(net472),
    .B(_09680_),
    .Y(_01062_));
 sg13g2_xnor2_1 _16747_ (.Y(_09681_),
    .A(\rbzero.texV[-7] ),
    .B(_09549_));
 sg13g2_xnor2_1 _16748_ (.Y(_09682_),
    .A(_09564_),
    .B(_09681_));
 sg13g2_nor2_1 _16749_ (.A(net472),
    .B(_09682_),
    .Y(_01063_));
 sg13g2_xor2_1 _16750_ (.B(_09548_),
    .A(\rbzero.texV[-6] ),
    .X(_09683_));
 sg13g2_xnor2_1 _16751_ (.Y(_09684_),
    .A(_09567_),
    .B(_09683_));
 sg13g2_nor2_1 _16752_ (.A(net472),
    .B(_09684_),
    .Y(_01064_));
 sg13g2_xnor2_1 _16753_ (.Y(_09685_),
    .A(\rbzero.texV[-5] ),
    .B(_09546_));
 sg13g2_xnor2_1 _16754_ (.Y(_09686_),
    .A(_09570_),
    .B(_09685_));
 sg13g2_nor2_1 _16755_ (.A(_09653_),
    .B(_09686_),
    .Y(_01065_));
 sg13g2_xor2_1 _16756_ (.B(_09545_),
    .A(\rbzero.texV[-4] ),
    .X(_09687_));
 sg13g2_xnor2_1 _16757_ (.Y(_09688_),
    .A(_09573_),
    .B(_09687_));
 sg13g2_nor2_1 _16758_ (.A(_09653_),
    .B(_09688_),
    .Y(_01066_));
 sg13g2_xnor2_1 _16759_ (.Y(_09689_),
    .A(\rbzero.texV[-3] ),
    .B(_09543_));
 sg13g2_xnor2_1 _16760_ (.Y(_09690_),
    .A(_09576_),
    .B(_09689_));
 sg13g2_nor2_1 _16761_ (.A(net472),
    .B(_09690_),
    .Y(_01067_));
 sg13g2_xor2_1 _16762_ (.B(_09542_),
    .A(\rbzero.texV[-2] ),
    .X(_09691_));
 sg13g2_xnor2_1 _16763_ (.Y(_09692_),
    .A(_09579_),
    .B(_09691_));
 sg13g2_nor2_1 _16764_ (.A(net490),
    .B(_09692_),
    .Y(_01068_));
 sg13g2_inv_1 _16765_ (.Y(_09693_),
    .A(\rbzero.debug_overlay.h[0] ));
 sg13g2_nand2_1 _16766_ (.Y(_09694_),
    .A(_08409_),
    .B(_08473_));
 sg13g2_buf_2 _16767_ (.A(_09694_),
    .X(_09695_));
 sg13g2_nor2_1 _16768_ (.A(_09693_),
    .B(_09695_),
    .Y(_01453_));
 sg13g2_inv_2 _16769_ (.Y(_09696_),
    .A(_08458_));
 sg13g2_nand2_1 _16770_ (.Y(_09697_),
    .A(_09696_),
    .B(net723));
 sg13g2_buf_1 _16771_ (.A(_08458_),
    .X(_09698_));
 sg13g2_nand2b_1 _16772_ (.Y(_09699_),
    .B(net754),
    .A_N(net783));
 sg13g2_a21oi_1 _16773_ (.A1(_09697_),
    .A2(_09699_),
    .Y(_01454_),
    .B1(_09695_));
 sg13g2_buf_1 _16774_ (.A(_08638_),
    .X(_09700_));
 sg13g2_buf_1 _16775_ (.A(_09700_),
    .X(_09701_));
 sg13g2_buf_1 _16776_ (.A(net675),
    .X(_09702_));
 sg13g2_nand2_1 _16777_ (.Y(_09703_),
    .A(net754),
    .B(net723));
 sg13g2_xor2_1 _16778_ (.B(_09703_),
    .A(net829),
    .X(_09704_));
 sg13g2_nor2_1 _16779_ (.A(net607),
    .B(_09704_),
    .Y(_01455_));
 sg13g2_xnor2_1 _16780_ (.Y(_09705_),
    .A(_00014_),
    .B(_08461_));
 sg13g2_nor2_1 _16781_ (.A(_09695_),
    .B(_09705_),
    .Y(_01456_));
 sg13g2_xnor2_1 _16782_ (.Y(_09706_),
    .A(_08453_),
    .B(_08462_));
 sg13g2_buf_1 _16783_ (.A(_09706_),
    .X(_09707_));
 sg13g2_nor2_1 _16784_ (.A(_09695_),
    .B(_09707_),
    .Y(_01457_));
 sg13g2_xnor2_1 _16785_ (.Y(_09708_),
    .A(net786),
    .B(_08464_));
 sg13g2_nor2_1 _16786_ (.A(_09695_),
    .B(_09708_),
    .Y(_01458_));
 sg13g2_inv_2 _16787_ (.Y(_09709_),
    .A(_08465_));
 sg13g2_nand2_1 _16788_ (.Y(_09710_),
    .A(net786),
    .B(_08464_));
 sg13g2_xnor2_1 _16789_ (.Y(_09711_),
    .A(_09709_),
    .B(_09710_));
 sg13g2_nor2_1 _16790_ (.A(_09695_),
    .B(_09711_),
    .Y(_01459_));
 sg13g2_nand3_1 _16791_ (.B(_08663_),
    .C(_08464_),
    .A(net786),
    .Y(_09712_));
 sg13g2_xor2_1 _16792_ (.B(_09712_),
    .A(net787),
    .X(_09713_));
 sg13g2_nor2_1 _16793_ (.A(net607),
    .B(_09713_),
    .Y(_01460_));
 sg13g2_nand4_1 _16794_ (.B(_08663_),
    .C(net787),
    .A(_08651_),
    .Y(_09714_),
    .D(_08464_));
 sg13g2_xnor2_1 _16795_ (.Y(_09715_),
    .A(_08655_),
    .B(_09714_));
 sg13g2_nor2_1 _16796_ (.A(_09695_),
    .B(_09715_),
    .Y(_01461_));
 sg13g2_or2_1 _16797_ (.X(_09716_),
    .B(_09714_),
    .A(_08655_));
 sg13g2_xnor2_1 _16798_ (.Y(_09717_),
    .A(_08470_),
    .B(_09716_));
 sg13g2_nor2_1 _16799_ (.A(_09695_),
    .B(_09717_),
    .Y(_01462_));
 sg13g2_nor3_1 _16800_ (.A(net829),
    .B(_09698_),
    .C(_08459_),
    .Y(_09718_));
 sg13g2_and4_1 _16801_ (.A(_08456_),
    .B(net787),
    .C(_08469_),
    .D(_08655_),
    .X(_09719_));
 sg13g2_nand3_1 _16802_ (.B(_09718_),
    .C(_09719_),
    .A(net796),
    .Y(_09720_));
 sg13g2_nor2_1 _16803_ (.A(net785),
    .B(_09720_),
    .Y(_09721_));
 sg13g2_o21ai_1 _16804_ (.B1(_08683_),
    .Y(_09722_),
    .A1(\rbzero.hsync ),
    .A2(_09721_));
 sg13g2_o21ai_1 _16805_ (.B1(\rbzero.hsync ),
    .Y(_09723_),
    .A1(_09709_),
    .A2(_09720_));
 sg13g2_buf_1 _16806_ (.A(_09700_),
    .X(_09724_));
 sg13g2_a21oi_1 _16807_ (.A1(_09722_),
    .A2(_09723_),
    .Y(_01463_),
    .B1(net674));
 sg13g2_inv_1 _16808_ (.Y(_09725_),
    .A(_09398_));
 sg13g2_buf_1 _16809_ (.A(_09402_),
    .X(_09726_));
 sg13g2_nor4_1 _16810_ (.A(_09725_),
    .B(net753),
    .C(_09399_),
    .D(_09414_),
    .Y(_09727_));
 sg13g2_inv_1 _16811_ (.Y(_09728_),
    .A(_09400_));
 sg13g2_nor4_1 _16812_ (.A(_09728_),
    .B(net816),
    .C(_09404_),
    .D(_09405_),
    .Y(_09729_));
 sg13g2_a21oi_1 _16813_ (.A1(_09727_),
    .A2(_09729_),
    .Y(_09730_),
    .B1(\rbzero.vga_sync.vsync ));
 sg13g2_nor2_1 _16814_ (.A(_09400_),
    .B(net816),
    .Y(_09731_));
 sg13g2_and3_1 _16815_ (.X(_09732_),
    .A(_09407_),
    .B(_09727_),
    .C(_09731_));
 sg13g2_nor3_1 _16816_ (.A(_09701_),
    .B(_09730_),
    .C(_09732_),
    .Y(_01474_));
 sg13g2_nor4_1 _16817_ (.A(_09398_),
    .B(_09399_),
    .C(_09410_),
    .D(_09414_),
    .Y(_09733_));
 sg13g2_and3_1 _16818_ (.X(_09734_),
    .A(\rbzero.pov.ready ),
    .B(_09733_),
    .C(_09417_));
 sg13g2_buf_1 _16819_ (.A(_09734_),
    .X(_09735_));
 sg13g2_buf_1 _16820_ (.A(_09735_),
    .X(_09736_));
 sg13g2_buf_1 _16821_ (.A(net388),
    .X(_09737_));
 sg13g2_nand2_1 _16822_ (.Y(_09738_),
    .A(\rbzero.pov.ready_buffer[33] ),
    .B(net358));
 sg13g2_buf_1 _16823_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .X(_09739_));
 sg13g2_buf_1 _16824_ (.A(_09733_),
    .X(_09740_));
 sg13g2_nand3_1 _16825_ (.B(net451),
    .C(_09417_),
    .A(\rbzero.pov.ready ),
    .Y(_09741_));
 sg13g2_buf_2 _16826_ (.A(_09741_),
    .X(_09742_));
 sg13g2_buf_1 _16827_ (.A(_09742_),
    .X(_09743_));
 sg13g2_nand2_1 _16828_ (.Y(_09744_),
    .A(_09739_),
    .B(_09743_));
 sg13g2_a21oi_1 _16829_ (.A1(_09738_),
    .A2(_09744_),
    .Y(_00476_),
    .B1(net674));
 sg13g2_buf_1 _16830_ (.A(net388),
    .X(_09745_));
 sg13g2_nand2_1 _16831_ (.Y(_09746_),
    .A(\rbzero.pov.ready_buffer[43] ),
    .B(net356));
 sg13g2_buf_2 _16832_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .X(_09747_));
 sg13g2_buf_1 _16833_ (.A(_09742_),
    .X(_09748_));
 sg13g2_nand2_1 _16834_ (.Y(_09749_),
    .A(_09747_),
    .B(_09748_));
 sg13g2_a21oi_1 _16835_ (.A1(_09746_),
    .A2(_09749_),
    .Y(_00477_),
    .B1(net674));
 sg13g2_nand2_1 _16836_ (.Y(_09750_),
    .A(\rbzero.pov.ready_buffer[34] ),
    .B(net356));
 sg13g2_buf_2 _16837_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .X(_09751_));
 sg13g2_nand2_1 _16838_ (.Y(_09752_),
    .A(_09751_),
    .B(net355));
 sg13g2_a21oi_1 _16839_ (.A1(_09750_),
    .A2(_09752_),
    .Y(_00478_),
    .B1(net674));
 sg13g2_nand2_1 _16840_ (.Y(_09753_),
    .A(\rbzero.pov.ready_buffer[35] ),
    .B(net356));
 sg13g2_buf_2 _16841_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .X(_09754_));
 sg13g2_nand2_1 _16842_ (.Y(_09755_),
    .A(_09754_),
    .B(net355));
 sg13g2_a21oi_1 _16843_ (.A1(_09753_),
    .A2(_09755_),
    .Y(_00479_),
    .B1(net674));
 sg13g2_nand2_1 _16844_ (.Y(_09756_),
    .A(\rbzero.pov.ready_buffer[36] ),
    .B(net356));
 sg13g2_buf_1 _16845_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .X(_09757_));
 sg13g2_nand2_1 _16846_ (.Y(_09758_),
    .A(_09757_),
    .B(net355));
 sg13g2_buf_1 _16847_ (.A(_09700_),
    .X(_09759_));
 sg13g2_buf_1 _16848_ (.A(_09759_),
    .X(_09760_));
 sg13g2_a21oi_1 _16849_ (.A1(_09756_),
    .A2(_09758_),
    .Y(_00480_),
    .B1(net606));
 sg13g2_buf_1 _16850_ (.A(_09424_),
    .X(_09761_));
 sg13g2_buf_1 _16851_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .X(_09762_));
 sg13g2_buf_1 _16852_ (.A(_09742_),
    .X(_09763_));
 sg13g2_nand2_1 _16853_ (.Y(_09764_),
    .A(_09762_),
    .B(net354));
 sg13g2_buf_1 _16854_ (.A(net388),
    .X(_09765_));
 sg13g2_nand2_1 _16855_ (.Y(_09766_),
    .A(\rbzero.pov.ready_buffer[37] ),
    .B(net353));
 sg13g2_nand3_1 _16856_ (.B(_09764_),
    .C(_09766_),
    .A(net752),
    .Y(_00481_));
 sg13g2_buf_1 _16857_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .X(_09767_));
 sg13g2_nand2_1 _16858_ (.Y(_09768_),
    .A(_09767_),
    .B(net354));
 sg13g2_nand2_1 _16859_ (.Y(_09769_),
    .A(\rbzero.pov.ready_buffer[38] ),
    .B(net353));
 sg13g2_nand3_1 _16860_ (.B(_09768_),
    .C(_09769_),
    .A(net752),
    .Y(_00482_));
 sg13g2_buf_1 _16861_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .X(_09770_));
 sg13g2_nand2_1 _16862_ (.Y(_09771_),
    .A(_09770_),
    .B(net354));
 sg13g2_nand2_1 _16863_ (.Y(_09772_),
    .A(\rbzero.pov.ready_buffer[39] ),
    .B(_09765_));
 sg13g2_nand3_1 _16864_ (.B(_09771_),
    .C(_09772_),
    .A(net752),
    .Y(_00483_));
 sg13g2_nand2_1 _16865_ (.Y(_09773_),
    .A(\rbzero.pov.ready_buffer[40] ),
    .B(_09745_));
 sg13g2_buf_2 _16866_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .X(_09774_));
 sg13g2_nand2_1 _16867_ (.Y(_09775_),
    .A(_09774_),
    .B(net355));
 sg13g2_a21oi_1 _16868_ (.A1(_09773_),
    .A2(_09775_),
    .Y(_00484_),
    .B1(net606));
 sg13g2_buf_1 _16869_ (.A(net758),
    .X(_09776_));
 sg13g2_buf_2 _16870_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .X(_09777_));
 sg13g2_nand2_1 _16871_ (.Y(_09778_),
    .A(_09777_),
    .B(net354));
 sg13g2_nand2_1 _16872_ (.Y(_09779_),
    .A(\rbzero.pov.ready_buffer[41] ),
    .B(_09765_));
 sg13g2_nand3_1 _16873_ (.B(_09778_),
    .C(_09779_),
    .A(net717),
    .Y(_00485_));
 sg13g2_nand2_1 _16874_ (.Y(_09780_),
    .A(\rbzero.pov.ready_buffer[42] ),
    .B(_09745_));
 sg13g2_buf_2 _16875_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .X(_09781_));
 sg13g2_nand2_1 _16876_ (.Y(_09782_),
    .A(_09781_),
    .B(net355));
 sg13g2_a21oi_1 _16877_ (.A1(_09780_),
    .A2(_09782_),
    .Y(_00486_),
    .B1(net606));
 sg13g2_buf_1 _16878_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .X(_09783_));
 sg13g2_nand2_1 _16879_ (.Y(_09784_),
    .A(_09783_),
    .B(net354));
 sg13g2_nand2_1 _16880_ (.Y(_09785_),
    .A(\rbzero.pov.ready_buffer[22] ),
    .B(net353));
 sg13g2_nand3_1 _16881_ (.B(_09784_),
    .C(_09785_),
    .A(net717),
    .Y(_00487_));
 sg13g2_buf_2 _16882_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .X(_09786_));
 sg13g2_nand2_1 _16883_ (.Y(_09787_),
    .A(_09786_),
    .B(net354));
 sg13g2_nand2_1 _16884_ (.Y(_09788_),
    .A(\rbzero.pov.ready_buffer[32] ),
    .B(net353));
 sg13g2_nand3_1 _16885_ (.B(_09787_),
    .C(_09788_),
    .A(net717),
    .Y(_00488_));
 sg13g2_nand2_1 _16886_ (.Y(_09789_),
    .A(\rbzero.pov.ready_buffer[23] ),
    .B(net356));
 sg13g2_buf_1 _16887_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .X(_09790_));
 sg13g2_nand2_1 _16888_ (.Y(_09791_),
    .A(_09790_),
    .B(net355));
 sg13g2_a21oi_1 _16889_ (.A1(_09789_),
    .A2(_09791_),
    .Y(_00489_),
    .B1(net606));
 sg13g2_buf_1 _16890_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .X(_09792_));
 sg13g2_nand2_1 _16891_ (.Y(_09793_),
    .A(_09792_),
    .B(_09763_));
 sg13g2_nand2_1 _16892_ (.Y(_09794_),
    .A(\rbzero.pov.ready_buffer[24] ),
    .B(net353));
 sg13g2_nand3_1 _16893_ (.B(_09793_),
    .C(_09794_),
    .A(net717),
    .Y(_00490_));
 sg13g2_buf_1 _16894_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .X(_09795_));
 sg13g2_nand2_1 _16895_ (.Y(_09796_),
    .A(_09795_),
    .B(net354));
 sg13g2_nand2_1 _16896_ (.Y(_09797_),
    .A(\rbzero.pov.ready_buffer[25] ),
    .B(net353));
 sg13g2_nand3_1 _16897_ (.B(_09796_),
    .C(_09797_),
    .A(net717),
    .Y(_00491_));
 sg13g2_buf_2 _16898_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .X(_09798_));
 sg13g2_nand2_1 _16899_ (.Y(_09799_),
    .A(_09798_),
    .B(net354));
 sg13g2_nand2_1 _16900_ (.Y(_09800_),
    .A(\rbzero.pov.ready_buffer[26] ),
    .B(net353));
 sg13g2_nand3_1 _16901_ (.B(_09799_),
    .C(_09800_),
    .A(_09776_),
    .Y(_00492_));
 sg13g2_nand2_1 _16902_ (.Y(_09801_),
    .A(\rbzero.pov.ready_buffer[27] ),
    .B(net356));
 sg13g2_buf_2 _16903_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .X(_09802_));
 sg13g2_nand2_1 _16904_ (.Y(_09803_),
    .A(_09802_),
    .B(net355));
 sg13g2_a21oi_1 _16905_ (.A1(_09801_),
    .A2(_09803_),
    .Y(_00493_),
    .B1(net606));
 sg13g2_nand2_1 _16906_ (.Y(_09804_),
    .A(\rbzero.pov.ready_buffer[28] ),
    .B(net356));
 sg13g2_buf_2 _16907_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .X(_09805_));
 sg13g2_nand2_1 _16908_ (.Y(_09806_),
    .A(_09805_),
    .B(net355));
 sg13g2_a21oi_1 _16909_ (.A1(_09804_),
    .A2(_09806_),
    .Y(_00494_),
    .B1(_09760_));
 sg13g2_buf_2 _16910_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .X(_09807_));
 sg13g2_nand2_1 _16911_ (.Y(_09808_),
    .A(_09807_),
    .B(_09763_));
 sg13g2_nand2_1 _16912_ (.Y(_09809_),
    .A(\rbzero.pov.ready_buffer[29] ),
    .B(net353));
 sg13g2_nand3_1 _16913_ (.B(_09808_),
    .C(_09809_),
    .A(_09776_),
    .Y(_00495_));
 sg13g2_nand2_1 _16914_ (.Y(_09810_),
    .A(\rbzero.pov.ready_buffer[30] ),
    .B(net356));
 sg13g2_buf_1 _16915_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .X(_09811_));
 sg13g2_nand2_1 _16916_ (.Y(_09812_),
    .A(_09811_),
    .B(_09748_));
 sg13g2_a21oi_1 _16917_ (.A1(_09810_),
    .A2(_09812_),
    .Y(_00496_),
    .B1(_09760_));
 sg13g2_buf_1 _16918_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .X(_09813_));
 sg13g2_nand2_1 _16919_ (.Y(_09814_),
    .A(_09813_),
    .B(_09743_));
 sg13g2_nand2_1 _16920_ (.Y(_09815_),
    .A(\rbzero.pov.ready_buffer[31] ),
    .B(_09737_));
 sg13g2_nand3_1 _16921_ (.B(_09814_),
    .C(_09815_),
    .A(net717),
    .Y(_00497_));
 sg13g2_buf_1 _16922_ (.A(_09424_),
    .X(_09816_));
 sg13g2_and2_1 _16923_ (.A(_09816_),
    .B(net2),
    .X(_00498_));
 sg13g2_and2_1 _16924_ (.A(_09816_),
    .B(\rbzero.pov.mosi_buffer[0] ),
    .X(_00499_));
 sg13g2_buf_1 _16925_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .X(_09817_));
 sg13g2_a21oi_1 _16926_ (.A1(net5),
    .A2(net451),
    .Y(_09818_),
    .B1(net388));
 sg13g2_buf_1 _16927_ (.A(_09818_),
    .X(_09819_));
 sg13g2_buf_1 _16928_ (.A(_00057_),
    .X(_09820_));
 sg13g2_buf_1 _16929_ (.A(_09419_),
    .X(_09821_));
 sg13g2_nand2_1 _16930_ (.Y(_09822_),
    .A(_09820_),
    .B(net352));
 sg13g2_nand2b_1 _16931_ (.Y(_09823_),
    .B(net451),
    .A_N(_09417_));
 sg13g2_buf_1 _16932_ (.A(_09823_),
    .X(_09824_));
 sg13g2_buf_1 _16933_ (.A(_09824_),
    .X(_09825_));
 sg13g2_nand2_1 _16934_ (.Y(_09826_),
    .A(\rbzero.pov.ready_buffer[59] ),
    .B(net351));
 sg13g2_a21oi_1 _16935_ (.A1(_09822_),
    .A2(_09826_),
    .Y(_09827_),
    .B1(_09819_));
 sg13g2_a21oi_1 _16936_ (.A1(_09817_),
    .A2(_09819_),
    .Y(_09828_),
    .B1(_09827_));
 sg13g2_nor2_1 _16937_ (.A(net607),
    .B(_09828_),
    .Y(_00500_));
 sg13g2_a21o_1 _16938_ (.A2(net451),
    .A1(net5),
    .B1(_09735_),
    .X(_09829_));
 sg13g2_buf_1 _16939_ (.A(_09829_),
    .X(_09830_));
 sg13g2_buf_1 _16940_ (.A(_09830_),
    .X(_09831_));
 sg13g2_buf_1 _16941_ (.A(_09419_),
    .X(_09832_));
 sg13g2_inv_1 _16942_ (.Y(_09833_),
    .A(_08494_));
 sg13g2_buf_1 _16943_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .X(_09834_));
 sg13g2_buf_1 _16944_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .X(_09835_));
 sg13g2_buf_2 _16945_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .X(_09836_));
 sg13g2_buf_1 _16946_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .X(_09837_));
 sg13g2_buf_1 _16947_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .X(_09838_));
 sg13g2_buf_2 _16948_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .X(_09839_));
 sg13g2_buf_2 _16949_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .X(_09840_));
 sg13g2_buf_1 _16950_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .X(_09841_));
 sg13g2_nor3_2 _16951_ (.A(_09840_),
    .B(_09841_),
    .C(_09817_),
    .Y(_09842_));
 sg13g2_nor2b_1 _16952_ (.A(_09839_),
    .B_N(_09842_),
    .Y(_09843_));
 sg13g2_buf_1 _16953_ (.A(_09843_),
    .X(_09844_));
 sg13g2_nand2b_1 _16954_ (.Y(_09845_),
    .B(_09844_),
    .A_N(_09838_));
 sg13g2_buf_1 _16955_ (.A(_09845_),
    .X(_09846_));
 sg13g2_nor3_2 _16956_ (.A(_09836_),
    .B(_09837_),
    .C(_09846_),
    .Y(_09847_));
 sg13g2_nand2b_1 _16957_ (.Y(_09848_),
    .B(_09847_),
    .A_N(_09835_));
 sg13g2_buf_1 _16958_ (.A(_09848_),
    .X(_09849_));
 sg13g2_nor2_1 _16959_ (.A(_09834_),
    .B(_09849_),
    .Y(_09850_));
 sg13g2_nand4_1 _16960_ (.B(_08511_),
    .C(net359),
    .A(_09833_),
    .Y(_09851_),
    .D(_09850_));
 sg13g2_o21ai_1 _16961_ (.B1(_09851_),
    .Y(_09852_),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .A2(net350));
 sg13g2_nor2b_1 _16962_ (.A(_09835_),
    .B_N(_09847_),
    .Y(_09853_));
 sg13g2_nand2b_1 _16963_ (.Y(_09854_),
    .B(_09853_),
    .A_N(_09834_));
 sg13g2_buf_1 _16964_ (.A(_09854_),
    .X(_09855_));
 sg13g2_o21ai_1 _16965_ (.B1(_09420_),
    .Y(_09856_),
    .A1(_08494_),
    .A2(_09855_));
 sg13g2_a21oi_1 _16966_ (.A1(_09830_),
    .A2(_09856_),
    .Y(_09857_),
    .B1(_08511_));
 sg13g2_a21oi_1 _16967_ (.A1(net339),
    .A2(_09852_),
    .Y(_09858_),
    .B1(_09857_));
 sg13g2_nand2b_1 _16968_ (.Y(_00501_),
    .B(net752),
    .A_N(_09858_));
 sg13g2_buf_1 _16969_ (.A(_09830_),
    .X(_09859_));
 sg13g2_buf_1 _16970_ (.A(_09824_),
    .X(_09860_));
 sg13g2_buf_1 _16971_ (.A(_09860_),
    .X(_09861_));
 sg13g2_nor3_1 _16972_ (.A(_08494_),
    .B(_08511_),
    .C(_09855_),
    .Y(_09862_));
 sg13g2_nand2b_1 _16973_ (.Y(_09863_),
    .B(_09862_),
    .A_N(_08501_));
 sg13g2_buf_1 _16974_ (.A(_09863_),
    .X(_09864_));
 sg13g2_nand2_1 _16975_ (.Y(_09865_),
    .A(\rbzero.pov.ready_buffer[70] ),
    .B(net351));
 sg13g2_o21ai_1 _16976_ (.B1(_09865_),
    .Y(_09866_),
    .A1(net337),
    .A2(_09864_));
 sg13g2_buf_1 _16977_ (.A(net349),
    .X(_09867_));
 sg13g2_o21ai_1 _16978_ (.B1(net339),
    .Y(_09868_),
    .A1(net336),
    .A2(_09862_));
 sg13g2_a22oi_1 _16979_ (.Y(_09869_),
    .B1(_09868_),
    .B2(_08501_),
    .A2(_09866_),
    .A1(net338));
 sg13g2_nor2_1 _16980_ (.A(net607),
    .B(_09869_),
    .Y(_00502_));
 sg13g2_a21oi_1 _16981_ (.A1(net340),
    .A2(_09864_),
    .Y(_09870_),
    .B1(_09819_));
 sg13g2_nor2_1 _16982_ (.A(\rbzero.pov.ready_buffer[71] ),
    .B(_09821_),
    .Y(_09871_));
 sg13g2_inv_1 _16983_ (.Y(_09872_),
    .A(_08483_));
 sg13g2_nor3_1 _16984_ (.A(_09872_),
    .B(net349),
    .C(_09864_),
    .Y(_09873_));
 sg13g2_o21ai_1 _16985_ (.B1(net339),
    .Y(_09874_),
    .A1(_09871_),
    .A2(_09873_));
 sg13g2_o21ai_1 _16986_ (.B1(_09874_),
    .Y(_09875_),
    .A1(_08483_),
    .A2(_09870_));
 sg13g2_nand2_1 _16987_ (.Y(_00503_),
    .A(net752),
    .B(_09875_));
 sg13g2_inv_1 _16988_ (.Y(_09876_),
    .A(\rbzero.pov.ready_buffer[72] ));
 sg13g2_nor3_1 _16989_ (.A(_08483_),
    .B(_08514_),
    .C(_09864_),
    .Y(_09877_));
 sg13g2_nand2_1 _16990_ (.Y(_09878_),
    .A(net359),
    .B(_09877_));
 sg13g2_o21ai_1 _16991_ (.B1(_09878_),
    .Y(_09879_),
    .A1(_09876_),
    .A2(net340));
 sg13g2_o21ai_1 _16992_ (.B1(net350),
    .Y(_09880_),
    .A1(_08483_),
    .A2(_09864_));
 sg13g2_nand2_1 _16993_ (.Y(_09881_),
    .A(net339),
    .B(_09880_));
 sg13g2_a22oi_1 _16994_ (.Y(_09882_),
    .B1(_09881_),
    .B2(_08514_),
    .A2(_09879_),
    .A1(net338));
 sg13g2_nor2_1 _16995_ (.A(net607),
    .B(_09882_),
    .Y(_00504_));
 sg13g2_nand2_1 _16996_ (.Y(_09883_),
    .A(\rbzero.pov.ready_buffer[73] ),
    .B(net351));
 sg13g2_o21ai_1 _16997_ (.B1(_09883_),
    .Y(_09884_),
    .A1(_08522_),
    .A2(_09878_));
 sg13g2_o21ai_1 _16998_ (.B1(net339),
    .Y(_09885_),
    .A1(net336),
    .A2(_09877_));
 sg13g2_a22oi_1 _16999_ (.Y(_09886_),
    .B1(_09885_),
    .B2(_08522_),
    .A2(_09884_),
    .A1(net338));
 sg13g2_nor2_1 _17000_ (.A(net607),
    .B(_09886_),
    .Y(_00505_));
 sg13g2_a21o_1 _17001_ (.A2(net350),
    .A1(_09817_),
    .B1(_09819_),
    .X(_09887_));
 sg13g2_nor2_1 _17002_ (.A(_09840_),
    .B(_09817_),
    .Y(_09888_));
 sg13g2_mux2_1 _17003_ (.A0(\rbzero.pov.ready_buffer[60] ),
    .A1(_09888_),
    .S(net350),
    .X(_09889_));
 sg13g2_a22oi_1 _17004_ (.Y(_09890_),
    .B1(_09889_),
    .B2(net338),
    .A2(_09887_),
    .A1(_09840_));
 sg13g2_nor2_1 _17005_ (.A(net607),
    .B(_09890_),
    .Y(_00506_));
 sg13g2_mux2_1 _17006_ (.A0(\rbzero.pov.ready_buffer[61] ),
    .A1(_09842_),
    .S(_09832_),
    .X(_09891_));
 sg13g2_o21ai_1 _17007_ (.B1(_09831_),
    .Y(_09892_),
    .A1(net336),
    .A2(_09888_));
 sg13g2_a22oi_1 _17008_ (.Y(_09893_),
    .B1(_09892_),
    .B2(_09841_),
    .A2(_09891_),
    .A1(net338));
 sg13g2_nor2_1 _17009_ (.A(net607),
    .B(_09893_),
    .Y(_00507_));
 sg13g2_mux2_1 _17010_ (.A0(\rbzero.pov.ready_buffer[62] ),
    .A1(_09844_),
    .S(_09832_),
    .X(_09894_));
 sg13g2_o21ai_1 _17011_ (.B1(_09831_),
    .Y(_09895_),
    .A1(net336),
    .A2(_09842_));
 sg13g2_a22oi_1 _17012_ (.Y(_09896_),
    .B1(_09895_),
    .B2(_09839_),
    .A2(_09894_),
    .A1(net338));
 sg13g2_nor2_1 _17013_ (.A(_09702_),
    .B(_09896_),
    .Y(_00508_));
 sg13g2_nand2_1 _17014_ (.Y(_09897_),
    .A(\rbzero.pov.ready_buffer[63] ),
    .B(_09825_));
 sg13g2_o21ai_1 _17015_ (.B1(_09897_),
    .Y(_09898_),
    .A1(net337),
    .A2(_09846_));
 sg13g2_o21ai_1 _17016_ (.B1(net339),
    .Y(_09899_),
    .A1(_09867_),
    .A2(_09844_));
 sg13g2_a22oi_1 _17017_ (.Y(_09900_),
    .B1(_09899_),
    .B2(_09838_),
    .A2(_09898_),
    .A1(net338));
 sg13g2_nor2_1 _17018_ (.A(_09702_),
    .B(_09900_),
    .Y(_00509_));
 sg13g2_buf_1 _17019_ (.A(_09759_),
    .X(_09901_));
 sg13g2_nor2_1 _17020_ (.A(_09836_),
    .B(_09846_),
    .Y(_09902_));
 sg13g2_mux2_1 _17021_ (.A0(\rbzero.pov.ready_buffer[64] ),
    .A1(_09902_),
    .S(net352),
    .X(_09903_));
 sg13g2_a21o_1 _17022_ (.A2(_09846_),
    .A1(net340),
    .B1(_09819_),
    .X(_09904_));
 sg13g2_a22oi_1 _17023_ (.Y(_09905_),
    .B1(_09904_),
    .B2(_09836_),
    .A2(_09903_),
    .A1(net338));
 sg13g2_nor2_1 _17024_ (.A(net605),
    .B(_09905_),
    .Y(_00510_));
 sg13g2_mux2_1 _17025_ (.A0(\rbzero.pov.ready_buffer[65] ),
    .A1(_09847_),
    .S(net352),
    .X(_09906_));
 sg13g2_o21ai_1 _17026_ (.B1(_09830_),
    .Y(_09907_),
    .A1(net336),
    .A2(_09902_));
 sg13g2_a22oi_1 _17027_ (.Y(_09908_),
    .B1(_09907_),
    .B2(_09837_),
    .A2(_09906_),
    .A1(_09859_));
 sg13g2_nor2_1 _17028_ (.A(net605),
    .B(_09908_),
    .Y(_00511_));
 sg13g2_nand2_1 _17029_ (.Y(_09909_),
    .A(\rbzero.pov.ready_buffer[66] ),
    .B(net351));
 sg13g2_o21ai_1 _17030_ (.B1(_09909_),
    .Y(_09910_),
    .A1(net337),
    .A2(_09849_));
 sg13g2_o21ai_1 _17031_ (.B1(_09830_),
    .Y(_09911_),
    .A1(net336),
    .A2(_09847_));
 sg13g2_a22oi_1 _17032_ (.Y(_09912_),
    .B1(_09911_),
    .B2(_09835_),
    .A2(_09910_),
    .A1(_09859_));
 sg13g2_nor2_1 _17033_ (.A(net605),
    .B(_09912_),
    .Y(_00512_));
 sg13g2_a21oi_1 _17034_ (.A1(net340),
    .A2(_09849_),
    .Y(_09913_),
    .B1(_09819_));
 sg13g2_nand3_1 _17035_ (.B(_09420_),
    .C(_09853_),
    .A(_09834_),
    .Y(_09914_));
 sg13g2_o21ai_1 _17036_ (.B1(_09914_),
    .Y(_09915_),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .A2(net352));
 sg13g2_nand2_1 _17037_ (.Y(_09916_),
    .A(net339),
    .B(_09915_));
 sg13g2_o21ai_1 _17038_ (.B1(_09916_),
    .Y(_09917_),
    .A1(_09834_),
    .A2(_09913_));
 sg13g2_nand2_1 _17039_ (.Y(_00513_),
    .A(net752),
    .B(_09917_));
 sg13g2_a21oi_1 _17040_ (.A1(_09421_),
    .A2(_09855_),
    .Y(_09918_),
    .B1(_09819_));
 sg13g2_nor2_1 _17041_ (.A(\rbzero.pov.ready_buffer[68] ),
    .B(net359),
    .Y(_09919_));
 sg13g2_nor3_1 _17042_ (.A(_09833_),
    .B(net349),
    .C(_09855_),
    .Y(_09920_));
 sg13g2_o21ai_1 _17043_ (.B1(net339),
    .Y(_09921_),
    .A1(_09919_),
    .A2(_09920_));
 sg13g2_o21ai_1 _17044_ (.B1(_09921_),
    .Y(_09922_),
    .A1(_08494_),
    .A2(_09918_));
 sg13g2_nand2_1 _17045_ (.Y(_00514_),
    .A(net752),
    .B(_09922_));
 sg13g2_buf_1 _17046_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .X(_09923_));
 sg13g2_a21oi_1 _17047_ (.A1(net6),
    .A2(_09740_),
    .Y(_09924_),
    .B1(_09736_));
 sg13g2_buf_1 _17048_ (.A(_09924_),
    .X(_09925_));
 sg13g2_buf_1 _17049_ (.A(_00059_),
    .X(_09926_));
 sg13g2_nand2_1 _17050_ (.Y(_09927_),
    .A(_09926_),
    .B(_09821_));
 sg13g2_nand2_1 _17051_ (.Y(_09928_),
    .A(\rbzero.pov.ready_buffer[44] ),
    .B(net351));
 sg13g2_a21oi_1 _17052_ (.A1(_09927_),
    .A2(_09928_),
    .Y(_09929_),
    .B1(_09925_));
 sg13g2_a21oi_1 _17053_ (.A1(_09923_),
    .A2(_09925_),
    .Y(_09930_),
    .B1(_09929_));
 sg13g2_nor2_1 _17054_ (.A(net605),
    .B(_09930_),
    .Y(_00515_));
 sg13g2_buf_1 _17055_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .X(_09931_));
 sg13g2_buf_1 _17056_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .X(_09932_));
 sg13g2_buf_2 _17057_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .X(_09933_));
 sg13g2_buf_1 _17058_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .X(_09934_));
 sg13g2_buf_1 _17059_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .X(_09935_));
 sg13g2_buf_1 _17060_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .X(_09936_));
 sg13g2_buf_2 _17061_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .X(_09937_));
 sg13g2_buf_1 _17062_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .X(_09938_));
 sg13g2_nor3_1 _17063_ (.A(_09937_),
    .B(_09938_),
    .C(_09923_),
    .Y(_09939_));
 sg13g2_nor2b_1 _17064_ (.A(_09936_),
    .B_N(_09939_),
    .Y(_09940_));
 sg13g2_buf_1 _17065_ (.A(_09940_),
    .X(_09941_));
 sg13g2_nand2b_1 _17066_ (.Y(_09942_),
    .B(_09941_),
    .A_N(_09935_));
 sg13g2_buf_1 _17067_ (.A(_09942_),
    .X(_09943_));
 sg13g2_nor3_1 _17068_ (.A(_09933_),
    .B(_09934_),
    .C(_09943_),
    .Y(_09944_));
 sg13g2_nand2b_1 _17069_ (.Y(_09945_),
    .B(_09944_),
    .A_N(_09932_));
 sg13g2_buf_1 _17070_ (.A(_09945_),
    .X(_09946_));
 sg13g2_nor2_1 _17071_ (.A(_09931_),
    .B(_09946_),
    .Y(_09947_));
 sg13g2_nand2b_1 _17072_ (.Y(_09948_),
    .B(_09947_),
    .A_N(_08485_));
 sg13g2_buf_1 _17073_ (.A(_09948_),
    .X(_09949_));
 sg13g2_a21oi_1 _17074_ (.A1(net340),
    .A2(_09949_),
    .Y(_09950_),
    .B1(_09925_));
 sg13g2_nor2_1 _17075_ (.A(\rbzero.pov.ready_buffer[54] ),
    .B(net359),
    .Y(_09951_));
 sg13g2_inv_1 _17076_ (.Y(_09952_),
    .A(_08507_));
 sg13g2_nor3_1 _17077_ (.A(_09952_),
    .B(net349),
    .C(_09949_),
    .Y(_09953_));
 sg13g2_a21o_1 _17078_ (.A2(_09740_),
    .A1(net6),
    .B1(_09735_),
    .X(_09954_));
 sg13g2_buf_1 _17079_ (.A(_09954_),
    .X(_09955_));
 sg13g2_buf_1 _17080_ (.A(_09955_),
    .X(_09956_));
 sg13g2_o21ai_1 _17081_ (.B1(net335),
    .Y(_09957_),
    .A1(_09951_),
    .A2(_09953_));
 sg13g2_o21ai_1 _17082_ (.B1(_09957_),
    .Y(_09958_),
    .A1(_08507_),
    .A2(_09950_));
 sg13g2_nand2_1 _17083_ (.Y(_00516_),
    .A(net752),
    .B(_09958_));
 sg13g2_buf_1 _17084_ (.A(_09955_),
    .X(_09959_));
 sg13g2_nor2_1 _17085_ (.A(_08507_),
    .B(_09949_),
    .Y(_09960_));
 sg13g2_nand2b_1 _17086_ (.Y(_09961_),
    .B(_09960_),
    .A_N(_08518_));
 sg13g2_buf_1 _17087_ (.A(_09961_),
    .X(_09962_));
 sg13g2_nand2_1 _17088_ (.Y(_09963_),
    .A(\rbzero.pov.ready_buffer[55] ),
    .B(net351));
 sg13g2_o21ai_1 _17089_ (.B1(_09963_),
    .Y(_09964_),
    .A1(net337),
    .A2(_09962_));
 sg13g2_o21ai_1 _17090_ (.B1(net335),
    .Y(_09965_),
    .A1(net336),
    .A2(_09960_));
 sg13g2_a22oi_1 _17091_ (.Y(_09966_),
    .B1(_09965_),
    .B2(_08518_),
    .A2(_09964_),
    .A1(net334));
 sg13g2_nor2_1 _17092_ (.A(net605),
    .B(_09966_),
    .Y(_00517_));
 sg13g2_a21oi_1 _17093_ (.A1(net340),
    .A2(_09962_),
    .Y(_09967_),
    .B1(_09925_));
 sg13g2_nor2_1 _17094_ (.A(\rbzero.pov.ready_buffer[56] ),
    .B(net359),
    .Y(_09968_));
 sg13g2_inv_1 _17095_ (.Y(_09969_),
    .A(_08489_));
 sg13g2_nor3_1 _17096_ (.A(_09969_),
    .B(net349),
    .C(_09962_),
    .Y(_09970_));
 sg13g2_o21ai_1 _17097_ (.B1(net335),
    .Y(_09971_),
    .A1(_09968_),
    .A2(_09970_));
 sg13g2_o21ai_1 _17098_ (.B1(_09971_),
    .Y(_09972_),
    .A1(_08489_),
    .A2(_09967_));
 sg13g2_nand2_1 _17099_ (.Y(_00518_),
    .A(_09761_),
    .B(_09972_));
 sg13g2_inv_1 _17100_ (.Y(_09973_),
    .A(\rbzero.pov.ready_buffer[57] ));
 sg13g2_nor3_1 _17101_ (.A(_08489_),
    .B(_08492_),
    .C(_09962_),
    .Y(_09974_));
 sg13g2_nand2_1 _17102_ (.Y(_09975_),
    .A(net359),
    .B(_09974_));
 sg13g2_o21ai_1 _17103_ (.B1(_09975_),
    .Y(_09976_),
    .A1(_09973_),
    .A2(net340));
 sg13g2_o21ai_1 _17104_ (.B1(net350),
    .Y(_09977_),
    .A1(_08489_),
    .A2(_09962_));
 sg13g2_nand2_1 _17105_ (.Y(_09978_),
    .A(net335),
    .B(_09977_));
 sg13g2_a22oi_1 _17106_ (.Y(_09979_),
    .B1(_09978_),
    .B2(_08492_),
    .A2(_09976_),
    .A1(net334));
 sg13g2_nor2_1 _17107_ (.A(net605),
    .B(_09979_),
    .Y(_00519_));
 sg13g2_nand2_1 _17108_ (.Y(_09980_),
    .A(\rbzero.pov.ready_buffer[58] ),
    .B(net351));
 sg13g2_o21ai_1 _17109_ (.B1(_09980_),
    .Y(_09981_),
    .A1(_08498_),
    .A2(_09975_));
 sg13g2_o21ai_1 _17110_ (.B1(net335),
    .Y(_09982_),
    .A1(net336),
    .A2(_09974_));
 sg13g2_a22oi_1 _17111_ (.Y(_09983_),
    .B1(_09982_),
    .B2(_08498_),
    .A2(_09981_),
    .A1(net334));
 sg13g2_nor2_1 _17112_ (.A(net605),
    .B(_09983_),
    .Y(_00520_));
 sg13g2_a21o_1 _17113_ (.A2(net350),
    .A1(_09923_),
    .B1(_09925_),
    .X(_09984_));
 sg13g2_nor2_1 _17114_ (.A(_09937_),
    .B(_09923_),
    .Y(_09985_));
 sg13g2_mux2_1 _17115_ (.A0(\rbzero.pov.ready_buffer[45] ),
    .A1(_09985_),
    .S(net350),
    .X(_09986_));
 sg13g2_a22oi_1 _17116_ (.Y(_09987_),
    .B1(_09986_),
    .B2(net334),
    .A2(_09984_),
    .A1(_09937_));
 sg13g2_nor2_1 _17117_ (.A(net605),
    .B(_09987_),
    .Y(_00521_));
 sg13g2_mux2_1 _17118_ (.A0(\rbzero.pov.ready_buffer[46] ),
    .A1(_09939_),
    .S(net352),
    .X(_09988_));
 sg13g2_o21ai_1 _17119_ (.B1(_09956_),
    .Y(_09989_),
    .A1(_09867_),
    .A2(_09985_));
 sg13g2_a22oi_1 _17120_ (.Y(_09990_),
    .B1(_09989_),
    .B2(_09938_),
    .A2(_09988_),
    .A1(net334));
 sg13g2_nor2_1 _17121_ (.A(_09901_),
    .B(_09990_),
    .Y(_00522_));
 sg13g2_mux2_1 _17122_ (.A0(\rbzero.pov.ready_buffer[47] ),
    .A1(_09941_),
    .S(net352),
    .X(_09991_));
 sg13g2_o21ai_1 _17123_ (.B1(net335),
    .Y(_09992_),
    .A1(net337),
    .A2(_09939_));
 sg13g2_a22oi_1 _17124_ (.Y(_09993_),
    .B1(_09992_),
    .B2(_09936_),
    .A2(_09991_),
    .A1(net334));
 sg13g2_nor2_1 _17125_ (.A(_09901_),
    .B(_09993_),
    .Y(_00523_));
 sg13g2_nand2_1 _17126_ (.Y(_09994_),
    .A(\rbzero.pov.ready_buffer[48] ),
    .B(net349));
 sg13g2_o21ai_1 _17127_ (.B1(_09994_),
    .Y(_09995_),
    .A1(net337),
    .A2(_09943_));
 sg13g2_o21ai_1 _17128_ (.B1(_09956_),
    .Y(_09996_),
    .A1(_09861_),
    .A2(_09941_));
 sg13g2_a22oi_1 _17129_ (.Y(_09997_),
    .B1(_09996_),
    .B2(_09935_),
    .A2(_09995_),
    .A1(net334));
 sg13g2_nor2_1 _17130_ (.A(net674),
    .B(_09997_),
    .Y(_00524_));
 sg13g2_nor2_1 _17131_ (.A(_09933_),
    .B(_09943_),
    .Y(_09998_));
 sg13g2_mux2_1 _17132_ (.A0(\rbzero.pov.ready_buffer[49] ),
    .A1(_09998_),
    .S(net352),
    .X(_09999_));
 sg13g2_a21o_1 _17133_ (.A2(_09943_),
    .A1(net350),
    .B1(_09925_),
    .X(_10000_));
 sg13g2_a22oi_1 _17134_ (.Y(_10001_),
    .B1(_10000_),
    .B2(_09933_),
    .A2(_09999_),
    .A1(net334));
 sg13g2_nor2_1 _17135_ (.A(net674),
    .B(_10001_),
    .Y(_00525_));
 sg13g2_mux2_1 _17136_ (.A0(\rbzero.pov.ready_buffer[50] ),
    .A1(_09944_),
    .S(net352),
    .X(_10002_));
 sg13g2_o21ai_1 _17137_ (.B1(_09955_),
    .Y(_10003_),
    .A1(_09861_),
    .A2(_09998_));
 sg13g2_a22oi_1 _17138_ (.Y(_10004_),
    .B1(_10003_),
    .B2(_09934_),
    .A2(_10002_),
    .A1(_09959_));
 sg13g2_nor2_1 _17139_ (.A(net674),
    .B(_10004_),
    .Y(_00526_));
 sg13g2_nand2_1 _17140_ (.Y(_10005_),
    .A(\rbzero.pov.ready_buffer[51] ),
    .B(net349));
 sg13g2_o21ai_1 _17141_ (.B1(_10005_),
    .Y(_10006_),
    .A1(net351),
    .A2(_09946_));
 sg13g2_o21ai_1 _17142_ (.B1(_09955_),
    .Y(_10007_),
    .A1(net337),
    .A2(_09944_));
 sg13g2_a22oi_1 _17143_ (.Y(_10008_),
    .B1(_10007_),
    .B2(_09932_),
    .A2(_10006_),
    .A1(_09959_));
 sg13g2_nor2_1 _17144_ (.A(_09724_),
    .B(_10008_),
    .Y(_00527_));
 sg13g2_a21oi_1 _17145_ (.A1(_09421_),
    .A2(_09946_),
    .Y(_10009_),
    .B1(_09925_));
 sg13g2_nor2_1 _17146_ (.A(\rbzero.pov.ready_buffer[52] ),
    .B(net359),
    .Y(_10010_));
 sg13g2_inv_1 _17147_ (.Y(_10011_),
    .A(_09931_));
 sg13g2_nor3_1 _17148_ (.A(_10011_),
    .B(net349),
    .C(_09946_),
    .Y(_10012_));
 sg13g2_o21ai_1 _17149_ (.B1(net335),
    .Y(_10013_),
    .A1(_10010_),
    .A2(_10012_));
 sg13g2_o21ai_1 _17150_ (.B1(_10013_),
    .Y(_10014_),
    .A1(_09931_),
    .A2(_10009_));
 sg13g2_nand2_1 _17151_ (.Y(_00528_),
    .A(_09761_),
    .B(_10014_));
 sg13g2_nand2_1 _17152_ (.Y(_10015_),
    .A(\rbzero.pov.ready_buffer[53] ),
    .B(_09860_));
 sg13g2_o21ai_1 _17153_ (.B1(_10015_),
    .Y(_10016_),
    .A1(_09825_),
    .A2(_09949_));
 sg13g2_o21ai_1 _17154_ (.B1(_09955_),
    .Y(_10017_),
    .A1(net337),
    .A2(_09947_));
 sg13g2_a22oi_1 _17155_ (.Y(_10018_),
    .B1(_10017_),
    .B2(_08485_),
    .A2(_10016_),
    .A1(net335));
 sg13g2_nor2_1 _17156_ (.A(_09724_),
    .B(_10018_),
    .Y(_00529_));
 sg13g2_nand2_1 _17157_ (.Y(_10019_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[0] ));
 sg13g2_nand2b_1 _17158_ (.Y(_10020_),
    .B(\rbzero.pov.ready_buffer[0] ),
    .A_N(net759));
 sg13g2_a21oi_1 _17159_ (.A1(_10019_),
    .A2(_10020_),
    .Y(_00531_),
    .B1(net606));
 sg13g2_nand2_1 _17160_ (.Y(_10021_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[10] ));
 sg13g2_nand2b_1 _17161_ (.Y(_10022_),
    .B(\rbzero.pov.ready_buffer[10] ),
    .A_N(net759));
 sg13g2_a21oi_1 _17162_ (.A1(_10021_),
    .A2(_10022_),
    .Y(_00532_),
    .B1(net606));
 sg13g2_nand2_1 _17163_ (.Y(_10023_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[11] ));
 sg13g2_nand2b_1 _17164_ (.Y(_10024_),
    .B(\rbzero.pov.ready_buffer[11] ),
    .A_N(net759));
 sg13g2_a21oi_1 _17165_ (.A1(_10023_),
    .A2(_10024_),
    .Y(_00533_),
    .B1(net606));
 sg13g2_nand2_1 _17166_ (.Y(_10025_),
    .A(_09457_),
    .B(\rbzero.pov.spi_buffer[12] ));
 sg13g2_nand2b_1 _17167_ (.Y(_10026_),
    .B(\rbzero.pov.ready_buffer[12] ),
    .A_N(net759));
 sg13g2_buf_1 _17168_ (.A(_09759_),
    .X(_10027_));
 sg13g2_a21oi_1 _17169_ (.A1(_10025_),
    .A2(_10026_),
    .Y(_00534_),
    .B1(net604));
 sg13g2_nand2_1 _17170_ (.Y(_10028_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[13] ));
 sg13g2_buf_1 _17171_ (.A(_09422_),
    .X(_10029_));
 sg13g2_buf_1 _17172_ (.A(_10029_),
    .X(_10030_));
 sg13g2_nand2b_1 _17173_ (.Y(_10031_),
    .B(\rbzero.pov.ready_buffer[13] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17174_ (.A1(_10028_),
    .A2(_10031_),
    .Y(_00535_),
    .B1(net604));
 sg13g2_nand2_1 _17175_ (.Y(_10032_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[14] ));
 sg13g2_nand2b_1 _17176_ (.Y(_10033_),
    .B(\rbzero.pov.ready_buffer[14] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17177_ (.A1(_10032_),
    .A2(_10033_),
    .Y(_00536_),
    .B1(net604));
 sg13g2_nand2_1 _17178_ (.Y(_10034_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[15] ));
 sg13g2_nand2b_1 _17179_ (.Y(_10035_),
    .B(\rbzero.pov.ready_buffer[15] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17180_ (.A1(_10034_),
    .A2(_10035_),
    .Y(_00537_),
    .B1(net604));
 sg13g2_nand2_1 _17181_ (.Y(_10036_),
    .A(net720),
    .B(\rbzero.pov.spi_buffer[16] ));
 sg13g2_nand2b_1 _17182_ (.Y(_10037_),
    .B(\rbzero.pov.ready_buffer[16] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17183_ (.A1(_10036_),
    .A2(_10037_),
    .Y(_00538_),
    .B1(net604));
 sg13g2_nand2_1 _17184_ (.Y(_10038_),
    .A(_09457_),
    .B(\rbzero.pov.spi_buffer[17] ));
 sg13g2_nand2b_1 _17185_ (.Y(_10039_),
    .B(\rbzero.pov.ready_buffer[17] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17186_ (.A1(_10038_),
    .A2(_10039_),
    .Y(_00539_),
    .B1(_10027_));
 sg13g2_buf_1 _17187_ (.A(_09456_),
    .X(_10040_));
 sg13g2_nand2_1 _17188_ (.Y(_10041_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[18] ));
 sg13g2_nand2b_1 _17189_ (.Y(_10042_),
    .B(\rbzero.pov.ready_buffer[18] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17190_ (.A1(_10041_),
    .A2(_10042_),
    .Y(_00540_),
    .B1(net604));
 sg13g2_nand2_1 _17191_ (.Y(_10043_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[19] ));
 sg13g2_nand2b_1 _17192_ (.Y(_10044_),
    .B(\rbzero.pov.ready_buffer[19] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17193_ (.A1(_10043_),
    .A2(_10044_),
    .Y(_00541_),
    .B1(net604));
 sg13g2_nand2_1 _17194_ (.Y(_10045_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[1] ));
 sg13g2_nand2b_1 _17195_ (.Y(_10046_),
    .B(\rbzero.pov.ready_buffer[1] ),
    .A_N(_10030_));
 sg13g2_a21oi_1 _17196_ (.A1(_10045_),
    .A2(_10046_),
    .Y(_00542_),
    .B1(_10027_));
 sg13g2_nand2_1 _17197_ (.Y(_10047_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[20] ));
 sg13g2_nand2b_1 _17198_ (.Y(_10048_),
    .B(\rbzero.pov.ready_buffer[20] ),
    .A_N(net716));
 sg13g2_a21oi_1 _17199_ (.A1(_10047_),
    .A2(_10048_),
    .Y(_00543_),
    .B1(net604));
 sg13g2_nand2_1 _17200_ (.Y(_10049_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[21] ));
 sg13g2_nand2b_1 _17201_ (.Y(_10050_),
    .B(\rbzero.pov.ready_buffer[21] ),
    .A_N(_10030_));
 sg13g2_buf_1 _17202_ (.A(_09759_),
    .X(_10051_));
 sg13g2_a21oi_1 _17203_ (.A1(_10049_),
    .A2(_10050_),
    .Y(_00544_),
    .B1(net603));
 sg13g2_nand2_1 _17204_ (.Y(_10052_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[22] ));
 sg13g2_buf_1 _17205_ (.A(_10029_),
    .X(_10053_));
 sg13g2_nand2b_1 _17206_ (.Y(_10054_),
    .B(\rbzero.pov.ready_buffer[22] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17207_ (.A1(_10052_),
    .A2(_10054_),
    .Y(_00545_),
    .B1(net603));
 sg13g2_nand2_1 _17208_ (.Y(_10055_),
    .A(_10040_),
    .B(\rbzero.pov.spi_buffer[23] ));
 sg13g2_nand2b_1 _17209_ (.Y(_10056_),
    .B(\rbzero.pov.ready_buffer[23] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17210_ (.A1(_10055_),
    .A2(_10056_),
    .Y(_00546_),
    .B1(net603));
 sg13g2_nand2_1 _17211_ (.Y(_10057_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[24] ));
 sg13g2_nand2b_1 _17212_ (.Y(_10058_),
    .B(\rbzero.pov.ready_buffer[24] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17213_ (.A1(_10057_),
    .A2(_10058_),
    .Y(_00547_),
    .B1(net603));
 sg13g2_nand2_1 _17214_ (.Y(_10059_),
    .A(net715),
    .B(\rbzero.pov.spi_buffer[25] ));
 sg13g2_nand2b_1 _17215_ (.Y(_10060_),
    .B(\rbzero.pov.ready_buffer[25] ),
    .A_N(_10053_));
 sg13g2_a21oi_1 _17216_ (.A1(_10059_),
    .A2(_10060_),
    .Y(_00548_),
    .B1(_10051_));
 sg13g2_nand2_1 _17217_ (.Y(_10061_),
    .A(_10040_),
    .B(\rbzero.pov.spi_buffer[26] ));
 sg13g2_nand2b_1 _17218_ (.Y(_10062_),
    .B(\rbzero.pov.ready_buffer[26] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17219_ (.A1(_10061_),
    .A2(_10062_),
    .Y(_00549_),
    .B1(net603));
 sg13g2_buf_1 _17220_ (.A(_09456_),
    .X(_10063_));
 sg13g2_nand2_1 _17221_ (.Y(_10064_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[27] ));
 sg13g2_nand2b_1 _17222_ (.Y(_10065_),
    .B(\rbzero.pov.ready_buffer[27] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17223_ (.A1(_10064_),
    .A2(_10065_),
    .Y(_00550_),
    .B1(net603));
 sg13g2_nand2_1 _17224_ (.Y(_10066_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[28] ));
 sg13g2_nand2b_1 _17225_ (.Y(_10067_),
    .B(\rbzero.pov.ready_buffer[28] ),
    .A_N(_10053_));
 sg13g2_a21oi_1 _17226_ (.A1(_10066_),
    .A2(_10067_),
    .Y(_00551_),
    .B1(net603));
 sg13g2_nand2_1 _17227_ (.Y(_10068_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[29] ));
 sg13g2_nand2b_1 _17228_ (.Y(_10069_),
    .B(\rbzero.pov.ready_buffer[29] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17229_ (.A1(_10068_),
    .A2(_10069_),
    .Y(_00552_),
    .B1(_10051_));
 sg13g2_nand2_1 _17230_ (.Y(_10070_),
    .A(_10063_),
    .B(\rbzero.pov.spi_buffer[2] ));
 sg13g2_nand2b_1 _17231_ (.Y(_10071_),
    .B(\rbzero.pov.ready_buffer[2] ),
    .A_N(net714));
 sg13g2_a21oi_1 _17232_ (.A1(_10070_),
    .A2(_10071_),
    .Y(_00553_),
    .B1(net603));
 sg13g2_nand2_1 _17233_ (.Y(_10072_),
    .A(_10063_),
    .B(\rbzero.pov.spi_buffer[30] ));
 sg13g2_nand2b_1 _17234_ (.Y(_10073_),
    .B(\rbzero.pov.ready_buffer[30] ),
    .A_N(net714));
 sg13g2_buf_1 _17235_ (.A(_09759_),
    .X(_10074_));
 sg13g2_a21oi_1 _17236_ (.A1(_10072_),
    .A2(_10073_),
    .Y(_00554_),
    .B1(net602));
 sg13g2_nand2_1 _17237_ (.Y(_10075_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[31] ));
 sg13g2_buf_1 _17238_ (.A(_10029_),
    .X(_10076_));
 sg13g2_nand2b_1 _17239_ (.Y(_10077_),
    .B(\rbzero.pov.ready_buffer[31] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17240_ (.A1(_10075_),
    .A2(_10077_),
    .Y(_00555_),
    .B1(net602));
 sg13g2_nand2_1 _17241_ (.Y(_10078_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[32] ));
 sg13g2_nand2b_1 _17242_ (.Y(_10079_),
    .B(\rbzero.pov.ready_buffer[32] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17243_ (.A1(_10078_),
    .A2(_10079_),
    .Y(_00556_),
    .B1(net602));
 sg13g2_nand2_1 _17244_ (.Y(_10080_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[33] ));
 sg13g2_nand2b_1 _17245_ (.Y(_10081_),
    .B(\rbzero.pov.ready_buffer[33] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17246_ (.A1(_10080_),
    .A2(_10081_),
    .Y(_00557_),
    .B1(net602));
 sg13g2_nand2_1 _17247_ (.Y(_10082_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[34] ));
 sg13g2_nand2b_1 _17248_ (.Y(_10083_),
    .B(\rbzero.pov.ready_buffer[34] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17249_ (.A1(_10082_),
    .A2(_10083_),
    .Y(_00558_),
    .B1(net602));
 sg13g2_nand2_1 _17250_ (.Y(_10084_),
    .A(net713),
    .B(\rbzero.pov.spi_buffer[35] ));
 sg13g2_nand2b_1 _17251_ (.Y(_10085_),
    .B(\rbzero.pov.ready_buffer[35] ),
    .A_N(_10076_));
 sg13g2_a21oi_1 _17252_ (.A1(_10084_),
    .A2(_10085_),
    .Y(_00559_),
    .B1(net602));
 sg13g2_buf_1 _17253_ (.A(_09456_),
    .X(_10086_));
 sg13g2_nand2_1 _17254_ (.Y(_10087_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[36] ));
 sg13g2_nand2b_1 _17255_ (.Y(_10088_),
    .B(\rbzero.pov.ready_buffer[36] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17256_ (.A1(_10087_),
    .A2(_10088_),
    .Y(_00560_),
    .B1(_10074_));
 sg13g2_nand2_1 _17257_ (.Y(_10089_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[37] ));
 sg13g2_nand2b_1 _17258_ (.Y(_10090_),
    .B(\rbzero.pov.ready_buffer[37] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17259_ (.A1(_10089_),
    .A2(_10090_),
    .Y(_00561_),
    .B1(_10074_));
 sg13g2_nand2_1 _17260_ (.Y(_10091_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[38] ));
 sg13g2_nand2b_1 _17261_ (.Y(_10092_),
    .B(\rbzero.pov.ready_buffer[38] ),
    .A_N(net712));
 sg13g2_a21oi_1 _17262_ (.A1(_10091_),
    .A2(_10092_),
    .Y(_00562_),
    .B1(net602));
 sg13g2_nand2_1 _17263_ (.Y(_10093_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[39] ));
 sg13g2_nand2b_1 _17264_ (.Y(_10094_),
    .B(\rbzero.pov.ready_buffer[39] ),
    .A_N(_10076_));
 sg13g2_a21oi_1 _17265_ (.A1(_10093_),
    .A2(_10094_),
    .Y(_00563_),
    .B1(net602));
 sg13g2_nand2_1 _17266_ (.Y(_10095_),
    .A(_10086_),
    .B(\rbzero.pov.spi_buffer[3] ));
 sg13g2_nand2b_1 _17267_ (.Y(_10096_),
    .B(\rbzero.pov.ready_buffer[3] ),
    .A_N(net712));
 sg13g2_buf_1 _17268_ (.A(_09759_),
    .X(_10097_));
 sg13g2_a21oi_1 _17269_ (.A1(_10095_),
    .A2(_10096_),
    .Y(_00564_),
    .B1(net601));
 sg13g2_nand2_1 _17270_ (.Y(_10098_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[40] ));
 sg13g2_buf_1 _17271_ (.A(_10029_),
    .X(_10099_));
 sg13g2_nand2b_1 _17272_ (.Y(_10100_),
    .B(\rbzero.pov.ready_buffer[40] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17273_ (.A1(_10098_),
    .A2(_10100_),
    .Y(_00565_),
    .B1(net601));
 sg13g2_nand2_1 _17274_ (.Y(_10101_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[41] ));
 sg13g2_nand2b_1 _17275_ (.Y(_10102_),
    .B(\rbzero.pov.ready_buffer[41] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17276_ (.A1(_10101_),
    .A2(_10102_),
    .Y(_00566_),
    .B1(net601));
 sg13g2_nand2_1 _17277_ (.Y(_10103_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[42] ));
 sg13g2_nand2b_1 _17278_ (.Y(_10104_),
    .B(\rbzero.pov.ready_buffer[42] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17279_ (.A1(_10103_),
    .A2(_10104_),
    .Y(_00567_),
    .B1(net601));
 sg13g2_nand2_1 _17280_ (.Y(_10105_),
    .A(_10086_),
    .B(\rbzero.pov.spi_buffer[43] ));
 sg13g2_nand2b_1 _17281_ (.Y(_10106_),
    .B(\rbzero.pov.ready_buffer[43] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17282_ (.A1(_10105_),
    .A2(_10106_),
    .Y(_00568_),
    .B1(net601));
 sg13g2_nand2_1 _17283_ (.Y(_10107_),
    .A(net711),
    .B(\rbzero.pov.spi_buffer[44] ));
 sg13g2_nand2b_1 _17284_ (.Y(_10108_),
    .B(\rbzero.pov.ready_buffer[44] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17285_ (.A1(_10107_),
    .A2(_10108_),
    .Y(_00569_),
    .B1(net601));
 sg13g2_buf_1 _17286_ (.A(_09456_),
    .X(_10109_));
 sg13g2_nand2_1 _17287_ (.Y(_10110_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[45] ));
 sg13g2_nand2b_1 _17288_ (.Y(_10111_),
    .B(\rbzero.pov.ready_buffer[45] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17289_ (.A1(_10110_),
    .A2(_10111_),
    .Y(_00570_),
    .B1(net601));
 sg13g2_nand2_1 _17290_ (.Y(_10112_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[46] ));
 sg13g2_nand2b_1 _17291_ (.Y(_10113_),
    .B(\rbzero.pov.ready_buffer[46] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17292_ (.A1(_10112_),
    .A2(_10113_),
    .Y(_00571_),
    .B1(net601));
 sg13g2_nand2_1 _17293_ (.Y(_10114_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[47] ));
 sg13g2_nand2b_1 _17294_ (.Y(_10115_),
    .B(\rbzero.pov.ready_buffer[47] ),
    .A_N(net710));
 sg13g2_a21oi_1 _17295_ (.A1(_10114_),
    .A2(_10115_),
    .Y(_00572_),
    .B1(_10097_));
 sg13g2_nand2_1 _17296_ (.Y(_10116_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[48] ));
 sg13g2_nand2b_1 _17297_ (.Y(_10117_),
    .B(\rbzero.pov.ready_buffer[48] ),
    .A_N(_10099_));
 sg13g2_a21oi_1 _17298_ (.A1(_10116_),
    .A2(_10117_),
    .Y(_00573_),
    .B1(_10097_));
 sg13g2_nand2_1 _17299_ (.Y(_10118_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[49] ));
 sg13g2_nand2b_1 _17300_ (.Y(_10119_),
    .B(\rbzero.pov.ready_buffer[49] ),
    .A_N(_10099_));
 sg13g2_buf_1 _17301_ (.A(_09759_),
    .X(_10120_));
 sg13g2_a21oi_1 _17302_ (.A1(_10118_),
    .A2(_10119_),
    .Y(_00574_),
    .B1(_10120_));
 sg13g2_nand2_1 _17303_ (.Y(_10121_),
    .A(_10109_),
    .B(\rbzero.pov.spi_buffer[4] ));
 sg13g2_buf_1 _17304_ (.A(_10029_),
    .X(_10122_));
 sg13g2_nand2b_1 _17305_ (.Y(_10123_),
    .B(\rbzero.pov.ready_buffer[4] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17306_ (.A1(_10121_),
    .A2(_10123_),
    .Y(_00575_),
    .B1(net600));
 sg13g2_nand2_1 _17307_ (.Y(_10124_),
    .A(_10109_),
    .B(\rbzero.pov.spi_buffer[50] ));
 sg13g2_nand2b_1 _17308_ (.Y(_10125_),
    .B(\rbzero.pov.ready_buffer[50] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17309_ (.A1(_10124_),
    .A2(_10125_),
    .Y(_00576_),
    .B1(net600));
 sg13g2_nand2_1 _17310_ (.Y(_10126_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[51] ));
 sg13g2_nand2b_1 _17311_ (.Y(_10127_),
    .B(\rbzero.pov.ready_buffer[51] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17312_ (.A1(_10126_),
    .A2(_10127_),
    .Y(_00577_),
    .B1(net600));
 sg13g2_nand2_1 _17313_ (.Y(_10128_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[52] ));
 sg13g2_nand2b_1 _17314_ (.Y(_10129_),
    .B(\rbzero.pov.ready_buffer[52] ),
    .A_N(_10122_));
 sg13g2_a21oi_1 _17315_ (.A1(_10128_),
    .A2(_10129_),
    .Y(_00578_),
    .B1(net600));
 sg13g2_nand2_1 _17316_ (.Y(_10130_),
    .A(net709),
    .B(\rbzero.pov.spi_buffer[53] ));
 sg13g2_nand2b_1 _17317_ (.Y(_10131_),
    .B(\rbzero.pov.ready_buffer[53] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17318_ (.A1(_10130_),
    .A2(_10131_),
    .Y(_00579_),
    .B1(_10120_));
 sg13g2_buf_1 _17319_ (.A(_09456_),
    .X(_10132_));
 sg13g2_nand2_1 _17320_ (.Y(_10133_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[54] ));
 sg13g2_nand2b_1 _17321_ (.Y(_10134_),
    .B(\rbzero.pov.ready_buffer[54] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17322_ (.A1(_10133_),
    .A2(_10134_),
    .Y(_00580_),
    .B1(net600));
 sg13g2_nand2_1 _17323_ (.Y(_10135_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[55] ));
 sg13g2_nand2b_1 _17324_ (.Y(_10136_),
    .B(\rbzero.pov.ready_buffer[55] ),
    .A_N(_10122_));
 sg13g2_a21oi_1 _17325_ (.A1(_10135_),
    .A2(_10136_),
    .Y(_00581_),
    .B1(net600));
 sg13g2_nand2_1 _17326_ (.Y(_10137_),
    .A(_10132_),
    .B(\rbzero.pov.spi_buffer[56] ));
 sg13g2_nand2b_1 _17327_ (.Y(_10138_),
    .B(\rbzero.pov.ready_buffer[56] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17328_ (.A1(_10137_),
    .A2(_10138_),
    .Y(_00582_),
    .B1(net600));
 sg13g2_nand2_1 _17329_ (.Y(_10139_),
    .A(_10132_),
    .B(\rbzero.pov.spi_buffer[57] ));
 sg13g2_nand2b_1 _17330_ (.Y(_10140_),
    .B(\rbzero.pov.ready_buffer[57] ),
    .A_N(net708));
 sg13g2_a21oi_1 _17331_ (.A1(_10139_),
    .A2(_10140_),
    .Y(_00583_),
    .B1(net600));
 sg13g2_nand2_1 _17332_ (.Y(_10141_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[58] ));
 sg13g2_nand2b_1 _17333_ (.Y(_10142_),
    .B(\rbzero.pov.ready_buffer[58] ),
    .A_N(net708));
 sg13g2_buf_1 _17334_ (.A(_09700_),
    .X(_10143_));
 sg13g2_buf_1 _17335_ (.A(_10143_),
    .X(_10144_));
 sg13g2_a21oi_1 _17336_ (.A1(_10141_),
    .A2(_10142_),
    .Y(_00584_),
    .B1(net599));
 sg13g2_nand2_1 _17337_ (.Y(_10145_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[59] ));
 sg13g2_buf_1 _17338_ (.A(_10029_),
    .X(_10146_));
 sg13g2_nand2b_1 _17339_ (.Y(_10147_),
    .B(\rbzero.pov.ready_buffer[59] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17340_ (.A1(_10145_),
    .A2(_10147_),
    .Y(_00585_),
    .B1(_10144_));
 sg13g2_nand2_1 _17341_ (.Y(_10148_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[5] ));
 sg13g2_nand2b_1 _17342_ (.Y(_10149_),
    .B(\rbzero.pov.ready_buffer[5] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17343_ (.A1(_10148_),
    .A2(_10149_),
    .Y(_00586_),
    .B1(net599));
 sg13g2_nand2_1 _17344_ (.Y(_10150_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[60] ));
 sg13g2_nand2b_1 _17345_ (.Y(_10151_),
    .B(\rbzero.pov.ready_buffer[60] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17346_ (.A1(_10150_),
    .A2(_10151_),
    .Y(_00587_),
    .B1(net599));
 sg13g2_nand2_1 _17347_ (.Y(_10152_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[61] ));
 sg13g2_nand2b_1 _17348_ (.Y(_10153_),
    .B(\rbzero.pov.ready_buffer[61] ),
    .A_N(_10146_));
 sg13g2_a21oi_1 _17349_ (.A1(_10152_),
    .A2(_10153_),
    .Y(_00588_),
    .B1(_10144_));
 sg13g2_nand2_1 _17350_ (.Y(_10154_),
    .A(net707),
    .B(\rbzero.pov.spi_buffer[62] ));
 sg13g2_nand2b_1 _17351_ (.Y(_10155_),
    .B(\rbzero.pov.ready_buffer[62] ),
    .A_N(_10146_));
 sg13g2_a21oi_1 _17352_ (.A1(_10154_),
    .A2(_10155_),
    .Y(_00589_),
    .B1(net599));
 sg13g2_buf_1 _17353_ (.A(_09456_),
    .X(_10156_));
 sg13g2_nand2_1 _17354_ (.Y(_10157_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[63] ));
 sg13g2_nand2b_1 _17355_ (.Y(_10158_),
    .B(\rbzero.pov.ready_buffer[63] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17356_ (.A1(_10157_),
    .A2(_10158_),
    .Y(_00590_),
    .B1(net599));
 sg13g2_nand2_1 _17357_ (.Y(_10159_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[64] ));
 sg13g2_nand2b_1 _17358_ (.Y(_10160_),
    .B(\rbzero.pov.ready_buffer[64] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17359_ (.A1(_10159_),
    .A2(_10160_),
    .Y(_00591_),
    .B1(net599));
 sg13g2_nand2_1 _17360_ (.Y(_10161_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[65] ));
 sg13g2_nand2b_1 _17361_ (.Y(_10162_),
    .B(\rbzero.pov.ready_buffer[65] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17362_ (.A1(_10161_),
    .A2(_10162_),
    .Y(_00592_),
    .B1(net599));
 sg13g2_nand2_1 _17363_ (.Y(_10163_),
    .A(_10156_),
    .B(\rbzero.pov.spi_buffer[66] ));
 sg13g2_nand2b_1 _17364_ (.Y(_10164_),
    .B(\rbzero.pov.ready_buffer[66] ),
    .A_N(net706));
 sg13g2_a21oi_1 _17365_ (.A1(_10163_),
    .A2(_10164_),
    .Y(_00593_),
    .B1(net599));
 sg13g2_nand2_1 _17366_ (.Y(_10165_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[67] ));
 sg13g2_nand2b_1 _17367_ (.Y(_10166_),
    .B(\rbzero.pov.ready_buffer[67] ),
    .A_N(net706));
 sg13g2_buf_1 _17368_ (.A(_10143_),
    .X(_10167_));
 sg13g2_a21oi_1 _17369_ (.A1(_10165_),
    .A2(_10166_),
    .Y(_00594_),
    .B1(net598));
 sg13g2_nand2_1 _17370_ (.Y(_10168_),
    .A(_10156_),
    .B(\rbzero.pov.spi_buffer[68] ));
 sg13g2_buf_1 _17371_ (.A(_10029_),
    .X(_10169_));
 sg13g2_nand2b_1 _17372_ (.Y(_10170_),
    .B(\rbzero.pov.ready_buffer[68] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17373_ (.A1(_10168_),
    .A2(_10170_),
    .Y(_00595_),
    .B1(net598));
 sg13g2_nand2_1 _17374_ (.Y(_10171_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[69] ));
 sg13g2_nand2b_1 _17375_ (.Y(_10172_),
    .B(\rbzero.pov.ready_buffer[69] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17376_ (.A1(_10171_),
    .A2(_10172_),
    .Y(_00596_),
    .B1(net598));
 sg13g2_nand2_1 _17377_ (.Y(_10173_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[6] ));
 sg13g2_nand2b_1 _17378_ (.Y(_10174_),
    .B(\rbzero.pov.ready_buffer[6] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17379_ (.A1(_10173_),
    .A2(_10174_),
    .Y(_00597_),
    .B1(net598));
 sg13g2_nand2_1 _17380_ (.Y(_10175_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[70] ));
 sg13g2_nand2b_1 _17381_ (.Y(_10176_),
    .B(\rbzero.pov.ready_buffer[70] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17382_ (.A1(_10175_),
    .A2(_10176_),
    .Y(_00598_),
    .B1(net598));
 sg13g2_nand2_1 _17383_ (.Y(_10177_),
    .A(net705),
    .B(\rbzero.pov.spi_buffer[71] ));
 sg13g2_nand2b_1 _17384_ (.Y(_10178_),
    .B(\rbzero.pov.ready_buffer[71] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17385_ (.A1(_10177_),
    .A2(_10178_),
    .Y(_00599_),
    .B1(net598));
 sg13g2_nand2_1 _17386_ (.Y(_10179_),
    .A(_09423_),
    .B(\rbzero.pov.spi_buffer[72] ));
 sg13g2_nand2b_1 _17387_ (.Y(_10180_),
    .B(\rbzero.pov.ready_buffer[72] ),
    .A_N(_10169_));
 sg13g2_a21oi_1 _17388_ (.A1(_10179_),
    .A2(_10180_),
    .Y(_00600_),
    .B1(_10167_));
 sg13g2_nand2_1 _17389_ (.Y(_10181_),
    .A(_09423_),
    .B(\rbzero.pov.spi_buffer[73] ));
 sg13g2_nand2b_1 _17390_ (.Y(_10182_),
    .B(\rbzero.pov.ready_buffer[73] ),
    .A_N(_10169_));
 sg13g2_a21oi_1 _17391_ (.A1(_10181_),
    .A2(_10182_),
    .Y(_00601_),
    .B1(_10167_));
 sg13g2_nand2_1 _17392_ (.Y(_10183_),
    .A(net759),
    .B(\rbzero.pov.spi_buffer[7] ));
 sg13g2_nand2b_1 _17393_ (.Y(_10184_),
    .B(\rbzero.pov.ready_buffer[7] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17394_ (.A1(_10183_),
    .A2(_10184_),
    .Y(_00602_),
    .B1(net598));
 sg13g2_nand2_1 _17395_ (.Y(_10185_),
    .A(net759),
    .B(\rbzero.pov.spi_buffer[8] ));
 sg13g2_nand2b_1 _17396_ (.Y(_10186_),
    .B(\rbzero.pov.ready_buffer[8] ),
    .A_N(net704));
 sg13g2_a21oi_1 _17397_ (.A1(_10185_),
    .A2(_10186_),
    .Y(_00603_),
    .B1(net598));
 sg13g2_nand2_1 _17398_ (.Y(_10187_),
    .A(net759),
    .B(\rbzero.pov.spi_buffer[9] ));
 sg13g2_nand2b_1 _17399_ (.Y(_10188_),
    .B(\rbzero.pov.ready_buffer[9] ),
    .A_N(net704));
 sg13g2_buf_1 _17400_ (.A(_10143_),
    .X(_10189_));
 sg13g2_a21oi_1 _17401_ (.A1(_10187_),
    .A2(_10188_),
    .Y(_00604_),
    .B1(_10189_));
 sg13g2_buf_1 _17402_ (.A(_09424_),
    .X(_10190_));
 sg13g2_and2_1 _17403_ (.A(net750),
    .B(net1),
    .X(_00605_));
 sg13g2_and2_1 _17404_ (.A(_10190_),
    .B(\rbzero.pov.sclk_buffer[0] ),
    .X(_00606_));
 sg13g2_and2_1 _17405_ (.A(net750),
    .B(\rbzero.pov.sclk_buffer[1] ),
    .X(_00607_));
 sg13g2_nor2b_1 _17406_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B_N(_09429_),
    .Y(_10191_));
 sg13g2_buf_1 _17407_ (.A(_10191_),
    .X(_10192_));
 sg13g2_buf_1 _17408_ (.A(_10192_),
    .X(_10193_));
 sg13g2_buf_1 _17409_ (.A(net596),
    .X(_10194_));
 sg13g2_nand2_1 _17410_ (.Y(_10195_),
    .A(\rbzero.pov.mosi ),
    .B(net542));
 sg13g2_buf_1 _17411_ (.A(_10192_),
    .X(_10196_));
 sg13g2_nand2b_1 _17412_ (.Y(_10197_),
    .B(\rbzero.pov.spi_buffer[0] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17413_ (.A1(_10195_),
    .A2(_10197_),
    .Y(_00608_),
    .B1(net597));
 sg13g2_nand2_1 _17414_ (.Y(_10198_),
    .A(\rbzero.pov.spi_buffer[9] ),
    .B(net542));
 sg13g2_nand2b_1 _17415_ (.Y(_10199_),
    .B(\rbzero.pov.spi_buffer[10] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17416_ (.A1(_10198_),
    .A2(_10199_),
    .Y(_00609_),
    .B1(net597));
 sg13g2_nand2_1 _17417_ (.Y(_10200_),
    .A(\rbzero.pov.spi_buffer[10] ),
    .B(net542));
 sg13g2_nand2b_1 _17418_ (.Y(_10201_),
    .B(\rbzero.pov.spi_buffer[11] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17419_ (.A1(_10200_),
    .A2(_10201_),
    .Y(_00610_),
    .B1(net597));
 sg13g2_nand2_1 _17420_ (.Y(_10202_),
    .A(\rbzero.pov.spi_buffer[11] ),
    .B(net542));
 sg13g2_nand2b_1 _17421_ (.Y(_10203_),
    .B(\rbzero.pov.spi_buffer[12] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17422_ (.A1(_10202_),
    .A2(_10203_),
    .Y(_00611_),
    .B1(net597));
 sg13g2_nand2_1 _17423_ (.Y(_10204_),
    .A(\rbzero.pov.spi_buffer[12] ),
    .B(net542));
 sg13g2_nand2b_1 _17424_ (.Y(_10205_),
    .B(\rbzero.pov.spi_buffer[13] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17425_ (.A1(_10204_),
    .A2(_10205_),
    .Y(_00612_),
    .B1(net597));
 sg13g2_nand2_1 _17426_ (.Y(_10206_),
    .A(\rbzero.pov.spi_buffer[13] ),
    .B(net542));
 sg13g2_nand2b_1 _17427_ (.Y(_10207_),
    .B(\rbzero.pov.spi_buffer[14] ),
    .A_N(net595));
 sg13g2_a21oi_1 _17428_ (.A1(_10206_),
    .A2(_10207_),
    .Y(_00613_),
    .B1(net597));
 sg13g2_nand2_1 _17429_ (.Y(_10208_),
    .A(\rbzero.pov.spi_buffer[14] ),
    .B(net542));
 sg13g2_buf_1 _17430_ (.A(_10192_),
    .X(_10209_));
 sg13g2_buf_1 _17431_ (.A(_10209_),
    .X(_10210_));
 sg13g2_nand2b_1 _17432_ (.Y(_10211_),
    .B(\rbzero.pov.spi_buffer[15] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17433_ (.A1(_10208_),
    .A2(_10211_),
    .Y(_00614_),
    .B1(net597));
 sg13g2_nand2_1 _17434_ (.Y(_10212_),
    .A(\rbzero.pov.spi_buffer[15] ),
    .B(net542));
 sg13g2_nand2b_1 _17435_ (.Y(_10213_),
    .B(\rbzero.pov.spi_buffer[16] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17436_ (.A1(_10212_),
    .A2(_10213_),
    .Y(_00615_),
    .B1(net597));
 sg13g2_nand2_1 _17437_ (.Y(_10214_),
    .A(\rbzero.pov.spi_buffer[16] ),
    .B(_10194_));
 sg13g2_nand2b_1 _17438_ (.Y(_10215_),
    .B(\rbzero.pov.spi_buffer[17] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17439_ (.A1(_10214_),
    .A2(_10215_),
    .Y(_00616_),
    .B1(_10189_));
 sg13g2_nand2_1 _17440_ (.Y(_10216_),
    .A(\rbzero.pov.spi_buffer[17] ),
    .B(_10194_));
 sg13g2_nand2b_1 _17441_ (.Y(_10217_),
    .B(\rbzero.pov.spi_buffer[18] ),
    .A_N(_10210_));
 sg13g2_buf_1 _17442_ (.A(_10143_),
    .X(_10218_));
 sg13g2_a21oi_1 _17443_ (.A1(_10216_),
    .A2(_10217_),
    .Y(_00617_),
    .B1(net594));
 sg13g2_buf_1 _17444_ (.A(net596),
    .X(_10219_));
 sg13g2_nand2_1 _17445_ (.Y(_10220_),
    .A(\rbzero.pov.spi_buffer[18] ),
    .B(net540));
 sg13g2_nand2b_1 _17446_ (.Y(_10221_),
    .B(\rbzero.pov.spi_buffer[19] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17447_ (.A1(_10220_),
    .A2(_10221_),
    .Y(_00618_),
    .B1(net594));
 sg13g2_nand2_1 _17448_ (.Y(_10222_),
    .A(\rbzero.pov.spi_buffer[0] ),
    .B(net540));
 sg13g2_nand2b_1 _17449_ (.Y(_10223_),
    .B(\rbzero.pov.spi_buffer[1] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17450_ (.A1(_10222_),
    .A2(_10223_),
    .Y(_00619_),
    .B1(net594));
 sg13g2_nand2_1 _17451_ (.Y(_10224_),
    .A(\rbzero.pov.spi_buffer[19] ),
    .B(net540));
 sg13g2_nand2b_1 _17452_ (.Y(_10225_),
    .B(\rbzero.pov.spi_buffer[20] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17453_ (.A1(_10224_),
    .A2(_10225_),
    .Y(_00620_),
    .B1(net594));
 sg13g2_nand2_1 _17454_ (.Y(_10226_),
    .A(\rbzero.pov.spi_buffer[20] ),
    .B(net540));
 sg13g2_nand2b_1 _17455_ (.Y(_10227_),
    .B(\rbzero.pov.spi_buffer[21] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17456_ (.A1(_10226_),
    .A2(_10227_),
    .Y(_00621_),
    .B1(net594));
 sg13g2_nand2_1 _17457_ (.Y(_10228_),
    .A(\rbzero.pov.spi_buffer[21] ),
    .B(net540));
 sg13g2_nand2b_1 _17458_ (.Y(_10229_),
    .B(\rbzero.pov.spi_buffer[22] ),
    .A_N(net541));
 sg13g2_a21oi_1 _17459_ (.A1(_10228_),
    .A2(_10229_),
    .Y(_00622_),
    .B1(net594));
 sg13g2_nand2_1 _17460_ (.Y(_10230_),
    .A(\rbzero.pov.spi_buffer[22] ),
    .B(_10219_));
 sg13g2_nand2b_1 _17461_ (.Y(_10231_),
    .B(\rbzero.pov.spi_buffer[23] ),
    .A_N(_10210_));
 sg13g2_a21oi_1 _17462_ (.A1(_10230_),
    .A2(_10231_),
    .Y(_00623_),
    .B1(net594));
 sg13g2_nand2_1 _17463_ (.Y(_10232_),
    .A(\rbzero.pov.spi_buffer[23] ),
    .B(net540));
 sg13g2_buf_1 _17464_ (.A(_10209_),
    .X(_10233_));
 sg13g2_nand2b_1 _17465_ (.Y(_10234_),
    .B(\rbzero.pov.spi_buffer[24] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17466_ (.A1(_10232_),
    .A2(_10234_),
    .Y(_00624_),
    .B1(_10218_));
 sg13g2_nand2_1 _17467_ (.Y(_10235_),
    .A(\rbzero.pov.spi_buffer[24] ),
    .B(net540));
 sg13g2_nand2b_1 _17468_ (.Y(_10236_),
    .B(\rbzero.pov.spi_buffer[25] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17469_ (.A1(_10235_),
    .A2(_10236_),
    .Y(_00625_),
    .B1(_10218_));
 sg13g2_nand2_1 _17470_ (.Y(_10237_),
    .A(\rbzero.pov.spi_buffer[25] ),
    .B(_10219_));
 sg13g2_nand2b_1 _17471_ (.Y(_10238_),
    .B(\rbzero.pov.spi_buffer[26] ),
    .A_N(_10233_));
 sg13g2_a21oi_1 _17472_ (.A1(_10237_),
    .A2(_10238_),
    .Y(_00626_),
    .B1(net594));
 sg13g2_nand2_1 _17473_ (.Y(_10239_),
    .A(\rbzero.pov.spi_buffer[26] ),
    .B(net540));
 sg13g2_nand2b_1 _17474_ (.Y(_10240_),
    .B(\rbzero.pov.spi_buffer[27] ),
    .A_N(net539));
 sg13g2_buf_1 _17475_ (.A(_10143_),
    .X(_10241_));
 sg13g2_a21oi_1 _17476_ (.A1(_10239_),
    .A2(_10240_),
    .Y(_00627_),
    .B1(_10241_));
 sg13g2_buf_1 _17477_ (.A(_10209_),
    .X(_10242_));
 sg13g2_nand2_1 _17478_ (.Y(_10243_),
    .A(\rbzero.pov.spi_buffer[27] ),
    .B(net538));
 sg13g2_nand2b_1 _17479_ (.Y(_10244_),
    .B(\rbzero.pov.spi_buffer[28] ),
    .A_N(_10233_));
 sg13g2_a21oi_1 _17480_ (.A1(_10243_),
    .A2(_10244_),
    .Y(_00628_),
    .B1(net593));
 sg13g2_nand2_1 _17481_ (.Y(_10245_),
    .A(\rbzero.pov.spi_buffer[28] ),
    .B(_10242_));
 sg13g2_nand2b_1 _17482_ (.Y(_10246_),
    .B(\rbzero.pov.spi_buffer[29] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17483_ (.A1(_10245_),
    .A2(_10246_),
    .Y(_00629_),
    .B1(net593));
 sg13g2_nand2_1 _17484_ (.Y(_10247_),
    .A(\rbzero.pov.spi_buffer[1] ),
    .B(_10242_));
 sg13g2_nand2b_1 _17485_ (.Y(_10248_),
    .B(\rbzero.pov.spi_buffer[2] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17486_ (.A1(_10247_),
    .A2(_10248_),
    .Y(_00630_),
    .B1(_10241_));
 sg13g2_nand2_1 _17487_ (.Y(_10249_),
    .A(\rbzero.pov.spi_buffer[29] ),
    .B(net538));
 sg13g2_nand2b_1 _17488_ (.Y(_10250_),
    .B(\rbzero.pov.spi_buffer[30] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17489_ (.A1(_10249_),
    .A2(_10250_),
    .Y(_00631_),
    .B1(net593));
 sg13g2_nand2_1 _17490_ (.Y(_10251_),
    .A(\rbzero.pov.spi_buffer[30] ),
    .B(net538));
 sg13g2_nand2b_1 _17491_ (.Y(_10252_),
    .B(\rbzero.pov.spi_buffer[31] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17492_ (.A1(_10251_),
    .A2(_10252_),
    .Y(_00632_),
    .B1(net593));
 sg13g2_nand2_1 _17493_ (.Y(_10253_),
    .A(\rbzero.pov.spi_buffer[31] ),
    .B(net538));
 sg13g2_nand2b_1 _17494_ (.Y(_10254_),
    .B(\rbzero.pov.spi_buffer[32] ),
    .A_N(net539));
 sg13g2_a21oi_1 _17495_ (.A1(_10253_),
    .A2(_10254_),
    .Y(_00633_),
    .B1(net593));
 sg13g2_nand2_1 _17496_ (.Y(_10255_),
    .A(\rbzero.pov.spi_buffer[32] ),
    .B(net538));
 sg13g2_buf_1 _17497_ (.A(_10192_),
    .X(_10256_));
 sg13g2_nand2b_1 _17498_ (.Y(_10257_),
    .B(\rbzero.pov.spi_buffer[33] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17499_ (.A1(_10255_),
    .A2(_10257_),
    .Y(_00634_),
    .B1(net593));
 sg13g2_nand2_1 _17500_ (.Y(_10258_),
    .A(\rbzero.pov.spi_buffer[33] ),
    .B(net538));
 sg13g2_nand2b_1 _17501_ (.Y(_10259_),
    .B(\rbzero.pov.spi_buffer[34] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17502_ (.A1(_10258_),
    .A2(_10259_),
    .Y(_00635_),
    .B1(net593));
 sg13g2_nand2_1 _17503_ (.Y(_10260_),
    .A(\rbzero.pov.spi_buffer[34] ),
    .B(net538));
 sg13g2_nand2b_1 _17504_ (.Y(_10261_),
    .B(\rbzero.pov.spi_buffer[35] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17505_ (.A1(_10260_),
    .A2(_10261_),
    .Y(_00636_),
    .B1(net593));
 sg13g2_nand2_1 _17506_ (.Y(_10262_),
    .A(\rbzero.pov.spi_buffer[35] ),
    .B(net538));
 sg13g2_nand2b_1 _17507_ (.Y(_10263_),
    .B(\rbzero.pov.spi_buffer[36] ),
    .A_N(net592));
 sg13g2_buf_1 _17508_ (.A(_10143_),
    .X(_10264_));
 sg13g2_a21oi_1 _17509_ (.A1(_10262_),
    .A2(_10263_),
    .Y(_00637_),
    .B1(net591));
 sg13g2_buf_1 _17510_ (.A(_10209_),
    .X(_10265_));
 sg13g2_nand2_1 _17511_ (.Y(_10266_),
    .A(\rbzero.pov.spi_buffer[36] ),
    .B(net537));
 sg13g2_nand2b_1 _17512_ (.Y(_10267_),
    .B(\rbzero.pov.spi_buffer[37] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17513_ (.A1(_10266_),
    .A2(_10267_),
    .Y(_00638_),
    .B1(net591));
 sg13g2_nand2_1 _17514_ (.Y(_10268_),
    .A(\rbzero.pov.spi_buffer[37] ),
    .B(net537));
 sg13g2_nand2b_1 _17515_ (.Y(_10269_),
    .B(\rbzero.pov.spi_buffer[38] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17516_ (.A1(_10268_),
    .A2(_10269_),
    .Y(_00639_),
    .B1(net591));
 sg13g2_nand2_1 _17517_ (.Y(_10270_),
    .A(\rbzero.pov.spi_buffer[38] ),
    .B(net537));
 sg13g2_nand2b_1 _17518_ (.Y(_10271_),
    .B(\rbzero.pov.spi_buffer[39] ),
    .A_N(_10256_));
 sg13g2_a21oi_1 _17519_ (.A1(_10270_),
    .A2(_10271_),
    .Y(_00640_),
    .B1(net591));
 sg13g2_nand2_1 _17520_ (.Y(_10272_),
    .A(\rbzero.pov.spi_buffer[2] ),
    .B(_10265_));
 sg13g2_nand2b_1 _17521_ (.Y(_10273_),
    .B(\rbzero.pov.spi_buffer[3] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17522_ (.A1(_10272_),
    .A2(_10273_),
    .Y(_00641_),
    .B1(_10264_));
 sg13g2_nand2_1 _17523_ (.Y(_10274_),
    .A(\rbzero.pov.spi_buffer[39] ),
    .B(net537));
 sg13g2_nand2b_1 _17524_ (.Y(_10275_),
    .B(\rbzero.pov.spi_buffer[40] ),
    .A_N(_10256_));
 sg13g2_a21oi_1 _17525_ (.A1(_10274_),
    .A2(_10275_),
    .Y(_00642_),
    .B1(net591));
 sg13g2_nand2_1 _17526_ (.Y(_10276_),
    .A(\rbzero.pov.spi_buffer[40] ),
    .B(_10265_));
 sg13g2_nand2b_1 _17527_ (.Y(_10277_),
    .B(\rbzero.pov.spi_buffer[41] ),
    .A_N(net592));
 sg13g2_a21oi_1 _17528_ (.A1(_10276_),
    .A2(_10277_),
    .Y(_00643_),
    .B1(net591));
 sg13g2_nand2_1 _17529_ (.Y(_10278_),
    .A(\rbzero.pov.spi_buffer[41] ),
    .B(net537));
 sg13g2_buf_1 _17530_ (.A(_10192_),
    .X(_10279_));
 sg13g2_nand2b_1 _17531_ (.Y(_10280_),
    .B(\rbzero.pov.spi_buffer[42] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17532_ (.A1(_10278_),
    .A2(_10280_),
    .Y(_00644_),
    .B1(net591));
 sg13g2_nand2_1 _17533_ (.Y(_10281_),
    .A(\rbzero.pov.spi_buffer[42] ),
    .B(net537));
 sg13g2_nand2b_1 _17534_ (.Y(_10282_),
    .B(\rbzero.pov.spi_buffer[43] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17535_ (.A1(_10281_),
    .A2(_10282_),
    .Y(_00645_),
    .B1(_10264_));
 sg13g2_nand2_1 _17536_ (.Y(_10283_),
    .A(\rbzero.pov.spi_buffer[43] ),
    .B(net537));
 sg13g2_nand2b_1 _17537_ (.Y(_10284_),
    .B(\rbzero.pov.spi_buffer[44] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17538_ (.A1(_10283_),
    .A2(_10284_),
    .Y(_00646_),
    .B1(net591));
 sg13g2_nand2_1 _17539_ (.Y(_10285_),
    .A(\rbzero.pov.spi_buffer[44] ),
    .B(net537));
 sg13g2_nand2b_1 _17540_ (.Y(_10286_),
    .B(\rbzero.pov.spi_buffer[45] ),
    .A_N(net590));
 sg13g2_buf_1 _17541_ (.A(_10143_),
    .X(_10287_));
 sg13g2_a21oi_1 _17542_ (.A1(_10285_),
    .A2(_10286_),
    .Y(_00647_),
    .B1(net589));
 sg13g2_buf_1 _17543_ (.A(_10209_),
    .X(_10288_));
 sg13g2_nand2_1 _17544_ (.Y(_10289_),
    .A(\rbzero.pov.spi_buffer[45] ),
    .B(net536));
 sg13g2_nand2b_1 _17545_ (.Y(_10290_),
    .B(\rbzero.pov.spi_buffer[46] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17546_ (.A1(_10289_),
    .A2(_10290_),
    .Y(_00648_),
    .B1(net589));
 sg13g2_nand2_1 _17547_ (.Y(_10291_),
    .A(\rbzero.pov.spi_buffer[46] ),
    .B(net536));
 sg13g2_nand2b_1 _17548_ (.Y(_10292_),
    .B(\rbzero.pov.spi_buffer[47] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17549_ (.A1(_10291_),
    .A2(_10292_),
    .Y(_00649_),
    .B1(net589));
 sg13g2_nand2_1 _17550_ (.Y(_10293_),
    .A(\rbzero.pov.spi_buffer[47] ),
    .B(net536));
 sg13g2_nand2b_1 _17551_ (.Y(_10294_),
    .B(\rbzero.pov.spi_buffer[48] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17552_ (.A1(_10293_),
    .A2(_10294_),
    .Y(_00650_),
    .B1(net589));
 sg13g2_nand2_1 _17553_ (.Y(_10295_),
    .A(\rbzero.pov.spi_buffer[48] ),
    .B(net536));
 sg13g2_nand2b_1 _17554_ (.Y(_10296_),
    .B(\rbzero.pov.spi_buffer[49] ),
    .A_N(_10279_));
 sg13g2_a21oi_1 _17555_ (.A1(_10295_),
    .A2(_10296_),
    .Y(_00651_),
    .B1(net589));
 sg13g2_nand2_1 _17556_ (.Y(_10297_),
    .A(\rbzero.pov.spi_buffer[3] ),
    .B(_10288_));
 sg13g2_nand2b_1 _17557_ (.Y(_10298_),
    .B(\rbzero.pov.spi_buffer[4] ),
    .A_N(net590));
 sg13g2_a21oi_1 _17558_ (.A1(_10297_),
    .A2(_10298_),
    .Y(_00652_),
    .B1(net589));
 sg13g2_nand2_1 _17559_ (.Y(_10299_),
    .A(\rbzero.pov.spi_buffer[49] ),
    .B(net536));
 sg13g2_nand2b_1 _17560_ (.Y(_10300_),
    .B(\rbzero.pov.spi_buffer[50] ),
    .A_N(_10279_));
 sg13g2_a21oi_1 _17561_ (.A1(_10299_),
    .A2(_10300_),
    .Y(_00653_),
    .B1(net589));
 sg13g2_nand2_1 _17562_ (.Y(_10301_),
    .A(\rbzero.pov.spi_buffer[50] ),
    .B(net536));
 sg13g2_buf_1 _17563_ (.A(_10192_),
    .X(_10302_));
 sg13g2_nand2b_1 _17564_ (.Y(_10303_),
    .B(\rbzero.pov.spi_buffer[51] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17565_ (.A1(_10301_),
    .A2(_10303_),
    .Y(_00654_),
    .B1(net589));
 sg13g2_nand2_1 _17566_ (.Y(_10304_),
    .A(\rbzero.pov.spi_buffer[51] ),
    .B(net536));
 sg13g2_nand2b_1 _17567_ (.Y(_10305_),
    .B(\rbzero.pov.spi_buffer[52] ),
    .A_N(_10302_));
 sg13g2_a21oi_1 _17568_ (.A1(_10304_),
    .A2(_10305_),
    .Y(_00655_),
    .B1(_10287_));
 sg13g2_nand2_1 _17569_ (.Y(_10306_),
    .A(\rbzero.pov.spi_buffer[52] ),
    .B(_10288_));
 sg13g2_nand2b_1 _17570_ (.Y(_10307_),
    .B(\rbzero.pov.spi_buffer[53] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17571_ (.A1(_10306_),
    .A2(_10307_),
    .Y(_00656_),
    .B1(_10287_));
 sg13g2_nand2_1 _17572_ (.Y(_10308_),
    .A(\rbzero.pov.spi_buffer[53] ),
    .B(net536));
 sg13g2_nand2b_1 _17573_ (.Y(_10309_),
    .B(\rbzero.pov.spi_buffer[54] ),
    .A_N(net588));
 sg13g2_buf_1 _17574_ (.A(_08638_),
    .X(_10310_));
 sg13g2_buf_1 _17575_ (.A(_10310_),
    .X(_10311_));
 sg13g2_a21oi_1 _17576_ (.A1(_10308_),
    .A2(_10309_),
    .Y(_00657_),
    .B1(net673));
 sg13g2_buf_1 _17577_ (.A(_10209_),
    .X(_10312_));
 sg13g2_nand2_1 _17578_ (.Y(_10313_),
    .A(\rbzero.pov.spi_buffer[54] ),
    .B(net535));
 sg13g2_nand2b_1 _17579_ (.Y(_10314_),
    .B(\rbzero.pov.spi_buffer[55] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17580_ (.A1(_10313_),
    .A2(_10314_),
    .Y(_00658_),
    .B1(net673));
 sg13g2_nand2_1 _17581_ (.Y(_10315_),
    .A(\rbzero.pov.spi_buffer[55] ),
    .B(net535));
 sg13g2_nand2b_1 _17582_ (.Y(_10316_),
    .B(\rbzero.pov.spi_buffer[56] ),
    .A_N(_10302_));
 sg13g2_a21oi_1 _17583_ (.A1(_10315_),
    .A2(_10316_),
    .Y(_00659_),
    .B1(net673));
 sg13g2_nand2_1 _17584_ (.Y(_10317_),
    .A(\rbzero.pov.spi_buffer[56] ),
    .B(_10312_));
 sg13g2_nand2b_1 _17585_ (.Y(_10318_),
    .B(\rbzero.pov.spi_buffer[57] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17586_ (.A1(_10317_),
    .A2(_10318_),
    .Y(_00660_),
    .B1(_10311_));
 sg13g2_nand2_1 _17587_ (.Y(_10319_),
    .A(\rbzero.pov.spi_buffer[57] ),
    .B(_10312_));
 sg13g2_nand2b_1 _17588_ (.Y(_10320_),
    .B(\rbzero.pov.spi_buffer[58] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17589_ (.A1(_10319_),
    .A2(_10320_),
    .Y(_00661_),
    .B1(_10311_));
 sg13g2_nand2_1 _17590_ (.Y(_10321_),
    .A(\rbzero.pov.spi_buffer[58] ),
    .B(net535));
 sg13g2_nand2b_1 _17591_ (.Y(_10322_),
    .B(\rbzero.pov.spi_buffer[59] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17592_ (.A1(_10321_),
    .A2(_10322_),
    .Y(_00662_),
    .B1(net673));
 sg13g2_nand2_1 _17593_ (.Y(_10323_),
    .A(\rbzero.pov.spi_buffer[4] ),
    .B(net535));
 sg13g2_nand2b_1 _17594_ (.Y(_10324_),
    .B(\rbzero.pov.spi_buffer[5] ),
    .A_N(net588));
 sg13g2_a21oi_1 _17595_ (.A1(_10323_),
    .A2(_10324_),
    .Y(_00663_),
    .B1(net673));
 sg13g2_nand2_1 _17596_ (.Y(_10325_),
    .A(\rbzero.pov.spi_buffer[59] ),
    .B(net535));
 sg13g2_buf_1 _17597_ (.A(_10192_),
    .X(_10326_));
 sg13g2_nand2b_1 _17598_ (.Y(_10327_),
    .B(\rbzero.pov.spi_buffer[60] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17599_ (.A1(_10325_),
    .A2(_10327_),
    .Y(_00664_),
    .B1(net673));
 sg13g2_nand2_1 _17600_ (.Y(_10328_),
    .A(\rbzero.pov.spi_buffer[60] ),
    .B(net535));
 sg13g2_nand2b_1 _17601_ (.Y(_10329_),
    .B(\rbzero.pov.spi_buffer[61] ),
    .A_N(_10326_));
 sg13g2_a21oi_1 _17602_ (.A1(_10328_),
    .A2(_10329_),
    .Y(_00665_),
    .B1(net673));
 sg13g2_nand2_1 _17603_ (.Y(_10330_),
    .A(\rbzero.pov.spi_buffer[61] ),
    .B(net535));
 sg13g2_nand2b_1 _17604_ (.Y(_10331_),
    .B(\rbzero.pov.spi_buffer[62] ),
    .A_N(_10326_));
 sg13g2_a21oi_1 _17605_ (.A1(_10330_),
    .A2(_10331_),
    .Y(_00666_),
    .B1(net673));
 sg13g2_nand2_1 _17606_ (.Y(_10332_),
    .A(\rbzero.pov.spi_buffer[62] ),
    .B(net535));
 sg13g2_nand2b_1 _17607_ (.Y(_10333_),
    .B(\rbzero.pov.spi_buffer[63] ),
    .A_N(net587));
 sg13g2_buf_1 _17608_ (.A(_10310_),
    .X(_10334_));
 sg13g2_a21oi_1 _17609_ (.A1(_10332_),
    .A2(_10333_),
    .Y(_00667_),
    .B1(net672));
 sg13g2_buf_1 _17610_ (.A(_10209_),
    .X(_10335_));
 sg13g2_nand2_1 _17611_ (.Y(_10336_),
    .A(\rbzero.pov.spi_buffer[63] ),
    .B(net534));
 sg13g2_nand2b_1 _17612_ (.Y(_10337_),
    .B(\rbzero.pov.spi_buffer[64] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17613_ (.A1(_10336_),
    .A2(_10337_),
    .Y(_00668_),
    .B1(net672));
 sg13g2_nand2_1 _17614_ (.Y(_10338_),
    .A(\rbzero.pov.spi_buffer[64] ),
    .B(net534));
 sg13g2_nand2b_1 _17615_ (.Y(_10339_),
    .B(\rbzero.pov.spi_buffer[65] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17616_ (.A1(_10338_),
    .A2(_10339_),
    .Y(_00669_),
    .B1(net672));
 sg13g2_nand2_1 _17617_ (.Y(_10340_),
    .A(\rbzero.pov.spi_buffer[65] ),
    .B(net534));
 sg13g2_nand2b_1 _17618_ (.Y(_10341_),
    .B(\rbzero.pov.spi_buffer[66] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17619_ (.A1(_10340_),
    .A2(_10341_),
    .Y(_00670_),
    .B1(_10334_));
 sg13g2_nand2_1 _17620_ (.Y(_10342_),
    .A(\rbzero.pov.spi_buffer[66] ),
    .B(_10335_));
 sg13g2_nand2b_1 _17621_ (.Y(_10343_),
    .B(\rbzero.pov.spi_buffer[67] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17622_ (.A1(_10342_),
    .A2(_10343_),
    .Y(_00671_),
    .B1(_10334_));
 sg13g2_nand2_1 _17623_ (.Y(_10344_),
    .A(\rbzero.pov.spi_buffer[67] ),
    .B(net534));
 sg13g2_nand2b_1 _17624_ (.Y(_10345_),
    .B(\rbzero.pov.spi_buffer[68] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17625_ (.A1(_10344_),
    .A2(_10345_),
    .Y(_00672_),
    .B1(net672));
 sg13g2_nand2_1 _17626_ (.Y(_10346_),
    .A(\rbzero.pov.spi_buffer[68] ),
    .B(_10335_));
 sg13g2_nand2b_1 _17627_ (.Y(_10347_),
    .B(\rbzero.pov.spi_buffer[69] ),
    .A_N(net587));
 sg13g2_a21oi_1 _17628_ (.A1(_10346_),
    .A2(_10347_),
    .Y(_00673_),
    .B1(net672));
 sg13g2_nand2_1 _17629_ (.Y(_10348_),
    .A(\rbzero.pov.spi_buffer[5] ),
    .B(net534));
 sg13g2_nand2b_1 _17630_ (.Y(_10349_),
    .B(\rbzero.pov.spi_buffer[6] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17631_ (.A1(_10348_),
    .A2(_10349_),
    .Y(_00674_),
    .B1(net672));
 sg13g2_nand2_1 _17632_ (.Y(_10350_),
    .A(\rbzero.pov.spi_buffer[69] ),
    .B(net534));
 sg13g2_nand2b_1 _17633_ (.Y(_10351_),
    .B(\rbzero.pov.spi_buffer[70] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17634_ (.A1(_10350_),
    .A2(_10351_),
    .Y(_00675_),
    .B1(net672));
 sg13g2_nand2_1 _17635_ (.Y(_10352_),
    .A(\rbzero.pov.spi_buffer[70] ),
    .B(net534));
 sg13g2_nand2b_1 _17636_ (.Y(_10353_),
    .B(\rbzero.pov.spi_buffer[71] ),
    .A_N(_10193_));
 sg13g2_a21oi_1 _17637_ (.A1(_10352_),
    .A2(_10353_),
    .Y(_00676_),
    .B1(net672));
 sg13g2_nand2_1 _17638_ (.Y(_10354_),
    .A(\rbzero.pov.spi_buffer[71] ),
    .B(net534));
 sg13g2_nand2b_1 _17639_ (.Y(_10355_),
    .B(\rbzero.pov.spi_buffer[72] ),
    .A_N(_10193_));
 sg13g2_buf_1 _17640_ (.A(_10310_),
    .X(_10356_));
 sg13g2_a21oi_1 _17641_ (.A1(_10354_),
    .A2(_10355_),
    .Y(_00677_),
    .B1(net671));
 sg13g2_nand2_1 _17642_ (.Y(_10357_),
    .A(\rbzero.pov.spi_buffer[72] ),
    .B(_10196_));
 sg13g2_nand2b_1 _17643_ (.Y(_10358_),
    .B(\rbzero.pov.spi_buffer[73] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17644_ (.A1(_10357_),
    .A2(_10358_),
    .Y(_00678_),
    .B1(net671));
 sg13g2_nand2_1 _17645_ (.Y(_10359_),
    .A(\rbzero.pov.spi_buffer[6] ),
    .B(_10196_));
 sg13g2_nand2b_1 _17646_ (.Y(_10360_),
    .B(\rbzero.pov.spi_buffer[7] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17647_ (.A1(_10359_),
    .A2(_10360_),
    .Y(_00679_),
    .B1(net671));
 sg13g2_nand2_1 _17648_ (.Y(_10361_),
    .A(\rbzero.pov.spi_buffer[7] ),
    .B(net595));
 sg13g2_nand2b_1 _17649_ (.Y(_10362_),
    .B(\rbzero.pov.spi_buffer[8] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17650_ (.A1(_10361_),
    .A2(_10362_),
    .Y(_00680_),
    .B1(net671));
 sg13g2_nand2_1 _17651_ (.Y(_10363_),
    .A(\rbzero.pov.spi_buffer[8] ),
    .B(net595));
 sg13g2_nand2b_1 _17652_ (.Y(_10364_),
    .B(\rbzero.pov.spi_buffer[9] ),
    .A_N(net596));
 sg13g2_a21oi_1 _17653_ (.A1(_10363_),
    .A2(_10364_),
    .Y(_00681_),
    .B1(net671));
 sg13g2_and2_1 _17654_ (.A(net750),
    .B(net3),
    .X(_00690_));
 sg13g2_and2_1 _17655_ (.A(_10190_),
    .B(\rbzero.pov.ss_buffer[0] ),
    .X(_00691_));
 sg13g2_nand2_1 _17656_ (.Y(_10365_),
    .A(_08815_),
    .B(net357));
 sg13g2_nand2_1 _17657_ (.Y(_10366_),
    .A(\rbzero.pov.ready_buffer[11] ),
    .B(net358));
 sg13g2_nand3_1 _17658_ (.B(_10365_),
    .C(_10366_),
    .A(net717),
    .Y(_00692_));
 sg13g2_buf_1 _17659_ (.A(net388),
    .X(_10367_));
 sg13g2_nand2_1 _17660_ (.Y(_10368_),
    .A(\rbzero.pov.ready_buffer[21] ),
    .B(net348));
 sg13g2_buf_1 _17661_ (.A(_09742_),
    .X(_10369_));
 sg13g2_nand2_1 _17662_ (.Y(_10370_),
    .A(_08831_),
    .B(_10369_));
 sg13g2_a21oi_1 _17663_ (.A1(_10368_),
    .A2(_10370_),
    .Y(_00693_),
    .B1(net671));
 sg13g2_nand2_1 _17664_ (.Y(_10371_),
    .A(\rbzero.pov.ready_buffer[12] ),
    .B(net348));
 sg13g2_nand2_1 _17665_ (.Y(_10372_),
    .A(net781),
    .B(net347));
 sg13g2_a21oi_1 _17666_ (.A1(_10371_),
    .A2(_10372_),
    .Y(_00694_),
    .B1(net671));
 sg13g2_nand2_1 _17667_ (.Y(_10373_),
    .A(\rbzero.pov.ready_buffer[13] ),
    .B(net348));
 sg13g2_nand2_1 _17668_ (.Y(_10374_),
    .A(net780),
    .B(net347));
 sg13g2_a21oi_1 _17669_ (.A1(_10373_),
    .A2(_10374_),
    .Y(_00695_),
    .B1(net671));
 sg13g2_nand2_1 _17670_ (.Y(_10375_),
    .A(\rbzero.pov.ready_buffer[14] ),
    .B(net348));
 sg13g2_nand2_1 _17671_ (.Y(_10376_),
    .A(net778),
    .B(net347));
 sg13g2_a21oi_1 _17672_ (.A1(_10375_),
    .A2(_10376_),
    .Y(_00696_),
    .B1(_10356_));
 sg13g2_nand2_1 _17673_ (.Y(_10377_),
    .A(net722),
    .B(net357));
 sg13g2_nand2_1 _17674_ (.Y(_10378_),
    .A(\rbzero.pov.ready_buffer[15] ),
    .B(net358));
 sg13g2_nand3_1 _17675_ (.B(_10377_),
    .C(_10378_),
    .A(net717),
    .Y(_00697_));
 sg13g2_buf_1 _17676_ (.A(_09424_),
    .X(_10379_));
 sg13g2_nand2_1 _17677_ (.Y(_10380_),
    .A(net779),
    .B(net357));
 sg13g2_nand2_1 _17678_ (.Y(_10381_),
    .A(\rbzero.pov.ready_buffer[16] ),
    .B(net358));
 sg13g2_nand3_1 _17679_ (.B(_10380_),
    .C(_10381_),
    .A(net749),
    .Y(_00698_));
 sg13g2_nand2_1 _17680_ (.Y(_10382_),
    .A(\rbzero.pov.ready_buffer[17] ),
    .B(net348));
 sg13g2_nand2_1 _17681_ (.Y(_10383_),
    .A(net775),
    .B(net347));
 sg13g2_a21oi_1 _17682_ (.A1(_10382_),
    .A2(_10383_),
    .Y(_00699_),
    .B1(_10356_));
 sg13g2_nand2_1 _17683_ (.Y(_10384_),
    .A(net773),
    .B(net357));
 sg13g2_nand2_1 _17684_ (.Y(_10385_),
    .A(\rbzero.pov.ready_buffer[18] ),
    .B(net358));
 sg13g2_nand3_1 _17685_ (.B(_10384_),
    .C(_10385_),
    .A(net749),
    .Y(_00700_));
 sg13g2_nand2_1 _17686_ (.Y(_10386_),
    .A(\rbzero.pov.ready_buffer[19] ),
    .B(net348));
 sg13g2_nand2_1 _17687_ (.Y(_10387_),
    .A(net772),
    .B(net347));
 sg13g2_buf_1 _17688_ (.A(_10310_),
    .X(_10388_));
 sg13g2_a21oi_1 _17689_ (.A1(_10386_),
    .A2(_10387_),
    .Y(_00701_),
    .B1(net670));
 sg13g2_nand2_1 _17690_ (.Y(_10389_),
    .A(\rbzero.pov.ready_buffer[20] ),
    .B(net348));
 sg13g2_nand2_1 _17691_ (.Y(_10390_),
    .A(net771),
    .B(net347));
 sg13g2_a21oi_1 _17692_ (.A1(_10389_),
    .A2(_10390_),
    .Y(_00702_),
    .B1(net670));
 sg13g2_nand2_1 _17693_ (.Y(_10391_),
    .A(\rbzero.pov.ready_buffer[0] ),
    .B(net348));
 sg13g2_nand2_1 _17694_ (.Y(_10392_),
    .A(net769),
    .B(net347));
 sg13g2_a21oi_1 _17695_ (.A1(_10391_),
    .A2(_10392_),
    .Y(_00703_),
    .B1(net670));
 sg13g2_nand2_1 _17696_ (.Y(_10393_),
    .A(\rbzero.pov.ready_buffer[10] ),
    .B(_10367_));
 sg13g2_nand2_1 _17697_ (.Y(_10394_),
    .A(net764),
    .B(net347));
 sg13g2_a21oi_1 _17698_ (.A1(_10393_),
    .A2(_10394_),
    .Y(_00704_),
    .B1(net670));
 sg13g2_nand2_1 _17699_ (.Y(_10395_),
    .A(\rbzero.pov.ready_buffer[1] ),
    .B(_10367_));
 sg13g2_nand2_1 _17700_ (.Y(_10396_),
    .A(net768),
    .B(_10369_));
 sg13g2_a21oi_1 _17701_ (.A1(_10395_),
    .A2(_10396_),
    .Y(_00705_),
    .B1(net670));
 sg13g2_nand2_1 _17702_ (.Y(_10397_),
    .A(\rbzero.pov.ready_buffer[2] ),
    .B(net388));
 sg13g2_nand2_1 _17703_ (.Y(_10398_),
    .A(net766),
    .B(_09742_));
 sg13g2_a21oi_1 _17704_ (.A1(_10397_),
    .A2(_10398_),
    .Y(_00706_),
    .B1(net670));
 sg13g2_nand2_1 _17705_ (.Y(_10399_),
    .A(net765),
    .B(net357));
 sg13g2_nand2_1 _17706_ (.Y(_10400_),
    .A(\rbzero.pov.ready_buffer[3] ),
    .B(net358));
 sg13g2_nand3_1 _17707_ (.B(_10399_),
    .C(_10400_),
    .A(net749),
    .Y(_00707_));
 sg13g2_nand2_1 _17708_ (.Y(_10401_),
    .A(net770),
    .B(net357));
 sg13g2_nand2_1 _17709_ (.Y(_10402_),
    .A(\rbzero.pov.ready_buffer[4] ),
    .B(net358));
 sg13g2_nand3_1 _17710_ (.B(_10401_),
    .C(_10402_),
    .A(net749),
    .Y(_00708_));
 sg13g2_nand2_1 _17711_ (.Y(_10403_),
    .A(net767),
    .B(net357));
 sg13g2_nand2_1 _17712_ (.Y(_10404_),
    .A(\rbzero.pov.ready_buffer[5] ),
    .B(_09737_));
 sg13g2_nand3_1 _17713_ (.B(_10403_),
    .C(_10404_),
    .A(_10379_),
    .Y(_00709_));
 sg13g2_nand2_1 _17714_ (.Y(_10405_),
    .A(\rbzero.pov.ready_buffer[6] ),
    .B(_09736_));
 sg13g2_nand2_1 _17715_ (.Y(_10406_),
    .A(net763),
    .B(_09742_));
 sg13g2_a21oi_1 _17716_ (.A1(_10405_),
    .A2(_10406_),
    .Y(_00710_),
    .B1(net670));
 sg13g2_nand2_1 _17717_ (.Y(_10407_),
    .A(_09292_),
    .B(net357));
 sg13g2_nand2_1 _17718_ (.Y(_10408_),
    .A(\rbzero.pov.ready_buffer[7] ),
    .B(net358));
 sg13g2_nand3_1 _17719_ (.B(_10407_),
    .C(_10408_),
    .A(_10379_),
    .Y(_00711_));
 sg13g2_nand2_1 _17720_ (.Y(_10409_),
    .A(\rbzero.pov.ready_buffer[8] ),
    .B(net388));
 sg13g2_nand2_1 _17721_ (.Y(_10410_),
    .A(net762),
    .B(_09742_));
 sg13g2_a21oi_1 _17722_ (.A1(_10409_),
    .A2(_10410_),
    .Y(_00712_),
    .B1(net670));
 sg13g2_nand2_1 _17723_ (.Y(_10411_),
    .A(\rbzero.pov.ready_buffer[9] ),
    .B(net388));
 sg13g2_nand2_1 _17724_ (.Y(_10412_),
    .A(net821),
    .B(_09742_));
 sg13g2_a21oi_1 _17725_ (.A1(_10411_),
    .A2(_10412_),
    .Y(_00713_),
    .B1(_10388_));
 sg13g2_buf_1 _17726_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(_10413_));
 sg13g2_buf_1 _17727_ (.A(_10413_),
    .X(_10414_));
 sg13g2_nand2b_1 _17728_ (.Y(_10415_),
    .B(_09461_),
    .A_N(net757));
 sg13g2_buf_2 _17729_ (.A(_10415_),
    .X(_10416_));
 sg13g2_nand2_1 _17730_ (.Y(_10417_),
    .A(_09536_),
    .B(_09505_));
 sg13g2_buf_2 _17731_ (.A(_10417_),
    .X(_10418_));
 sg13g2_nor2_1 _17732_ (.A(_10416_),
    .B(_10418_),
    .Y(_10419_));
 sg13g2_buf_1 _17733_ (.A(_10419_),
    .X(_10420_));
 sg13g2_nand2_1 _17734_ (.Y(_10421_),
    .A(net748),
    .B(_10420_));
 sg13g2_buf_1 _17735_ (.A(_10416_),
    .X(_10422_));
 sg13g2_buf_1 _17736_ (.A(_10418_),
    .X(_10423_));
 sg13g2_o21ai_1 _17737_ (.B1(\rbzero.spi_registers.buf_floor[0] ),
    .Y(_10424_),
    .A1(net586),
    .A2(_10423_));
 sg13g2_a21oi_1 _17738_ (.A1(_10421_),
    .A2(_10424_),
    .Y(_00714_),
    .B1(_10388_));
 sg13g2_o21ai_1 _17739_ (.B1(\rbzero.spi_registers.buf_floor[1] ),
    .Y(_10425_),
    .A1(net586),
    .A2(net585));
 sg13g2_buf_1 _17740_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(_10426_));
 sg13g2_buf_1 _17741_ (.A(_10426_),
    .X(_10427_));
 sg13g2_nand2_1 _17742_ (.Y(_10428_),
    .A(net747),
    .B(_10420_));
 sg13g2_nand3_1 _17743_ (.B(_10425_),
    .C(_10428_),
    .A(net749),
    .Y(_00715_));
 sg13g2_buf_1 _17744_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(_10429_));
 sg13g2_buf_1 _17745_ (.A(_10429_),
    .X(_10430_));
 sg13g2_nand2_1 _17746_ (.Y(_10431_),
    .A(net746),
    .B(_10420_));
 sg13g2_o21ai_1 _17747_ (.B1(\rbzero.spi_registers.buf_floor[2] ),
    .Y(_10432_),
    .A1(net586),
    .A2(net585));
 sg13g2_buf_1 _17748_ (.A(_10310_),
    .X(_10433_));
 sg13g2_a21oi_1 _17749_ (.A1(_10431_),
    .A2(_10432_),
    .Y(_00716_),
    .B1(net669));
 sg13g2_o21ai_1 _17750_ (.B1(\rbzero.spi_registers.buf_floor[3] ),
    .Y(_10434_),
    .A1(net586),
    .A2(net585));
 sg13g2_buf_1 _17751_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(_10435_));
 sg13g2_buf_1 _17752_ (.A(_10435_),
    .X(_10436_));
 sg13g2_nand2_1 _17753_ (.Y(_10437_),
    .A(net745),
    .B(_10420_));
 sg13g2_nand3_1 _17754_ (.B(_10434_),
    .C(_10437_),
    .A(net749),
    .Y(_00717_));
 sg13g2_buf_1 _17755_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(_10438_));
 sg13g2_buf_1 _17756_ (.A(_10438_),
    .X(_10439_));
 sg13g2_nand2_1 _17757_ (.Y(_10440_),
    .A(net744),
    .B(_10420_));
 sg13g2_o21ai_1 _17758_ (.B1(\rbzero.spi_registers.buf_floor[4] ),
    .Y(_10441_),
    .A1(_10422_),
    .A2(net585));
 sg13g2_a21oi_1 _17759_ (.A1(_10440_),
    .A2(_10441_),
    .Y(_00718_),
    .B1(net669));
 sg13g2_o21ai_1 _17760_ (.B1(\rbzero.spi_registers.buf_floor[5] ),
    .Y(_10442_),
    .A1(_10422_),
    .A2(_10423_));
 sg13g2_buf_1 _17761_ (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(_10443_));
 sg13g2_nand2_1 _17762_ (.Y(_10444_),
    .A(net814),
    .B(_10420_));
 sg13g2_nand3_1 _17763_ (.B(_10442_),
    .C(_10444_),
    .A(net749),
    .Y(_00719_));
 sg13g2_nand2_1 _17764_ (.Y(_10445_),
    .A(_09474_),
    .B(net757));
 sg13g2_buf_1 _17765_ (.A(_10445_),
    .X(_10446_));
 sg13g2_nor2_1 _17766_ (.A(_10418_),
    .B(net668),
    .Y(_10447_));
 sg13g2_buf_1 _17767_ (.A(_10447_),
    .X(_10448_));
 sg13g2_nand2_1 _17768_ (.Y(_10449_),
    .A(net748),
    .B(_10448_));
 sg13g2_buf_1 _17769_ (.A(_10418_),
    .X(_10450_));
 sg13g2_buf_1 _17770_ (.A(net668),
    .X(_10451_));
 sg13g2_o21ai_1 _17771_ (.B1(\rbzero.spi_registers.buf_leak[0] ),
    .Y(_10452_),
    .A1(net584),
    .A2(net583));
 sg13g2_a21oi_1 _17772_ (.A1(_10449_),
    .A2(_10452_),
    .Y(_00720_),
    .B1(net669));
 sg13g2_nand2_1 _17773_ (.Y(_10453_),
    .A(net747),
    .B(_10448_));
 sg13g2_o21ai_1 _17774_ (.B1(\rbzero.spi_registers.buf_leak[1] ),
    .Y(_10454_),
    .A1(net584),
    .A2(net583));
 sg13g2_a21oi_1 _17775_ (.A1(_10453_),
    .A2(_10454_),
    .Y(_00721_),
    .B1(net669));
 sg13g2_nand2_1 _17776_ (.Y(_10455_),
    .A(net746),
    .B(_10448_));
 sg13g2_o21ai_1 _17777_ (.B1(\rbzero.spi_registers.buf_leak[2] ),
    .Y(_10456_),
    .A1(_10450_),
    .A2(_10451_));
 sg13g2_a21oi_1 _17778_ (.A1(_10455_),
    .A2(_10456_),
    .Y(_00722_),
    .B1(net669));
 sg13g2_nand2_1 _17779_ (.Y(_10457_),
    .A(net745),
    .B(_10448_));
 sg13g2_o21ai_1 _17780_ (.B1(\rbzero.spi_registers.buf_leak[3] ),
    .Y(_10458_),
    .A1(_10450_),
    .A2(_10451_));
 sg13g2_a21oi_1 _17781_ (.A1(_10457_),
    .A2(_10458_),
    .Y(_00723_),
    .B1(_10433_));
 sg13g2_nand2_1 _17782_ (.Y(_10459_),
    .A(net744),
    .B(_10448_));
 sg13g2_o21ai_1 _17783_ (.B1(\rbzero.spi_registers.buf_leak[4] ),
    .Y(_10460_),
    .A1(_10418_),
    .A2(net583));
 sg13g2_a21oi_1 _17784_ (.A1(_10459_),
    .A2(_10460_),
    .Y(_00724_),
    .B1(_10433_));
 sg13g2_nand2_1 _17785_ (.Y(_10461_),
    .A(net814),
    .B(_10448_));
 sg13g2_o21ai_1 _17786_ (.B1(\rbzero.spi_registers.buf_leak[5] ),
    .Y(_10462_),
    .A1(_10418_),
    .A2(net583));
 sg13g2_a21oi_1 _17787_ (.A1(_10461_),
    .A2(_10462_),
    .Y(_00725_),
    .B1(net669));
 sg13g2_buf_2 _17788_ (.A(\rbzero.spi_registers.spi_buffer[10] ),
    .X(_10463_));
 sg13g2_nand3_1 _17789_ (.B(_09487_),
    .C(_09536_),
    .A(net756),
    .Y(_10464_));
 sg13g2_buf_2 _17790_ (.A(_10464_),
    .X(_10465_));
 sg13g2_nor2_1 _17791_ (.A(net668),
    .B(_10465_),
    .Y(_10466_));
 sg13g2_buf_1 _17792_ (.A(_10466_),
    .X(_10467_));
 sg13g2_buf_1 _17793_ (.A(_10467_),
    .X(_10468_));
 sg13g2_nand2_1 _17794_ (.Y(_10469_),
    .A(_10463_),
    .B(net511));
 sg13g2_buf_1 _17795_ (.A(_10465_),
    .X(_10470_));
 sg13g2_o21ai_1 _17796_ (.B1(\rbzero.spi_registers.buf_mapdx[0] ),
    .Y(_10471_),
    .A1(net583),
    .A2(_10470_));
 sg13g2_a21oi_1 _17797_ (.A1(_10469_),
    .A2(_10471_),
    .Y(_00726_),
    .B1(net669));
 sg13g2_buf_2 _17798_ (.A(\rbzero.spi_registers.spi_buffer[11] ),
    .X(_10472_));
 sg13g2_nand2_1 _17799_ (.Y(_10473_),
    .A(_10472_),
    .B(net511));
 sg13g2_o21ai_1 _17800_ (.B1(\rbzero.spi_registers.buf_mapdx[1] ),
    .Y(_10474_),
    .A1(net583),
    .A2(net582));
 sg13g2_a21oi_1 _17801_ (.A1(_10473_),
    .A2(_10474_),
    .Y(_00727_),
    .B1(net669));
 sg13g2_buf_2 _17802_ (.A(\rbzero.spi_registers.spi_buffer[12] ),
    .X(_10475_));
 sg13g2_nand2_1 _17803_ (.Y(_10476_),
    .A(_10475_),
    .B(net511));
 sg13g2_o21ai_1 _17804_ (.B1(\rbzero.spi_registers.buf_mapdx[2] ),
    .Y(_10477_),
    .A1(net583),
    .A2(net582));
 sg13g2_buf_1 _17805_ (.A(_10310_),
    .X(_10478_));
 sg13g2_a21oi_1 _17806_ (.A1(_10476_),
    .A2(_10477_),
    .Y(_00728_),
    .B1(net667));
 sg13g2_buf_2 _17807_ (.A(\rbzero.spi_registers.spi_buffer[13] ),
    .X(_10479_));
 sg13g2_nand2_1 _17808_ (.Y(_10480_),
    .A(_10479_),
    .B(net511));
 sg13g2_o21ai_1 _17809_ (.B1(\rbzero.spi_registers.buf_mapdx[3] ),
    .Y(_10481_),
    .A1(net583),
    .A2(net582));
 sg13g2_a21oi_1 _17810_ (.A1(_10480_),
    .A2(_10481_),
    .Y(_00729_),
    .B1(net667));
 sg13g2_buf_2 _17811_ (.A(\rbzero.spi_registers.spi_buffer[14] ),
    .X(_10482_));
 sg13g2_nand2_1 _17812_ (.Y(_10483_),
    .A(_10482_),
    .B(net511));
 sg13g2_buf_1 _17813_ (.A(net668),
    .X(_10484_));
 sg13g2_o21ai_1 _17814_ (.B1(\rbzero.spi_registers.buf_mapdx[4] ),
    .Y(_10485_),
    .A1(_10484_),
    .A2(net582));
 sg13g2_a21oi_1 _17815_ (.A1(_10483_),
    .A2(_10485_),
    .Y(_00730_),
    .B1(net667));
 sg13g2_nand2_1 _17816_ (.Y(_10486_),
    .A(net746),
    .B(net511));
 sg13g2_o21ai_1 _17817_ (.B1(\rbzero.spi_registers.buf_mapdxw[0] ),
    .Y(_10487_),
    .A1(net581),
    .A2(_10470_));
 sg13g2_a21oi_1 _17818_ (.A1(_10486_),
    .A2(_10487_),
    .Y(_00731_),
    .B1(net667));
 sg13g2_nand2_1 _17819_ (.Y(_10488_),
    .A(net745),
    .B(net511));
 sg13g2_o21ai_1 _17820_ (.B1(\rbzero.spi_registers.buf_mapdxw[1] ),
    .Y(_10489_),
    .A1(net581),
    .A2(net582));
 sg13g2_a21oi_1 _17821_ (.A1(_10488_),
    .A2(_10489_),
    .Y(_00732_),
    .B1(_10478_));
 sg13g2_nand2_1 _17822_ (.Y(_10490_),
    .A(net744),
    .B(net511));
 sg13g2_o21ai_1 _17823_ (.B1(\rbzero.spi_registers.buf_mapdy[0] ),
    .Y(_10491_),
    .A1(net581),
    .A2(net582));
 sg13g2_a21oi_1 _17824_ (.A1(_10490_),
    .A2(_10491_),
    .Y(_00733_),
    .B1(net667));
 sg13g2_nand2_1 _17825_ (.Y(_10492_),
    .A(net814),
    .B(_10468_));
 sg13g2_o21ai_1 _17826_ (.B1(\rbzero.spi_registers.buf_mapdy[1] ),
    .Y(_10493_),
    .A1(_10484_),
    .A2(net582));
 sg13g2_a21oi_1 _17827_ (.A1(_10492_),
    .A2(_10493_),
    .Y(_00734_),
    .B1(_10478_));
 sg13g2_buf_2 _17828_ (.A(\rbzero.spi_registers.spi_buffer[6] ),
    .X(_10494_));
 sg13g2_nand2_1 _17829_ (.Y(_10495_),
    .A(_10494_),
    .B(_10468_));
 sg13g2_o21ai_1 _17830_ (.B1(\rbzero.spi_registers.buf_mapdy[2] ),
    .Y(_10496_),
    .A1(net581),
    .A2(net582));
 sg13g2_a21oi_1 _17831_ (.A1(_10495_),
    .A2(_10496_),
    .Y(_00735_),
    .B1(net667));
 sg13g2_buf_2 _17832_ (.A(\rbzero.spi_registers.spi_buffer[7] ),
    .X(_10497_));
 sg13g2_nand2_1 _17833_ (.Y(_10498_),
    .A(_10497_),
    .B(_10467_));
 sg13g2_buf_1 _17834_ (.A(_10465_),
    .X(_10499_));
 sg13g2_o21ai_1 _17835_ (.B1(\rbzero.spi_registers.buf_mapdy[3] ),
    .Y(_10500_),
    .A1(net581),
    .A2(net580));
 sg13g2_a21oi_1 _17836_ (.A1(_10498_),
    .A2(_10500_),
    .Y(_00736_),
    .B1(net667));
 sg13g2_buf_2 _17837_ (.A(\rbzero.spi_registers.spi_buffer[8] ),
    .X(_10501_));
 sg13g2_nand2_1 _17838_ (.Y(_10502_),
    .A(_10501_),
    .B(_10467_));
 sg13g2_o21ai_1 _17839_ (.B1(\rbzero.spi_registers.buf_mapdy[4] ),
    .Y(_10503_),
    .A1(net581),
    .A2(net580));
 sg13g2_a21oi_1 _17840_ (.A1(_10502_),
    .A2(_10503_),
    .Y(_00737_),
    .B1(net667));
 sg13g2_nand2_1 _17841_ (.Y(_10504_),
    .A(_10414_),
    .B(_10467_));
 sg13g2_o21ai_1 _17842_ (.B1(\rbzero.spi_registers.buf_mapdyw[0] ),
    .Y(_10505_),
    .A1(net581),
    .A2(_10499_));
 sg13g2_buf_1 _17843_ (.A(_10310_),
    .X(_10506_));
 sg13g2_a21oi_1 _17844_ (.A1(_10504_),
    .A2(_10505_),
    .Y(_00738_),
    .B1(_10506_));
 sg13g2_nand2_1 _17845_ (.Y(_10507_),
    .A(net747),
    .B(_10467_));
 sg13g2_o21ai_1 _17846_ (.B1(\rbzero.spi_registers.buf_mapdyw[1] ),
    .Y(_10508_),
    .A1(net581),
    .A2(_10499_));
 sg13g2_a21oi_1 _17847_ (.A1(_10507_),
    .A2(_10508_),
    .Y(_00739_),
    .B1(net666));
 sg13g2_nor2_1 _17848_ (.A(net718),
    .B(_10418_),
    .Y(_10509_));
 sg13g2_buf_1 _17849_ (.A(_10509_),
    .X(_10510_));
 sg13g2_nand2_1 _17850_ (.Y(_10511_),
    .A(_10494_),
    .B(net533));
 sg13g2_buf_1 _17851_ (.A(net718),
    .X(_10512_));
 sg13g2_o21ai_1 _17852_ (.B1(\rbzero.spi_registers.buf_otherx[0] ),
    .Y(_10513_),
    .A1(net665),
    .A2(net585));
 sg13g2_a21oi_1 _17853_ (.A1(_10511_),
    .A2(_10513_),
    .Y(_00740_),
    .B1(_10506_));
 sg13g2_nand2_1 _17854_ (.Y(_10514_),
    .A(_10497_),
    .B(net533));
 sg13g2_o21ai_1 _17855_ (.B1(\rbzero.spi_registers.buf_otherx[1] ),
    .Y(_10515_),
    .A1(_10512_),
    .A2(net585));
 sg13g2_a21oi_1 _17856_ (.A1(_10514_),
    .A2(_10515_),
    .Y(_00741_),
    .B1(net666));
 sg13g2_nand2_1 _17857_ (.Y(_10516_),
    .A(_10501_),
    .B(net533));
 sg13g2_o21ai_1 _17858_ (.B1(\rbzero.spi_registers.buf_otherx[2] ),
    .Y(_10517_),
    .A1(net665),
    .A2(net585));
 sg13g2_a21oi_1 _17859_ (.A1(_10516_),
    .A2(_10517_),
    .Y(_00742_),
    .B1(net666));
 sg13g2_buf_2 _17860_ (.A(\rbzero.spi_registers.spi_buffer[9] ),
    .X(_10518_));
 sg13g2_nand2_1 _17861_ (.Y(_10519_),
    .A(_10518_),
    .B(_10510_));
 sg13g2_o21ai_1 _17862_ (.B1(\rbzero.spi_registers.buf_otherx[3] ),
    .Y(_10520_),
    .A1(net665),
    .A2(net585));
 sg13g2_a21oi_1 _17863_ (.A1(_10519_),
    .A2(_10520_),
    .Y(_00743_),
    .B1(net666));
 sg13g2_nand2_1 _17864_ (.Y(_10521_),
    .A(_10463_),
    .B(net533));
 sg13g2_o21ai_1 _17865_ (.B1(\rbzero.spi_registers.buf_otherx[4] ),
    .Y(_10522_),
    .A1(net665),
    .A2(net584));
 sg13g2_a21oi_1 _17866_ (.A1(_10521_),
    .A2(_10522_),
    .Y(_00744_),
    .B1(net666));
 sg13g2_nand2_1 _17867_ (.Y(_10523_),
    .A(net748),
    .B(net533));
 sg13g2_o21ai_1 _17868_ (.B1(\rbzero.spi_registers.buf_othery[0] ),
    .Y(_10524_),
    .A1(net665),
    .A2(net584));
 sg13g2_a21oi_1 _17869_ (.A1(_10523_),
    .A2(_10524_),
    .Y(_00745_),
    .B1(net666));
 sg13g2_nand2_1 _17870_ (.Y(_10525_),
    .A(net747),
    .B(net533));
 sg13g2_o21ai_1 _17871_ (.B1(\rbzero.spi_registers.buf_othery[1] ),
    .Y(_10526_),
    .A1(net665),
    .A2(net584));
 sg13g2_a21oi_1 _17872_ (.A1(_10525_),
    .A2(_10526_),
    .Y(_00746_),
    .B1(net666));
 sg13g2_nand2_1 _17873_ (.Y(_10527_),
    .A(net746),
    .B(_10510_));
 sg13g2_o21ai_1 _17874_ (.B1(\rbzero.spi_registers.buf_othery[2] ),
    .Y(_10528_),
    .A1(_10512_),
    .A2(net584));
 sg13g2_a21oi_1 _17875_ (.A1(_10527_),
    .A2(_10528_),
    .Y(_00747_),
    .B1(net666));
 sg13g2_nand2_1 _17876_ (.Y(_10529_),
    .A(net745),
    .B(net533));
 sg13g2_o21ai_1 _17877_ (.B1(\rbzero.spi_registers.buf_othery[3] ),
    .Y(_10530_),
    .A1(net665),
    .A2(net584));
 sg13g2_buf_1 _17878_ (.A(_08638_),
    .X(_10531_));
 sg13g2_buf_1 _17879_ (.A(_10531_),
    .X(_10532_));
 sg13g2_a21oi_1 _17880_ (.A1(_10529_),
    .A2(_10530_),
    .Y(_00748_),
    .B1(net664));
 sg13g2_nand2_1 _17881_ (.Y(_10533_),
    .A(net744),
    .B(net533));
 sg13g2_o21ai_1 _17882_ (.B1(\rbzero.spi_registers.buf_othery[4] ),
    .Y(_10534_),
    .A1(net665),
    .A2(net584));
 sg13g2_a21oi_1 _17883_ (.A1(_10533_),
    .A2(_10534_),
    .Y(_00749_),
    .B1(_10532_));
 sg13g2_nor3_1 _17884_ (.A(net815),
    .B(_09476_),
    .C(_10418_),
    .Y(_10535_));
 sg13g2_buf_1 _17885_ (.A(_10535_),
    .X(_10536_));
 sg13g2_nand2_1 _17886_ (.Y(_10537_),
    .A(_10414_),
    .B(net532));
 sg13g2_nand2b_1 _17887_ (.Y(_10538_),
    .B(\rbzero.spi_registers.buf_sky[0] ),
    .A_N(net532));
 sg13g2_nand3_1 _17888_ (.B(_10537_),
    .C(_10538_),
    .A(net749),
    .Y(_00750_));
 sg13g2_nand2_1 _17889_ (.Y(_10539_),
    .A(_10427_),
    .B(net532));
 sg13g2_nand2b_1 _17890_ (.Y(_10540_),
    .B(\rbzero.spi_registers.buf_sky[1] ),
    .A_N(net532));
 sg13g2_a21oi_1 _17891_ (.A1(_10539_),
    .A2(_10540_),
    .Y(_00751_),
    .B1(_10532_));
 sg13g2_nand2_1 _17892_ (.Y(_10541_),
    .A(_10430_),
    .B(_10536_));
 sg13g2_nand2b_1 _17893_ (.Y(_10542_),
    .B(\rbzero.spi_registers.buf_sky[2] ),
    .A_N(net532));
 sg13g2_nand3_1 _17894_ (.B(_10541_),
    .C(_10542_),
    .A(net751),
    .Y(_00752_));
 sg13g2_nand2_1 _17895_ (.Y(_10543_),
    .A(_10436_),
    .B(net532));
 sg13g2_nand2b_1 _17896_ (.Y(_10544_),
    .B(\rbzero.spi_registers.buf_sky[3] ),
    .A_N(_10535_));
 sg13g2_a21oi_1 _17897_ (.A1(_10543_),
    .A2(_10544_),
    .Y(_00753_),
    .B1(net664));
 sg13g2_nand2_1 _17898_ (.Y(_10545_),
    .A(_10439_),
    .B(_10536_));
 sg13g2_nand2b_1 _17899_ (.Y(_10546_),
    .B(\rbzero.spi_registers.buf_sky[4] ),
    .A_N(net532));
 sg13g2_nand3_1 _17900_ (.B(_10545_),
    .C(_10546_),
    .A(net751),
    .Y(_00754_));
 sg13g2_nand2_1 _17901_ (.Y(_10547_),
    .A(net814),
    .B(net532));
 sg13g2_nand2b_1 _17902_ (.Y(_10548_),
    .B(\rbzero.spi_registers.buf_sky[5] ),
    .A_N(_10535_));
 sg13g2_a21oi_1 _17903_ (.A1(_10547_),
    .A2(_10548_),
    .Y(_00755_),
    .B1(net664));
 sg13g2_nor2_1 _17904_ (.A(net718),
    .B(_10465_),
    .Y(_10549_));
 sg13g2_buf_1 _17905_ (.A(_10549_),
    .X(_10550_));
 sg13g2_buf_1 _17906_ (.A(_10550_),
    .X(_10551_));
 sg13g2_nand2_1 _17907_ (.Y(_10552_),
    .A(net748),
    .B(net510));
 sg13g2_buf_1 _17908_ (.A(_09513_),
    .X(_10553_));
 sg13g2_o21ai_1 _17909_ (.B1(\rbzero.spi_registers.buf_texadd0[0] ),
    .Y(_10554_),
    .A1(net663),
    .A2(net580));
 sg13g2_a21oi_1 _17910_ (.A1(_10552_),
    .A2(_10554_),
    .Y(_00756_),
    .B1(net664));
 sg13g2_nand2_1 _17911_ (.Y(_10555_),
    .A(_10463_),
    .B(net510));
 sg13g2_o21ai_1 _17912_ (.B1(\rbzero.spi_registers.buf_texadd0[10] ),
    .Y(_10556_),
    .A1(net663),
    .A2(net580));
 sg13g2_a21oi_1 _17913_ (.A1(_10555_),
    .A2(_10556_),
    .Y(_00757_),
    .B1(net664));
 sg13g2_nand2_1 _17914_ (.Y(_10557_),
    .A(_10472_),
    .B(net510));
 sg13g2_o21ai_1 _17915_ (.B1(\rbzero.spi_registers.buf_texadd0[11] ),
    .Y(_10558_),
    .A1(net663),
    .A2(net580));
 sg13g2_a21oi_1 _17916_ (.A1(_10557_),
    .A2(_10558_),
    .Y(_00758_),
    .B1(net664));
 sg13g2_nand2_1 _17917_ (.Y(_10559_),
    .A(_10475_),
    .B(_10551_));
 sg13g2_o21ai_1 _17918_ (.B1(\rbzero.spi_registers.buf_texadd0[12] ),
    .Y(_10560_),
    .A1(_10553_),
    .A2(net580));
 sg13g2_a21oi_1 _17919_ (.A1(_10559_),
    .A2(_10560_),
    .Y(_00759_),
    .B1(net664));
 sg13g2_nand2_1 _17920_ (.Y(_10561_),
    .A(_10479_),
    .B(_10551_));
 sg13g2_o21ai_1 _17921_ (.B1(\rbzero.spi_registers.buf_texadd0[13] ),
    .Y(_10562_),
    .A1(_10553_),
    .A2(net580));
 sg13g2_a21oi_1 _17922_ (.A1(_10561_),
    .A2(_10562_),
    .Y(_00760_),
    .B1(net664));
 sg13g2_nand2_1 _17923_ (.Y(_10563_),
    .A(_10482_),
    .B(net510));
 sg13g2_o21ai_1 _17924_ (.B1(\rbzero.spi_registers.buf_texadd0[14] ),
    .Y(_10564_),
    .A1(net663),
    .A2(net580));
 sg13g2_buf_1 _17925_ (.A(_10531_),
    .X(_10565_));
 sg13g2_a21oi_1 _17926_ (.A1(_10563_),
    .A2(_10564_),
    .Y(_00761_),
    .B1(_10565_));
 sg13g2_buf_1 _17927_ (.A(\rbzero.spi_registers.spi_buffer[15] ),
    .X(_10566_));
 sg13g2_nand2_1 _17928_ (.Y(_10567_),
    .A(_10566_),
    .B(net510));
 sg13g2_buf_1 _17929_ (.A(_10465_),
    .X(_10568_));
 sg13g2_o21ai_1 _17930_ (.B1(\rbzero.spi_registers.buf_texadd0[15] ),
    .Y(_10569_),
    .A1(net663),
    .A2(net579));
 sg13g2_a21oi_1 _17931_ (.A1(_10567_),
    .A2(_10569_),
    .Y(_00762_),
    .B1(_10565_));
 sg13g2_buf_1 _17932_ (.A(\rbzero.spi_registers.spi_buffer[16] ),
    .X(_10570_));
 sg13g2_nand2_1 _17933_ (.Y(_10571_),
    .A(_10570_),
    .B(net510));
 sg13g2_o21ai_1 _17934_ (.B1(\rbzero.spi_registers.buf_texadd0[16] ),
    .Y(_10572_),
    .A1(net663),
    .A2(net579));
 sg13g2_a21oi_1 _17935_ (.A1(_10571_),
    .A2(_10572_),
    .Y(_00763_),
    .B1(net662));
 sg13g2_buf_1 _17936_ (.A(\rbzero.spi_registers.spi_buffer[17] ),
    .X(_10573_));
 sg13g2_nand2_1 _17937_ (.Y(_10574_),
    .A(_10573_),
    .B(net510));
 sg13g2_o21ai_1 _17938_ (.B1(\rbzero.spi_registers.buf_texadd0[17] ),
    .Y(_10575_),
    .A1(net663),
    .A2(_10568_));
 sg13g2_a21oi_1 _17939_ (.A1(_10574_),
    .A2(_10575_),
    .Y(_00764_),
    .B1(net662));
 sg13g2_buf_1 _17940_ (.A(\rbzero.spi_registers.spi_buffer[18] ),
    .X(_10576_));
 sg13g2_nand2_1 _17941_ (.Y(_10577_),
    .A(_10576_),
    .B(net510));
 sg13g2_o21ai_1 _17942_ (.B1(\rbzero.spi_registers.buf_texadd0[18] ),
    .Y(_10578_),
    .A1(net663),
    .A2(_10568_));
 sg13g2_a21oi_1 _17943_ (.A1(_10577_),
    .A2(_10578_),
    .Y(_00765_),
    .B1(net662));
 sg13g2_buf_1 _17944_ (.A(\rbzero.spi_registers.spi_buffer[19] ),
    .X(_10579_));
 sg13g2_buf_1 _17945_ (.A(_10550_),
    .X(_10580_));
 sg13g2_nand2_1 _17946_ (.Y(_10581_),
    .A(_10579_),
    .B(net509));
 sg13g2_buf_1 _17947_ (.A(net718),
    .X(_10582_));
 sg13g2_o21ai_1 _17948_ (.B1(\rbzero.spi_registers.buf_texadd0[19] ),
    .Y(_10583_),
    .A1(net661),
    .A2(net579));
 sg13g2_a21oi_1 _17949_ (.A1(_10581_),
    .A2(_10583_),
    .Y(_00766_),
    .B1(net662));
 sg13g2_nand2_1 _17950_ (.Y(_10584_),
    .A(net747),
    .B(net509));
 sg13g2_o21ai_1 _17951_ (.B1(\rbzero.spi_registers.buf_texadd0[1] ),
    .Y(_10585_),
    .A1(net661),
    .A2(net579));
 sg13g2_a21oi_1 _17952_ (.A1(_10584_),
    .A2(_10585_),
    .Y(_00767_),
    .B1(net662));
 sg13g2_buf_1 _17953_ (.A(\rbzero.spi_registers.spi_buffer[20] ),
    .X(_10586_));
 sg13g2_nand2_1 _17954_ (.Y(_10587_),
    .A(_10586_),
    .B(net509));
 sg13g2_o21ai_1 _17955_ (.B1(\rbzero.spi_registers.buf_texadd0[20] ),
    .Y(_10588_),
    .A1(net661),
    .A2(net579));
 sg13g2_a21oi_1 _17956_ (.A1(_10587_),
    .A2(_10588_),
    .Y(_00768_),
    .B1(net662));
 sg13g2_buf_1 _17957_ (.A(\rbzero.spi_registers.spi_buffer[21] ),
    .X(_10589_));
 sg13g2_nand2_1 _17958_ (.Y(_10590_),
    .A(_10589_),
    .B(net509));
 sg13g2_o21ai_1 _17959_ (.B1(\rbzero.spi_registers.buf_texadd0[21] ),
    .Y(_10591_),
    .A1(net661),
    .A2(net579));
 sg13g2_a21oi_1 _17960_ (.A1(_10590_),
    .A2(_10591_),
    .Y(_00769_),
    .B1(net662));
 sg13g2_buf_1 _17961_ (.A(\rbzero.spi_registers.spi_buffer[22] ),
    .X(_10592_));
 sg13g2_nand2_1 _17962_ (.Y(_10593_),
    .A(_10592_),
    .B(net509));
 sg13g2_o21ai_1 _17963_ (.B1(\rbzero.spi_registers.buf_texadd0[22] ),
    .Y(_10594_),
    .A1(net661),
    .A2(net579));
 sg13g2_a21oi_1 _17964_ (.A1(_10593_),
    .A2(_10594_),
    .Y(_00770_),
    .B1(net662));
 sg13g2_buf_1 _17965_ (.A(\rbzero.spi_registers.spi_buffer[23] ),
    .X(_10595_));
 sg13g2_nand2_1 _17966_ (.Y(_10596_),
    .A(_10595_),
    .B(net509));
 sg13g2_o21ai_1 _17967_ (.B1(\rbzero.spi_registers.buf_texadd0[23] ),
    .Y(_10597_),
    .A1(net661),
    .A2(net579));
 sg13g2_buf_1 _17968_ (.A(_10531_),
    .X(_10598_));
 sg13g2_a21oi_1 _17969_ (.A1(_10596_),
    .A2(_10597_),
    .Y(_00771_),
    .B1(_10598_));
 sg13g2_nand2_1 _17970_ (.Y(_10599_),
    .A(net746),
    .B(net509));
 sg13g2_buf_1 _17971_ (.A(_10465_),
    .X(_10600_));
 sg13g2_o21ai_1 _17972_ (.B1(\rbzero.spi_registers.buf_texadd0[2] ),
    .Y(_10601_),
    .A1(net661),
    .A2(net578));
 sg13g2_a21oi_1 _17973_ (.A1(_10599_),
    .A2(_10601_),
    .Y(_00772_),
    .B1(net660));
 sg13g2_nand2_1 _17974_ (.Y(_10602_),
    .A(net745),
    .B(net509));
 sg13g2_o21ai_1 _17975_ (.B1(\rbzero.spi_registers.buf_texadd0[3] ),
    .Y(_10603_),
    .A1(net661),
    .A2(net578));
 sg13g2_a21oi_1 _17976_ (.A1(_10602_),
    .A2(_10603_),
    .Y(_00773_),
    .B1(net660));
 sg13g2_nand2_1 _17977_ (.Y(_10604_),
    .A(net744),
    .B(_10580_));
 sg13g2_o21ai_1 _17978_ (.B1(\rbzero.spi_registers.buf_texadd0[4] ),
    .Y(_10605_),
    .A1(_10582_),
    .A2(net578));
 sg13g2_a21oi_1 _17979_ (.A1(_10604_),
    .A2(_10605_),
    .Y(_00774_),
    .B1(net660));
 sg13g2_nand2_1 _17980_ (.Y(_10606_),
    .A(net814),
    .B(_10580_));
 sg13g2_o21ai_1 _17981_ (.B1(\rbzero.spi_registers.buf_texadd0[5] ),
    .Y(_10607_),
    .A1(_10582_),
    .A2(net578));
 sg13g2_a21oi_1 _17982_ (.A1(_10606_),
    .A2(_10607_),
    .Y(_00775_),
    .B1(net660));
 sg13g2_nand2_1 _17983_ (.Y(_10608_),
    .A(_10494_),
    .B(_10550_));
 sg13g2_o21ai_1 _17984_ (.B1(\rbzero.spi_registers.buf_texadd0[6] ),
    .Y(_10609_),
    .A1(net718),
    .A2(net578));
 sg13g2_a21oi_1 _17985_ (.A1(_10608_),
    .A2(_10609_),
    .Y(_00776_),
    .B1(net660));
 sg13g2_nand2_1 _17986_ (.Y(_10610_),
    .A(_10497_),
    .B(_10550_));
 sg13g2_o21ai_1 _17987_ (.B1(\rbzero.spi_registers.buf_texadd0[7] ),
    .Y(_10611_),
    .A1(net718),
    .A2(net578));
 sg13g2_a21oi_1 _17988_ (.A1(_10610_),
    .A2(_10611_),
    .Y(_00777_),
    .B1(net660));
 sg13g2_nand2_1 _17989_ (.Y(_10612_),
    .A(_10501_),
    .B(_10550_));
 sg13g2_o21ai_1 _17990_ (.B1(\rbzero.spi_registers.buf_texadd0[8] ),
    .Y(_10613_),
    .A1(net718),
    .A2(net578));
 sg13g2_a21oi_1 _17991_ (.A1(_10612_),
    .A2(_10613_),
    .Y(_00778_),
    .B1(net660));
 sg13g2_nand2_1 _17992_ (.Y(_10614_),
    .A(_10518_),
    .B(_10550_));
 sg13g2_o21ai_1 _17993_ (.B1(\rbzero.spi_registers.buf_texadd0[9] ),
    .Y(_10615_),
    .A1(net718),
    .A2(net578));
 sg13g2_a21oi_1 _17994_ (.A1(_10614_),
    .A2(_10615_),
    .Y(_00779_),
    .B1(net660));
 sg13g2_nand2_1 _17995_ (.Y(_10616_),
    .A(_09536_),
    .B(_09514_));
 sg13g2_buf_1 _17996_ (.A(_10616_),
    .X(_10617_));
 sg13g2_nor3_1 _17997_ (.A(net815),
    .B(net757),
    .C(_10617_),
    .Y(_10618_));
 sg13g2_buf_1 _17998_ (.A(_10618_),
    .X(_10619_));
 sg13g2_buf_1 _17999_ (.A(_10619_),
    .X(_10620_));
 sg13g2_buf_1 _18000_ (.A(net489),
    .X(_10621_));
 sg13g2_nand2_1 _18001_ (.Y(_10622_),
    .A(net748),
    .B(net471));
 sg13g2_buf_1 _18002_ (.A(_10619_),
    .X(_10623_));
 sg13g2_nand2b_1 _18003_ (.Y(_10624_),
    .B(\rbzero.spi_registers.buf_texadd1[0] ),
    .A_N(net488));
 sg13g2_a21oi_1 _18004_ (.A1(_10622_),
    .A2(_10624_),
    .Y(_00780_),
    .B1(_10598_));
 sg13g2_nand2_1 _18005_ (.Y(_10625_),
    .A(_10463_),
    .B(net471));
 sg13g2_nand2b_1 _18006_ (.Y(_10626_),
    .B(\rbzero.spi_registers.buf_texadd1[10] ),
    .A_N(net488));
 sg13g2_buf_1 _18007_ (.A(_10531_),
    .X(_10627_));
 sg13g2_a21oi_1 _18008_ (.A1(_10625_),
    .A2(_10626_),
    .Y(_00781_),
    .B1(net659));
 sg13g2_nand2_1 _18009_ (.Y(_10628_),
    .A(_10472_),
    .B(net471));
 sg13g2_nand2b_1 _18010_ (.Y(_10629_),
    .B(\rbzero.spi_registers.buf_texadd1[11] ),
    .A_N(net488));
 sg13g2_a21oi_1 _18011_ (.A1(_10628_),
    .A2(_10629_),
    .Y(_00782_),
    .B1(_10627_));
 sg13g2_nand2_1 _18012_ (.Y(_10630_),
    .A(_10475_),
    .B(net471));
 sg13g2_nand2b_1 _18013_ (.Y(_10631_),
    .B(\rbzero.spi_registers.buf_texadd1[12] ),
    .A_N(net488));
 sg13g2_a21oi_1 _18014_ (.A1(_10630_),
    .A2(_10631_),
    .Y(_00783_),
    .B1(_10627_));
 sg13g2_nand2_1 _18015_ (.Y(_10632_),
    .A(_10479_),
    .B(_10621_));
 sg13g2_nand2b_1 _18016_ (.Y(_10633_),
    .B(\rbzero.spi_registers.buf_texadd1[13] ),
    .A_N(net488));
 sg13g2_a21oi_1 _18017_ (.A1(_10632_),
    .A2(_10633_),
    .Y(_00784_),
    .B1(net659));
 sg13g2_nand2_1 _18018_ (.Y(_10634_),
    .A(_10482_),
    .B(_10621_));
 sg13g2_nand2b_1 _18019_ (.Y(_10635_),
    .B(\rbzero.spi_registers.buf_texadd1[14] ),
    .A_N(net488));
 sg13g2_a21oi_1 _18020_ (.A1(_10634_),
    .A2(_10635_),
    .Y(_00785_),
    .B1(net659));
 sg13g2_nand2_1 _18021_ (.Y(_10636_),
    .A(_10566_),
    .B(net471));
 sg13g2_buf_1 _18022_ (.A(_10619_),
    .X(_10637_));
 sg13g2_nand2b_1 _18023_ (.Y(_10638_),
    .B(\rbzero.spi_registers.buf_texadd1[15] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18024_ (.A1(_10636_),
    .A2(_10638_),
    .Y(_00786_),
    .B1(net659));
 sg13g2_nand2_1 _18025_ (.Y(_10639_),
    .A(_10570_),
    .B(net471));
 sg13g2_nand2b_1 _18026_ (.Y(_10640_),
    .B(\rbzero.spi_registers.buf_texadd1[16] ),
    .A_N(_10637_));
 sg13g2_a21oi_1 _18027_ (.A1(_10639_),
    .A2(_10640_),
    .Y(_00787_),
    .B1(net659));
 sg13g2_nand2_1 _18028_ (.Y(_10641_),
    .A(_10573_),
    .B(net471));
 sg13g2_nand2b_1 _18029_ (.Y(_10642_),
    .B(\rbzero.spi_registers.buf_texadd1[17] ),
    .A_N(_10637_));
 sg13g2_a21oi_1 _18030_ (.A1(_10641_),
    .A2(_10642_),
    .Y(_00788_),
    .B1(net659));
 sg13g2_nand2_1 _18031_ (.Y(_10643_),
    .A(_10576_),
    .B(net471));
 sg13g2_nand2b_1 _18032_ (.Y(_10644_),
    .B(\rbzero.spi_registers.buf_texadd1[18] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18033_ (.A1(_10643_),
    .A2(_10644_),
    .Y(_00789_),
    .B1(net659));
 sg13g2_buf_1 _18034_ (.A(net489),
    .X(_10645_));
 sg13g2_nand2_1 _18035_ (.Y(_10646_),
    .A(_10579_),
    .B(net470));
 sg13g2_nand2b_1 _18036_ (.Y(_10647_),
    .B(\rbzero.spi_registers.buf_texadd1[19] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18037_ (.A1(_10646_),
    .A2(_10647_),
    .Y(_00790_),
    .B1(net659));
 sg13g2_nand2_1 _18038_ (.Y(_10648_),
    .A(net747),
    .B(net470));
 sg13g2_nand2b_1 _18039_ (.Y(_10649_),
    .B(\rbzero.spi_registers.buf_texadd1[1] ),
    .A_N(net487));
 sg13g2_buf_1 _18040_ (.A(_10531_),
    .X(_10650_));
 sg13g2_a21oi_1 _18041_ (.A1(_10648_),
    .A2(_10649_),
    .Y(_00791_),
    .B1(net658));
 sg13g2_nand2_1 _18042_ (.Y(_10651_),
    .A(_10586_),
    .B(net470));
 sg13g2_nand2b_1 _18043_ (.Y(_10652_),
    .B(\rbzero.spi_registers.buf_texadd1[20] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18044_ (.A1(_10651_),
    .A2(_10652_),
    .Y(_00792_),
    .B1(net658));
 sg13g2_nand2_1 _18045_ (.Y(_10653_),
    .A(_10589_),
    .B(net470));
 sg13g2_nand2b_1 _18046_ (.Y(_10654_),
    .B(\rbzero.spi_registers.buf_texadd1[21] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18047_ (.A1(_10653_),
    .A2(_10654_),
    .Y(_00793_),
    .B1(net658));
 sg13g2_nand2_1 _18048_ (.Y(_10655_),
    .A(_10592_),
    .B(net470));
 sg13g2_nand2b_1 _18049_ (.Y(_10656_),
    .B(\rbzero.spi_registers.buf_texadd1[22] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18050_ (.A1(_10655_),
    .A2(_10656_),
    .Y(_00794_),
    .B1(net658));
 sg13g2_nand2_1 _18051_ (.Y(_10657_),
    .A(_10595_),
    .B(net470));
 sg13g2_nand2b_1 _18052_ (.Y(_10658_),
    .B(\rbzero.spi_registers.buf_texadd1[23] ),
    .A_N(net487));
 sg13g2_a21oi_1 _18053_ (.A1(_10657_),
    .A2(_10658_),
    .Y(_00795_),
    .B1(net658));
 sg13g2_nand2_1 _18054_ (.Y(_10659_),
    .A(net746),
    .B(net470));
 sg13g2_nand2b_1 _18055_ (.Y(_10660_),
    .B(\rbzero.spi_registers.buf_texadd1[2] ),
    .A_N(net489));
 sg13g2_a21oi_1 _18056_ (.A1(_10659_),
    .A2(_10660_),
    .Y(_00796_),
    .B1(_10650_));
 sg13g2_nand2_1 _18057_ (.Y(_10661_),
    .A(net745),
    .B(net470));
 sg13g2_nand2b_1 _18058_ (.Y(_10662_),
    .B(\rbzero.spi_registers.buf_texadd1[3] ),
    .A_N(net489));
 sg13g2_a21oi_1 _18059_ (.A1(_10661_),
    .A2(_10662_),
    .Y(_00797_),
    .B1(net658));
 sg13g2_nand2_1 _18060_ (.Y(_10663_),
    .A(net744),
    .B(_10645_));
 sg13g2_nand2b_1 _18061_ (.Y(_10664_),
    .B(\rbzero.spi_registers.buf_texadd1[4] ),
    .A_N(net489));
 sg13g2_a21oi_1 _18062_ (.A1(_10663_),
    .A2(_10664_),
    .Y(_00798_),
    .B1(net658));
 sg13g2_nand2_1 _18063_ (.Y(_10665_),
    .A(net814),
    .B(_10645_));
 sg13g2_nand2b_1 _18064_ (.Y(_10666_),
    .B(\rbzero.spi_registers.buf_texadd1[5] ),
    .A_N(net489));
 sg13g2_a21oi_1 _18065_ (.A1(_10665_),
    .A2(_10666_),
    .Y(_00799_),
    .B1(net658));
 sg13g2_nand2_1 _18066_ (.Y(_10667_),
    .A(_10494_),
    .B(net488));
 sg13g2_nand2b_1 _18067_ (.Y(_10668_),
    .B(\rbzero.spi_registers.buf_texadd1[6] ),
    .A_N(net489));
 sg13g2_a21oi_1 _18068_ (.A1(_10667_),
    .A2(_10668_),
    .Y(_00800_),
    .B1(_10650_));
 sg13g2_nand2_1 _18069_ (.Y(_10669_),
    .A(_10497_),
    .B(net488));
 sg13g2_nand2b_1 _18070_ (.Y(_10670_),
    .B(\rbzero.spi_registers.buf_texadd1[7] ),
    .A_N(net489));
 sg13g2_buf_1 _18071_ (.A(_10531_),
    .X(_10671_));
 sg13g2_a21oi_1 _18072_ (.A1(_10669_),
    .A2(_10670_),
    .Y(_00801_),
    .B1(_10671_));
 sg13g2_nand2_1 _18073_ (.Y(_10672_),
    .A(_10501_),
    .B(_10623_));
 sg13g2_nand2b_1 _18074_ (.Y(_10673_),
    .B(\rbzero.spi_registers.buf_texadd1[8] ),
    .A_N(_10620_));
 sg13g2_a21oi_1 _18075_ (.A1(_10672_),
    .A2(_10673_),
    .Y(_00802_),
    .B1(net657));
 sg13g2_nand2_1 _18076_ (.Y(_10674_),
    .A(_10518_),
    .B(_10623_));
 sg13g2_nand2b_1 _18077_ (.Y(_10675_),
    .B(\rbzero.spi_registers.buf_texadd1[9] ),
    .A_N(_10620_));
 sg13g2_a21oi_1 _18078_ (.A1(_10674_),
    .A2(_10675_),
    .Y(_00803_),
    .B1(_10671_));
 sg13g2_nor2_1 _18079_ (.A(_10416_),
    .B(_10617_),
    .Y(_10676_));
 sg13g2_buf_1 _18080_ (.A(_10676_),
    .X(_10677_));
 sg13g2_buf_1 _18081_ (.A(_10677_),
    .X(_10678_));
 sg13g2_nand2_1 _18082_ (.Y(_10679_),
    .A(net748),
    .B(net486));
 sg13g2_buf_1 _18083_ (.A(_10617_),
    .X(_10680_));
 sg13g2_buf_1 _18084_ (.A(net531),
    .X(_10681_));
 sg13g2_o21ai_1 _18085_ (.B1(\rbzero.spi_registers.buf_texadd2[0] ),
    .Y(_10682_),
    .A1(net586),
    .A2(net508));
 sg13g2_a21oi_1 _18086_ (.A1(_10679_),
    .A2(_10682_),
    .Y(_00804_),
    .B1(net657));
 sg13g2_nand2_1 _18087_ (.Y(_10683_),
    .A(_10463_),
    .B(net486));
 sg13g2_o21ai_1 _18088_ (.B1(\rbzero.spi_registers.buf_texadd2[10] ),
    .Y(_10684_),
    .A1(net586),
    .A2(net508));
 sg13g2_a21oi_1 _18089_ (.A1(_10683_),
    .A2(_10684_),
    .Y(_00805_),
    .B1(net657));
 sg13g2_nand2_1 _18090_ (.Y(_10685_),
    .A(_10472_),
    .B(_10678_));
 sg13g2_o21ai_1 _18091_ (.B1(\rbzero.spi_registers.buf_texadd2[11] ),
    .Y(_10686_),
    .A1(net586),
    .A2(_10681_));
 sg13g2_a21oi_1 _18092_ (.A1(_10685_),
    .A2(_10686_),
    .Y(_00806_),
    .B1(net657));
 sg13g2_nand2_1 _18093_ (.Y(_10687_),
    .A(_10475_),
    .B(net486));
 sg13g2_o21ai_1 _18094_ (.B1(\rbzero.spi_registers.buf_texadd2[12] ),
    .Y(_10688_),
    .A1(net586),
    .A2(net508));
 sg13g2_a21oi_1 _18095_ (.A1(_10687_),
    .A2(_10688_),
    .Y(_00807_),
    .B1(net657));
 sg13g2_nand2_1 _18096_ (.Y(_10689_),
    .A(_10479_),
    .B(net486));
 sg13g2_buf_1 _18097_ (.A(_10416_),
    .X(_10690_));
 sg13g2_o21ai_1 _18098_ (.B1(\rbzero.spi_registers.buf_texadd2[13] ),
    .Y(_10691_),
    .A1(net577),
    .A2(net508));
 sg13g2_a21oi_1 _18099_ (.A1(_10689_),
    .A2(_10691_),
    .Y(_00808_),
    .B1(net657));
 sg13g2_nand2_1 _18100_ (.Y(_10692_),
    .A(_10482_),
    .B(net486));
 sg13g2_o21ai_1 _18101_ (.B1(\rbzero.spi_registers.buf_texadd2[14] ),
    .Y(_10693_),
    .A1(net577),
    .A2(net508));
 sg13g2_a21oi_1 _18102_ (.A1(_10692_),
    .A2(_10693_),
    .Y(_00809_),
    .B1(net657));
 sg13g2_nand2_1 _18103_ (.Y(_10694_),
    .A(_10566_),
    .B(_10678_));
 sg13g2_o21ai_1 _18104_ (.B1(\rbzero.spi_registers.buf_texadd2[15] ),
    .Y(_10695_),
    .A1(net577),
    .A2(_10681_));
 sg13g2_a21oi_1 _18105_ (.A1(_10694_),
    .A2(_10695_),
    .Y(_00810_),
    .B1(net657));
 sg13g2_nand2_1 _18106_ (.Y(_10696_),
    .A(_10570_),
    .B(net486));
 sg13g2_o21ai_1 _18107_ (.B1(\rbzero.spi_registers.buf_texadd2[16] ),
    .Y(_10697_),
    .A1(net577),
    .A2(net508));
 sg13g2_buf_1 _18108_ (.A(_10531_),
    .X(_10698_));
 sg13g2_a21oi_1 _18109_ (.A1(_10696_),
    .A2(_10697_),
    .Y(_00811_),
    .B1(net656));
 sg13g2_nand2_1 _18110_ (.Y(_10699_),
    .A(_10573_),
    .B(net486));
 sg13g2_o21ai_1 _18111_ (.B1(\rbzero.spi_registers.buf_texadd2[17] ),
    .Y(_10700_),
    .A1(_10690_),
    .A2(net508));
 sg13g2_a21oi_1 _18112_ (.A1(_10699_),
    .A2(_10700_),
    .Y(_00812_),
    .B1(net656));
 sg13g2_nand2_1 _18113_ (.Y(_10701_),
    .A(_10576_),
    .B(net486));
 sg13g2_o21ai_1 _18114_ (.B1(\rbzero.spi_registers.buf_texadd2[18] ),
    .Y(_10702_),
    .A1(_10690_),
    .A2(net508));
 sg13g2_a21oi_1 _18115_ (.A1(_10701_),
    .A2(_10702_),
    .Y(_00813_),
    .B1(_10698_));
 sg13g2_buf_1 _18116_ (.A(_10677_),
    .X(_10703_));
 sg13g2_nand2_1 _18117_ (.Y(_10704_),
    .A(_10579_),
    .B(net485));
 sg13g2_buf_1 _18118_ (.A(net531),
    .X(_10705_));
 sg13g2_o21ai_1 _18119_ (.B1(\rbzero.spi_registers.buf_texadd2[19] ),
    .Y(_10706_),
    .A1(net577),
    .A2(net507));
 sg13g2_a21oi_1 _18120_ (.A1(_10704_),
    .A2(_10706_),
    .Y(_00814_),
    .B1(net656));
 sg13g2_nand2_1 _18121_ (.Y(_10707_),
    .A(net747),
    .B(net485));
 sg13g2_o21ai_1 _18122_ (.B1(\rbzero.spi_registers.buf_texadd2[1] ),
    .Y(_10708_),
    .A1(net577),
    .A2(net507));
 sg13g2_a21oi_1 _18123_ (.A1(_10707_),
    .A2(_10708_),
    .Y(_00815_),
    .B1(net656));
 sg13g2_nand2_1 _18124_ (.Y(_10709_),
    .A(_10586_),
    .B(net485));
 sg13g2_o21ai_1 _18125_ (.B1(\rbzero.spi_registers.buf_texadd2[20] ),
    .Y(_10710_),
    .A1(net577),
    .A2(net507));
 sg13g2_a21oi_1 _18126_ (.A1(_10709_),
    .A2(_10710_),
    .Y(_00816_),
    .B1(net656));
 sg13g2_nand2_1 _18127_ (.Y(_10711_),
    .A(_10589_),
    .B(net485));
 sg13g2_o21ai_1 _18128_ (.B1(\rbzero.spi_registers.buf_texadd2[21] ),
    .Y(_10712_),
    .A1(net577),
    .A2(net507));
 sg13g2_a21oi_1 _18129_ (.A1(_10711_),
    .A2(_10712_),
    .Y(_00817_),
    .B1(net656));
 sg13g2_nand2_1 _18130_ (.Y(_10713_),
    .A(_10592_),
    .B(net485));
 sg13g2_buf_1 _18131_ (.A(_10416_),
    .X(_10714_));
 sg13g2_o21ai_1 _18132_ (.B1(\rbzero.spi_registers.buf_texadd2[22] ),
    .Y(_10715_),
    .A1(net576),
    .A2(net507));
 sg13g2_a21oi_1 _18133_ (.A1(_10713_),
    .A2(_10715_),
    .Y(_00818_),
    .B1(net656));
 sg13g2_nand2_1 _18134_ (.Y(_10716_),
    .A(_10595_),
    .B(net485));
 sg13g2_o21ai_1 _18135_ (.B1(\rbzero.spi_registers.buf_texadd2[23] ),
    .Y(_10717_),
    .A1(net576),
    .A2(net507));
 sg13g2_a21oi_1 _18136_ (.A1(_10716_),
    .A2(_10717_),
    .Y(_00819_),
    .B1(net656));
 sg13g2_nand2_1 _18137_ (.Y(_10718_),
    .A(net746),
    .B(net485));
 sg13g2_o21ai_1 _18138_ (.B1(\rbzero.spi_registers.buf_texadd2[2] ),
    .Y(_10719_),
    .A1(net576),
    .A2(net507));
 sg13g2_a21oi_1 _18139_ (.A1(_10718_),
    .A2(_10719_),
    .Y(_00820_),
    .B1(_10698_));
 sg13g2_nand2_1 _18140_ (.Y(_10720_),
    .A(net745),
    .B(net485));
 sg13g2_o21ai_1 _18141_ (.B1(\rbzero.spi_registers.buf_texadd2[3] ),
    .Y(_10721_),
    .A1(net576),
    .A2(net507));
 sg13g2_buf_1 _18142_ (.A(_08638_),
    .X(_10722_));
 sg13g2_buf_1 _18143_ (.A(_10722_),
    .X(_10723_));
 sg13g2_a21oi_1 _18144_ (.A1(_10720_),
    .A2(_10721_),
    .Y(_00821_),
    .B1(net655));
 sg13g2_nand2_1 _18145_ (.Y(_10724_),
    .A(net744),
    .B(_10703_));
 sg13g2_o21ai_1 _18146_ (.B1(\rbzero.spi_registers.buf_texadd2[4] ),
    .Y(_10725_),
    .A1(net576),
    .A2(_10705_));
 sg13g2_a21oi_1 _18147_ (.A1(_10724_),
    .A2(_10725_),
    .Y(_00822_),
    .B1(net655));
 sg13g2_nand2_1 _18148_ (.Y(_10726_),
    .A(net814),
    .B(_10703_));
 sg13g2_o21ai_1 _18149_ (.B1(\rbzero.spi_registers.buf_texadd2[5] ),
    .Y(_10727_),
    .A1(_10714_),
    .A2(_10705_));
 sg13g2_a21oi_1 _18150_ (.A1(_10726_),
    .A2(_10727_),
    .Y(_00823_),
    .B1(net655));
 sg13g2_nand2_1 _18151_ (.Y(_10728_),
    .A(_10494_),
    .B(_10677_));
 sg13g2_buf_1 _18152_ (.A(_10617_),
    .X(_10729_));
 sg13g2_o21ai_1 _18153_ (.B1(\rbzero.spi_registers.buf_texadd2[6] ),
    .Y(_10730_),
    .A1(net576),
    .A2(net530));
 sg13g2_a21oi_1 _18154_ (.A1(_10728_),
    .A2(_10730_),
    .Y(_00824_),
    .B1(net655));
 sg13g2_nand2_1 _18155_ (.Y(_10731_),
    .A(_10497_),
    .B(_10677_));
 sg13g2_o21ai_1 _18156_ (.B1(\rbzero.spi_registers.buf_texadd2[7] ),
    .Y(_10732_),
    .A1(net576),
    .A2(net530));
 sg13g2_a21oi_1 _18157_ (.A1(_10731_),
    .A2(_10732_),
    .Y(_00825_),
    .B1(net655));
 sg13g2_nand2_1 _18158_ (.Y(_10733_),
    .A(_10501_),
    .B(_10677_));
 sg13g2_o21ai_1 _18159_ (.B1(\rbzero.spi_registers.buf_texadd2[8] ),
    .Y(_10734_),
    .A1(net576),
    .A2(_10729_));
 sg13g2_a21oi_1 _18160_ (.A1(_10733_),
    .A2(_10734_),
    .Y(_00826_),
    .B1(net655));
 sg13g2_nand2_1 _18161_ (.Y(_10735_),
    .A(_10518_),
    .B(_10677_));
 sg13g2_o21ai_1 _18162_ (.B1(\rbzero.spi_registers.buf_texadd2[9] ),
    .Y(_10736_),
    .A1(_10714_),
    .A2(_10729_));
 sg13g2_a21oi_1 _18163_ (.A1(_10735_),
    .A2(_10736_),
    .Y(_00827_),
    .B1(net655));
 sg13g2_nor2_1 _18164_ (.A(_10445_),
    .B(_10617_),
    .Y(_10737_));
 sg13g2_buf_1 _18165_ (.A(_10737_),
    .X(_10738_));
 sg13g2_buf_1 _18166_ (.A(_10738_),
    .X(_10739_));
 sg13g2_nand2_1 _18167_ (.Y(_10740_),
    .A(net748),
    .B(net484));
 sg13g2_buf_1 _18168_ (.A(net668),
    .X(_10741_));
 sg13g2_o21ai_1 _18169_ (.B1(\rbzero.spi_registers.buf_texadd3[0] ),
    .Y(_10742_),
    .A1(net575),
    .A2(net530));
 sg13g2_a21oi_1 _18170_ (.A1(_10740_),
    .A2(_10742_),
    .Y(_00828_),
    .B1(net655));
 sg13g2_nand2_1 _18171_ (.Y(_10743_),
    .A(_10463_),
    .B(net484));
 sg13g2_o21ai_1 _18172_ (.B1(\rbzero.spi_registers.buf_texadd3[10] ),
    .Y(_10744_),
    .A1(net575),
    .A2(net530));
 sg13g2_a21oi_1 _18173_ (.A1(_10743_),
    .A2(_10744_),
    .Y(_00829_),
    .B1(_10723_));
 sg13g2_nand2_1 _18174_ (.Y(_10745_),
    .A(_10472_),
    .B(_10739_));
 sg13g2_o21ai_1 _18175_ (.B1(\rbzero.spi_registers.buf_texadd3[11] ),
    .Y(_10746_),
    .A1(net575),
    .A2(net530));
 sg13g2_a21oi_1 _18176_ (.A1(_10745_),
    .A2(_10746_),
    .Y(_00830_),
    .B1(_10723_));
 sg13g2_nand2_1 _18177_ (.Y(_10747_),
    .A(_10475_),
    .B(_10739_));
 sg13g2_o21ai_1 _18178_ (.B1(\rbzero.spi_registers.buf_texadd3[12] ),
    .Y(_10748_),
    .A1(net575),
    .A2(net530));
 sg13g2_buf_1 _18179_ (.A(_10722_),
    .X(_10749_));
 sg13g2_a21oi_1 _18180_ (.A1(_10747_),
    .A2(_10748_),
    .Y(_00831_),
    .B1(net654));
 sg13g2_nand2_1 _18181_ (.Y(_10750_),
    .A(_10479_),
    .B(net484));
 sg13g2_o21ai_1 _18182_ (.B1(\rbzero.spi_registers.buf_texadd3[13] ),
    .Y(_10751_),
    .A1(_10741_),
    .A2(net530));
 sg13g2_a21oi_1 _18183_ (.A1(_10750_),
    .A2(_10751_),
    .Y(_00832_),
    .B1(_10749_));
 sg13g2_nand2_1 _18184_ (.Y(_10752_),
    .A(_10482_),
    .B(net484));
 sg13g2_o21ai_1 _18185_ (.B1(\rbzero.spi_registers.buf_texadd3[14] ),
    .Y(_10753_),
    .A1(_10741_),
    .A2(net530));
 sg13g2_a21oi_1 _18186_ (.A1(_10752_),
    .A2(_10753_),
    .Y(_00833_),
    .B1(net654));
 sg13g2_nand2_1 _18187_ (.Y(_10754_),
    .A(_10566_),
    .B(net484));
 sg13g2_buf_1 _18188_ (.A(_10617_),
    .X(_10755_));
 sg13g2_o21ai_1 _18189_ (.B1(\rbzero.spi_registers.buf_texadd3[15] ),
    .Y(_10756_),
    .A1(net575),
    .A2(_10755_));
 sg13g2_a21oi_1 _18190_ (.A1(_10754_),
    .A2(_10756_),
    .Y(_00834_),
    .B1(_10749_));
 sg13g2_nand2_1 _18191_ (.Y(_10757_),
    .A(_10570_),
    .B(net484));
 sg13g2_o21ai_1 _18192_ (.B1(\rbzero.spi_registers.buf_texadd3[16] ),
    .Y(_10758_),
    .A1(net575),
    .A2(_10755_));
 sg13g2_a21oi_1 _18193_ (.A1(_10757_),
    .A2(_10758_),
    .Y(_00835_),
    .B1(net654));
 sg13g2_nand2_1 _18194_ (.Y(_10759_),
    .A(_10573_),
    .B(net484));
 sg13g2_o21ai_1 _18195_ (.B1(\rbzero.spi_registers.buf_texadd3[17] ),
    .Y(_10760_),
    .A1(net575),
    .A2(net529));
 sg13g2_a21oi_1 _18196_ (.A1(_10759_),
    .A2(_10760_),
    .Y(_00836_),
    .B1(net654));
 sg13g2_nand2_1 _18197_ (.Y(_10761_),
    .A(_10576_),
    .B(net484));
 sg13g2_o21ai_1 _18198_ (.B1(\rbzero.spi_registers.buf_texadd3[18] ),
    .Y(_10762_),
    .A1(net575),
    .A2(net529));
 sg13g2_a21oi_1 _18199_ (.A1(_10761_),
    .A2(_10762_),
    .Y(_00837_),
    .B1(net654));
 sg13g2_buf_1 _18200_ (.A(_10738_),
    .X(_10763_));
 sg13g2_nand2_1 _18201_ (.Y(_10764_),
    .A(_10579_),
    .B(net483));
 sg13g2_buf_1 _18202_ (.A(net668),
    .X(_10765_));
 sg13g2_o21ai_1 _18203_ (.B1(\rbzero.spi_registers.buf_texadd3[19] ),
    .Y(_10766_),
    .A1(net574),
    .A2(net529));
 sg13g2_a21oi_1 _18204_ (.A1(_10764_),
    .A2(_10766_),
    .Y(_00838_),
    .B1(net654));
 sg13g2_nand2_1 _18205_ (.Y(_10767_),
    .A(net747),
    .B(net483));
 sg13g2_o21ai_1 _18206_ (.B1(\rbzero.spi_registers.buf_texadd3[1] ),
    .Y(_10768_),
    .A1(net574),
    .A2(net529));
 sg13g2_a21oi_1 _18207_ (.A1(_10767_),
    .A2(_10768_),
    .Y(_00839_),
    .B1(net654));
 sg13g2_nand2_1 _18208_ (.Y(_10769_),
    .A(_10586_),
    .B(net483));
 sg13g2_o21ai_1 _18209_ (.B1(\rbzero.spi_registers.buf_texadd3[20] ),
    .Y(_10770_),
    .A1(net574),
    .A2(net529));
 sg13g2_a21oi_1 _18210_ (.A1(_10769_),
    .A2(_10770_),
    .Y(_00840_),
    .B1(net654));
 sg13g2_nand2_1 _18211_ (.Y(_10771_),
    .A(_10589_),
    .B(net483));
 sg13g2_o21ai_1 _18212_ (.B1(\rbzero.spi_registers.buf_texadd3[21] ),
    .Y(_10772_),
    .A1(net574),
    .A2(net529));
 sg13g2_buf_1 _18213_ (.A(_10722_),
    .X(_10773_));
 sg13g2_a21oi_1 _18214_ (.A1(_10771_),
    .A2(_10772_),
    .Y(_00841_),
    .B1(net653));
 sg13g2_nand2_1 _18215_ (.Y(_10774_),
    .A(_10592_),
    .B(net483));
 sg13g2_o21ai_1 _18216_ (.B1(\rbzero.spi_registers.buf_texadd3[22] ),
    .Y(_10775_),
    .A1(net574),
    .A2(net529));
 sg13g2_a21oi_1 _18217_ (.A1(_10774_),
    .A2(_10775_),
    .Y(_00842_),
    .B1(net653));
 sg13g2_nand2_1 _18218_ (.Y(_10776_),
    .A(_10595_),
    .B(net483));
 sg13g2_o21ai_1 _18219_ (.B1(\rbzero.spi_registers.buf_texadd3[23] ),
    .Y(_10777_),
    .A1(net574),
    .A2(net529));
 sg13g2_a21oi_1 _18220_ (.A1(_10776_),
    .A2(_10777_),
    .Y(_00843_),
    .B1(net653));
 sg13g2_nand2_1 _18221_ (.Y(_10778_),
    .A(net746),
    .B(net483));
 sg13g2_o21ai_1 _18222_ (.B1(\rbzero.spi_registers.buf_texadd3[2] ),
    .Y(_10779_),
    .A1(net574),
    .A2(net531));
 sg13g2_a21oi_1 _18223_ (.A1(_10778_),
    .A2(_10779_),
    .Y(_00844_),
    .B1(net653));
 sg13g2_nand2_1 _18224_ (.Y(_10780_),
    .A(net745),
    .B(net483));
 sg13g2_o21ai_1 _18225_ (.B1(\rbzero.spi_registers.buf_texadd3[3] ),
    .Y(_10781_),
    .A1(net574),
    .A2(net531));
 sg13g2_a21oi_1 _18226_ (.A1(_10780_),
    .A2(_10781_),
    .Y(_00845_),
    .B1(net653));
 sg13g2_nand2_1 _18227_ (.Y(_10782_),
    .A(net744),
    .B(_10763_));
 sg13g2_o21ai_1 _18228_ (.B1(\rbzero.spi_registers.buf_texadd3[4] ),
    .Y(_10783_),
    .A1(_10765_),
    .A2(net531));
 sg13g2_a21oi_1 _18229_ (.A1(_10782_),
    .A2(_10783_),
    .Y(_00846_),
    .B1(net653));
 sg13g2_nand2_1 _18230_ (.Y(_10784_),
    .A(net814),
    .B(_10763_));
 sg13g2_o21ai_1 _18231_ (.B1(\rbzero.spi_registers.buf_texadd3[5] ),
    .Y(_10785_),
    .A1(_10765_),
    .A2(net531));
 sg13g2_a21oi_1 _18232_ (.A1(_10784_),
    .A2(_10785_),
    .Y(_00847_),
    .B1(net653));
 sg13g2_nand2_1 _18233_ (.Y(_10786_),
    .A(_10494_),
    .B(_10738_));
 sg13g2_o21ai_1 _18234_ (.B1(\rbzero.spi_registers.buf_texadd3[6] ),
    .Y(_10787_),
    .A1(net668),
    .A2(net531));
 sg13g2_a21oi_1 _18235_ (.A1(_10786_),
    .A2(_10787_),
    .Y(_00848_),
    .B1(_10773_));
 sg13g2_nand2_1 _18236_ (.Y(_10788_),
    .A(_10497_),
    .B(_10738_));
 sg13g2_o21ai_1 _18237_ (.B1(\rbzero.spi_registers.buf_texadd3[7] ),
    .Y(_10789_),
    .A1(_10446_),
    .A2(net531));
 sg13g2_a21oi_1 _18238_ (.A1(_10788_),
    .A2(_10789_),
    .Y(_00849_),
    .B1(_10773_));
 sg13g2_nand2_1 _18239_ (.Y(_10790_),
    .A(_10501_),
    .B(_10738_));
 sg13g2_o21ai_1 _18240_ (.B1(\rbzero.spi_registers.buf_texadd3[8] ),
    .Y(_10791_),
    .A1(net668),
    .A2(_10680_));
 sg13g2_a21oi_1 _18241_ (.A1(_10790_),
    .A2(_10791_),
    .Y(_00850_),
    .B1(net653));
 sg13g2_nand2_1 _18242_ (.Y(_10792_),
    .A(_10518_),
    .B(_10738_));
 sg13g2_o21ai_1 _18243_ (.B1(\rbzero.spi_registers.buf_texadd3[9] ),
    .Y(_10793_),
    .A1(_10446_),
    .A2(_10680_));
 sg13g2_buf_1 _18244_ (.A(_10722_),
    .X(_10794_));
 sg13g2_a21oi_1 _18245_ (.A1(_10792_),
    .A2(_10793_),
    .Y(_00851_),
    .B1(net652));
 sg13g2_nor2_1 _18246_ (.A(_10416_),
    .B(_10600_),
    .Y(_10795_));
 sg13g2_nand2_1 _18247_ (.Y(_10796_),
    .A(net748),
    .B(_10795_));
 sg13g2_o21ai_1 _18248_ (.B1(\rbzero.spi_registers.buf_vinf ),
    .Y(_10797_),
    .A1(_10416_),
    .A2(_10600_));
 sg13g2_a21oi_1 _18249_ (.A1(_10796_),
    .A2(_10797_),
    .Y(_00852_),
    .B1(net652));
 sg13g2_nor3_1 _18250_ (.A(_09461_),
    .B(_09476_),
    .C(_10465_),
    .Y(_10798_));
 sg13g2_buf_1 _18251_ (.A(_10798_),
    .X(_10799_));
 sg13g2_nand2_1 _18252_ (.Y(_10800_),
    .A(_10413_),
    .B(net528));
 sg13g2_nand2b_1 _18253_ (.Y(_10801_),
    .B(\rbzero.spi_registers.buf_vshift[0] ),
    .A_N(net528));
 sg13g2_a21oi_1 _18254_ (.A1(_10800_),
    .A2(_10801_),
    .Y(_00853_),
    .B1(net652));
 sg13g2_nand2_1 _18255_ (.Y(_10802_),
    .A(_10427_),
    .B(net528));
 sg13g2_nand2b_1 _18256_ (.Y(_10803_),
    .B(\rbzero.spi_registers.buf_vshift[1] ),
    .A_N(net528));
 sg13g2_a21oi_1 _18257_ (.A1(_10802_),
    .A2(_10803_),
    .Y(_00854_),
    .B1(net652));
 sg13g2_nand2_1 _18258_ (.Y(_10804_),
    .A(_10430_),
    .B(net528));
 sg13g2_nand2b_1 _18259_ (.Y(_10805_),
    .B(\rbzero.spi_registers.buf_vshift[2] ),
    .A_N(net528));
 sg13g2_a21oi_1 _18260_ (.A1(_10804_),
    .A2(_10805_),
    .Y(_00855_),
    .B1(net652));
 sg13g2_nand2_1 _18261_ (.Y(_10806_),
    .A(_10436_),
    .B(net528));
 sg13g2_nand2b_1 _18262_ (.Y(_10807_),
    .B(\rbzero.spi_registers.buf_vshift[3] ),
    .A_N(net528));
 sg13g2_a21oi_1 _18263_ (.A1(_10806_),
    .A2(_10807_),
    .Y(_00856_),
    .B1(net652));
 sg13g2_nand2_1 _18264_ (.Y(_10808_),
    .A(_10439_),
    .B(_10799_));
 sg13g2_nand2b_1 _18265_ (.Y(_10809_),
    .B(\rbzero.spi_registers.buf_vshift[4] ),
    .A_N(_10798_));
 sg13g2_a21oi_1 _18266_ (.A1(_10808_),
    .A2(_10809_),
    .Y(_00857_),
    .B1(net652));
 sg13g2_nand2_1 _18267_ (.Y(_10810_),
    .A(_10443_),
    .B(_10799_));
 sg13g2_nand2b_1 _18268_ (.Y(_10811_),
    .B(\rbzero.spi_registers.buf_vshift[5] ),
    .A_N(_10798_));
 sg13g2_a21oi_1 _18269_ (.A1(_10810_),
    .A2(_10811_),
    .Y(_00858_),
    .B1(net652));
 sg13g2_buf_1 _18270_ (.A(net451),
    .X(_10812_));
 sg13g2_buf_1 _18271_ (.A(net413),
    .X(_10813_));
 sg13g2_nand2_1 _18272_ (.Y(_10814_),
    .A(\rbzero.spi_registers.buf_floor[0] ),
    .B(net387));
 sg13g2_buf_1 _18273_ (.A(_09416_),
    .X(_10815_));
 sg13g2_buf_1 _18274_ (.A(net412),
    .X(_10816_));
 sg13g2_nand2_1 _18275_ (.Y(_10817_),
    .A(\rbzero.color_floor[0] ),
    .B(net386));
 sg13g2_a21oi_1 _18276_ (.A1(_10814_),
    .A2(_10817_),
    .Y(_00859_),
    .B1(_10794_));
 sg13g2_nand2_1 _18277_ (.Y(_10818_),
    .A(\rbzero.color_floor[1] ),
    .B(net386));
 sg13g2_nand2_1 _18278_ (.Y(_10819_),
    .A(\rbzero.spi_registers.buf_floor[1] ),
    .B(net387));
 sg13g2_nand3_1 _18279_ (.B(_10818_),
    .C(_10819_),
    .A(net751),
    .Y(_00860_));
 sg13g2_nand2_1 _18280_ (.Y(_10820_),
    .A(\rbzero.spi_registers.buf_floor[2] ),
    .B(net387));
 sg13g2_nand2_1 _18281_ (.Y(_10821_),
    .A(\rbzero.color_floor[2] ),
    .B(_10816_));
 sg13g2_a21oi_1 _18282_ (.A1(_10820_),
    .A2(_10821_),
    .Y(_00861_),
    .B1(_10794_));
 sg13g2_nand2_1 _18283_ (.Y(_10822_),
    .A(\rbzero.spi_registers.buf_floor[3] ),
    .B(net387));
 sg13g2_nand2_1 _18284_ (.Y(_10823_),
    .A(\rbzero.color_floor[3] ),
    .B(net386));
 sg13g2_nand3_1 _18285_ (.B(_10822_),
    .C(_10823_),
    .A(net751),
    .Y(_00862_));
 sg13g2_nand2_1 _18286_ (.Y(_10824_),
    .A(\rbzero.spi_registers.buf_floor[4] ),
    .B(_10813_));
 sg13g2_nand2_1 _18287_ (.Y(_10825_),
    .A(\rbzero.color_floor[4] ),
    .B(net386));
 sg13g2_buf_1 _18288_ (.A(_10722_),
    .X(_10826_));
 sg13g2_a21oi_1 _18289_ (.A1(_10824_),
    .A2(_10825_),
    .Y(_00863_),
    .B1(net651));
 sg13g2_nand2_1 _18290_ (.Y(_10827_),
    .A(\rbzero.spi_registers.buf_floor[5] ),
    .B(net387));
 sg13g2_nand2_1 _18291_ (.Y(_10828_),
    .A(\rbzero.color_floor[5] ),
    .B(net386));
 sg13g2_nand3_1 _18292_ (.B(_10827_),
    .C(_10828_),
    .A(net751),
    .Y(_00864_));
 sg13g2_nand2_1 _18293_ (.Y(_10829_),
    .A(\rbzero.spi_registers.buf_leak[0] ),
    .B(_10813_));
 sg13g2_nand2_1 _18294_ (.Y(_10830_),
    .A(\rbzero.floor_leak[0] ),
    .B(_10816_));
 sg13g2_a21oi_1 _18295_ (.A1(_10829_),
    .A2(_10830_),
    .Y(_00865_),
    .B1(net651));
 sg13g2_buf_1 _18296_ (.A(net413),
    .X(_10831_));
 sg13g2_nand2_1 _18297_ (.Y(_10832_),
    .A(\rbzero.spi_registers.buf_leak[1] ),
    .B(net385));
 sg13g2_buf_1 _18298_ (.A(net412),
    .X(_10833_));
 sg13g2_nand2_1 _18299_ (.Y(_10834_),
    .A(\rbzero.floor_leak[1] ),
    .B(net384));
 sg13g2_a21oi_1 _18300_ (.A1(_10832_),
    .A2(_10834_),
    .Y(_00866_),
    .B1(net651));
 sg13g2_nand2_1 _18301_ (.Y(_10835_),
    .A(\rbzero.spi_registers.buf_leak[2] ),
    .B(net385));
 sg13g2_nand2_1 _18302_ (.Y(_10836_),
    .A(\rbzero.floor_leak[2] ),
    .B(net384));
 sg13g2_a21oi_1 _18303_ (.A1(_10835_),
    .A2(_10836_),
    .Y(_00867_),
    .B1(net651));
 sg13g2_nand2_1 _18304_ (.Y(_10837_),
    .A(\rbzero.spi_registers.buf_leak[3] ),
    .B(net385));
 sg13g2_nand2_1 _18305_ (.Y(_10838_),
    .A(\rbzero.floor_leak[3] ),
    .B(net384));
 sg13g2_a21oi_1 _18306_ (.A1(_10837_),
    .A2(_10838_),
    .Y(_00868_),
    .B1(_10826_));
 sg13g2_nand2_1 _18307_ (.Y(_10839_),
    .A(\rbzero.spi_registers.buf_leak[4] ),
    .B(_10831_));
 sg13g2_nand2_1 _18308_ (.Y(_10840_),
    .A(\rbzero.floor_leak[4] ),
    .B(_10833_));
 sg13g2_a21oi_1 _18309_ (.A1(_10839_),
    .A2(_10840_),
    .Y(_00869_),
    .B1(net651));
 sg13g2_nand2_1 _18310_ (.Y(_10841_),
    .A(\rbzero.spi_registers.buf_leak[5] ),
    .B(_10831_));
 sg13g2_nand2_1 _18311_ (.Y(_10842_),
    .A(\rbzero.floor_leak[5] ),
    .B(_10833_));
 sg13g2_a21oi_1 _18312_ (.A1(_10841_),
    .A2(_10842_),
    .Y(_00870_),
    .B1(_10826_));
 sg13g2_nand2_1 _18313_ (.Y(_10843_),
    .A(\rbzero.spi_registers.buf_mapdx[0] ),
    .B(net385));
 sg13g2_nand2_1 _18314_ (.Y(_10844_),
    .A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(net384));
 sg13g2_a21oi_1 _18315_ (.A1(_10843_),
    .A2(_10844_),
    .Y(_00871_),
    .B1(net651));
 sg13g2_nand2_1 _18316_ (.Y(_10845_),
    .A(\rbzero.spi_registers.buf_mapdx[1] ),
    .B(net385));
 sg13g2_nand2_1 _18317_ (.Y(_10846_),
    .A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(net384));
 sg13g2_a21oi_1 _18318_ (.A1(_10845_),
    .A2(_10846_),
    .Y(_00872_),
    .B1(net651));
 sg13g2_nand2_1 _18319_ (.Y(_10847_),
    .A(\rbzero.spi_registers.buf_mapdx[2] ),
    .B(net385));
 sg13g2_nand2_1 _18320_ (.Y(_10848_),
    .A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(net384));
 sg13g2_a21oi_1 _18321_ (.A1(_10847_),
    .A2(_10848_),
    .Y(_00873_),
    .B1(net651));
 sg13g2_nand2_1 _18322_ (.Y(_10849_),
    .A(\rbzero.spi_registers.buf_mapdx[3] ),
    .B(net385));
 sg13g2_nand2_1 _18323_ (.Y(_10850_),
    .A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(net384));
 sg13g2_buf_1 _18324_ (.A(_10722_),
    .X(_10851_));
 sg13g2_a21oi_1 _18325_ (.A1(_10849_),
    .A2(_10850_),
    .Y(_00874_),
    .B1(_10851_));
 sg13g2_nand2_1 _18326_ (.Y(_10852_),
    .A(\rbzero.spi_registers.buf_mapdx[4] ),
    .B(net385));
 sg13g2_nand2_1 _18327_ (.Y(_10853_),
    .A(\rbzero.map_overlay.i_mapdx[4] ),
    .B(net384));
 sg13g2_a21oi_1 _18328_ (.A1(_10852_),
    .A2(_10853_),
    .Y(_00875_),
    .B1(net650));
 sg13g2_buf_1 _18329_ (.A(net413),
    .X(_10854_));
 sg13g2_nand2_1 _18330_ (.Y(_10855_),
    .A(\rbzero.spi_registers.buf_mapdxw[0] ),
    .B(net383));
 sg13g2_buf_1 _18331_ (.A(net412),
    .X(_10856_));
 sg13g2_nand2_1 _18332_ (.Y(_10857_),
    .A(\rbzero.mapdxw[0] ),
    .B(net382));
 sg13g2_a21oi_1 _18333_ (.A1(_10855_),
    .A2(_10857_),
    .Y(_00876_),
    .B1(net650));
 sg13g2_nand2_1 _18334_ (.Y(_10858_),
    .A(\rbzero.spi_registers.buf_mapdxw[1] ),
    .B(_10854_));
 sg13g2_nand2_1 _18335_ (.Y(_10859_),
    .A(\rbzero.mapdxw[1] ),
    .B(net382));
 sg13g2_a21oi_1 _18336_ (.A1(_10858_),
    .A2(_10859_),
    .Y(_00877_),
    .B1(_10851_));
 sg13g2_nand2_1 _18337_ (.Y(_10860_),
    .A(\rbzero.spi_registers.buf_mapdy[0] ),
    .B(net383));
 sg13g2_nand2_1 _18338_ (.Y(_10861_),
    .A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(net382));
 sg13g2_a21oi_1 _18339_ (.A1(_10860_),
    .A2(_10861_),
    .Y(_00878_),
    .B1(net650));
 sg13g2_nand2_1 _18340_ (.Y(_10862_),
    .A(\rbzero.spi_registers.buf_mapdy[1] ),
    .B(net383));
 sg13g2_nand2_1 _18341_ (.Y(_10863_),
    .A(\rbzero.map_overlay.i_mapdy[1] ),
    .B(net382));
 sg13g2_a21oi_1 _18342_ (.A1(_10862_),
    .A2(_10863_),
    .Y(_00879_),
    .B1(net650));
 sg13g2_nand2_1 _18343_ (.Y(_10864_),
    .A(\rbzero.spi_registers.buf_mapdy[2] ),
    .B(net383));
 sg13g2_nand2_1 _18344_ (.Y(_10865_),
    .A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(net382));
 sg13g2_a21oi_1 _18345_ (.A1(_10864_),
    .A2(_10865_),
    .Y(_00880_),
    .B1(net650));
 sg13g2_nand2_1 _18346_ (.Y(_10866_),
    .A(\rbzero.spi_registers.buf_mapdy[3] ),
    .B(net383));
 sg13g2_nand2_1 _18347_ (.Y(_10867_),
    .A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(net382));
 sg13g2_a21oi_1 _18348_ (.A1(_10866_),
    .A2(_10867_),
    .Y(_00881_),
    .B1(net650));
 sg13g2_nand2_1 _18349_ (.Y(_10868_),
    .A(\rbzero.spi_registers.buf_mapdy[4] ),
    .B(net383));
 sg13g2_nand2_1 _18350_ (.Y(_10869_),
    .A(\rbzero.map_overlay.i_mapdy[4] ),
    .B(_10856_));
 sg13g2_a21oi_1 _18351_ (.A1(_10868_),
    .A2(_10869_),
    .Y(_00882_),
    .B1(net650));
 sg13g2_nand2_1 _18352_ (.Y(_10870_),
    .A(\rbzero.spi_registers.buf_mapdyw[0] ),
    .B(net383));
 sg13g2_nand2_1 _18353_ (.Y(_10871_),
    .A(\rbzero.mapdyw[0] ),
    .B(_10856_));
 sg13g2_a21oi_1 _18354_ (.A1(_10870_),
    .A2(_10871_),
    .Y(_00883_),
    .B1(net650));
 sg13g2_nand2_1 _18355_ (.Y(_10872_),
    .A(\rbzero.spi_registers.buf_mapdyw[1] ),
    .B(net383));
 sg13g2_nand2_1 _18356_ (.Y(_10873_),
    .A(\rbzero.mapdyw[1] ),
    .B(net382));
 sg13g2_buf_1 _18357_ (.A(_10722_),
    .X(_10874_));
 sg13g2_a21oi_1 _18358_ (.A1(_10872_),
    .A2(_10873_),
    .Y(_00884_),
    .B1(_10874_));
 sg13g2_and2_1 _18359_ (.A(net750),
    .B(net8),
    .X(_00885_));
 sg13g2_and2_1 _18360_ (.A(net750),
    .B(\rbzero.spi_registers.mosi_buffer[0] ),
    .X(_00886_));
 sg13g2_nand2_1 _18361_ (.Y(_10875_),
    .A(\rbzero.spi_registers.buf_otherx[0] ),
    .B(_10854_));
 sg13g2_nand2_1 _18362_ (.Y(_10876_),
    .A(\rbzero.map_overlay.i_otherx[0] ),
    .B(net382));
 sg13g2_a21oi_1 _18363_ (.A1(_10875_),
    .A2(_10876_),
    .Y(_00887_),
    .B1(_10874_));
 sg13g2_buf_1 _18364_ (.A(net413),
    .X(_10877_));
 sg13g2_nand2_1 _18365_ (.Y(_10878_),
    .A(\rbzero.spi_registers.buf_otherx[1] ),
    .B(net381));
 sg13g2_buf_1 _18366_ (.A(net412),
    .X(_10879_));
 sg13g2_nand2_1 _18367_ (.Y(_10880_),
    .A(\rbzero.map_overlay.i_otherx[1] ),
    .B(net380));
 sg13g2_a21oi_1 _18368_ (.A1(_10878_),
    .A2(_10880_),
    .Y(_00888_),
    .B1(net649));
 sg13g2_nand2_1 _18369_ (.Y(_10881_),
    .A(\rbzero.spi_registers.buf_otherx[2] ),
    .B(_10877_));
 sg13g2_nand2_1 _18370_ (.Y(_10882_),
    .A(\rbzero.map_overlay.i_otherx[2] ),
    .B(net380));
 sg13g2_a21oi_1 _18371_ (.A1(_10881_),
    .A2(_10882_),
    .Y(_00889_),
    .B1(net649));
 sg13g2_nand2_1 _18372_ (.Y(_10883_),
    .A(\rbzero.spi_registers.buf_otherx[3] ),
    .B(net381));
 sg13g2_nand2_1 _18373_ (.Y(_10884_),
    .A(\rbzero.map_overlay.i_otherx[3] ),
    .B(net380));
 sg13g2_a21oi_1 _18374_ (.A1(_10883_),
    .A2(_10884_),
    .Y(_00890_),
    .B1(net649));
 sg13g2_nand2_1 _18375_ (.Y(_10885_),
    .A(\rbzero.spi_registers.buf_otherx[4] ),
    .B(net381));
 sg13g2_nand2_1 _18376_ (.Y(_10886_),
    .A(\rbzero.map_overlay.i_otherx[4] ),
    .B(net380));
 sg13g2_a21oi_1 _18377_ (.A1(_10885_),
    .A2(_10886_),
    .Y(_00891_),
    .B1(net649));
 sg13g2_nand2_1 _18378_ (.Y(_10887_),
    .A(\rbzero.spi_registers.buf_othery[0] ),
    .B(net381));
 sg13g2_nand2_1 _18379_ (.Y(_10888_),
    .A(\rbzero.map_overlay.i_othery[0] ),
    .B(net380));
 sg13g2_a21oi_1 _18380_ (.A1(_10887_),
    .A2(_10888_),
    .Y(_00892_),
    .B1(net649));
 sg13g2_nand2_1 _18381_ (.Y(_10889_),
    .A(\rbzero.spi_registers.buf_othery[1] ),
    .B(_10877_));
 sg13g2_nand2_1 _18382_ (.Y(_10890_),
    .A(\rbzero.map_overlay.i_othery[1] ),
    .B(_10879_));
 sg13g2_a21oi_1 _18383_ (.A1(_10889_),
    .A2(_10890_),
    .Y(_00893_),
    .B1(net649));
 sg13g2_nand2_1 _18384_ (.Y(_10891_),
    .A(\rbzero.spi_registers.buf_othery[2] ),
    .B(net381));
 sg13g2_nand2_1 _18385_ (.Y(_10892_),
    .A(\rbzero.map_overlay.i_othery[2] ),
    .B(_10879_));
 sg13g2_a21oi_1 _18386_ (.A1(_10891_),
    .A2(_10892_),
    .Y(_00894_),
    .B1(net649));
 sg13g2_nand2_1 _18387_ (.Y(_10893_),
    .A(\rbzero.spi_registers.buf_othery[3] ),
    .B(net381));
 sg13g2_nand2_1 _18388_ (.Y(_10894_),
    .A(\rbzero.map_overlay.i_othery[3] ),
    .B(net380));
 sg13g2_a21oi_1 _18389_ (.A1(_10893_),
    .A2(_10894_),
    .Y(_00895_),
    .B1(net649));
 sg13g2_nand2_1 _18390_ (.Y(_10895_),
    .A(\rbzero.spi_registers.buf_othery[4] ),
    .B(net381));
 sg13g2_nand2_1 _18391_ (.Y(_10896_),
    .A(\rbzero.map_overlay.i_othery[4] ),
    .B(net380));
 sg13g2_buf_1 _18392_ (.A(_08638_),
    .X(_10897_));
 sg13g2_buf_1 _18393_ (.A(_10897_),
    .X(_10898_));
 sg13g2_a21oi_1 _18394_ (.A1(_10895_),
    .A2(_10896_),
    .Y(_00896_),
    .B1(net648));
 sg13g2_and2_1 _18395_ (.A(net750),
    .B(net7),
    .X(_00897_));
 sg13g2_and2_1 _18396_ (.A(net750),
    .B(\rbzero.spi_registers.sclk_buffer[0] ),
    .X(_00898_));
 sg13g2_and2_1 _18397_ (.A(net750),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(_00899_));
 sg13g2_nand2_1 _18398_ (.Y(_10899_),
    .A(\rbzero.spi_registers.buf_sky[0] ),
    .B(net387));
 sg13g2_nand2_1 _18399_ (.Y(_10900_),
    .A(\rbzero.color_sky[0] ),
    .B(net386));
 sg13g2_nand3_1 _18400_ (.B(_10899_),
    .C(_10900_),
    .A(net751),
    .Y(_00900_));
 sg13g2_nand2_1 _18401_ (.Y(_10901_),
    .A(\rbzero.spi_registers.buf_sky[1] ),
    .B(net381));
 sg13g2_nand2_1 _18402_ (.Y(_10902_),
    .A(\rbzero.color_sky[1] ),
    .B(net380));
 sg13g2_a21oi_1 _18403_ (.A1(_10901_),
    .A2(_10902_),
    .Y(_00901_),
    .B1(net648));
 sg13g2_nand2_1 _18404_ (.Y(_10903_),
    .A(\rbzero.spi_registers.buf_sky[2] ),
    .B(net387));
 sg13g2_nand2_1 _18405_ (.Y(_10904_),
    .A(\rbzero.color_sky[2] ),
    .B(net386));
 sg13g2_nand3_1 _18406_ (.B(_10903_),
    .C(_10904_),
    .A(net751),
    .Y(_00902_));
 sg13g2_buf_1 _18407_ (.A(net413),
    .X(_10905_));
 sg13g2_nand2_1 _18408_ (.Y(_10906_),
    .A(\rbzero.spi_registers.buf_sky[3] ),
    .B(net379));
 sg13g2_buf_1 _18409_ (.A(net412),
    .X(_10907_));
 sg13g2_nand2_1 _18410_ (.Y(_10908_),
    .A(\rbzero.color_sky[3] ),
    .B(net378));
 sg13g2_a21oi_1 _18411_ (.A1(_10906_),
    .A2(_10908_),
    .Y(_00903_),
    .B1(_10898_));
 sg13g2_nand2_1 _18412_ (.Y(_10909_),
    .A(\rbzero.spi_registers.buf_sky[4] ),
    .B(net387));
 sg13g2_nand2_1 _18413_ (.Y(_10910_),
    .A(\rbzero.color_sky[4] ),
    .B(net386));
 sg13g2_nand3_1 _18414_ (.B(_10909_),
    .C(_10910_),
    .A(net751),
    .Y(_00904_));
 sg13g2_nand2_1 _18415_ (.Y(_10911_),
    .A(\rbzero.spi_registers.buf_sky[5] ),
    .B(_10905_));
 sg13g2_nand2_1 _18416_ (.Y(_10912_),
    .A(\rbzero.color_sky[5] ),
    .B(_10907_));
 sg13g2_a21oi_1 _18417_ (.A1(_10911_),
    .A2(_10912_),
    .Y(_00905_),
    .B1(net648));
 sg13g2_buf_1 _18418_ (.A(_09424_),
    .X(_10913_));
 sg13g2_or3_1 _18419_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_09469_),
    .C(_09537_),
    .X(_10914_));
 sg13g2_buf_2 _18420_ (.A(_10914_),
    .X(_10915_));
 sg13g2_buf_1 _18421_ (.A(_10915_),
    .X(_10916_));
 sg13g2_mux2_1 _18422_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(_10413_),
    .S(_10916_),
    .X(_10917_));
 sg13g2_and2_1 _18423_ (.A(_10913_),
    .B(_10917_),
    .X(_00906_));
 sg13g2_mux2_1 _18424_ (.A0(_10518_),
    .A1(_10463_),
    .S(net527),
    .X(_10918_));
 sg13g2_and2_1 _18425_ (.A(net743),
    .B(_10918_),
    .X(_00907_));
 sg13g2_mux2_1 _18426_ (.A0(_10463_),
    .A1(_10472_),
    .S(net527),
    .X(_10919_));
 sg13g2_and2_1 _18427_ (.A(net743),
    .B(_10919_),
    .X(_00908_));
 sg13g2_mux2_1 _18428_ (.A0(_10472_),
    .A1(_10475_),
    .S(_10916_),
    .X(_10920_));
 sg13g2_and2_1 _18429_ (.A(net743),
    .B(_10920_),
    .X(_00909_));
 sg13g2_mux2_1 _18430_ (.A0(_10475_),
    .A1(_10479_),
    .S(net527),
    .X(_10921_));
 sg13g2_and2_1 _18431_ (.A(_10913_),
    .B(_10921_),
    .X(_00910_));
 sg13g2_mux2_1 _18432_ (.A0(_10479_),
    .A1(_10482_),
    .S(net527),
    .X(_10922_));
 sg13g2_and2_1 _18433_ (.A(net743),
    .B(_10922_),
    .X(_00911_));
 sg13g2_mux2_1 _18434_ (.A0(_10482_),
    .A1(_10566_),
    .S(net527),
    .X(_10923_));
 sg13g2_and2_1 _18435_ (.A(net743),
    .B(_10923_),
    .X(_00912_));
 sg13g2_mux2_1 _18436_ (.A0(_10566_),
    .A1(_10570_),
    .S(net527),
    .X(_10924_));
 sg13g2_and2_1 _18437_ (.A(net743),
    .B(_10924_),
    .X(_00913_));
 sg13g2_mux2_1 _18438_ (.A0(_10570_),
    .A1(_10573_),
    .S(net527),
    .X(_10925_));
 sg13g2_and2_1 _18439_ (.A(net743),
    .B(_10925_),
    .X(_00914_));
 sg13g2_mux2_1 _18440_ (.A0(_10573_),
    .A1(_10576_),
    .S(net527),
    .X(_10926_));
 sg13g2_and2_1 _18441_ (.A(net743),
    .B(_10926_),
    .X(_00915_));
 sg13g2_buf_1 _18442_ (.A(_09424_),
    .X(_10927_));
 sg13g2_buf_1 _18443_ (.A(_10915_),
    .X(_10928_));
 sg13g2_mux2_1 _18444_ (.A0(_10576_),
    .A1(_10579_),
    .S(net526),
    .X(_10929_));
 sg13g2_and2_1 _18445_ (.A(net742),
    .B(_10929_),
    .X(_00916_));
 sg13g2_mux2_1 _18446_ (.A0(_10413_),
    .A1(_10426_),
    .S(net526),
    .X(_10930_));
 sg13g2_and2_1 _18447_ (.A(net742),
    .B(_10930_),
    .X(_00917_));
 sg13g2_mux2_1 _18448_ (.A0(_10579_),
    .A1(_10586_),
    .S(net526),
    .X(_10931_));
 sg13g2_and2_1 _18449_ (.A(net742),
    .B(_10931_),
    .X(_00918_));
 sg13g2_mux2_1 _18450_ (.A0(_10586_),
    .A1(_10589_),
    .S(net526),
    .X(_10932_));
 sg13g2_and2_1 _18451_ (.A(net742),
    .B(_10932_),
    .X(_00919_));
 sg13g2_mux2_1 _18452_ (.A0(_10589_),
    .A1(_10592_),
    .S(net526),
    .X(_10933_));
 sg13g2_and2_1 _18453_ (.A(net742),
    .B(_10933_),
    .X(_00920_));
 sg13g2_mux2_1 _18454_ (.A0(_10592_),
    .A1(_10595_),
    .S(net526),
    .X(_10934_));
 sg13g2_and2_1 _18455_ (.A(net742),
    .B(_10934_),
    .X(_00921_));
 sg13g2_mux2_1 _18456_ (.A0(_10426_),
    .A1(_10429_),
    .S(net526),
    .X(_10935_));
 sg13g2_and2_1 _18457_ (.A(net742),
    .B(_10935_),
    .X(_00922_));
 sg13g2_mux2_1 _18458_ (.A0(_10429_),
    .A1(_10435_),
    .S(net526),
    .X(_10936_));
 sg13g2_and2_1 _18459_ (.A(net742),
    .B(_10936_),
    .X(_00923_));
 sg13g2_mux2_1 _18460_ (.A0(_10435_),
    .A1(_10438_),
    .S(_10928_),
    .X(_10937_));
 sg13g2_and2_1 _18461_ (.A(_10927_),
    .B(_10937_),
    .X(_00924_));
 sg13g2_mux2_1 _18462_ (.A0(_10438_),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_10928_),
    .X(_10938_));
 sg13g2_and2_1 _18463_ (.A(_10927_),
    .B(_10938_),
    .X(_00925_));
 sg13g2_mux2_1 _18464_ (.A0(_10443_),
    .A1(_10494_),
    .S(_10915_),
    .X(_10939_));
 sg13g2_and2_1 _18465_ (.A(net758),
    .B(_10939_),
    .X(_00926_));
 sg13g2_mux2_1 _18466_ (.A0(_10494_),
    .A1(_10497_),
    .S(_10915_),
    .X(_10940_));
 sg13g2_and2_1 _18467_ (.A(net758),
    .B(_10940_),
    .X(_00927_));
 sg13g2_mux2_1 _18468_ (.A0(_10497_),
    .A1(_10501_),
    .S(_10915_),
    .X(_10941_));
 sg13g2_and2_1 _18469_ (.A(net758),
    .B(_10941_),
    .X(_00928_));
 sg13g2_mux2_1 _18470_ (.A0(_10501_),
    .A1(_10518_),
    .S(_10915_),
    .X(_10942_));
 sg13g2_and2_1 _18471_ (.A(net758),
    .B(_10942_),
    .X(_00929_));
 sg13g2_and2_1 _18472_ (.A(net758),
    .B(net9),
    .X(_00942_));
 sg13g2_and2_1 _18473_ (.A(net758),
    .B(\rbzero.spi_registers.ss_buffer[0] ),
    .X(_00943_));
 sg13g2_nand2_1 _18474_ (.Y(_10943_),
    .A(\rbzero.spi_registers.buf_texadd0[0] ),
    .B(net379));
 sg13g2_nand2_1 _18475_ (.Y(_10944_),
    .A(\rbzero.spi_registers.texadd0[0] ),
    .B(_10907_));
 sg13g2_a21oi_1 _18476_ (.A1(_10943_),
    .A2(_10944_),
    .Y(_00944_),
    .B1(net648));
 sg13g2_nand2_1 _18477_ (.Y(_10945_),
    .A(\rbzero.spi_registers.buf_texadd0[10] ),
    .B(net379));
 sg13g2_nand2_1 _18478_ (.Y(_10946_),
    .A(\rbzero.spi_registers.texadd0[10] ),
    .B(net378));
 sg13g2_a21oi_1 _18479_ (.A1(_10945_),
    .A2(_10946_),
    .Y(_00945_),
    .B1(net648));
 sg13g2_nand2_1 _18480_ (.Y(_10947_),
    .A(\rbzero.spi_registers.buf_texadd0[11] ),
    .B(net379));
 sg13g2_nand2_1 _18481_ (.Y(_10948_),
    .A(\rbzero.spi_registers.texadd0[11] ),
    .B(net378));
 sg13g2_a21oi_1 _18482_ (.A1(_10947_),
    .A2(_10948_),
    .Y(_00946_),
    .B1(_10898_));
 sg13g2_nand2_1 _18483_ (.Y(_10949_),
    .A(\rbzero.spi_registers.buf_texadd0[12] ),
    .B(net379));
 sg13g2_nand2_1 _18484_ (.Y(_10950_),
    .A(\rbzero.spi_registers.texadd0[12] ),
    .B(net378));
 sg13g2_a21oi_1 _18485_ (.A1(_10949_),
    .A2(_10950_),
    .Y(_00947_),
    .B1(net648));
 sg13g2_nand2_1 _18486_ (.Y(_10951_),
    .A(\rbzero.spi_registers.buf_texadd0[13] ),
    .B(_10905_));
 sg13g2_nand2_1 _18487_ (.Y(_10952_),
    .A(\rbzero.spi_registers.texadd0[13] ),
    .B(net378));
 sg13g2_a21oi_1 _18488_ (.A1(_10951_),
    .A2(_10952_),
    .Y(_00948_),
    .B1(net648));
 sg13g2_nand2_1 _18489_ (.Y(_10953_),
    .A(\rbzero.spi_registers.buf_texadd0[14] ),
    .B(net379));
 sg13g2_nand2_1 _18490_ (.Y(_10954_),
    .A(\rbzero.spi_registers.texadd0[14] ),
    .B(net378));
 sg13g2_a21oi_1 _18491_ (.A1(_10953_),
    .A2(_10954_),
    .Y(_00949_),
    .B1(net648));
 sg13g2_nand2_1 _18492_ (.Y(_10955_),
    .A(\rbzero.spi_registers.buf_texadd0[15] ),
    .B(net379));
 sg13g2_nand2_1 _18493_ (.Y(_10956_),
    .A(\rbzero.spi_registers.texadd0[15] ),
    .B(net378));
 sg13g2_buf_1 _18494_ (.A(_10897_),
    .X(_10957_));
 sg13g2_a21oi_1 _18495_ (.A1(_10955_),
    .A2(_10956_),
    .Y(_00950_),
    .B1(_10957_));
 sg13g2_nand2_1 _18496_ (.Y(_10958_),
    .A(\rbzero.spi_registers.buf_texadd0[16] ),
    .B(net379));
 sg13g2_nand2_1 _18497_ (.Y(_10959_),
    .A(\rbzero.spi_registers.texadd0[16] ),
    .B(net378));
 sg13g2_a21oi_1 _18498_ (.A1(_10958_),
    .A2(_10959_),
    .Y(_00951_),
    .B1(_10957_));
 sg13g2_buf_1 _18499_ (.A(net451),
    .X(_10960_));
 sg13g2_buf_1 _18500_ (.A(_10960_),
    .X(_10961_));
 sg13g2_nand2_1 _18501_ (.Y(_10962_),
    .A(\rbzero.spi_registers.buf_texadd0[17] ),
    .B(_10961_));
 sg13g2_buf_1 _18502_ (.A(_09416_),
    .X(_10963_));
 sg13g2_buf_1 _18503_ (.A(_10963_),
    .X(_10964_));
 sg13g2_nand2_1 _18504_ (.Y(_10965_),
    .A(\rbzero.spi_registers.texadd0[17] ),
    .B(_10964_));
 sg13g2_a21oi_1 _18505_ (.A1(_10962_),
    .A2(_10965_),
    .Y(_00952_),
    .B1(net647));
 sg13g2_nand2_1 _18506_ (.Y(_10966_),
    .A(\rbzero.spi_registers.buf_texadd0[18] ),
    .B(net377));
 sg13g2_nand2_1 _18507_ (.Y(_10967_),
    .A(\rbzero.spi_registers.texadd0[18] ),
    .B(net376));
 sg13g2_a21oi_1 _18508_ (.A1(_10966_),
    .A2(_10967_),
    .Y(_00953_),
    .B1(net647));
 sg13g2_nand2_1 _18509_ (.Y(_10968_),
    .A(\rbzero.spi_registers.buf_texadd0[19] ),
    .B(net377));
 sg13g2_nand2_1 _18510_ (.Y(_10969_),
    .A(\rbzero.spi_registers.texadd0[19] ),
    .B(net376));
 sg13g2_a21oi_1 _18511_ (.A1(_10968_),
    .A2(_10969_),
    .Y(_00954_),
    .B1(net647));
 sg13g2_nand2_1 _18512_ (.Y(_10970_),
    .A(\rbzero.spi_registers.buf_texadd0[1] ),
    .B(net377));
 sg13g2_nand2_1 _18513_ (.Y(_10971_),
    .A(\rbzero.spi_registers.texadd0[1] ),
    .B(net376));
 sg13g2_a21oi_1 _18514_ (.A1(_10970_),
    .A2(_10971_),
    .Y(_00955_),
    .B1(net647));
 sg13g2_nand2_1 _18515_ (.Y(_10972_),
    .A(\rbzero.spi_registers.buf_texadd0[20] ),
    .B(net377));
 sg13g2_nand2_1 _18516_ (.Y(_10973_),
    .A(\rbzero.spi_registers.texadd0[20] ),
    .B(net376));
 sg13g2_a21oi_1 _18517_ (.A1(_10972_),
    .A2(_10973_),
    .Y(_00956_),
    .B1(net647));
 sg13g2_nand2_1 _18518_ (.Y(_10974_),
    .A(\rbzero.spi_registers.buf_texadd0[21] ),
    .B(net377));
 sg13g2_nand2_1 _18519_ (.Y(_10975_),
    .A(\rbzero.spi_registers.texadd0[21] ),
    .B(net376));
 sg13g2_a21oi_1 _18520_ (.A1(_10974_),
    .A2(_10975_),
    .Y(_00957_),
    .B1(net647));
 sg13g2_nand2_1 _18521_ (.Y(_10976_),
    .A(\rbzero.spi_registers.buf_texadd0[22] ),
    .B(net377));
 sg13g2_nand2_1 _18522_ (.Y(_10977_),
    .A(\rbzero.spi_registers.texadd0[22] ),
    .B(net376));
 sg13g2_a21oi_1 _18523_ (.A1(_10976_),
    .A2(_10977_),
    .Y(_00958_),
    .B1(net647));
 sg13g2_nand2_1 _18524_ (.Y(_10978_),
    .A(\rbzero.spi_registers.buf_texadd0[23] ),
    .B(net377));
 sg13g2_nand2_1 _18525_ (.Y(_10979_),
    .A(\rbzero.spi_registers.texadd0[23] ),
    .B(net376));
 sg13g2_a21oi_1 _18526_ (.A1(_10978_),
    .A2(_10979_),
    .Y(_00959_),
    .B1(net647));
 sg13g2_nand2_1 _18527_ (.Y(_10980_),
    .A(\rbzero.spi_registers.buf_texadd0[2] ),
    .B(net377));
 sg13g2_nand2_1 _18528_ (.Y(_10981_),
    .A(\rbzero.spi_registers.texadd0[2] ),
    .B(net376));
 sg13g2_buf_1 _18529_ (.A(_10897_),
    .X(_10982_));
 sg13g2_a21oi_1 _18530_ (.A1(_10980_),
    .A2(_10981_),
    .Y(_00960_),
    .B1(net646));
 sg13g2_nand2_1 _18531_ (.Y(_10983_),
    .A(\rbzero.spi_registers.buf_texadd0[3] ),
    .B(_10961_));
 sg13g2_nand2_1 _18532_ (.Y(_10984_),
    .A(\rbzero.spi_registers.texadd0[3] ),
    .B(_10964_));
 sg13g2_a21oi_1 _18533_ (.A1(_10983_),
    .A2(_10984_),
    .Y(_00961_),
    .B1(net646));
 sg13g2_buf_1 _18534_ (.A(_10960_),
    .X(_10985_));
 sg13g2_nand2_1 _18535_ (.Y(_10986_),
    .A(\rbzero.spi_registers.buf_texadd0[4] ),
    .B(net375));
 sg13g2_buf_1 _18536_ (.A(_10963_),
    .X(_10987_));
 sg13g2_nand2_1 _18537_ (.Y(_10988_),
    .A(\rbzero.spi_registers.texadd0[4] ),
    .B(net374));
 sg13g2_a21oi_1 _18538_ (.A1(_10986_),
    .A2(_10988_),
    .Y(_00962_),
    .B1(net646));
 sg13g2_nand2_1 _18539_ (.Y(_10989_),
    .A(\rbzero.spi_registers.buf_texadd0[5] ),
    .B(net375));
 sg13g2_nand2_1 _18540_ (.Y(_10990_),
    .A(\rbzero.spi_registers.texadd0[5] ),
    .B(net374));
 sg13g2_a21oi_1 _18541_ (.A1(_10989_),
    .A2(_10990_),
    .Y(_00963_),
    .B1(net646));
 sg13g2_nand2_1 _18542_ (.Y(_10991_),
    .A(\rbzero.spi_registers.buf_texadd0[6] ),
    .B(net375));
 sg13g2_nand2_1 _18543_ (.Y(_10992_),
    .A(\rbzero.spi_registers.texadd0[6] ),
    .B(net374));
 sg13g2_a21oi_1 _18544_ (.A1(_10991_),
    .A2(_10992_),
    .Y(_00964_),
    .B1(net646));
 sg13g2_nand2_1 _18545_ (.Y(_10993_),
    .A(\rbzero.spi_registers.buf_texadd0[7] ),
    .B(net375));
 sg13g2_nand2_1 _18546_ (.Y(_10994_),
    .A(\rbzero.spi_registers.texadd0[7] ),
    .B(net374));
 sg13g2_a21oi_1 _18547_ (.A1(_10993_),
    .A2(_10994_),
    .Y(_00965_),
    .B1(net646));
 sg13g2_nand2_1 _18548_ (.Y(_10995_),
    .A(\rbzero.spi_registers.buf_texadd0[8] ),
    .B(net375));
 sg13g2_nand2_1 _18549_ (.Y(_10996_),
    .A(\rbzero.spi_registers.texadd0[8] ),
    .B(net374));
 sg13g2_a21oi_1 _18550_ (.A1(_10995_),
    .A2(_10996_),
    .Y(_00966_),
    .B1(net646));
 sg13g2_nand2_1 _18551_ (.Y(_10997_),
    .A(\rbzero.spi_registers.buf_texadd0[9] ),
    .B(net375));
 sg13g2_nand2_1 _18552_ (.Y(_10998_),
    .A(\rbzero.spi_registers.texadd0[9] ),
    .B(net374));
 sg13g2_a21oi_1 _18553_ (.A1(_10997_),
    .A2(_10998_),
    .Y(_00967_),
    .B1(net646));
 sg13g2_nand2_1 _18554_ (.Y(_10999_),
    .A(\rbzero.spi_registers.buf_texadd1[0] ),
    .B(_10985_));
 sg13g2_nand2_1 _18555_ (.Y(_11000_),
    .A(\rbzero.spi_registers.texadd1[0] ),
    .B(net374));
 sg13g2_a21oi_1 _18556_ (.A1(_10999_),
    .A2(_11000_),
    .Y(_00968_),
    .B1(_10982_));
 sg13g2_nand2_1 _18557_ (.Y(_11001_),
    .A(\rbzero.spi_registers.buf_texadd1[10] ),
    .B(net375));
 sg13g2_nand2_1 _18558_ (.Y(_11002_),
    .A(\rbzero.spi_registers.texadd1[10] ),
    .B(_10987_));
 sg13g2_a21oi_1 _18559_ (.A1(_11001_),
    .A2(_11002_),
    .Y(_00969_),
    .B1(_10982_));
 sg13g2_nand2_1 _18560_ (.Y(_11003_),
    .A(\rbzero.spi_registers.buf_texadd1[11] ),
    .B(net375));
 sg13g2_nand2_1 _18561_ (.Y(_11004_),
    .A(\rbzero.spi_registers.texadd1[11] ),
    .B(_10987_));
 sg13g2_buf_1 _18562_ (.A(_10897_),
    .X(_11005_));
 sg13g2_a21oi_1 _18563_ (.A1(_11003_),
    .A2(_11004_),
    .Y(_00970_),
    .B1(net645));
 sg13g2_nand2_1 _18564_ (.Y(_11006_),
    .A(\rbzero.spi_registers.buf_texadd1[12] ),
    .B(_10985_));
 sg13g2_nand2_1 _18565_ (.Y(_11007_),
    .A(\rbzero.spi_registers.texadd1[12] ),
    .B(net374));
 sg13g2_a21oi_1 _18566_ (.A1(_11006_),
    .A2(_11007_),
    .Y(_00971_),
    .B1(net645));
 sg13g2_buf_1 _18567_ (.A(_10960_),
    .X(_11008_));
 sg13g2_nand2_1 _18568_ (.Y(_11009_),
    .A(\rbzero.spi_registers.buf_texadd1[13] ),
    .B(_11008_));
 sg13g2_buf_1 _18569_ (.A(_10963_),
    .X(_11010_));
 sg13g2_nand2_1 _18570_ (.Y(_11011_),
    .A(\rbzero.spi_registers.texadd1[13] ),
    .B(_11010_));
 sg13g2_a21oi_1 _18571_ (.A1(_11009_),
    .A2(_11011_),
    .Y(_00972_),
    .B1(_11005_));
 sg13g2_nand2_1 _18572_ (.Y(_11012_),
    .A(\rbzero.spi_registers.buf_texadd1[14] ),
    .B(_11008_));
 sg13g2_nand2_1 _18573_ (.Y(_11013_),
    .A(\rbzero.spi_registers.texadd1[14] ),
    .B(net372));
 sg13g2_a21oi_1 _18574_ (.A1(_11012_),
    .A2(_11013_),
    .Y(_00973_),
    .B1(_11005_));
 sg13g2_nand2_1 _18575_ (.Y(_11014_),
    .A(\rbzero.spi_registers.buf_texadd1[15] ),
    .B(net373));
 sg13g2_nand2_1 _18576_ (.Y(_11015_),
    .A(\rbzero.spi_registers.texadd1[15] ),
    .B(_11010_));
 sg13g2_a21oi_1 _18577_ (.A1(_11014_),
    .A2(_11015_),
    .Y(_00974_),
    .B1(net645));
 sg13g2_nand2_1 _18578_ (.Y(_11016_),
    .A(\rbzero.spi_registers.buf_texadd1[16] ),
    .B(net373));
 sg13g2_nand2_1 _18579_ (.Y(_11017_),
    .A(\rbzero.spi_registers.texadd1[16] ),
    .B(net372));
 sg13g2_a21oi_1 _18580_ (.A1(_11016_),
    .A2(_11017_),
    .Y(_00975_),
    .B1(net645));
 sg13g2_nand2_1 _18581_ (.Y(_11018_),
    .A(\rbzero.spi_registers.buf_texadd1[17] ),
    .B(net373));
 sg13g2_nand2_1 _18582_ (.Y(_11019_),
    .A(\rbzero.spi_registers.texadd1[17] ),
    .B(net372));
 sg13g2_a21oi_1 _18583_ (.A1(_11018_),
    .A2(_11019_),
    .Y(_00976_),
    .B1(net645));
 sg13g2_nand2_1 _18584_ (.Y(_11020_),
    .A(\rbzero.spi_registers.buf_texadd1[18] ),
    .B(net373));
 sg13g2_nand2_1 _18585_ (.Y(_11021_),
    .A(\rbzero.spi_registers.texadd1[18] ),
    .B(net372));
 sg13g2_a21oi_1 _18586_ (.A1(_11020_),
    .A2(_11021_),
    .Y(_00977_),
    .B1(net645));
 sg13g2_nand2_1 _18587_ (.Y(_11022_),
    .A(\rbzero.spi_registers.buf_texadd1[19] ),
    .B(net373));
 sg13g2_nand2_1 _18588_ (.Y(_11023_),
    .A(\rbzero.spi_registers.texadd1[19] ),
    .B(net372));
 sg13g2_a21oi_1 _18589_ (.A1(_11022_),
    .A2(_11023_),
    .Y(_00978_),
    .B1(net645));
 sg13g2_nand2_1 _18590_ (.Y(_11024_),
    .A(\rbzero.spi_registers.buf_texadd1[1] ),
    .B(net373));
 sg13g2_nand2_1 _18591_ (.Y(_11025_),
    .A(\rbzero.spi_registers.texadd1[1] ),
    .B(net372));
 sg13g2_a21oi_1 _18592_ (.A1(_11024_),
    .A2(_11025_),
    .Y(_00979_),
    .B1(net645));
 sg13g2_nand2_1 _18593_ (.Y(_11026_),
    .A(\rbzero.spi_registers.buf_texadd1[20] ),
    .B(net373));
 sg13g2_nand2_1 _18594_ (.Y(_11027_),
    .A(\rbzero.spi_registers.texadd1[20] ),
    .B(net372));
 sg13g2_buf_1 _18595_ (.A(_10897_),
    .X(_11028_));
 sg13g2_a21oi_1 _18596_ (.A1(_11026_),
    .A2(_11027_),
    .Y(_00980_),
    .B1(net644));
 sg13g2_nand2_1 _18597_ (.Y(_11029_),
    .A(\rbzero.spi_registers.buf_texadd1[21] ),
    .B(net373));
 sg13g2_nand2_1 _18598_ (.Y(_11030_),
    .A(\rbzero.spi_registers.texadd1[21] ),
    .B(net372));
 sg13g2_a21oi_1 _18599_ (.A1(_11029_),
    .A2(_11030_),
    .Y(_00981_),
    .B1(net644));
 sg13g2_buf_1 _18600_ (.A(_10960_),
    .X(_11031_));
 sg13g2_nand2_1 _18601_ (.Y(_11032_),
    .A(\rbzero.spi_registers.buf_texadd1[22] ),
    .B(net371));
 sg13g2_buf_1 _18602_ (.A(_10963_),
    .X(_11033_));
 sg13g2_nand2_1 _18603_ (.Y(_11034_),
    .A(\rbzero.spi_registers.texadd1[22] ),
    .B(net370));
 sg13g2_a21oi_1 _18604_ (.A1(_11032_),
    .A2(_11034_),
    .Y(_00982_),
    .B1(net644));
 sg13g2_nand2_1 _18605_ (.Y(_11035_),
    .A(\rbzero.spi_registers.buf_texadd1[23] ),
    .B(net371));
 sg13g2_nand2_1 _18606_ (.Y(_11036_),
    .A(\rbzero.spi_registers.texadd1[23] ),
    .B(net370));
 sg13g2_a21oi_1 _18607_ (.A1(_11035_),
    .A2(_11036_),
    .Y(_00983_),
    .B1(net644));
 sg13g2_nand2_1 _18608_ (.Y(_11037_),
    .A(\rbzero.spi_registers.buf_texadd1[2] ),
    .B(net371));
 sg13g2_nand2_1 _18609_ (.Y(_11038_),
    .A(\rbzero.spi_registers.texadd1[2] ),
    .B(net370));
 sg13g2_a21oi_1 _18610_ (.A1(_11037_),
    .A2(_11038_),
    .Y(_00984_),
    .B1(net644));
 sg13g2_nand2_1 _18611_ (.Y(_11039_),
    .A(\rbzero.spi_registers.buf_texadd1[3] ),
    .B(net371));
 sg13g2_nand2_1 _18612_ (.Y(_11040_),
    .A(\rbzero.spi_registers.texadd1[3] ),
    .B(net370));
 sg13g2_a21oi_1 _18613_ (.A1(_11039_),
    .A2(_11040_),
    .Y(_00985_),
    .B1(net644));
 sg13g2_nand2_1 _18614_ (.Y(_11041_),
    .A(\rbzero.spi_registers.buf_texadd1[4] ),
    .B(net371));
 sg13g2_nand2_1 _18615_ (.Y(_11042_),
    .A(\rbzero.spi_registers.texadd1[4] ),
    .B(net370));
 sg13g2_a21oi_1 _18616_ (.A1(_11041_),
    .A2(_11042_),
    .Y(_00986_),
    .B1(net644));
 sg13g2_nand2_1 _18617_ (.Y(_11043_),
    .A(\rbzero.spi_registers.buf_texadd1[5] ),
    .B(net371));
 sg13g2_nand2_1 _18618_ (.Y(_11044_),
    .A(\rbzero.spi_registers.texadd1[5] ),
    .B(net370));
 sg13g2_a21oi_1 _18619_ (.A1(_11043_),
    .A2(_11044_),
    .Y(_00987_),
    .B1(net644));
 sg13g2_nand2_1 _18620_ (.Y(_11045_),
    .A(\rbzero.spi_registers.buf_texadd1[6] ),
    .B(net371));
 sg13g2_nand2_1 _18621_ (.Y(_11046_),
    .A(\rbzero.spi_registers.texadd1[6] ),
    .B(net370));
 sg13g2_a21oi_1 _18622_ (.A1(_11045_),
    .A2(_11046_),
    .Y(_00988_),
    .B1(_11028_));
 sg13g2_nand2_1 _18623_ (.Y(_11047_),
    .A(\rbzero.spi_registers.buf_texadd1[7] ),
    .B(net371));
 sg13g2_nand2_1 _18624_ (.Y(_11048_),
    .A(\rbzero.spi_registers.texadd1[7] ),
    .B(net370));
 sg13g2_a21oi_1 _18625_ (.A1(_11047_),
    .A2(_11048_),
    .Y(_00989_),
    .B1(_11028_));
 sg13g2_nand2_1 _18626_ (.Y(_11049_),
    .A(\rbzero.spi_registers.buf_texadd1[8] ),
    .B(_11031_));
 sg13g2_nand2_1 _18627_ (.Y(_11050_),
    .A(\rbzero.spi_registers.texadd1[8] ),
    .B(_11033_));
 sg13g2_buf_1 _18628_ (.A(_10897_),
    .X(_11051_));
 sg13g2_a21oi_1 _18629_ (.A1(_11049_),
    .A2(_11050_),
    .Y(_00990_),
    .B1(_11051_));
 sg13g2_nand2_1 _18630_ (.Y(_11052_),
    .A(\rbzero.spi_registers.buf_texadd1[9] ),
    .B(_11031_));
 sg13g2_nand2_1 _18631_ (.Y(_11053_),
    .A(\rbzero.spi_registers.texadd1[9] ),
    .B(_11033_));
 sg13g2_a21oi_1 _18632_ (.A1(_11052_),
    .A2(_11053_),
    .Y(_00991_),
    .B1(_11051_));
 sg13g2_buf_1 _18633_ (.A(_10960_),
    .X(_11054_));
 sg13g2_nand2_1 _18634_ (.Y(_11055_),
    .A(\rbzero.spi_registers.buf_texadd2[0] ),
    .B(net369));
 sg13g2_buf_1 _18635_ (.A(_10963_),
    .X(_11056_));
 sg13g2_nand2_1 _18636_ (.Y(_11057_),
    .A(\rbzero.spi_registers.texadd2[0] ),
    .B(net368));
 sg13g2_a21oi_1 _18637_ (.A1(_11055_),
    .A2(_11057_),
    .Y(_00992_),
    .B1(net643));
 sg13g2_nand2_1 _18638_ (.Y(_11058_),
    .A(\rbzero.spi_registers.buf_texadd2[10] ),
    .B(net369));
 sg13g2_nand2_1 _18639_ (.Y(_11059_),
    .A(\rbzero.spi_registers.texadd2[10] ),
    .B(net368));
 sg13g2_a21oi_1 _18640_ (.A1(_11058_),
    .A2(_11059_),
    .Y(_00993_),
    .B1(net643));
 sg13g2_nand2_1 _18641_ (.Y(_11060_),
    .A(\rbzero.spi_registers.buf_texadd2[11] ),
    .B(net369));
 sg13g2_nand2_1 _18642_ (.Y(_11061_),
    .A(\rbzero.spi_registers.texadd2[11] ),
    .B(net368));
 sg13g2_a21oi_1 _18643_ (.A1(_11060_),
    .A2(_11061_),
    .Y(_00994_),
    .B1(net643));
 sg13g2_nand2_1 _18644_ (.Y(_11062_),
    .A(\rbzero.spi_registers.buf_texadd2[12] ),
    .B(_11054_));
 sg13g2_nand2_1 _18645_ (.Y(_11063_),
    .A(\rbzero.spi_registers.texadd2[12] ),
    .B(_11056_));
 sg13g2_a21oi_1 _18646_ (.A1(_11062_),
    .A2(_11063_),
    .Y(_00995_),
    .B1(net643));
 sg13g2_nand2_1 _18647_ (.Y(_11064_),
    .A(\rbzero.spi_registers.buf_texadd2[13] ),
    .B(_11054_));
 sg13g2_nand2_1 _18648_ (.Y(_11065_),
    .A(\rbzero.spi_registers.texadd2[13] ),
    .B(_11056_));
 sg13g2_a21oi_1 _18649_ (.A1(_11064_),
    .A2(_11065_),
    .Y(_00996_),
    .B1(net643));
 sg13g2_nand2_1 _18650_ (.Y(_11066_),
    .A(\rbzero.spi_registers.buf_texadd2[14] ),
    .B(net369));
 sg13g2_nand2_1 _18651_ (.Y(_11067_),
    .A(\rbzero.spi_registers.texadd2[14] ),
    .B(net368));
 sg13g2_a21oi_1 _18652_ (.A1(_11066_),
    .A2(_11067_),
    .Y(_00997_),
    .B1(net643));
 sg13g2_nand2_1 _18653_ (.Y(_11068_),
    .A(\rbzero.spi_registers.buf_texadd2[15] ),
    .B(net369));
 sg13g2_nand2_1 _18654_ (.Y(_11069_),
    .A(\rbzero.spi_registers.texadd2[15] ),
    .B(net368));
 sg13g2_a21oi_1 _18655_ (.A1(_11068_),
    .A2(_11069_),
    .Y(_00998_),
    .B1(net643));
 sg13g2_nand2_1 _18656_ (.Y(_11070_),
    .A(\rbzero.spi_registers.buf_texadd2[16] ),
    .B(net369));
 sg13g2_nand2_1 _18657_ (.Y(_11071_),
    .A(\rbzero.spi_registers.texadd2[16] ),
    .B(net368));
 sg13g2_a21oi_1 _18658_ (.A1(_11070_),
    .A2(_11071_),
    .Y(_00999_),
    .B1(net643));
 sg13g2_nand2_1 _18659_ (.Y(_11072_),
    .A(\rbzero.spi_registers.buf_texadd2[17] ),
    .B(net369));
 sg13g2_nand2_1 _18660_ (.Y(_11073_),
    .A(\rbzero.spi_registers.texadd2[17] ),
    .B(net368));
 sg13g2_buf_1 _18661_ (.A(_10897_),
    .X(_11074_));
 sg13g2_a21oi_1 _18662_ (.A1(_11072_),
    .A2(_11073_),
    .Y(_01000_),
    .B1(net642));
 sg13g2_nand2_1 _18663_ (.Y(_11075_),
    .A(\rbzero.spi_registers.buf_texadd2[18] ),
    .B(net369));
 sg13g2_nand2_1 _18664_ (.Y(_11076_),
    .A(\rbzero.spi_registers.texadd2[18] ),
    .B(net368));
 sg13g2_a21oi_1 _18665_ (.A1(_11075_),
    .A2(_11076_),
    .Y(_01001_),
    .B1(net642));
 sg13g2_buf_1 _18666_ (.A(_10960_),
    .X(_11077_));
 sg13g2_nand2_1 _18667_ (.Y(_11078_),
    .A(\rbzero.spi_registers.buf_texadd2[19] ),
    .B(net367));
 sg13g2_buf_1 _18668_ (.A(_10963_),
    .X(_11079_));
 sg13g2_nand2_1 _18669_ (.Y(_11080_),
    .A(\rbzero.spi_registers.texadd2[19] ),
    .B(net366));
 sg13g2_a21oi_1 _18670_ (.A1(_11078_),
    .A2(_11080_),
    .Y(_01002_),
    .B1(net642));
 sg13g2_nand2_1 _18671_ (.Y(_11081_),
    .A(\rbzero.spi_registers.buf_texadd2[1] ),
    .B(net367));
 sg13g2_nand2_1 _18672_ (.Y(_11082_),
    .A(\rbzero.spi_registers.texadd2[1] ),
    .B(net366));
 sg13g2_a21oi_1 _18673_ (.A1(_11081_),
    .A2(_11082_),
    .Y(_01003_),
    .B1(net642));
 sg13g2_nand2_1 _18674_ (.Y(_11083_),
    .A(\rbzero.spi_registers.buf_texadd2[20] ),
    .B(net367));
 sg13g2_nand2_1 _18675_ (.Y(_11084_),
    .A(\rbzero.spi_registers.texadd2[20] ),
    .B(net366));
 sg13g2_a21oi_1 _18676_ (.A1(_11083_),
    .A2(_11084_),
    .Y(_01004_),
    .B1(net642));
 sg13g2_nand2_1 _18677_ (.Y(_11085_),
    .A(\rbzero.spi_registers.buf_texadd2[21] ),
    .B(net367));
 sg13g2_nand2_1 _18678_ (.Y(_11086_),
    .A(\rbzero.spi_registers.texadd2[21] ),
    .B(net366));
 sg13g2_a21oi_1 _18679_ (.A1(_11085_),
    .A2(_11086_),
    .Y(_01005_),
    .B1(_11074_));
 sg13g2_nand2_1 _18680_ (.Y(_11087_),
    .A(\rbzero.spi_registers.buf_texadd2[22] ),
    .B(net367));
 sg13g2_nand2_1 _18681_ (.Y(_11088_),
    .A(\rbzero.spi_registers.texadd2[22] ),
    .B(_11079_));
 sg13g2_a21oi_1 _18682_ (.A1(_11087_),
    .A2(_11088_),
    .Y(_01006_),
    .B1(net642));
 sg13g2_nand2_1 _18683_ (.Y(_11089_),
    .A(\rbzero.spi_registers.buf_texadd2[23] ),
    .B(net367));
 sg13g2_nand2_1 _18684_ (.Y(_11090_),
    .A(\rbzero.spi_registers.texadd2[23] ),
    .B(_11079_));
 sg13g2_a21oi_1 _18685_ (.A1(_11089_),
    .A2(_11090_),
    .Y(_01007_),
    .B1(_11074_));
 sg13g2_nand2_1 _18686_ (.Y(_11091_),
    .A(\rbzero.spi_registers.buf_texadd2[2] ),
    .B(net367));
 sg13g2_nand2_1 _18687_ (.Y(_11092_),
    .A(\rbzero.spi_registers.texadd2[2] ),
    .B(net366));
 sg13g2_a21oi_1 _18688_ (.A1(_11091_),
    .A2(_11092_),
    .Y(_01008_),
    .B1(net642));
 sg13g2_nand2_1 _18689_ (.Y(_11093_),
    .A(\rbzero.spi_registers.buf_texadd2[3] ),
    .B(net367));
 sg13g2_nand2_1 _18690_ (.Y(_11094_),
    .A(\rbzero.spi_registers.texadd2[3] ),
    .B(net366));
 sg13g2_a21oi_1 _18691_ (.A1(_11093_),
    .A2(_11094_),
    .Y(_01009_),
    .B1(net642));
 sg13g2_nand2_1 _18692_ (.Y(_11095_),
    .A(\rbzero.spi_registers.buf_texadd2[4] ),
    .B(_11077_));
 sg13g2_nand2_1 _18693_ (.Y(_11096_),
    .A(\rbzero.spi_registers.texadd2[4] ),
    .B(net366));
 sg13g2_buf_1 _18694_ (.A(_09700_),
    .X(_11097_));
 sg13g2_a21oi_1 _18695_ (.A1(_11095_),
    .A2(_11096_),
    .Y(_01010_),
    .B1(net641));
 sg13g2_nand2_1 _18696_ (.Y(_11098_),
    .A(\rbzero.spi_registers.buf_texadd2[5] ),
    .B(_11077_));
 sg13g2_nand2_1 _18697_ (.Y(_11099_),
    .A(\rbzero.spi_registers.texadd2[5] ),
    .B(net366));
 sg13g2_a21oi_1 _18698_ (.A1(_11098_),
    .A2(_11099_),
    .Y(_01011_),
    .B1(net641));
 sg13g2_buf_1 _18699_ (.A(_10960_),
    .X(_11100_));
 sg13g2_nand2_1 _18700_ (.Y(_11101_),
    .A(\rbzero.spi_registers.buf_texadd2[6] ),
    .B(net365));
 sg13g2_buf_1 _18701_ (.A(_10963_),
    .X(_11102_));
 sg13g2_nand2_1 _18702_ (.Y(_11103_),
    .A(\rbzero.spi_registers.texadd2[6] ),
    .B(net364));
 sg13g2_a21oi_1 _18703_ (.A1(_11101_),
    .A2(_11103_),
    .Y(_01012_),
    .B1(_11097_));
 sg13g2_nand2_1 _18704_ (.Y(_11104_),
    .A(\rbzero.spi_registers.buf_texadd2[7] ),
    .B(net365));
 sg13g2_nand2_1 _18705_ (.Y(_11105_),
    .A(\rbzero.spi_registers.texadd2[7] ),
    .B(net364));
 sg13g2_a21oi_1 _18706_ (.A1(_11104_),
    .A2(_11105_),
    .Y(_01013_),
    .B1(_11097_));
 sg13g2_nand2_1 _18707_ (.Y(_11106_),
    .A(\rbzero.spi_registers.buf_texadd2[8] ),
    .B(_11100_));
 sg13g2_nand2_1 _18708_ (.Y(_11107_),
    .A(\rbzero.spi_registers.texadd2[8] ),
    .B(_11102_));
 sg13g2_a21oi_1 _18709_ (.A1(_11106_),
    .A2(_11107_),
    .Y(_01014_),
    .B1(net641));
 sg13g2_nand2_1 _18710_ (.Y(_11108_),
    .A(\rbzero.spi_registers.buf_texadd2[9] ),
    .B(net365));
 sg13g2_nand2_1 _18711_ (.Y(_11109_),
    .A(\rbzero.spi_registers.texadd2[9] ),
    .B(_11102_));
 sg13g2_a21oi_1 _18712_ (.A1(_11108_),
    .A2(_11109_),
    .Y(_01015_),
    .B1(net641));
 sg13g2_nand2_1 _18713_ (.Y(_11110_),
    .A(\rbzero.spi_registers.buf_texadd3[0] ),
    .B(net365));
 sg13g2_nand2_1 _18714_ (.Y(_11111_),
    .A(\rbzero.spi_registers.texadd3[0] ),
    .B(net364));
 sg13g2_a21oi_1 _18715_ (.A1(_11110_),
    .A2(_11111_),
    .Y(_01016_),
    .B1(net641));
 sg13g2_nand2_1 _18716_ (.Y(_11112_),
    .A(\rbzero.spi_registers.buf_texadd3[10] ),
    .B(net365));
 sg13g2_nand2_1 _18717_ (.Y(_11113_),
    .A(\rbzero.spi_registers.texadd3[10] ),
    .B(net364));
 sg13g2_a21oi_1 _18718_ (.A1(_11112_),
    .A2(_11113_),
    .Y(_01017_),
    .B1(net641));
 sg13g2_nand2_1 _18719_ (.Y(_11114_),
    .A(\rbzero.spi_registers.buf_texadd3[11] ),
    .B(net365));
 sg13g2_nand2_1 _18720_ (.Y(_11115_),
    .A(\rbzero.spi_registers.texadd3[11] ),
    .B(net364));
 sg13g2_a21oi_1 _18721_ (.A1(_11114_),
    .A2(_11115_),
    .Y(_01018_),
    .B1(net641));
 sg13g2_nand2_1 _18722_ (.Y(_11116_),
    .A(\rbzero.spi_registers.buf_texadd3[12] ),
    .B(net365));
 sg13g2_nand2_1 _18723_ (.Y(_11117_),
    .A(\rbzero.spi_registers.texadd3[12] ),
    .B(net364));
 sg13g2_a21oi_1 _18724_ (.A1(_11116_),
    .A2(_11117_),
    .Y(_01019_),
    .B1(net641));
 sg13g2_nand2_1 _18725_ (.Y(_11118_),
    .A(\rbzero.spi_registers.buf_texadd3[13] ),
    .B(net365));
 sg13g2_nand2_1 _18726_ (.Y(_11119_),
    .A(\rbzero.spi_registers.texadd3[13] ),
    .B(net364));
 sg13g2_buf_1 _18727_ (.A(_09700_),
    .X(_11120_));
 sg13g2_a21oi_1 _18728_ (.A1(_11118_),
    .A2(_11119_),
    .Y(_01020_),
    .B1(_11120_));
 sg13g2_nand2_1 _18729_ (.Y(_11121_),
    .A(\rbzero.spi_registers.buf_texadd3[14] ),
    .B(_11100_));
 sg13g2_nand2_1 _18730_ (.Y(_11122_),
    .A(\rbzero.spi_registers.texadd3[14] ),
    .B(net364));
 sg13g2_a21oi_1 _18731_ (.A1(_11121_),
    .A2(_11122_),
    .Y(_01021_),
    .B1(net640));
 sg13g2_buf_1 _18732_ (.A(net451),
    .X(_11123_));
 sg13g2_nand2_1 _18733_ (.Y(_11124_),
    .A(\rbzero.spi_registers.buf_texadd3[15] ),
    .B(_11123_));
 sg13g2_buf_1 _18734_ (.A(_09416_),
    .X(_11125_));
 sg13g2_nand2_1 _18735_ (.Y(_11126_),
    .A(\rbzero.spi_registers.texadd3[15] ),
    .B(net410));
 sg13g2_a21oi_1 _18736_ (.A1(_11124_),
    .A2(_11126_),
    .Y(_01022_),
    .B1(net640));
 sg13g2_nand2_1 _18737_ (.Y(_11127_),
    .A(\rbzero.spi_registers.buf_texadd3[16] ),
    .B(_11123_));
 sg13g2_nand2_1 _18738_ (.Y(_11128_),
    .A(\rbzero.spi_registers.texadd3[16] ),
    .B(net410));
 sg13g2_a21oi_1 _18739_ (.A1(_11127_),
    .A2(_11128_),
    .Y(_01023_),
    .B1(_11120_));
 sg13g2_nand2_1 _18740_ (.Y(_11129_),
    .A(\rbzero.spi_registers.buf_texadd3[17] ),
    .B(net411));
 sg13g2_nand2_1 _18741_ (.Y(_11130_),
    .A(\rbzero.spi_registers.texadd3[17] ),
    .B(net410));
 sg13g2_a21oi_1 _18742_ (.A1(_11129_),
    .A2(_11130_),
    .Y(_01024_),
    .B1(net640));
 sg13g2_nand2_1 _18743_ (.Y(_11131_),
    .A(\rbzero.spi_registers.buf_texadd3[18] ),
    .B(net411));
 sg13g2_nand2_1 _18744_ (.Y(_11132_),
    .A(\rbzero.spi_registers.texadd3[18] ),
    .B(net410));
 sg13g2_a21oi_1 _18745_ (.A1(_11131_),
    .A2(_11132_),
    .Y(_01025_),
    .B1(net640));
 sg13g2_nand2_1 _18746_ (.Y(_11133_),
    .A(\rbzero.spi_registers.buf_texadd3[19] ),
    .B(net411));
 sg13g2_nand2_1 _18747_ (.Y(_11134_),
    .A(\rbzero.spi_registers.texadd3[19] ),
    .B(net410));
 sg13g2_a21oi_1 _18748_ (.A1(_11133_),
    .A2(_11134_),
    .Y(_01026_),
    .B1(net640));
 sg13g2_nand2_1 _18749_ (.Y(_11135_),
    .A(\rbzero.spi_registers.buf_texadd3[1] ),
    .B(net411));
 sg13g2_nand2_1 _18750_ (.Y(_11136_),
    .A(\rbzero.spi_registers.texadd3[1] ),
    .B(net410));
 sg13g2_a21oi_1 _18751_ (.A1(_11135_),
    .A2(_11136_),
    .Y(_01027_),
    .B1(net640));
 sg13g2_nand2_1 _18752_ (.Y(_11137_),
    .A(\rbzero.spi_registers.buf_texadd3[20] ),
    .B(net411));
 sg13g2_nand2_1 _18753_ (.Y(_11138_),
    .A(\rbzero.spi_registers.texadd3[20] ),
    .B(net410));
 sg13g2_a21oi_1 _18754_ (.A1(_11137_),
    .A2(_11138_),
    .Y(_01028_),
    .B1(net640));
 sg13g2_nand2_1 _18755_ (.Y(_11139_),
    .A(\rbzero.spi_registers.buf_texadd3[21] ),
    .B(net411));
 sg13g2_nand2_1 _18756_ (.Y(_11140_),
    .A(\rbzero.spi_registers.texadd3[21] ),
    .B(net410));
 sg13g2_a21oi_1 _18757_ (.A1(_11139_),
    .A2(_11140_),
    .Y(_01029_),
    .B1(net640));
 sg13g2_nand2_1 _18758_ (.Y(_11141_),
    .A(\rbzero.spi_registers.buf_texadd3[22] ),
    .B(net411));
 sg13g2_nand2_1 _18759_ (.Y(_11142_),
    .A(\rbzero.spi_registers.texadd3[22] ),
    .B(_11125_));
 sg13g2_buf_1 _18760_ (.A(_09700_),
    .X(_11143_));
 sg13g2_a21oi_1 _18761_ (.A1(_11141_),
    .A2(_11142_),
    .Y(_01030_),
    .B1(net639));
 sg13g2_nand2_1 _18762_ (.Y(_11144_),
    .A(\rbzero.spi_registers.buf_texadd3[23] ),
    .B(net411));
 sg13g2_nand2_1 _18763_ (.Y(_11145_),
    .A(\rbzero.spi_registers.texadd3[23] ),
    .B(_11125_));
 sg13g2_a21oi_1 _18764_ (.A1(_11144_),
    .A2(_11145_),
    .Y(_01031_),
    .B1(net639));
 sg13g2_buf_1 _18765_ (.A(net451),
    .X(_11146_));
 sg13g2_nand2_1 _18766_ (.Y(_11147_),
    .A(\rbzero.spi_registers.buf_texadd3[2] ),
    .B(net409));
 sg13g2_buf_1 _18767_ (.A(_09416_),
    .X(_11148_));
 sg13g2_nand2_1 _18768_ (.Y(_11149_),
    .A(\rbzero.spi_registers.texadd3[2] ),
    .B(net408));
 sg13g2_a21oi_1 _18769_ (.A1(_11147_),
    .A2(_11149_),
    .Y(_01032_),
    .B1(net639));
 sg13g2_nand2_1 _18770_ (.Y(_11150_),
    .A(\rbzero.spi_registers.buf_texadd3[3] ),
    .B(net409));
 sg13g2_nand2_1 _18771_ (.Y(_11151_),
    .A(\rbzero.spi_registers.texadd3[3] ),
    .B(net408));
 sg13g2_a21oi_1 _18772_ (.A1(_11150_),
    .A2(_11151_),
    .Y(_01033_),
    .B1(net639));
 sg13g2_nand2_1 _18773_ (.Y(_11152_),
    .A(\rbzero.spi_registers.buf_texadd3[4] ),
    .B(net409));
 sg13g2_nand2_1 _18774_ (.Y(_11153_),
    .A(\rbzero.spi_registers.texadd3[4] ),
    .B(net408));
 sg13g2_a21oi_1 _18775_ (.A1(_11152_),
    .A2(_11153_),
    .Y(_01034_),
    .B1(net639));
 sg13g2_nand2_1 _18776_ (.Y(_11154_),
    .A(\rbzero.spi_registers.buf_texadd3[5] ),
    .B(net409));
 sg13g2_nand2_1 _18777_ (.Y(_11155_),
    .A(\rbzero.spi_registers.texadd3[5] ),
    .B(net408));
 sg13g2_a21oi_1 _18778_ (.A1(_11154_),
    .A2(_11155_),
    .Y(_01035_),
    .B1(net639));
 sg13g2_nand2_1 _18779_ (.Y(_11156_),
    .A(\rbzero.spi_registers.buf_texadd3[6] ),
    .B(net409));
 sg13g2_nand2_1 _18780_ (.Y(_11157_),
    .A(\rbzero.spi_registers.texadd3[6] ),
    .B(net408));
 sg13g2_a21oi_1 _18781_ (.A1(_11156_),
    .A2(_11157_),
    .Y(_01036_),
    .B1(net639));
 sg13g2_nand2_1 _18782_ (.Y(_11158_),
    .A(\rbzero.spi_registers.buf_texadd3[7] ),
    .B(net409));
 sg13g2_nand2_1 _18783_ (.Y(_11159_),
    .A(\rbzero.spi_registers.texadd3[7] ),
    .B(net408));
 sg13g2_a21oi_1 _18784_ (.A1(_11158_),
    .A2(_11159_),
    .Y(_01037_),
    .B1(net639));
 sg13g2_nand2_1 _18785_ (.Y(_11160_),
    .A(\rbzero.spi_registers.buf_texadd3[8] ),
    .B(net409));
 sg13g2_nand2_1 _18786_ (.Y(_11161_),
    .A(\rbzero.spi_registers.texadd3[8] ),
    .B(net408));
 sg13g2_a21oi_1 _18787_ (.A1(_11160_),
    .A2(_11161_),
    .Y(_01038_),
    .B1(_11143_));
 sg13g2_nand2_1 _18788_ (.Y(_11162_),
    .A(\rbzero.spi_registers.buf_texadd3[9] ),
    .B(net409));
 sg13g2_nand2_1 _18789_ (.Y(_11163_),
    .A(\rbzero.spi_registers.texadd3[9] ),
    .B(net408));
 sg13g2_a21oi_1 _18790_ (.A1(_11162_),
    .A2(_11163_),
    .Y(_01039_),
    .B1(_11143_));
 sg13g2_nand2_1 _18791_ (.Y(_11164_),
    .A(\rbzero.spi_registers.buf_vinf ),
    .B(_11146_));
 sg13g2_nand2_1 _18792_ (.Y(_11165_),
    .A(\rbzero.o_vinf ),
    .B(_11148_));
 sg13g2_a21oi_1 _18793_ (.A1(_11164_),
    .A2(_11165_),
    .Y(_01040_),
    .B1(net675));
 sg13g2_nand2_1 _18794_ (.Y(_11166_),
    .A(\rbzero.spi_registers.buf_vshift[0] ),
    .B(_11146_));
 sg13g2_buf_1 _18795_ (.A(\rbzero.spi_registers.vshift[0] ),
    .X(_11167_));
 sg13g2_nand2_1 _18796_ (.Y(_11168_),
    .A(_11167_),
    .B(_11148_));
 sg13g2_a21oi_1 _18797_ (.A1(_11166_),
    .A2(_11168_),
    .Y(_01041_),
    .B1(net675));
 sg13g2_nand2_1 _18798_ (.Y(_11169_),
    .A(\rbzero.spi_registers.buf_vshift[1] ),
    .B(net413));
 sg13g2_nand2_1 _18799_ (.Y(_11170_),
    .A(\rbzero.spi_registers.vshift[1] ),
    .B(net412));
 sg13g2_a21oi_1 _18800_ (.A1(_11169_),
    .A2(_11170_),
    .Y(_01042_),
    .B1(net675));
 sg13g2_nand2_1 _18801_ (.Y(_11171_),
    .A(\rbzero.spi_registers.buf_vshift[2] ),
    .B(net413));
 sg13g2_buf_2 _18802_ (.A(\rbzero.spi_registers.vshift[2] ),
    .X(_11172_));
 sg13g2_nand2_1 _18803_ (.Y(_11173_),
    .A(_11172_),
    .B(net412));
 sg13g2_a21oi_1 _18804_ (.A1(_11171_),
    .A2(_11173_),
    .Y(_01043_),
    .B1(net675));
 sg13g2_nand2_1 _18805_ (.Y(_11174_),
    .A(\rbzero.spi_registers.buf_vshift[3] ),
    .B(net413));
 sg13g2_nand2_1 _18806_ (.Y(_11175_),
    .A(\rbzero.spi_registers.vshift[3] ),
    .B(net412));
 sg13g2_a21oi_1 _18807_ (.A1(_11174_),
    .A2(_11175_),
    .Y(_01044_),
    .B1(net675));
 sg13g2_nand2_1 _18808_ (.Y(_11176_),
    .A(\rbzero.spi_registers.buf_vshift[4] ),
    .B(_10812_));
 sg13g2_nand2_1 _18809_ (.Y(_11177_),
    .A(\rbzero.spi_registers.vshift[4] ),
    .B(_10815_));
 sg13g2_a21oi_1 _18810_ (.A1(_11176_),
    .A2(_11177_),
    .Y(_01045_),
    .B1(net675));
 sg13g2_nand2_1 _18811_ (.Y(_11178_),
    .A(\rbzero.spi_registers.buf_vshift[5] ),
    .B(_10812_));
 sg13g2_buf_1 _18812_ (.A(\rbzero.spi_registers.vshift[5] ),
    .X(_11179_));
 sg13g2_nand2_1 _18813_ (.Y(_11180_),
    .A(_11179_),
    .B(_10815_));
 sg13g2_a21oi_1 _18814_ (.A1(_11178_),
    .A2(_11180_),
    .Y(_01046_),
    .B1(net675));
 sg13g2_nor2b_1 _18815_ (.A(_09412_),
    .B_N(_09399_),
    .Y(_11181_));
 sg13g2_nor2_1 _18816_ (.A(_09411_),
    .B(\rbzero.debug_overlay.vpos[8] ),
    .Y(_11182_));
 sg13g2_or2_1 _18817_ (.X(_11183_),
    .B(net816),
    .A(_09400_));
 sg13g2_buf_1 _18818_ (.A(_11183_),
    .X(_11184_));
 sg13g2_nor3_1 _18819_ (.A(_09398_),
    .B(net753),
    .C(_11184_),
    .Y(_11185_));
 sg13g2_nand4_1 _18820_ (.B(_11181_),
    .C(_11182_),
    .A(_09407_),
    .Y(_11186_),
    .D(_11185_));
 sg13g2_buf_1 _18821_ (.A(_11186_),
    .X(_11187_));
 sg13g2_nand3b_1 _18822_ (.B(net490),
    .C(_11187_),
    .Y(_11188_),
    .A_N(net816));
 sg13g2_nand2_1 _18823_ (.Y(_11189_),
    .A(net816),
    .B(_08473_));
 sg13g2_a21oi_1 _18824_ (.A1(_11188_),
    .A2(_11189_),
    .Y(_01464_),
    .B1(_09701_));
 sg13g2_nand2_1 _18825_ (.Y(_11190_),
    .A(net816),
    .B(net490));
 sg13g2_xnor2_1 _18826_ (.Y(_11191_),
    .A(_09400_),
    .B(_11190_));
 sg13g2_and2_1 _18827_ (.A(_09425_),
    .B(_11191_),
    .X(_01465_));
 sg13g2_o21ai_1 _18828_ (.B1(_09424_),
    .Y(_11192_),
    .A1(_08473_),
    .A2(_11187_));
 sg13g2_buf_2 _18829_ (.A(_11192_),
    .X(_11193_));
 sg13g2_nand3_1 _18830_ (.B(_09401_),
    .C(net490),
    .A(_09400_),
    .Y(_11194_));
 sg13g2_xnor2_1 _18831_ (.Y(_11195_),
    .A(_09406_),
    .B(_11194_));
 sg13g2_nor2_1 _18832_ (.A(_11193_),
    .B(_11195_),
    .Y(_01466_));
 sg13g2_or2_1 _18833_ (.X(_11196_),
    .B(_11194_),
    .A(_09406_));
 sg13g2_xnor2_1 _18834_ (.Y(_11197_),
    .A(_09404_),
    .B(_11196_));
 sg13g2_nor2_1 _18835_ (.A(_11193_),
    .B(_11197_),
    .Y(_01467_));
 sg13g2_nand4_1 _18836_ (.B(net816),
    .C(net490),
    .A(_09400_),
    .Y(_11198_),
    .D(_09407_));
 sg13g2_xor2_1 _18837_ (.B(_11198_),
    .A(net753),
    .X(_11199_));
 sg13g2_nor2_1 _18838_ (.A(_11193_),
    .B(_11199_),
    .Y(_01468_));
 sg13g2_buf_1 _18839_ (.A(_00058_),
    .X(_11200_));
 sg13g2_xnor2_1 _18840_ (.Y(_11201_),
    .A(_11200_),
    .B(_09408_));
 sg13g2_nor2_1 _18841_ (.A(_08473_),
    .B(_11201_),
    .Y(_11202_));
 sg13g2_a22oi_1 _18842_ (.Y(_11203_),
    .B1(_11187_),
    .B2(_11202_),
    .A2(_08473_),
    .A1(_09398_));
 sg13g2_nor2b_1 _18843_ (.A(_11203_),
    .B_N(_09425_),
    .Y(_01469_));
 sg13g2_nor2_1 _18844_ (.A(_09725_),
    .B(_09410_),
    .Y(_11204_));
 sg13g2_xnor2_1 _18845_ (.Y(_11205_),
    .A(_09412_),
    .B(_11204_));
 sg13g2_nor2_1 _18846_ (.A(_11193_),
    .B(_11205_),
    .Y(_01470_));
 sg13g2_nand2_1 _18847_ (.Y(_11206_),
    .A(_09412_),
    .B(_11204_));
 sg13g2_xor2_1 _18848_ (.B(_11206_),
    .A(_09411_),
    .X(_11207_));
 sg13g2_nor2_1 _18849_ (.A(_11193_),
    .B(_11207_),
    .Y(_01471_));
 sg13g2_nand3_1 _18850_ (.B(_09412_),
    .C(_11204_),
    .A(_09411_),
    .Y(_11208_));
 sg13g2_xor2_1 _18851_ (.B(_11208_),
    .A(\rbzero.debug_overlay.vpos[8] ),
    .X(_11209_));
 sg13g2_nor2_1 _18852_ (.A(_11193_),
    .B(_11209_),
    .Y(_01472_));
 sg13g2_nor3_1 _18853_ (.A(_09725_),
    .B(_09410_),
    .C(_09414_),
    .Y(_11210_));
 sg13g2_xnor2_1 _18854_ (.Y(_11211_),
    .A(_09399_),
    .B(_11210_));
 sg13g2_nor2_1 _18855_ (.A(_11193_),
    .B(_11211_),
    .Y(_01473_));
 sg13g2_buf_1 _18856_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .X(_11212_));
 sg13g2_inv_1 _18857_ (.Y(_11213_),
    .A(_11212_));
 sg13g2_buf_1 _18858_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_11214_));
 sg13g2_inv_1 _18859_ (.Y(_11215_),
    .A(_11214_));
 sg13g2_buf_1 _18860_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .X(_11216_));
 sg13g2_inv_1 _18861_ (.Y(_11217_),
    .A(_11216_));
 sg13g2_buf_2 _18862_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_11218_));
 sg13g2_buf_1 _18863_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .X(_11219_));
 sg13g2_nor2b_1 _18864_ (.A(_11218_),
    .B_N(_11219_),
    .Y(_11220_));
 sg13g2_buf_2 _18865_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .X(_11221_));
 sg13g2_buf_1 _18866_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .X(_11222_));
 sg13g2_inv_1 _18867_ (.Y(_11223_),
    .A(_11222_));
 sg13g2_buf_1 _18868_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .X(_11224_));
 sg13g2_inv_1 _18869_ (.Y(_11225_),
    .A(_11224_));
 sg13g2_buf_1 _18870_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .X(_11226_));
 sg13g2_buf_1 _18871_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .X(_11227_));
 sg13g2_buf_2 _18872_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .X(_11228_));
 sg13g2_buf_1 _18873_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .X(_11229_));
 sg13g2_nor2b_1 _18874_ (.A(_11228_),
    .B_N(_11229_),
    .Y(_11230_));
 sg13g2_buf_1 _18875_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .X(_11231_));
 sg13g2_buf_2 _18876_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .X(_11232_));
 sg13g2_buf_1 _18877_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .X(_11233_));
 sg13g2_buf_2 _18878_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .X(_11234_));
 sg13g2_nand2b_1 _18879_ (.Y(_11235_),
    .B(_11234_),
    .A_N(_11233_));
 sg13g2_buf_1 _18880_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .X(_11236_));
 sg13g2_buf_1 _18881_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .X(_11237_));
 sg13g2_buf_1 _18882_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .X(_11238_));
 sg13g2_buf_2 _18883_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .X(_11239_));
 sg13g2_inv_1 _18884_ (.Y(_11240_),
    .A(_11239_));
 sg13g2_inv_1 _18885_ (.Y(_11241_),
    .A(_11238_));
 sg13g2_buf_2 _18886_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .X(_11242_));
 sg13g2_buf_1 _18887_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(_11243_));
 sg13g2_buf_2 _18888_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_11244_));
 sg13g2_nand2b_1 _18889_ (.Y(_11245_),
    .B(_11244_),
    .A_N(_11243_));
 sg13g2_buf_1 _18890_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .X(_11246_));
 sg13g2_buf_1 _18891_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .X(_11247_));
 sg13g2_buf_1 _18892_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(_11248_));
 sg13g2_buf_2 _18893_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .X(_11249_));
 sg13g2_inv_1 _18894_ (.Y(_11250_),
    .A(_11249_));
 sg13g2_inv_1 _18895_ (.Y(_11251_),
    .A(_11248_));
 sg13g2_buf_1 _18896_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .X(_11252_));
 sg13g2_inv_1 _18897_ (.Y(_11253_),
    .A(_11252_));
 sg13g2_buf_1 _18898_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .X(_11254_));
 sg13g2_inv_1 _18899_ (.Y(_11255_),
    .A(_11254_));
 sg13g2_buf_1 _18900_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .X(_11256_));
 sg13g2_buf_1 _18901_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(_11257_));
 sg13g2_buf_1 _18902_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .X(_11258_));
 sg13g2_inv_1 _18903_ (.Y(_11259_),
    .A(_11258_));
 sg13g2_inv_1 _18904_ (.Y(_11260_),
    .A(_11257_));
 sg13g2_buf_1 _18905_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .X(_11261_));
 sg13g2_buf_2 _18906_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .X(_11262_));
 sg13g2_inv_1 _18907_ (.Y(_11263_),
    .A(_11262_));
 sg13g2_buf_1 _18908_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_11264_));
 sg13g2_inv_1 _18909_ (.Y(_11265_),
    .A(_11264_));
 sg13g2_inv_1 _18910_ (.Y(_11266_),
    .A(\rbzero.wall_tracer.trackDistX[-10] ));
 sg13g2_buf_2 _18911_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .X(_11267_));
 sg13g2_buf_2 _18912_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(_11268_));
 sg13g2_nor2b_1 _18913_ (.A(_11267_),
    .B_N(_11268_),
    .Y(_11269_));
 sg13g2_nand2_1 _18914_ (.Y(_11270_),
    .A(_11266_),
    .B(_11269_));
 sg13g2_o21ai_1 _18915_ (.B1(\rbzero.wall_tracer.trackDistY[-10] ),
    .Y(_11271_),
    .A1(_11266_),
    .A2(_11269_));
 sg13g2_a22oi_1 _18916_ (.Y(_11272_),
    .B1(_11270_),
    .B2(_11271_),
    .A2(_11265_),
    .A1(_11262_));
 sg13g2_a21oi_1 _18917_ (.A1(_11263_),
    .A2(_11264_),
    .Y(_11273_),
    .B1(_11272_));
 sg13g2_buf_1 _18918_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .X(_11274_));
 sg13g2_nor2_1 _18919_ (.A(_11261_),
    .B(_11273_),
    .Y(_11275_));
 sg13g2_nor2_1 _18920_ (.A(_11274_),
    .B(_11275_),
    .Y(_11276_));
 sg13g2_a221oi_1 _18921_ (.B2(_11273_),
    .C1(_11276_),
    .B1(_11261_),
    .A1(_11260_),
    .Y(_11277_),
    .A2(_11258_));
 sg13g2_a21oi_1 _18922_ (.A1(_11257_),
    .A2(_11259_),
    .Y(_11278_),
    .B1(_11277_));
 sg13g2_buf_1 _18923_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_11279_));
 sg13g2_nor2_1 _18924_ (.A(_11256_),
    .B(_11278_),
    .Y(_11280_));
 sg13g2_nor2_1 _18925_ (.A(_11279_),
    .B(_11280_),
    .Y(_11281_));
 sg13g2_a221oi_1 _18926_ (.B2(_11278_),
    .C1(_11281_),
    .B1(_11256_),
    .A1(_11252_),
    .Y(_11282_),
    .A2(_11255_));
 sg13g2_a21oi_1 _18927_ (.A1(_11253_),
    .A2(_11254_),
    .Y(_11283_),
    .B1(_11282_));
 sg13g2_o21ai_1 _18928_ (.B1(_11283_),
    .Y(_11284_),
    .A1(_11251_),
    .A2(_11249_));
 sg13g2_o21ai_1 _18929_ (.B1(_11284_),
    .Y(_11285_),
    .A1(_11248_),
    .A2(_11250_));
 sg13g2_nor2_1 _18930_ (.A(_11247_),
    .B(_11285_),
    .Y(_11286_));
 sg13g2_nand2_1 _18931_ (.Y(_11287_),
    .A(_11247_),
    .B(_11285_));
 sg13g2_o21ai_1 _18932_ (.B1(_11287_),
    .Y(_11288_),
    .A1(_11246_),
    .A2(_11286_));
 sg13g2_nor2b_1 _18933_ (.A(_11244_),
    .B_N(_11243_),
    .Y(_11289_));
 sg13g2_a21oi_1 _18934_ (.A1(_11245_),
    .A2(_11288_),
    .Y(_11290_),
    .B1(_11289_));
 sg13g2_buf_1 _18935_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(_11291_));
 sg13g2_nand2_1 _18936_ (.Y(_11292_),
    .A(_11242_),
    .B(_11290_));
 sg13g2_nand2_1 _18937_ (.Y(_11293_),
    .A(_11291_),
    .B(_11292_));
 sg13g2_o21ai_1 _18938_ (.B1(_11293_),
    .Y(_11294_),
    .A1(_11242_),
    .A2(_11290_));
 sg13g2_o21ai_1 _18939_ (.B1(_11294_),
    .Y(_11295_),
    .A1(_11241_),
    .A2(_11239_));
 sg13g2_o21ai_1 _18940_ (.B1(_11295_),
    .Y(_11296_),
    .A1(_11238_),
    .A2(_11240_));
 sg13g2_nor2_1 _18941_ (.A(_11237_),
    .B(_11296_),
    .Y(_11297_));
 sg13g2_nand2_1 _18942_ (.Y(_11298_),
    .A(_11237_),
    .B(_11296_));
 sg13g2_o21ai_1 _18943_ (.B1(_11298_),
    .Y(_11299_),
    .A1(_11236_),
    .A2(_11297_));
 sg13g2_nor2b_1 _18944_ (.A(_11234_),
    .B_N(_11233_),
    .Y(_11300_));
 sg13g2_a21oi_1 _18945_ (.A1(_11235_),
    .A2(_11299_),
    .Y(_11301_),
    .B1(_11300_));
 sg13g2_nand2_1 _18946_ (.Y(_11302_),
    .A(_11232_),
    .B(_11301_));
 sg13g2_nor2_1 _18947_ (.A(_11232_),
    .B(_11301_),
    .Y(_11303_));
 sg13g2_a21oi_1 _18948_ (.A1(_11231_),
    .A2(_11302_),
    .Y(_11304_),
    .B1(_11303_));
 sg13g2_nand2b_1 _18949_ (.Y(_11305_),
    .B(_11228_),
    .A_N(_11229_));
 sg13g2_o21ai_1 _18950_ (.B1(_11305_),
    .Y(_11306_),
    .A1(_11230_),
    .A2(_11304_));
 sg13g2_nand2_1 _18951_ (.Y(_11307_),
    .A(_11227_),
    .B(_11306_));
 sg13g2_nor2_1 _18952_ (.A(_11227_),
    .B(_11306_),
    .Y(_11308_));
 sg13g2_a221oi_1 _18953_ (.B2(_11307_),
    .C1(_11308_),
    .B1(_11226_),
    .A1(_11222_),
    .Y(_11309_),
    .A2(_11225_));
 sg13g2_a21oi_1 _18954_ (.A1(_11223_),
    .A2(_11224_),
    .Y(_11310_),
    .B1(_11309_));
 sg13g2_buf_1 _18955_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .X(_11311_));
 sg13g2_nor2_1 _18956_ (.A(_11221_),
    .B(_11310_),
    .Y(_11312_));
 sg13g2_nor2_1 _18957_ (.A(_11311_),
    .B(_11312_),
    .Y(_11313_));
 sg13g2_a21oi_1 _18958_ (.A1(_11221_),
    .A2(_11310_),
    .Y(_11314_),
    .B1(_11313_));
 sg13g2_nand2b_1 _18959_ (.Y(_11315_),
    .B(_11218_),
    .A_N(_11219_));
 sg13g2_o21ai_1 _18960_ (.B1(_11315_),
    .Y(_11316_),
    .A1(_11220_),
    .A2(_11314_));
 sg13g2_buf_2 _18961_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_11317_));
 sg13g2_o21ai_1 _18962_ (.B1(_11317_),
    .Y(_11318_),
    .A1(_11217_),
    .A2(_11316_));
 sg13g2_nand2_1 _18963_ (.Y(_11319_),
    .A(_11217_),
    .B(_11316_));
 sg13g2_a22oi_1 _18964_ (.Y(_11320_),
    .B1(_11318_),
    .B2(_11319_),
    .A2(_11215_),
    .A1(_11212_));
 sg13g2_a21o_1 _18965_ (.A2(_11214_),
    .A1(_11213_),
    .B1(_11320_),
    .X(_11321_));
 sg13g2_buf_1 _18966_ (.A(_11321_),
    .X(_11322_));
 sg13g2_buf_1 _18967_ (.A(_00017_),
    .X(_11323_));
 sg13g2_or2_1 _18968_ (.X(_11324_),
    .B(_08631_),
    .A(_11323_));
 sg13g2_buf_1 _18969_ (.A(_11324_),
    .X(_11325_));
 sg13g2_nor2_1 _18970_ (.A(_11323_),
    .B(_08629_),
    .Y(_11326_));
 sg13g2_nand2_1 _18971_ (.Y(_11327_),
    .A(_08550_),
    .B(_08562_));
 sg13g2_nor2_1 _18972_ (.A(_11323_),
    .B(_08585_),
    .Y(_11328_));
 sg13g2_nand2_1 _18973_ (.Y(_11329_),
    .A(_08572_),
    .B(_11328_));
 sg13g2_o21ai_1 _18974_ (.B1(_11329_),
    .Y(_11330_),
    .A1(_08672_),
    .A2(_08572_));
 sg13g2_nor2b_1 _18975_ (.A(_11327_),
    .B_N(_11330_),
    .Y(_11331_));
 sg13g2_inv_1 _18976_ (.Y(_11332_),
    .A(_08550_));
 sg13g2_nor2_1 _18977_ (.A(_11332_),
    .B(_08562_),
    .Y(_11333_));
 sg13g2_inv_1 _18978_ (.Y(_11334_),
    .A(_11333_));
 sg13g2_nor2_1 _18979_ (.A(_08672_),
    .B(_11334_),
    .Y(_11335_));
 sg13g2_nor3_1 _18980_ (.A(_08423_),
    .B(net832),
    .C(_00023_),
    .Y(_11336_));
 sg13g2_a22oi_1 _18981_ (.Y(_11337_),
    .B1(_00023_),
    .B2(_08672_),
    .A2(net611),
    .A1(_08435_));
 sg13g2_nand2b_1 _18982_ (.Y(_11338_),
    .B(_11337_),
    .A_N(_11336_));
 sg13g2_nor4_1 _18983_ (.A(_11326_),
    .B(_11331_),
    .C(_11335_),
    .D(_11338_),
    .Y(_11339_));
 sg13g2_o21ai_1 _18984_ (.B1(_11339_),
    .Y(_11340_),
    .A1(_11322_),
    .A2(_11325_));
 sg13g2_buf_1 _18985_ (.A(_11340_),
    .X(_11341_));
 sg13g2_buf_1 _18986_ (.A(_11341_),
    .X(_11342_));
 sg13g2_buf_1 _18987_ (.A(_11342_),
    .X(_11343_));
 sg13g2_buf_1 _18988_ (.A(_11343_),
    .X(_11344_));
 sg13g2_buf_1 _18989_ (.A(_11341_),
    .X(_11345_));
 sg13g2_buf_1 _18990_ (.A(net71),
    .X(_11346_));
 sg13g2_buf_1 _18991_ (.A(_08672_),
    .X(_11347_));
 sg13g2_and2_1 _18992_ (.A(net795),
    .B(_00394_),
    .X(_11348_));
 sg13g2_a21oi_1 _18993_ (.A1(_08494_),
    .A2(net703),
    .Y(_11349_),
    .B1(_11348_));
 sg13g2_nor2_1 _18994_ (.A(net68),
    .B(_11349_),
    .Y(_11350_));
 sg13g2_a21oi_1 _18995_ (.A1(net827),
    .A2(net64),
    .Y(_11351_),
    .B1(_11350_));
 sg13g2_nor2_1 _18996_ (.A(net678),
    .B(_11351_),
    .Y(_01475_));
 sg13g2_buf_1 _18997_ (.A(_08672_),
    .X(_11352_));
 sg13g2_buf_1 _18998_ (.A(net702),
    .X(_11353_));
 sg13g2_buf_1 _18999_ (.A(_00396_),
    .X(_11354_));
 sg13g2_inv_1 _19000_ (.Y(_11355_),
    .A(_08933_));
 sg13g2_inv_1 _19001_ (.Y(_11356_),
    .A(_09762_));
 sg13g2_inv_1 _19002_ (.Y(_11357_),
    .A(_09767_));
 sg13g2_inv_1 _19003_ (.Y(_11358_),
    .A(_09757_));
 sg13g2_nand2_1 _19004_ (.Y(_11359_),
    .A(_08826_),
    .B(_09754_));
 sg13g2_nor2_1 _19005_ (.A(_08826_),
    .B(_09754_),
    .Y(_11360_));
 sg13g2_nor2_1 _19006_ (.A(_08800_),
    .B(_09751_),
    .Y(_11361_));
 sg13g2_a22oi_1 _19007_ (.Y(_11362_),
    .B1(_08800_),
    .B2(_09751_),
    .A2(_09739_),
    .A1(_08748_));
 sg13g2_or3_1 _19008_ (.A(_11360_),
    .B(_11361_),
    .C(_11362_),
    .X(_11363_));
 sg13g2_buf_1 _19009_ (.A(_11363_),
    .X(_11364_));
 sg13g2_nand3_1 _19010_ (.B(_11359_),
    .C(_11364_),
    .A(_11358_),
    .Y(_11365_));
 sg13g2_a21oi_1 _19011_ (.A1(_11359_),
    .A2(_11364_),
    .Y(_11366_),
    .B1(_11358_));
 sg13g2_a21oi_2 _19012_ (.B1(_11366_),
    .Y(_11367_),
    .A2(_11365_),
    .A1(_08846_));
 sg13g2_a221oi_1 _19013_ (.B2(_11357_),
    .C1(_11367_),
    .B1(_08899_),
    .A1(_08902_),
    .Y(_11368_),
    .A2(_11356_));
 sg13g2_buf_1 _19014_ (.A(_11368_),
    .X(_11369_));
 sg13g2_nor2_1 _19015_ (.A(_08902_),
    .B(_11356_),
    .Y(_11370_));
 sg13g2_o21ai_1 _19016_ (.B1(_11370_),
    .Y(_11371_),
    .A1(net824),
    .A2(_09767_));
 sg13g2_o21ai_1 _19017_ (.B1(_11371_),
    .Y(_11372_),
    .A1(_08899_),
    .A2(_11357_));
 sg13g2_o21ai_1 _19018_ (.B1(_09770_),
    .Y(_11373_),
    .A1(_11369_),
    .A2(_11372_));
 sg13g2_nor3_1 _19019_ (.A(_09770_),
    .B(_11369_),
    .C(_11372_),
    .Y(_11374_));
 sg13g2_a21o_1 _19020_ (.A2(_11373_),
    .A1(_11355_),
    .B1(_11374_),
    .X(_11375_));
 sg13g2_buf_1 _19021_ (.A(_11375_),
    .X(_11376_));
 sg13g2_nand2_1 _19022_ (.Y(_11377_),
    .A(_08953_),
    .B(_09774_));
 sg13g2_nand2_1 _19023_ (.Y(_11378_),
    .A(_09777_),
    .B(net823));
 sg13g2_nand2_1 _19024_ (.Y(_11379_),
    .A(_08980_),
    .B(net823));
 sg13g2_nor2_1 _19025_ (.A(_08953_),
    .B(_09774_),
    .Y(_11380_));
 sg13g2_a221oi_1 _19026_ (.B2(_11379_),
    .C1(_11380_),
    .B1(_11378_),
    .A1(_11376_),
    .Y(_11381_),
    .A2(_11377_));
 sg13g2_nand2_1 _19027_ (.Y(_11382_),
    .A(_09777_),
    .B(_09781_));
 sg13g2_nand2_1 _19028_ (.Y(_11383_),
    .A(_08980_),
    .B(_09781_));
 sg13g2_a221oi_1 _19029_ (.B2(_11383_),
    .C1(_11380_),
    .B1(_11382_),
    .A1(_11376_),
    .Y(_11384_),
    .A2(_11377_));
 sg13g2_nand2_1 _19030_ (.Y(_11385_),
    .A(net823),
    .B(_09781_));
 sg13g2_and2_1 _19031_ (.A(_08980_),
    .B(_09777_),
    .X(_11386_));
 sg13g2_o21ai_1 _19032_ (.B1(_11386_),
    .Y(_11387_),
    .A1(net823),
    .A2(_09781_));
 sg13g2_nand2_1 _19033_ (.Y(_11388_),
    .A(_11385_),
    .B(_11387_));
 sg13g2_nor3_1 _19034_ (.A(_11381_),
    .B(_11384_),
    .C(_11388_),
    .Y(_11389_));
 sg13g2_buf_2 _19035_ (.A(_11389_),
    .X(_11390_));
 sg13g2_or2_1 _19036_ (.X(_11391_),
    .B(_11390_),
    .A(_09037_));
 sg13g2_or2_1 _19037_ (.X(_11392_),
    .B(_09037_),
    .A(_09747_));
 sg13g2_a21oi_2 _19038_ (.B1(_11380_),
    .Y(_11393_),
    .A2(_11377_),
    .A1(_11376_));
 sg13g2_a21oi_1 _19039_ (.A1(_09777_),
    .A2(_11393_),
    .Y(_11394_),
    .B1(_08980_));
 sg13g2_nor2_1 _19040_ (.A(_09777_),
    .B(_11393_),
    .Y(_11395_));
 sg13g2_xnor2_1 _19041_ (.Y(_11396_),
    .A(_08997_),
    .B(_09781_));
 sg13g2_o21ai_1 _19042_ (.B1(_11396_),
    .Y(_11397_),
    .A1(_11394_),
    .A2(_11395_));
 sg13g2_or3_1 _19043_ (.A(_11396_),
    .B(_11394_),
    .C(_11395_),
    .X(_11398_));
 sg13g2_xnor2_1 _19044_ (.Y(_11399_),
    .A(_08980_),
    .B(_09777_));
 sg13g2_xnor2_1 _19045_ (.Y(_11400_),
    .A(_11393_),
    .B(_11399_));
 sg13g2_xnor2_1 _19046_ (.Y(_11401_),
    .A(_08953_),
    .B(_09774_));
 sg13g2_xnor2_1 _19047_ (.Y(_11402_),
    .A(_11376_),
    .B(_11401_));
 sg13g2_nor2_1 _19048_ (.A(_11369_),
    .B(_11372_),
    .Y(_11403_));
 sg13g2_xnor2_1 _19049_ (.Y(_11404_),
    .A(_08933_),
    .B(_09770_));
 sg13g2_xnor2_1 _19050_ (.Y(_11405_),
    .A(_11403_),
    .B(_11404_));
 sg13g2_nand2_1 _19051_ (.Y(_11406_),
    .A(_11356_),
    .B(_11367_));
 sg13g2_o21ai_1 _19052_ (.B1(_08902_),
    .Y(_11407_),
    .A1(_11356_),
    .A2(_11367_));
 sg13g2_nand2_1 _19053_ (.Y(_11408_),
    .A(_11406_),
    .B(_11407_));
 sg13g2_xor2_1 _19054_ (.B(_09767_),
    .A(net824),
    .X(_11409_));
 sg13g2_xnor2_1 _19055_ (.Y(_11410_),
    .A(_11408_),
    .B(_11409_));
 sg13g2_xnor2_1 _19056_ (.Y(_11411_),
    .A(_08872_),
    .B(_09762_));
 sg13g2_xnor2_1 _19057_ (.Y(_11412_),
    .A(_11367_),
    .B(_11411_));
 sg13g2_inv_1 _19058_ (.Y(_11413_),
    .A(_11412_));
 sg13g2_nand2_1 _19059_ (.Y(_11414_),
    .A(_11359_),
    .B(_11364_));
 sg13g2_xnor2_1 _19060_ (.Y(_11415_),
    .A(_08846_),
    .B(_09757_));
 sg13g2_xnor2_1 _19061_ (.Y(_11416_),
    .A(_11414_),
    .B(_11415_));
 sg13g2_nor2_1 _19062_ (.A(_11361_),
    .B(_11362_),
    .Y(_11417_));
 sg13g2_xor2_1 _19063_ (.B(_09754_),
    .A(_08826_),
    .X(_11418_));
 sg13g2_xnor2_1 _19064_ (.Y(_11419_),
    .A(_11417_),
    .B(_11418_));
 sg13g2_nand2_1 _19065_ (.Y(_11420_),
    .A(_08748_),
    .B(_09739_));
 sg13g2_xnor2_1 _19066_ (.Y(_11421_),
    .A(_08800_),
    .B(_09751_));
 sg13g2_xnor2_1 _19067_ (.Y(_11422_),
    .A(_11420_),
    .B(_11421_));
 sg13g2_xnor2_1 _19068_ (.Y(_11423_),
    .A(_08748_),
    .B(_09739_));
 sg13g2_nor2_1 _19069_ (.A(_08781_),
    .B(_08784_),
    .Y(_11424_));
 sg13g2_nand4_1 _19070_ (.B(_11422_),
    .C(_11423_),
    .A(_11419_),
    .Y(_11425_),
    .D(_11424_));
 sg13g2_nor4_1 _19071_ (.A(_11410_),
    .B(_11413_),
    .C(_11416_),
    .D(_11425_),
    .Y(_11426_));
 sg13g2_nand3_1 _19072_ (.B(_11405_),
    .C(_11426_),
    .A(_11402_),
    .Y(_11427_));
 sg13g2_or2_1 _19073_ (.X(_11428_),
    .B(_11427_),
    .A(_11400_));
 sg13g2_a21oi_1 _19074_ (.A1(_11397_),
    .A2(_11398_),
    .Y(_11429_),
    .B1(_11428_));
 sg13g2_a21oi_1 _19075_ (.A1(_11391_),
    .A2(_11392_),
    .Y(_11430_),
    .B1(_11429_));
 sg13g2_nand2b_1 _19076_ (.Y(_11431_),
    .B(_09023_),
    .A_N(_09037_));
 sg13g2_a21o_1 _19077_ (.A2(_11431_),
    .A1(_11392_),
    .B1(_11390_),
    .X(_11432_));
 sg13g2_o21ai_1 _19078_ (.B1(_11432_),
    .Y(_11433_),
    .A1(_11429_),
    .A2(_11431_));
 sg13g2_nand2b_1 _19079_ (.Y(_11434_),
    .B(_09023_),
    .A_N(_09747_));
 sg13g2_nor2_1 _19080_ (.A(_09037_),
    .B(_11434_),
    .Y(_11435_));
 sg13g2_nor3_1 _19081_ (.A(_11429_),
    .B(_11390_),
    .C(_11434_),
    .Y(_11436_));
 sg13g2_nor4_1 _19082_ (.A(_11430_),
    .B(_11433_),
    .C(_11435_),
    .D(_11436_),
    .Y(_11437_));
 sg13g2_buf_1 _19083_ (.A(_11437_),
    .X(_11438_));
 sg13g2_buf_1 _19084_ (.A(_11438_),
    .X(_11439_));
 sg13g2_buf_1 _19085_ (.A(net308),
    .X(_11440_));
 sg13g2_nor2_1 _19086_ (.A(_08604_),
    .B(_08593_),
    .Y(_11441_));
 sg13g2_nand3b_1 _19087_ (.B(_11441_),
    .C(_08623_),
    .Y(_11442_),
    .A_N(net302));
 sg13g2_buf_1 _19088_ (.A(_11442_),
    .X(_11443_));
 sg13g2_nor2_1 _19089_ (.A(_00395_),
    .B(_11443_),
    .Y(_11444_));
 sg13g2_nand2_1 _19090_ (.Y(_11445_),
    .A(_08521_),
    .B(_11444_));
 sg13g2_nor3_1 _19091_ (.A(_11354_),
    .B(_00397_),
    .C(_11445_),
    .Y(_11446_));
 sg13g2_buf_1 _19092_ (.A(_11440_),
    .X(_11447_));
 sg13g2_and2_1 _19093_ (.A(_00395_),
    .B(net302),
    .X(_11448_));
 sg13g2_or2_1 _19094_ (.X(_11449_),
    .B(_11448_),
    .A(_11444_));
 sg13g2_nor3_1 _19095_ (.A(_08604_),
    .B(_08622_),
    .C(net302),
    .Y(_11450_));
 sg13g2_a21o_1 _19096_ (.A2(net302),
    .A1(_08604_),
    .B1(_11450_),
    .X(_11451_));
 sg13g2_o21ai_1 _19097_ (.B1(_08604_),
    .Y(_11452_),
    .A1(net793),
    .A2(net791));
 sg13g2_nand2_1 _19098_ (.Y(_11453_),
    .A(_08589_),
    .B(_11452_));
 sg13g2_a22oi_1 _19099_ (.Y(_11454_),
    .B1(_11453_),
    .B2(net302),
    .A2(_11451_),
    .A1(net827));
 sg13g2_nand2b_1 _19100_ (.Y(_11455_),
    .B(_08593_),
    .A_N(_11454_));
 sg13g2_nand3b_1 _19101_ (.B(net302),
    .C(_11455_),
    .Y(_11456_),
    .A_N(_08513_));
 sg13g2_buf_1 _19102_ (.A(_11456_),
    .X(_11457_));
 sg13g2_a221oi_1 _19103_ (.B2(_11448_),
    .C1(\rbzero.wall_tracer.mapX[6] ),
    .B1(_11457_),
    .A1(_08521_),
    .Y(_11458_),
    .A2(_11449_));
 sg13g2_nand2b_1 _19104_ (.Y(_11459_),
    .B(_11354_),
    .A_N(_11458_));
 sg13g2_nand2b_1 _19105_ (.Y(_11460_),
    .B(_11459_),
    .A_N(\rbzero.wall_tracer.mapX[7] ));
 sg13g2_nand3_1 _19106_ (.B(net294),
    .C(_11460_),
    .A(_00397_),
    .Y(_11461_));
 sg13g2_nor2b_1 _19107_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B_N(_11461_),
    .Y(_11462_));
 sg13g2_nand2b_1 _19108_ (.Y(_11463_),
    .B(_11462_),
    .A_N(_11446_));
 sg13g2_inv_1 _19109_ (.Y(_11464_),
    .A(\rbzero.wall_tracer.mapX[9] ));
 sg13g2_a21oi_1 _19110_ (.A1(_11464_),
    .A2(net294),
    .Y(_11465_),
    .B1(_11446_));
 sg13g2_a21oi_1 _19111_ (.A1(_00398_),
    .A2(_11463_),
    .Y(_11466_),
    .B1(_11465_));
 sg13g2_nor2_1 _19112_ (.A(net638),
    .B(_11466_),
    .Y(_11467_));
 sg13g2_o21ai_1 _19113_ (.B1(\rbzero.wall_tracer.mapX[10] ),
    .Y(_11468_),
    .A1(net64),
    .A2(_11467_));
 sg13g2_inv_1 _19114_ (.Y(_11469_),
    .A(\rbzero.wall_tracer.mapX[10] ));
 sg13g2_buf_1 _19115_ (.A(net795),
    .X(_11470_));
 sg13g2_buf_1 _19116_ (.A(net701),
    .X(_11471_));
 sg13g2_inv_1 _19117_ (.Y(_11472_),
    .A(_11341_));
 sg13g2_nand4_1 _19118_ (.B(net637),
    .C(_11472_),
    .A(_11469_),
    .Y(_11473_),
    .D(_11466_));
 sg13g2_a21oi_1 _19119_ (.A1(_11468_),
    .A2(_11473_),
    .Y(_01476_),
    .B1(net682));
 sg13g2_xnor2_1 _19120_ (.Y(_11474_),
    .A(_00394_),
    .B(net294));
 sg13g2_nor2_1 _19121_ (.A(net793),
    .B(net702),
    .Y(_11475_));
 sg13g2_a22oi_1 _19122_ (.Y(_11476_),
    .B1(_11474_),
    .B2(_11475_),
    .A2(net703),
    .A1(_08511_));
 sg13g2_or2_1 _19123_ (.X(_11477_),
    .B(_11476_),
    .A(net68));
 sg13g2_buf_1 _19124_ (.A(net69),
    .X(_11478_));
 sg13g2_nor2_1 _19125_ (.A(net703),
    .B(_11474_),
    .Y(_11479_));
 sg13g2_o21ai_1 _19126_ (.B1(net793),
    .Y(_11480_),
    .A1(net63),
    .A2(_11479_));
 sg13g2_a21oi_1 _19127_ (.A1(_11477_),
    .A2(_11480_),
    .Y(_01477_),
    .B1(net682));
 sg13g2_nor2_1 _19128_ (.A(_08495_),
    .B(_08510_),
    .Y(_11481_));
 sg13g2_nor2b_1 _19129_ (.A(net294),
    .B_N(_08510_),
    .Y(_11482_));
 sg13g2_a22oi_1 _19130_ (.Y(_11483_),
    .B1(_11482_),
    .B2(_08495_),
    .A2(net294),
    .A1(_11481_));
 sg13g2_nor3_1 _19131_ (.A(_08558_),
    .B(net702),
    .C(_11483_),
    .Y(_11484_));
 sg13g2_a21o_1 _19132_ (.A2(net703),
    .A1(_08501_),
    .B1(_11484_),
    .X(_11485_));
 sg13g2_buf_1 _19133_ (.A(net795),
    .X(_11486_));
 sg13g2_a21o_1 _19134_ (.A2(_11483_),
    .A1(net700),
    .B1(net69),
    .X(_11487_));
 sg13g2_a22oi_1 _19135_ (.Y(_11488_),
    .B1(_11487_),
    .B2(net791),
    .A2(_11485_),
    .A1(_11472_));
 sg13g2_nor2_1 _19136_ (.A(net678),
    .B(_11488_),
    .Y(_01478_));
 sg13g2_mux2_1 _19137_ (.A0(_08623_),
    .A1(_08551_),
    .S(net294),
    .X(_11489_));
 sg13g2_xor2_1 _19138_ (.B(_11489_),
    .A(_08604_),
    .X(_11490_));
 sg13g2_nor2_1 _19139_ (.A(_11352_),
    .B(_11490_),
    .Y(_11491_));
 sg13g2_a21oi_1 _19140_ (.A1(_08483_),
    .A2(_11352_),
    .Y(_11492_),
    .B1(_11491_));
 sg13g2_nor2_1 _19141_ (.A(net68),
    .B(_11492_),
    .Y(_11493_));
 sg13g2_a21oi_1 _19142_ (.A1(_08482_),
    .A2(net64),
    .Y(_11494_),
    .B1(_11493_));
 sg13g2_nor2_1 _19143_ (.A(_09051_),
    .B(_11494_),
    .Y(_01479_));
 sg13g2_xnor2_1 _19144_ (.Y(_11495_),
    .A(_08593_),
    .B(net294));
 sg13g2_xnor2_1 _19145_ (.Y(_11496_),
    .A(_11454_),
    .B(_11495_));
 sg13g2_nor2b_1 _19146_ (.A(net795),
    .B_N(_08514_),
    .Y(_11497_));
 sg13g2_a21oi_1 _19147_ (.A1(net701),
    .A2(_11496_),
    .Y(_11498_),
    .B1(_11497_));
 sg13g2_nor2_1 _19148_ (.A(net68),
    .B(_11498_),
    .Y(_11499_));
 sg13g2_a21oi_1 _19149_ (.A1(_08513_),
    .A2(net64),
    .Y(_11500_),
    .B1(_11499_));
 sg13g2_nor2_1 _19150_ (.A(_09051_),
    .B(_11500_),
    .Y(_01480_));
 sg13g2_nand2_1 _19151_ (.Y(_11501_),
    .A(_11443_),
    .B(_11457_));
 sg13g2_nor2_1 _19152_ (.A(_08521_),
    .B(net702),
    .Y(_11502_));
 sg13g2_a22oi_1 _19153_ (.Y(_11503_),
    .B1(_11501_),
    .B2(_11502_),
    .A2(net703),
    .A1(_08522_));
 sg13g2_or2_1 _19154_ (.X(_11504_),
    .B(_11503_),
    .A(net68));
 sg13g2_nor2_1 _19155_ (.A(net703),
    .B(_11501_),
    .Y(_11505_));
 sg13g2_o21ai_1 _19156_ (.B1(_08521_),
    .Y(_11506_),
    .A1(net63),
    .A2(_11505_));
 sg13g2_a21oi_1 _19157_ (.A1(_11504_),
    .A2(_11506_),
    .Y(_01481_),
    .B1(net682));
 sg13g2_buf_1 _19158_ (.A(net729),
    .X(_11507_));
 sg13g2_mux2_1 _19159_ (.A0(_11457_),
    .A1(_11443_),
    .S(_08521_),
    .X(_11508_));
 sg13g2_xnor2_1 _19160_ (.Y(_11509_),
    .A(_00395_),
    .B(_11508_));
 sg13g2_nor3_1 _19161_ (.A(net638),
    .B(net69),
    .C(_11509_),
    .Y(_11510_));
 sg13g2_a21oi_1 _19162_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(net64),
    .Y(_11511_),
    .B1(_11510_));
 sg13g2_nor2_1 _19163_ (.A(net636),
    .B(_11511_),
    .Y(_01482_));
 sg13g2_nand2_1 _19164_ (.Y(_11512_),
    .A(net294),
    .B(_11458_));
 sg13g2_nand2_1 _19165_ (.Y(_11513_),
    .A(_11445_),
    .B(_11512_));
 sg13g2_xor2_1 _19166_ (.B(_11513_),
    .A(_11354_),
    .X(_11514_));
 sg13g2_nor3_1 _19167_ (.A(net638),
    .B(net69),
    .C(_11514_),
    .Y(_11515_));
 sg13g2_a21oi_1 _19168_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(net64),
    .Y(_11516_),
    .B1(_11515_));
 sg13g2_nor2_1 _19169_ (.A(net636),
    .B(_11516_),
    .Y(_01483_));
 sg13g2_inv_1 _19170_ (.Y(_11517_),
    .A(_11460_));
 sg13g2_nor2_1 _19171_ (.A(_11354_),
    .B(_11445_),
    .Y(_11518_));
 sg13g2_a21oi_1 _19172_ (.A1(_11447_),
    .A2(_11517_),
    .Y(_11519_),
    .B1(_11518_));
 sg13g2_xnor2_1 _19173_ (.Y(_11520_),
    .A(_00397_),
    .B(_11519_));
 sg13g2_nor3_1 _19174_ (.A(net638),
    .B(net69),
    .C(_11520_),
    .Y(_11521_));
 sg13g2_a21oi_1 _19175_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(net64),
    .Y(_11522_),
    .B1(_11521_));
 sg13g2_nor2_1 _19176_ (.A(_11507_),
    .B(_11522_),
    .Y(_01484_));
 sg13g2_a21oi_1 _19177_ (.A1(_11447_),
    .A2(_11462_),
    .Y(_11523_),
    .B1(_11446_));
 sg13g2_xnor2_1 _19178_ (.Y(_11524_),
    .A(_00398_),
    .B(_11523_));
 sg13g2_nor3_1 _19179_ (.A(net638),
    .B(net69),
    .C(_11524_),
    .Y(_11525_));
 sg13g2_a21oi_1 _19180_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(net64),
    .Y(_11526_),
    .B1(_11525_));
 sg13g2_nor2_1 _19181_ (.A(_11507_),
    .B(_11526_),
    .Y(_01485_));
 sg13g2_buf_1 _19182_ (.A(_08675_),
    .X(_11527_));
 sg13g2_nand2b_1 _19183_ (.Y(_11528_),
    .B(_11322_),
    .A_N(_08673_));
 sg13g2_and2_1 _19184_ (.A(_11339_),
    .B(_11528_),
    .X(_11529_));
 sg13g2_buf_2 _19185_ (.A(_11529_),
    .X(_11530_));
 sg13g2_buf_1 _19186_ (.A(_11530_),
    .X(_11531_));
 sg13g2_nor2_1 _19187_ (.A(net790),
    .B(net67),
    .Y(_11532_));
 sg13g2_and2_1 _19188_ (.A(net795),
    .B(_00393_),
    .X(_11533_));
 sg13g2_a21oi_1 _19189_ (.A1(_08485_),
    .A2(net703),
    .Y(_11534_),
    .B1(_11533_));
 sg13g2_and2_1 _19190_ (.A(net67),
    .B(_11534_),
    .X(_11535_));
 sg13g2_nor3_1 _19191_ (.A(net635),
    .B(_11532_),
    .C(_11535_),
    .Y(_01486_));
 sg13g2_inv_1 _19192_ (.Y(_11536_),
    .A(_09811_));
 sg13g2_inv_1 _19193_ (.Y(_11537_),
    .A(_09802_));
 sg13g2_nand2_1 _19194_ (.Y(_11538_),
    .A(_09805_),
    .B(_09271_));
 sg13g2_nand2_1 _19195_ (.Y(_11539_),
    .A(_09247_),
    .B(_09271_));
 sg13g2_inv_1 _19196_ (.Y(_11540_),
    .A(\rbzero.wall_tracer.rayAddendY[2] ));
 sg13g2_and2_1 _19197_ (.A(_09156_),
    .B(_09792_),
    .X(_11541_));
 sg13g2_buf_1 _19198_ (.A(_11541_),
    .X(_11542_));
 sg13g2_nor2_1 _19199_ (.A(_09156_),
    .B(_09792_),
    .Y(_11543_));
 sg13g2_nor2_1 _19200_ (.A(_09132_),
    .B(_09790_),
    .Y(_11544_));
 sg13g2_a22oi_1 _19201_ (.Y(_11545_),
    .B1(_09132_),
    .B2(_09790_),
    .A2(_09783_),
    .A1(_09083_));
 sg13g2_nor3_1 _19202_ (.A(_11543_),
    .B(_11544_),
    .C(_11545_),
    .Y(_11546_));
 sg13g2_nor3_1 _19203_ (.A(_09795_),
    .B(_11542_),
    .C(_11546_),
    .Y(_11547_));
 sg13g2_o21ai_1 _19204_ (.B1(_09795_),
    .Y(_11548_),
    .A1(_11542_),
    .A2(_11546_));
 sg13g2_o21ai_1 _19205_ (.B1(_11548_),
    .Y(_11549_),
    .A1(_11540_),
    .A2(_11547_));
 sg13g2_buf_1 _19206_ (.A(_11549_),
    .X(_11550_));
 sg13g2_a21o_1 _19207_ (.A2(_11550_),
    .A1(_09798_),
    .B1(net818),
    .X(_11551_));
 sg13g2_or2_1 _19208_ (.X(_11552_),
    .B(_11550_),
    .A(_09798_));
 sg13g2_a22oi_1 _19209_ (.Y(_11553_),
    .B1(_11551_),
    .B2(_11552_),
    .A2(_09802_),
    .A1(net817));
 sg13g2_a221oi_1 _19210_ (.B2(_11539_),
    .C1(_11553_),
    .B1(_11538_),
    .A1(_09208_),
    .Y(_11554_),
    .A2(_11537_));
 sg13g2_nand2_1 _19211_ (.Y(_11555_),
    .A(_09805_),
    .B(_09807_));
 sg13g2_nand2_1 _19212_ (.Y(_11556_),
    .A(_09248_),
    .B(_09807_));
 sg13g2_a221oi_1 _19213_ (.B2(_11556_),
    .C1(_11553_),
    .B1(_11555_),
    .A1(_09208_),
    .Y(_11557_),
    .A2(_11537_));
 sg13g2_nand2_1 _19214_ (.Y(_11558_),
    .A(_09271_),
    .B(_09807_));
 sg13g2_and2_1 _19215_ (.A(_09247_),
    .B(_09805_),
    .X(_11559_));
 sg13g2_o21ai_1 _19216_ (.B1(_11559_),
    .Y(_11560_),
    .A1(_09271_),
    .A2(_09807_));
 sg13g2_nand2_1 _19217_ (.Y(_11561_),
    .A(_11558_),
    .B(_11560_));
 sg13g2_nor3_2 _19218_ (.A(_11554_),
    .B(_11557_),
    .C(_11561_),
    .Y(_11562_));
 sg13g2_o21ai_1 _19219_ (.B1(_09320_),
    .Y(_11563_),
    .A1(_11536_),
    .A2(_11562_));
 sg13g2_nand2_1 _19220_ (.Y(_11564_),
    .A(_11536_),
    .B(_11562_));
 sg13g2_xnor2_1 _19221_ (.Y(_11565_),
    .A(_09319_),
    .B(_09813_));
 sg13g2_a21oi_1 _19222_ (.A1(_11563_),
    .A2(_11564_),
    .Y(_11566_),
    .B1(_11565_));
 sg13g2_and3_1 _19223_ (.X(_11567_),
    .A(_11565_),
    .B(_11563_),
    .C(_11564_));
 sg13g2_xnor2_1 _19224_ (.Y(_11568_),
    .A(_09297_),
    .B(_09811_));
 sg13g2_xnor2_1 _19225_ (.Y(_11569_),
    .A(_11562_),
    .B(_11568_));
 sg13g2_inv_1 _19226_ (.Y(_11570_),
    .A(_11569_));
 sg13g2_inv_1 _19227_ (.Y(_11571_),
    .A(_09248_));
 sg13g2_a21oi_1 _19228_ (.A1(_09798_),
    .A2(_11550_),
    .Y(_11572_),
    .B1(net818));
 sg13g2_nor2_1 _19229_ (.A(_09798_),
    .B(_11550_),
    .Y(_11573_));
 sg13g2_nand2_1 _19230_ (.Y(_11574_),
    .A(net817),
    .B(_09802_));
 sg13g2_o21ai_1 _19231_ (.B1(_11574_),
    .Y(_11575_),
    .A1(_11572_),
    .A2(_11573_));
 sg13g2_nand2_1 _19232_ (.Y(_11576_),
    .A(_09208_),
    .B(_11537_));
 sg13g2_nand3_1 _19233_ (.B(_11575_),
    .C(_11576_),
    .A(_09805_),
    .Y(_11577_));
 sg13g2_a21oi_1 _19234_ (.A1(_11575_),
    .A2(_11576_),
    .Y(_11578_),
    .B1(_09805_));
 sg13g2_a21oi_1 _19235_ (.A1(_11571_),
    .A2(_11577_),
    .Y(_11579_),
    .B1(_11578_));
 sg13g2_xnor2_1 _19236_ (.Y(_11580_),
    .A(_09271_),
    .B(_09807_));
 sg13g2_xnor2_1 _19237_ (.Y(_11581_),
    .A(_11579_),
    .B(_11580_));
 sg13g2_nand2_1 _19238_ (.Y(_11582_),
    .A(_11575_),
    .B(_11576_));
 sg13g2_xnor2_1 _19239_ (.Y(_11583_),
    .A(net761),
    .B(_09805_));
 sg13g2_xnor2_1 _19240_ (.Y(_11584_),
    .A(_11582_),
    .B(_11583_));
 sg13g2_nor2_1 _19241_ (.A(_11572_),
    .B(_11573_),
    .Y(_11585_));
 sg13g2_xnor2_1 _19242_ (.Y(_11586_),
    .A(_09207_),
    .B(_09802_));
 sg13g2_xnor2_1 _19243_ (.Y(_11587_),
    .A(_11585_),
    .B(_11586_));
 sg13g2_xnor2_1 _19244_ (.Y(_11588_),
    .A(_09190_),
    .B(_09798_));
 sg13g2_xnor2_1 _19245_ (.Y(_11589_),
    .A(_11550_),
    .B(_11588_));
 sg13g2_nor2_1 _19246_ (.A(_11542_),
    .B(_11546_),
    .Y(_11590_));
 sg13g2_xor2_1 _19247_ (.B(_09795_),
    .A(net819),
    .X(_11591_));
 sg13g2_xnor2_1 _19248_ (.Y(_11592_),
    .A(_11590_),
    .B(_11591_));
 sg13g2_nor2_1 _19249_ (.A(_11544_),
    .B(_11545_),
    .Y(_11593_));
 sg13g2_xor2_1 _19250_ (.B(_09792_),
    .A(_09156_),
    .X(_11594_));
 sg13g2_xnor2_1 _19251_ (.Y(_11595_),
    .A(_11593_),
    .B(_11594_));
 sg13g2_nand2_1 _19252_ (.Y(_11596_),
    .A(_09083_),
    .B(_09783_));
 sg13g2_xor2_1 _19253_ (.B(_09790_),
    .A(_09132_),
    .X(_11597_));
 sg13g2_xnor2_1 _19254_ (.Y(_11598_),
    .A(_11596_),
    .B(_11597_));
 sg13g2_xor2_1 _19255_ (.B(_09783_),
    .A(_09083_),
    .X(_11599_));
 sg13g2_nor4_1 _19256_ (.A(_09115_),
    .B(_09118_),
    .C(_11598_),
    .D(_11599_),
    .Y(_11600_));
 sg13g2_nand2_1 _19257_ (.Y(_11601_),
    .A(_11595_),
    .B(_11600_));
 sg13g2_nor4_1 _19258_ (.A(_11587_),
    .B(_11589_),
    .C(_11592_),
    .D(_11601_),
    .Y(_11602_));
 sg13g2_nand3b_1 _19259_ (.B(_11584_),
    .C(_11602_),
    .Y(_11603_),
    .A_N(_11581_));
 sg13g2_or4_1 _19260_ (.A(_11566_),
    .B(_11567_),
    .C(_11570_),
    .D(_11603_),
    .X(_11604_));
 sg13g2_buf_1 _19261_ (.A(_11604_),
    .X(_11605_));
 sg13g2_inv_1 _19262_ (.Y(_11606_),
    .A(_09786_));
 sg13g2_nand2_1 _19263_ (.Y(_11607_),
    .A(_09343_),
    .B(_11606_));
 sg13g2_inv_1 _19264_ (.Y(_11608_),
    .A(_09813_));
 sg13g2_a221oi_1 _19265_ (.B2(_11608_),
    .C1(_11562_),
    .B1(_09344_),
    .A1(_09320_),
    .Y(_11609_),
    .A2(_11536_));
 sg13g2_buf_1 _19266_ (.A(_11609_),
    .X(_11610_));
 sg13g2_nor2_1 _19267_ (.A(_09320_),
    .B(_11536_),
    .Y(_11611_));
 sg13g2_o21ai_1 _19268_ (.B1(_11611_),
    .Y(_11612_),
    .A1(_09319_),
    .A2(_09813_));
 sg13g2_o21ai_1 _19269_ (.B1(_11612_),
    .Y(_11613_),
    .A1(_09344_),
    .A2(_11608_));
 sg13g2_buf_1 _19270_ (.A(_11613_),
    .X(_11614_));
 sg13g2_nor2_2 _19271_ (.A(_11610_),
    .B(_11614_),
    .Y(_11615_));
 sg13g2_nor2_1 _19272_ (.A(_11607_),
    .B(_11615_),
    .Y(_11616_));
 sg13g2_nor2_1 _19273_ (.A(_09357_),
    .B(_11607_),
    .Y(_11617_));
 sg13g2_a21oi_1 _19274_ (.A1(_11605_),
    .A2(_11616_),
    .Y(_11618_),
    .B1(_11617_));
 sg13g2_nor2_1 _19275_ (.A(_09357_),
    .B(_11615_),
    .Y(_11619_));
 sg13g2_nor2_1 _19276_ (.A(_09786_),
    .B(_09357_),
    .Y(_11620_));
 sg13g2_o21ai_1 _19277_ (.B1(_11605_),
    .Y(_11621_),
    .A1(_11619_),
    .A2(_11620_));
 sg13g2_nor2b_1 _19278_ (.A(_09357_),
    .B_N(_09343_),
    .Y(_11622_));
 sg13g2_o21ai_1 _19279_ (.B1(_11620_),
    .Y(_11623_),
    .A1(_11610_),
    .A2(_11614_));
 sg13g2_o21ai_1 _19280_ (.B1(_11622_),
    .Y(_11624_),
    .A1(_11610_),
    .A2(_11614_));
 sg13g2_nand2_1 _19281_ (.Y(_11625_),
    .A(_11623_),
    .B(_11624_));
 sg13g2_a21oi_1 _19282_ (.A1(_11605_),
    .A2(_11622_),
    .Y(_11626_),
    .B1(_11625_));
 sg13g2_nand3_1 _19283_ (.B(_11621_),
    .C(_11626_),
    .A(_11618_),
    .Y(_11627_));
 sg13g2_buf_2 _19284_ (.A(_11627_),
    .X(_11628_));
 sg13g2_buf_1 _19285_ (.A(_11628_),
    .X(_11629_));
 sg13g2_or2_1 _19286_ (.X(_11630_),
    .B(net794),
    .A(net790));
 sg13g2_a21o_1 _19287_ (.A2(_11630_),
    .A1(_08614_),
    .B1(net792),
    .X(_11631_));
 sg13g2_buf_1 _19288_ (.A(_11631_),
    .X(_11632_));
 sg13g2_and2_1 _19289_ (.A(_08619_),
    .B(_11632_),
    .X(_11633_));
 sg13g2_or4_1 _19290_ (.A(_08491_),
    .B(_08497_),
    .C(net314),
    .D(_11633_),
    .X(_11634_));
 sg13g2_buf_1 _19291_ (.A(_11634_),
    .X(_11635_));
 sg13g2_a21oi_1 _19292_ (.A1(_08591_),
    .A2(_08619_),
    .Y(_11636_),
    .B1(_11635_));
 sg13g2_inv_1 _19293_ (.Y(_11637_),
    .A(\rbzero.wall_tracer.mapY[6] ));
 sg13g2_inv_1 _19294_ (.Y(_11638_),
    .A(_11629_));
 sg13g2_nand2_1 _19295_ (.Y(_11639_),
    .A(_08590_),
    .B(net794));
 sg13g2_nor3_2 _19296_ (.A(_08614_),
    .B(_11638_),
    .C(_11639_),
    .Y(_11640_));
 sg13g2_nand3_1 _19297_ (.B(_08497_),
    .C(_11640_),
    .A(net789),
    .Y(_11641_));
 sg13g2_nor3_1 _19298_ (.A(_11637_),
    .B(_08619_),
    .C(_11641_),
    .Y(_11642_));
 sg13g2_and3_1 _19299_ (.X(_11643_),
    .A(_08524_),
    .B(_08526_),
    .C(_11642_));
 sg13g2_a22oi_1 _19300_ (.Y(_11644_),
    .B1(_11643_),
    .B2(_08525_),
    .A2(_11636_),
    .A1(_08527_));
 sg13g2_nand2_1 _19301_ (.Y(_11645_),
    .A(net701),
    .B(_11644_));
 sg13g2_nand2_1 _19302_ (.Y(_11646_),
    .A(_11531_),
    .B(_11645_));
 sg13g2_nand2_2 _19303_ (.Y(_11647_),
    .A(net795),
    .B(_11530_));
 sg13g2_nor3_1 _19304_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_11644_),
    .C(_11647_),
    .Y(_11648_));
 sg13g2_a21oi_1 _19305_ (.A1(\rbzero.wall_tracer.mapY[10] ),
    .A2(_11646_),
    .Y(_11649_),
    .B1(_11648_));
 sg13g2_nor2_1 _19306_ (.A(net636),
    .B(_11649_),
    .Y(_01487_));
 sg13g2_xor2_1 _19307_ (.B(net314),
    .A(_00393_),
    .X(_11650_));
 sg13g2_nand3b_1 _19308_ (.B(net795),
    .C(_11650_),
    .Y(_11651_),
    .A_N(net794));
 sg13g2_o21ai_1 _19309_ (.B1(_11651_),
    .Y(_11652_),
    .A1(_09952_),
    .A2(net700));
 sg13g2_o21ai_1 _19310_ (.B1(net67),
    .Y(_11653_),
    .A1(net638),
    .A2(_11650_));
 sg13g2_a22oi_1 _19311_ (.Y(_11654_),
    .B1(_11653_),
    .B2(net794),
    .A2(_11652_),
    .A1(net67));
 sg13g2_nor2_1 _19312_ (.A(net636),
    .B(_11654_),
    .Y(_01488_));
 sg13g2_mux2_1 _19313_ (.A0(_11630_),
    .A1(_11639_),
    .S(net314),
    .X(_11655_));
 sg13g2_xnor2_1 _19314_ (.Y(_11656_),
    .A(_08614_),
    .B(_11655_));
 sg13g2_nor2_1 _19315_ (.A(_08518_),
    .B(net701),
    .Y(_11657_));
 sg13g2_a21oi_1 _19316_ (.A1(net700),
    .A2(_11656_),
    .Y(_11658_),
    .B1(_11657_));
 sg13g2_nand2_1 _19317_ (.Y(_11659_),
    .A(net67),
    .B(_11658_));
 sg13g2_nand2b_1 _19318_ (.Y(_11660_),
    .B(_08517_),
    .A_N(net67));
 sg13g2_a21oi_1 _19319_ (.A1(_11659_),
    .A2(_11660_),
    .Y(_01489_),
    .B1(net682));
 sg13g2_inv_1 _19320_ (.Y(_11661_),
    .A(_11640_));
 sg13g2_o21ai_1 _19321_ (.B1(_11661_),
    .Y(_11662_),
    .A1(net314),
    .A2(_11632_));
 sg13g2_o21ai_1 _19322_ (.B1(_11530_),
    .Y(_11663_),
    .A1(net638),
    .A2(_11662_));
 sg13g2_nor2_1 _19323_ (.A(net789),
    .B(net702),
    .Y(_11664_));
 sg13g2_a22oi_1 _19324_ (.Y(_11665_),
    .B1(_11662_),
    .B2(_11664_),
    .A2(net702),
    .A1(_08489_));
 sg13g2_nor2b_1 _19325_ (.A(_11665_),
    .B_N(_11530_),
    .Y(_11666_));
 sg13g2_a21oi_1 _19326_ (.A1(net789),
    .A2(_11663_),
    .Y(_11667_),
    .B1(_11666_));
 sg13g2_nor2_1 _19327_ (.A(net636),
    .B(_11667_),
    .Y(_01490_));
 sg13g2_o21ai_1 _19328_ (.B1(_08603_),
    .Y(_11668_),
    .A1(net314),
    .A2(_11632_));
 sg13g2_o21ai_1 _19329_ (.B1(_11668_),
    .Y(_11669_),
    .A1(_08603_),
    .A2(_11640_));
 sg13g2_xnor2_1 _19330_ (.Y(_11670_),
    .A(_08619_),
    .B(_11669_));
 sg13g2_nand2_1 _19331_ (.Y(_11671_),
    .A(net795),
    .B(_11670_));
 sg13g2_o21ai_1 _19332_ (.B1(_11671_),
    .Y(_11672_),
    .A1(_08492_),
    .A2(net701));
 sg13g2_mux2_1 _19333_ (.A0(_08592_),
    .A1(_11672_),
    .S(net67),
    .X(_11673_));
 sg13g2_nor2_1 _19334_ (.A(net636),
    .B(_11673_),
    .Y(_01491_));
 sg13g2_o21ai_1 _19335_ (.B1(_08619_),
    .Y(_11674_),
    .A1(net789),
    .A2(_11632_));
 sg13g2_nand2_1 _19336_ (.Y(_11675_),
    .A(_08592_),
    .B(_11674_));
 sg13g2_nand3b_1 _19337_ (.B(_11640_),
    .C(net789),
    .Y(_11676_),
    .A_N(_08619_));
 sg13g2_o21ai_1 _19338_ (.B1(_11676_),
    .Y(_11677_),
    .A1(net314),
    .A2(_11675_));
 sg13g2_o21ai_1 _19339_ (.B1(_11530_),
    .Y(_11678_),
    .A1(net703),
    .A2(_11677_));
 sg13g2_nor2_1 _19340_ (.A(_08497_),
    .B(net702),
    .Y(_11679_));
 sg13g2_a22oi_1 _19341_ (.Y(_11680_),
    .B1(_11677_),
    .B2(_11679_),
    .A2(net702),
    .A1(_08498_));
 sg13g2_nor2b_1 _19342_ (.A(_11680_),
    .B_N(_11530_),
    .Y(_11681_));
 sg13g2_a21oi_1 _19343_ (.A1(_08497_),
    .A2(_11678_),
    .Y(_11682_),
    .B1(_11681_));
 sg13g2_nor2_1 _19344_ (.A(net636),
    .B(_11682_),
    .Y(_01492_));
 sg13g2_a21oi_1 _19345_ (.A1(_11635_),
    .A2(_11641_),
    .Y(_11683_),
    .B1(_08619_));
 sg13g2_nor2_1 _19346_ (.A(_08591_),
    .B(_11635_),
    .Y(_11684_));
 sg13g2_nor2_1 _19347_ (.A(_11683_),
    .B(_11684_),
    .Y(_11685_));
 sg13g2_nand2_1 _19348_ (.Y(_11686_),
    .A(net701),
    .B(_11685_));
 sg13g2_a21oi_1 _19349_ (.A1(_11530_),
    .A2(_11686_),
    .Y(_11687_),
    .B1(_11637_));
 sg13g2_nor3_1 _19350_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_11647_),
    .C(_11685_),
    .Y(_11688_));
 sg13g2_nor2_1 _19351_ (.A(_11687_),
    .B(_11688_),
    .Y(_11689_));
 sg13g2_nor2_1 _19352_ (.A(net636),
    .B(_11689_),
    .Y(_01493_));
 sg13g2_buf_1 _19353_ (.A(net729),
    .X(_11690_));
 sg13g2_nand2_1 _19354_ (.Y(_11691_),
    .A(_11637_),
    .B(_11636_));
 sg13g2_nor2b_1 _19355_ (.A(_11642_),
    .B_N(_11691_),
    .Y(_11692_));
 sg13g2_nand2_1 _19356_ (.Y(_11693_),
    .A(net701),
    .B(_11692_));
 sg13g2_nand2_1 _19357_ (.Y(_11694_),
    .A(_11531_),
    .B(_11693_));
 sg13g2_nor3_1 _19358_ (.A(_08524_),
    .B(_11647_),
    .C(_11692_),
    .Y(_11695_));
 sg13g2_a21oi_1 _19359_ (.A1(_08524_),
    .A2(_11694_),
    .Y(_11696_),
    .B1(_11695_));
 sg13g2_nor2_1 _19360_ (.A(net634),
    .B(_11696_),
    .Y(_01494_));
 sg13g2_nand2_1 _19361_ (.Y(_11697_),
    .A(_08524_),
    .B(_11642_));
 sg13g2_o21ai_1 _19362_ (.B1(_11697_),
    .Y(_11698_),
    .A1(_08524_),
    .A2(_11691_));
 sg13g2_o21ai_1 _19363_ (.B1(_11530_),
    .Y(_11699_),
    .A1(_11347_),
    .A2(_11698_));
 sg13g2_inv_1 _19364_ (.Y(_11700_),
    .A(_11698_));
 sg13g2_nor3_1 _19365_ (.A(_08526_),
    .B(_11647_),
    .C(_11700_),
    .Y(_11701_));
 sg13g2_a21oi_1 _19366_ (.A1(_08526_),
    .A2(_11699_),
    .Y(_11702_),
    .B1(_11701_));
 sg13g2_nor2_1 _19367_ (.A(net634),
    .B(_11702_),
    .Y(_01495_));
 sg13g2_nor3_1 _19368_ (.A(_08524_),
    .B(_08526_),
    .C(_11691_),
    .Y(_11703_));
 sg13g2_nor2_1 _19369_ (.A(_11643_),
    .B(_11703_),
    .Y(_11704_));
 sg13g2_nand2_1 _19370_ (.Y(_11705_),
    .A(net701),
    .B(_11704_));
 sg13g2_nand2_1 _19371_ (.Y(_11706_),
    .A(net67),
    .B(_11705_));
 sg13g2_nor3_1 _19372_ (.A(_08525_),
    .B(_11647_),
    .C(_11704_),
    .Y(_11707_));
 sg13g2_a21oi_1 _19373_ (.A1(_08525_),
    .A2(_11706_),
    .Y(_11708_),
    .B1(_11707_));
 sg13g2_nor2_1 _19374_ (.A(net634),
    .B(_11708_),
    .Y(_01496_));
 sg13g2_buf_1 _19375_ (.A(\rbzero.wall_tracer.side ),
    .X(_11709_));
 sg13g2_buf_1 _19376_ (.A(_11709_),
    .X(_11710_));
 sg13g2_buf_1 _19377_ (.A(_11710_),
    .X(_11711_));
 sg13g2_buf_1 _19378_ (.A(net699),
    .X(_11712_));
 sg13g2_buf_1 _19379_ (.A(net633),
    .X(_11713_));
 sg13g2_buf_1 _19380_ (.A(_08807_),
    .X(_11714_));
 sg13g2_buf_1 _19381_ (.A(net459),
    .X(_11715_));
 sg13g2_nand2_1 _19382_ (.Y(_11716_),
    .A(net573),
    .B(net450));
 sg13g2_buf_1 _19383_ (.A(\rbzero.row_render.side ),
    .X(_11717_));
 sg13g2_nand2_1 _19384_ (.Y(_11718_),
    .A(net812),
    .B(net452));
 sg13g2_a21oi_1 _19385_ (.A1(_11716_),
    .A2(_11718_),
    .Y(_01497_),
    .B1(net682));
 sg13g2_nand2_1 _19386_ (.Y(_11719_),
    .A(net573),
    .B(net547));
 sg13g2_nand2_1 _19387_ (.Y(_11720_),
    .A(_08414_),
    .B(_08475_));
 sg13g2_buf_1 _19388_ (.A(_11720_),
    .X(_11721_));
 sg13g2_nand2_1 _19389_ (.Y(_11722_),
    .A(\rbzero.side_hot ),
    .B(_11721_));
 sg13g2_a21oi_1 _19390_ (.A1(_11719_),
    .A2(_11722_),
    .Y(_01498_),
    .B1(net682));
 sg13g2_nand2_1 _19391_ (.Y(_11723_),
    .A(\rbzero.wall_tracer.size[0] ),
    .B(net450));
 sg13g2_buf_1 _19392_ (.A(\rbzero.row_render.size[0] ),
    .X(_11724_));
 sg13g2_nand2_1 _19393_ (.Y(_11725_),
    .A(_11724_),
    .B(net452));
 sg13g2_buf_1 _19394_ (.A(net729),
    .X(_11726_));
 sg13g2_a21oi_1 _19395_ (.A1(_11723_),
    .A2(_11725_),
    .Y(_01499_),
    .B1(net632));
 sg13g2_buf_2 _19396_ (.A(\rbzero.wall_tracer.size[10] ),
    .X(_11727_));
 sg13g2_nand2_1 _19397_ (.Y(_11728_),
    .A(_11727_),
    .B(_11715_));
 sg13g2_buf_1 _19398_ (.A(\rbzero.row_render.size[10] ),
    .X(_11729_));
 sg13g2_nand2_1 _19399_ (.Y(_11730_),
    .A(_11729_),
    .B(net452));
 sg13g2_a21oi_1 _19400_ (.A1(_11728_),
    .A2(_11730_),
    .Y(_01500_),
    .B1(net632));
 sg13g2_nand2_1 _19401_ (.Y(_11731_),
    .A(\rbzero.wall_tracer.size[1] ),
    .B(net450));
 sg13g2_buf_1 _19402_ (.A(\rbzero.row_render.size[1] ),
    .X(_11732_));
 sg13g2_nand2_1 _19403_ (.Y(_11733_),
    .A(net811),
    .B(net452));
 sg13g2_a21oi_1 _19404_ (.A1(_11731_),
    .A2(_11733_),
    .Y(_01501_),
    .B1(net632));
 sg13g2_buf_1 _19405_ (.A(net462),
    .X(_11734_));
 sg13g2_nand2_1 _19406_ (.Y(_11735_),
    .A(\rbzero.wall_tracer.size[2] ),
    .B(net449));
 sg13g2_buf_2 _19407_ (.A(\rbzero.row_render.size[2] ),
    .X(_11736_));
 sg13g2_nand2_1 _19408_ (.Y(_11737_),
    .A(_11736_),
    .B(net452));
 sg13g2_a21oi_1 _19409_ (.A1(_11735_),
    .A2(_11737_),
    .Y(_01502_),
    .B1(net632));
 sg13g2_nand2_1 _19410_ (.Y(_11738_),
    .A(\rbzero.wall_tracer.size[3] ),
    .B(net449));
 sg13g2_buf_2 _19411_ (.A(\rbzero.row_render.size[3] ),
    .X(_11739_));
 sg13g2_nand2_1 _19412_ (.Y(_11740_),
    .A(_11739_),
    .B(net452));
 sg13g2_a21oi_1 _19413_ (.A1(_11738_),
    .A2(_11740_),
    .Y(_01503_),
    .B1(net632));
 sg13g2_nand2_1 _19414_ (.Y(_11741_),
    .A(\rbzero.wall_tracer.size[4] ),
    .B(net449));
 sg13g2_buf_2 _19415_ (.A(\rbzero.row_render.size[4] ),
    .X(_11742_));
 sg13g2_buf_1 _19416_ (.A(net464),
    .X(_11743_));
 sg13g2_nand2_1 _19417_ (.Y(_11744_),
    .A(_11742_),
    .B(net448));
 sg13g2_a21oi_1 _19418_ (.A1(_11741_),
    .A2(_11744_),
    .Y(_01504_),
    .B1(_11726_));
 sg13g2_nand2_1 _19419_ (.Y(_11745_),
    .A(\rbzero.wall_tracer.size[5] ),
    .B(net449));
 sg13g2_buf_1 _19420_ (.A(\rbzero.row_render.size[5] ),
    .X(_11746_));
 sg13g2_nand2_1 _19421_ (.Y(_11747_),
    .A(_11746_),
    .B(net448));
 sg13g2_a21oi_1 _19422_ (.A1(_11745_),
    .A2(_11747_),
    .Y(_01505_),
    .B1(net632));
 sg13g2_buf_2 _19423_ (.A(\rbzero.wall_tracer.size[6] ),
    .X(_11748_));
 sg13g2_nand2_1 _19424_ (.Y(_11749_),
    .A(_11748_),
    .B(_11734_));
 sg13g2_buf_2 _19425_ (.A(\rbzero.row_render.size[6] ),
    .X(_11750_));
 sg13g2_nand2_1 _19426_ (.Y(_11751_),
    .A(_11750_),
    .B(net448));
 sg13g2_a21oi_1 _19427_ (.A1(_11749_),
    .A2(_11751_),
    .Y(_01506_),
    .B1(net632));
 sg13g2_buf_1 _19428_ (.A(\rbzero.wall_tracer.size[7] ),
    .X(_11752_));
 sg13g2_nand2_1 _19429_ (.Y(_11753_),
    .A(_11752_),
    .B(net449));
 sg13g2_buf_2 _19430_ (.A(\rbzero.row_render.size[7] ),
    .X(_11754_));
 sg13g2_nand2_1 _19431_ (.Y(_11755_),
    .A(_11754_),
    .B(net448));
 sg13g2_a21oi_1 _19432_ (.A1(_11753_),
    .A2(_11755_),
    .Y(_01507_),
    .B1(_11726_));
 sg13g2_buf_1 _19433_ (.A(\rbzero.wall_tracer.size[8] ),
    .X(_11756_));
 sg13g2_nand2_1 _19434_ (.Y(_11757_),
    .A(_11756_),
    .B(net449));
 sg13g2_buf_1 _19435_ (.A(\rbzero.row_render.size[8] ),
    .X(_11758_));
 sg13g2_nand2_1 _19436_ (.Y(_11759_),
    .A(_11758_),
    .B(net448));
 sg13g2_a21oi_1 _19437_ (.A1(_11757_),
    .A2(_11759_),
    .Y(_01508_),
    .B1(net632));
 sg13g2_buf_1 _19438_ (.A(\rbzero.wall_tracer.size[9] ),
    .X(_11760_));
 sg13g2_nand2_1 _19439_ (.Y(_11761_),
    .A(_11760_),
    .B(_11734_));
 sg13g2_buf_2 _19440_ (.A(\rbzero.row_render.size[9] ),
    .X(_11762_));
 sg13g2_nand2_1 _19441_ (.Y(_11763_),
    .A(_11762_),
    .B(net448));
 sg13g2_buf_2 _19442_ (.A(_08746_),
    .X(_11764_));
 sg13g2_buf_1 _19443_ (.A(_11764_),
    .X(_11765_));
 sg13g2_a21oi_1 _19444_ (.A1(_11761_),
    .A2(_11763_),
    .Y(_01509_),
    .B1(_11765_));
 sg13g2_inv_2 _19445_ (.Y(_11766_),
    .A(_08443_));
 sg13g2_buf_1 _19446_ (.A(_11766_),
    .X(_11767_));
 sg13g2_buf_1 _19447_ (.A(net698),
    .X(_11768_));
 sg13g2_xnor2_1 _19448_ (.Y(_11769_),
    .A(_09937_),
    .B(_09923_));
 sg13g2_mux2_1 _19449_ (.A0(_00442_),
    .A1(_11769_),
    .S(_11628_),
    .X(_11770_));
 sg13g2_buf_1 _19450_ (.A(_08439_),
    .X(_11771_));
 sg13g2_mux2_1 _19451_ (.A0(_00441_),
    .A1(_11770_),
    .S(net740),
    .X(_11772_));
 sg13g2_buf_2 _19452_ (.A(_11772_),
    .X(_11773_));
 sg13g2_nand2_1 _19453_ (.Y(_11774_),
    .A(_00443_),
    .B(_11438_));
 sg13g2_xnor2_1 _19454_ (.Y(_11775_),
    .A(_09840_),
    .B(_09817_));
 sg13g2_nand2b_1 _19455_ (.Y(_11776_),
    .B(_11775_),
    .A_N(_11438_));
 sg13g2_a21oi_1 _19456_ (.A1(_11774_),
    .A2(_11776_),
    .Y(_11777_),
    .B1(_11766_));
 sg13g2_buf_2 _19457_ (.A(_11777_),
    .X(_11778_));
 sg13g2_a21oi_1 _19458_ (.A1(net631),
    .A2(_11773_),
    .Y(_11779_),
    .B1(_11778_));
 sg13g2_buf_1 _19459_ (.A(_11779_),
    .X(_11780_));
 sg13g2_buf_1 _19460_ (.A(net283),
    .X(_11781_));
 sg13g2_nand2b_1 _19461_ (.Y(_11782_),
    .B(net797),
    .A_N(_00438_));
 sg13g2_inv_2 _19462_ (.Y(_11783_),
    .A(_08439_));
 sg13g2_nor2_1 _19463_ (.A(_11783_),
    .B(_00439_),
    .Y(_11784_));
 sg13g2_inv_1 _19464_ (.Y(_11785_),
    .A(_11584_));
 sg13g2_nand2_1 _19465_ (.Y(_11786_),
    .A(net741),
    .B(_11405_));
 sg13g2_o21ai_1 _19466_ (.B1(_11786_),
    .Y(_11787_),
    .A1(net741),
    .A2(_11785_));
 sg13g2_mux2_1 _19467_ (.A0(_00440_),
    .A1(_11787_),
    .S(net833),
    .X(_11788_));
 sg13g2_nor2_1 _19468_ (.A(net740),
    .B(_11788_),
    .Y(_11789_));
 sg13g2_o21ai_1 _19469_ (.B1(_11766_),
    .Y(_11790_),
    .A1(_11784_),
    .A2(_11789_));
 sg13g2_buf_1 _19470_ (.A(_11790_),
    .X(_11791_));
 sg13g2_nand2_1 _19471_ (.Y(_11792_),
    .A(_11782_),
    .B(_11791_));
 sg13g2_buf_2 _19472_ (.A(_11792_),
    .X(_11793_));
 sg13g2_buf_1 _19473_ (.A(_11793_),
    .X(_11794_));
 sg13g2_nand2_1 _19474_ (.Y(_11795_),
    .A(net268),
    .B(net307));
 sg13g2_buf_2 _19475_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_11796_));
 sg13g2_nor2_1 _19476_ (.A(_11771_),
    .B(_08443_),
    .Y(_11797_));
 sg13g2_buf_1 _19477_ (.A(_11797_),
    .X(_11798_));
 sg13g2_and2_1 _19478_ (.A(_11796_),
    .B(net630),
    .X(_11799_));
 sg13g2_buf_1 _19479_ (.A(_11799_),
    .X(_11800_));
 sg13g2_nor2_1 _19480_ (.A(net813),
    .B(_11569_),
    .Y(_11801_));
 sg13g2_a21oi_1 _19481_ (.A1(net741),
    .A2(_11400_),
    .Y(_11802_),
    .B1(_11801_));
 sg13g2_xnor2_1 _19482_ (.Y(_11803_),
    .A(_11748_),
    .B(_11752_));
 sg13g2_nor2_1 _19483_ (.A(net833),
    .B(_11803_),
    .Y(_11804_));
 sg13g2_a21oi_1 _19484_ (.A1(_08419_),
    .A2(_11802_),
    .Y(_11805_),
    .B1(_11804_));
 sg13g2_nand2_1 _19485_ (.Y(_11806_),
    .A(net740),
    .B(_00448_));
 sg13g2_o21ai_1 _19486_ (.B1(_11806_),
    .Y(_11807_),
    .A1(net740),
    .A2(_11805_));
 sg13g2_and2_1 _19487_ (.A(_08443_),
    .B(_00447_),
    .X(_11808_));
 sg13g2_a21oi_1 _19488_ (.A1(_11766_),
    .A2(_11807_),
    .Y(_11809_),
    .B1(_11808_));
 sg13g2_buf_1 _19489_ (.A(_11809_),
    .X(_11810_));
 sg13g2_nand2_1 _19490_ (.Y(_11811_),
    .A(_11800_),
    .B(_11810_));
 sg13g2_mux2_1 _19491_ (.A0(_00446_),
    .A1(_09926_),
    .S(_08439_),
    .X(_11812_));
 sg13g2_and2_1 _19492_ (.A(_08443_),
    .B(_09820_),
    .X(_11813_));
 sg13g2_a21oi_1 _19493_ (.A1(_11766_),
    .A2(_11812_),
    .Y(_11814_),
    .B1(_11813_));
 sg13g2_buf_1 _19494_ (.A(_11814_),
    .X(_11815_));
 sg13g2_nand2b_1 _19495_ (.Y(_11816_),
    .B(net797),
    .A_N(_00444_));
 sg13g2_nor2_1 _19496_ (.A(_11783_),
    .B(_00445_),
    .Y(_11817_));
 sg13g2_nand2_1 _19497_ (.Y(_11818_),
    .A(net813),
    .B(_11402_));
 sg13g2_o21ai_1 _19498_ (.B1(_11818_),
    .Y(_11819_),
    .A1(net813),
    .A2(_11581_));
 sg13g2_mux2_1 _19499_ (.A0(_11748_),
    .A1(_11819_),
    .S(net833),
    .X(_11820_));
 sg13g2_nor2_1 _19500_ (.A(_08439_),
    .B(_11820_),
    .Y(_11821_));
 sg13g2_o21ai_1 _19501_ (.B1(_11766_),
    .Y(_11822_),
    .A1(_11817_),
    .A2(_11821_));
 sg13g2_buf_1 _19502_ (.A(_11822_),
    .X(_11823_));
 sg13g2_nand2_1 _19503_ (.Y(_11824_),
    .A(_11816_),
    .B(_11823_));
 sg13g2_buf_1 _19504_ (.A(_11824_),
    .X(_11825_));
 sg13g2_nand2_1 _19505_ (.Y(_11826_),
    .A(_11815_),
    .B(_11825_));
 sg13g2_xor2_1 _19506_ (.B(_11826_),
    .A(_11811_),
    .X(_11827_));
 sg13g2_xnor2_1 _19507_ (.Y(_11828_),
    .A(_11795_),
    .B(_11827_));
 sg13g2_nand2b_1 _19508_ (.Y(_11829_),
    .B(net797),
    .A_N(_00432_));
 sg13g2_nor2b_1 _19509_ (.A(net741),
    .B_N(_11587_),
    .Y(_11830_));
 sg13g2_a21oi_1 _19510_ (.A1(net741),
    .A2(_11410_),
    .Y(_11831_),
    .B1(_11830_));
 sg13g2_mux2_1 _19511_ (.A0(_00434_),
    .A1(_11831_),
    .S(net800),
    .X(_11832_));
 sg13g2_nand2b_1 _19512_ (.Y(_11833_),
    .B(net740),
    .A_N(_00433_));
 sg13g2_o21ai_1 _19513_ (.B1(_11833_),
    .Y(_11834_),
    .A1(_08440_),
    .A2(_11832_));
 sg13g2_nand2_1 _19514_ (.Y(_11835_),
    .A(net698),
    .B(_11834_));
 sg13g2_nand2_1 _19515_ (.Y(_11836_),
    .A(_11829_),
    .B(_11835_));
 sg13g2_buf_1 _19516_ (.A(_11836_),
    .X(_11837_));
 sg13g2_nand2_1 _19517_ (.Y(_11838_),
    .A(net283),
    .B(net333));
 sg13g2_buf_1 _19518_ (.A(_11815_),
    .X(_11839_));
 sg13g2_nand2_1 _19519_ (.Y(_11840_),
    .A(_11793_),
    .B(net571));
 sg13g2_buf_1 _19520_ (.A(_11800_),
    .X(_11841_));
 sg13g2_nand2_1 _19521_ (.Y(_11842_),
    .A(net506),
    .B(_11825_));
 sg13g2_or2_1 _19522_ (.X(_11843_),
    .B(_11842_),
    .A(_11840_));
 sg13g2_and2_1 _19523_ (.A(_11840_),
    .B(_11842_),
    .X(_11844_));
 sg13g2_a21oi_2 _19524_ (.B1(_11844_),
    .Y(_11845_),
    .A2(_11843_),
    .A1(_11838_));
 sg13g2_buf_1 _19525_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_11846_));
 sg13g2_and2_1 _19526_ (.A(_11846_),
    .B(net630),
    .X(_11847_));
 sg13g2_buf_1 _19527_ (.A(_11847_),
    .X(_11848_));
 sg13g2_or2_1 _19528_ (.X(_11849_),
    .B(_11567_),
    .A(_11566_));
 sg13g2_and2_1 _19529_ (.A(_11397_),
    .B(_11398_),
    .X(_11850_));
 sg13g2_mux2_1 _19530_ (.A0(_11849_),
    .A1(_11850_),
    .S(_11711_),
    .X(_11851_));
 sg13g2_o21ai_1 _19531_ (.B1(_11756_),
    .Y(_11852_),
    .A1(_11748_),
    .A2(_11752_));
 sg13g2_buf_1 _19532_ (.A(_11852_),
    .X(_11853_));
 sg13g2_inv_1 _19533_ (.Y(_11854_),
    .A(_11853_));
 sg13g2_nor3_1 _19534_ (.A(_11748_),
    .B(_11752_),
    .C(_11756_),
    .Y(_11855_));
 sg13g2_nor3_1 _19535_ (.A(net800),
    .B(_11854_),
    .C(_11855_),
    .Y(_11856_));
 sg13g2_a21o_1 _19536_ (.A2(_11851_),
    .A1(net728),
    .B1(_11856_),
    .X(_11857_));
 sg13g2_nand2_1 _19537_ (.Y(_11858_),
    .A(net726),
    .B(_00450_));
 sg13g2_o21ai_1 _19538_ (.B1(_11858_),
    .Y(_11859_),
    .A1(net726),
    .A2(_11857_));
 sg13g2_and2_1 _19539_ (.A(net797),
    .B(_00449_),
    .X(_11860_));
 sg13g2_a21oi_1 _19540_ (.A1(net631),
    .A2(_11859_),
    .Y(_11861_),
    .B1(_11860_));
 sg13g2_buf_1 _19541_ (.A(_11861_),
    .X(_11862_));
 sg13g2_and2_1 _19542_ (.A(net524),
    .B(_11862_),
    .X(_11863_));
 sg13g2_xnor2_1 _19543_ (.Y(_11864_),
    .A(_11845_),
    .B(_11863_));
 sg13g2_xnor2_1 _19544_ (.Y(_11865_),
    .A(_11828_),
    .B(_11864_));
 sg13g2_buf_1 _19545_ (.A(net631),
    .X(_11866_));
 sg13g2_xor2_1 _19546_ (.B(_09985_),
    .A(_09938_),
    .X(_11867_));
 sg13g2_mux2_1 _19547_ (.A0(_00436_),
    .A1(_11867_),
    .S(_11628_),
    .X(_11868_));
 sg13g2_mux2_1 _19548_ (.A0(_00435_),
    .A1(_11868_),
    .S(net798),
    .X(_11869_));
 sg13g2_buf_1 _19549_ (.A(_11869_),
    .X(_11870_));
 sg13g2_nor2b_1 _19550_ (.A(_00437_),
    .B_N(net308),
    .Y(_11871_));
 sg13g2_nor2b_1 _19551_ (.A(_09888_),
    .B_N(_09841_),
    .Y(_11872_));
 sg13g2_nor3_1 _19552_ (.A(_09842_),
    .B(net308),
    .C(_11872_),
    .Y(_11873_));
 sg13g2_nor3_2 _19553_ (.A(net698),
    .B(_11871_),
    .C(_11873_),
    .Y(_11874_));
 sg13g2_a21oi_1 _19554_ (.A1(net570),
    .A2(_11870_),
    .Y(_11875_),
    .B1(_11874_));
 sg13g2_buf_2 _19555_ (.A(_11875_),
    .X(_11876_));
 sg13g2_nand2b_1 _19556_ (.Y(_11877_),
    .B(_08443_),
    .A_N(_00426_));
 sg13g2_buf_1 _19557_ (.A(_11877_),
    .X(_11878_));
 sg13g2_nand2_1 _19558_ (.Y(_11879_),
    .A(net813),
    .B(_11412_));
 sg13g2_o21ai_1 _19559_ (.B1(_11879_),
    .Y(_11880_),
    .A1(net813),
    .A2(_11589_));
 sg13g2_nor2b_1 _19560_ (.A(net833),
    .B_N(_00428_),
    .Y(_11881_));
 sg13g2_a21oi_1 _19561_ (.A1(net833),
    .A2(_11880_),
    .Y(_11882_),
    .B1(_11881_));
 sg13g2_nor2_1 _19562_ (.A(net740),
    .B(_11882_),
    .Y(_11883_));
 sg13g2_a21oi_1 _19563_ (.A1(net740),
    .A2(_00427_),
    .Y(_11884_),
    .B1(_11883_));
 sg13g2_nand2_1 _19564_ (.Y(_11885_),
    .A(_11766_),
    .B(_11884_));
 sg13g2_nand2_1 _19565_ (.Y(_11886_),
    .A(_11878_),
    .B(_11885_));
 sg13g2_buf_2 _19566_ (.A(_11886_),
    .X(_11887_));
 sg13g2_nand2_1 _19567_ (.Y(_11888_),
    .A(_11876_),
    .B(_11887_));
 sg13g2_inv_1 _19568_ (.Y(_11889_),
    .A(_09926_));
 sg13g2_nor3_1 _19569_ (.A(_11889_),
    .B(_09937_),
    .C(_09938_),
    .Y(_11890_));
 sg13g2_xor2_1 _19570_ (.B(_11890_),
    .A(_09936_),
    .X(_11891_));
 sg13g2_mux2_1 _19571_ (.A0(_00430_),
    .A1(_11891_),
    .S(_11628_),
    .X(_11892_));
 sg13g2_nor2b_1 _19572_ (.A(net798),
    .B_N(_00429_),
    .Y(_11893_));
 sg13g2_a21oi_1 _19573_ (.A1(net726),
    .A2(_11892_),
    .Y(_11894_),
    .B1(_11893_));
 sg13g2_nand2b_1 _19574_ (.Y(_11895_),
    .B(net308),
    .A_N(_00431_));
 sg13g2_nor2_1 _19575_ (.A(_09840_),
    .B(_09841_),
    .Y(_11896_));
 sg13g2_nand2_1 _19576_ (.Y(_11897_),
    .A(_09820_),
    .B(_11896_));
 sg13g2_xor2_1 _19577_ (.B(_11897_),
    .A(_09839_),
    .X(_11898_));
 sg13g2_nand2b_1 _19578_ (.Y(_11899_),
    .B(_11898_),
    .A_N(_11438_));
 sg13g2_a21oi_1 _19579_ (.A1(_11895_),
    .A2(_11899_),
    .Y(_11900_),
    .B1(net698));
 sg13g2_a21oi_1 _19580_ (.A1(net570),
    .A2(_11894_),
    .Y(_11901_),
    .B1(_11900_));
 sg13g2_buf_1 _19581_ (.A(_11901_),
    .X(_11902_));
 sg13g2_nand2b_1 _19582_ (.Y(_11903_),
    .B(net797),
    .A_N(_00420_));
 sg13g2_buf_1 _19583_ (.A(_11903_),
    .X(_11904_));
 sg13g2_nor2b_1 _19584_ (.A(net741),
    .B_N(_11592_),
    .Y(_11905_));
 sg13g2_a21oi_1 _19585_ (.A1(net741),
    .A2(_11416_),
    .Y(_11906_),
    .B1(_11905_));
 sg13g2_nor2b_1 _19586_ (.A(net833),
    .B_N(_00422_),
    .Y(_11907_));
 sg13g2_a21oi_1 _19587_ (.A1(net800),
    .A2(_11906_),
    .Y(_11908_),
    .B1(_11907_));
 sg13g2_nor2_1 _19588_ (.A(net798),
    .B(_11908_),
    .Y(_11909_));
 sg13g2_a21oi_1 _19589_ (.A1(net798),
    .A2(_00421_),
    .Y(_11910_),
    .B1(_11909_));
 sg13g2_nand2_1 _19590_ (.Y(_11911_),
    .A(net698),
    .B(_11910_));
 sg13g2_and2_1 _19591_ (.A(_11904_),
    .B(_11911_),
    .X(_11912_));
 sg13g2_buf_2 _19592_ (.A(_11912_),
    .X(_11913_));
 sg13g2_nand2b_1 _19593_ (.Y(_11914_),
    .B(_08444_),
    .A_N(_00414_));
 sg13g2_buf_1 _19594_ (.A(_11914_),
    .X(_11915_));
 sg13g2_inv_1 _19595_ (.Y(_11916_),
    .A(_11419_));
 sg13g2_nor2_1 _19596_ (.A(_11710_),
    .B(_11595_),
    .Y(_11917_));
 sg13g2_a21oi_1 _19597_ (.A1(net699),
    .A2(_11916_),
    .Y(_11918_),
    .B1(_11917_));
 sg13g2_nor2b_1 _19598_ (.A(net800),
    .B_N(_00416_),
    .Y(_11919_));
 sg13g2_a21oi_1 _19599_ (.A1(net800),
    .A2(_11918_),
    .Y(_11920_),
    .B1(_11919_));
 sg13g2_nand2_1 _19600_ (.Y(_11921_),
    .A(_11783_),
    .B(_11920_));
 sg13g2_o21ai_1 _19601_ (.B1(_11921_),
    .Y(_11922_),
    .A1(_11783_),
    .A2(_00415_));
 sg13g2_nand2_2 _19602_ (.Y(_11923_),
    .A(net698),
    .B(_11922_));
 sg13g2_xor2_1 _19603_ (.B(_09941_),
    .A(_09935_),
    .X(_11924_));
 sg13g2_mux2_1 _19604_ (.A0(_00424_),
    .A1(_11924_),
    .S(_11628_),
    .X(_11925_));
 sg13g2_mux2_1 _19605_ (.A0(_00423_),
    .A1(_11925_),
    .S(net798),
    .X(_11926_));
 sg13g2_buf_1 _19606_ (.A(_11926_),
    .X(_11927_));
 sg13g2_buf_1 _19607_ (.A(_11768_),
    .X(_11928_));
 sg13g2_nor2b_1 _19608_ (.A(_00425_),
    .B_N(_11438_),
    .Y(_11929_));
 sg13g2_xor2_1 _19609_ (.B(_09844_),
    .A(_09838_),
    .X(_11930_));
 sg13g2_nor2_1 _19610_ (.A(_11438_),
    .B(_11930_),
    .Y(_11931_));
 sg13g2_nor3_1 _19611_ (.A(net698),
    .B(_11929_),
    .C(_11931_),
    .Y(_11932_));
 sg13g2_buf_1 _19612_ (.A(_11932_),
    .X(_11933_));
 sg13g2_a221oi_1 _19613_ (.B2(net569),
    .C1(_11933_),
    .B1(_11927_),
    .A1(_11915_),
    .Y(_11934_),
    .A2(_11923_));
 sg13g2_o21ai_1 _19614_ (.B1(_11934_),
    .Y(_11935_),
    .A1(_11902_),
    .A2(_11913_));
 sg13g2_a21o_1 _19615_ (.A2(_11894_),
    .A1(net631),
    .B1(_11900_),
    .X(_11936_));
 sg13g2_buf_1 _19616_ (.A(_11936_),
    .X(_11937_));
 sg13g2_buf_1 _19617_ (.A(_11937_),
    .X(_11938_));
 sg13g2_nand2_1 _19618_ (.Y(_11939_),
    .A(_11904_),
    .B(_11911_));
 sg13g2_buf_1 _19619_ (.A(_11939_),
    .X(_11940_));
 sg13g2_nand3b_1 _19620_ (.B(net267),
    .C(net407),
    .Y(_11941_),
    .A_N(_11934_));
 sg13g2_and3_1 _19621_ (.X(_11942_),
    .A(_11888_),
    .B(_11935_),
    .C(_11941_));
 sg13g2_buf_1 _19622_ (.A(_11942_),
    .X(_11943_));
 sg13g2_a21oi_1 _19623_ (.A1(_11935_),
    .A2(_11941_),
    .Y(_11944_),
    .B1(_11888_));
 sg13g2_nand2_1 _19624_ (.Y(_11945_),
    .A(_11915_),
    .B(_11923_));
 sg13g2_buf_2 _19625_ (.A(_11945_),
    .X(_11946_));
 sg13g2_nand2_1 _19626_ (.Y(_11947_),
    .A(_11946_),
    .B(net267));
 sg13g2_nand2b_1 _19627_ (.Y(_11948_),
    .B(_08444_),
    .A_N(_00409_));
 sg13g2_buf_4 _19628_ (.X(_11949_),
    .A(_11948_));
 sg13g2_nor2_1 _19629_ (.A(_11783_),
    .B(_00410_),
    .Y(_11950_));
 sg13g2_nand2_1 _19630_ (.Y(_11951_),
    .A(net813),
    .B(_11422_));
 sg13g2_o21ai_1 _19631_ (.B1(_11951_),
    .Y(_11952_),
    .A1(net741),
    .A2(_11598_));
 sg13g2_mux2_1 _19632_ (.A0(_00411_),
    .A1(_11952_),
    .S(net833),
    .X(_11953_));
 sg13g2_nor2_1 _19633_ (.A(net740),
    .B(_11953_),
    .Y(_11954_));
 sg13g2_o21ai_1 _19634_ (.B1(_11766_),
    .Y(_11955_),
    .A1(_11950_),
    .A2(_11954_));
 sg13g2_buf_4 _19635_ (.X(_11956_),
    .A(_11955_));
 sg13g2_nand2_1 _19636_ (.Y(_11957_),
    .A(_11949_),
    .B(_11956_));
 sg13g2_buf_1 _19637_ (.A(_11957_),
    .X(_11958_));
 sg13g2_a21oi_1 _19638_ (.A1(net570),
    .A2(_11927_),
    .Y(_11959_),
    .B1(_11933_));
 sg13g2_buf_2 _19639_ (.A(_11959_),
    .X(_11960_));
 sg13g2_nand4_1 _19640_ (.B(_11876_),
    .C(_11960_),
    .A(net458),
    .Y(_11961_),
    .D(net407));
 sg13g2_a22oi_1 _19641_ (.Y(_11962_),
    .B1(net407),
    .B2(_11876_),
    .A2(_11960_),
    .A1(net458));
 sg13g2_a21o_1 _19642_ (.A2(_11961_),
    .A1(_11947_),
    .B1(_11962_),
    .X(_11963_));
 sg13g2_buf_1 _19643_ (.A(_11963_),
    .X(_11964_));
 sg13g2_nor3_1 _19644_ (.A(_11943_),
    .B(_11944_),
    .C(_11964_),
    .Y(_11965_));
 sg13g2_nor2_1 _19645_ (.A(_09936_),
    .B(_09935_),
    .Y(_11966_));
 sg13g2_and2_1 _19646_ (.A(_11890_),
    .B(_11966_),
    .X(_11967_));
 sg13g2_xor2_1 _19647_ (.B(_11967_),
    .A(_09933_),
    .X(_11968_));
 sg13g2_mux2_1 _19648_ (.A0(_00418_),
    .A1(_11968_),
    .S(_11628_),
    .X(_11969_));
 sg13g2_mux2_1 _19649_ (.A0(_00417_),
    .A1(_11969_),
    .S(net726),
    .X(_11970_));
 sg13g2_nor2b_1 _19650_ (.A(_00419_),
    .B_N(_11439_),
    .Y(_11971_));
 sg13g2_nor3_1 _19651_ (.A(_09839_),
    .B(_09838_),
    .C(_11897_),
    .Y(_11972_));
 sg13g2_xor2_1 _19652_ (.B(_11972_),
    .A(_09836_),
    .X(_11973_));
 sg13g2_nor2_1 _19653_ (.A(_11439_),
    .B(_11973_),
    .Y(_11974_));
 sg13g2_o21ai_1 _19654_ (.B1(net797),
    .Y(_11975_),
    .A1(_11971_),
    .A2(_11974_));
 sg13g2_o21ai_1 _19655_ (.B1(_11975_),
    .Y(_11976_),
    .A1(net725),
    .A2(_11970_));
 sg13g2_buf_1 _19656_ (.A(_11976_),
    .X(_11977_));
 sg13g2_nand2b_1 _19657_ (.Y(_11978_),
    .B(net797),
    .A_N(_00403_));
 sg13g2_buf_1 _19658_ (.A(_11978_),
    .X(_11979_));
 sg13g2_nor2_1 _19659_ (.A(net813),
    .B(_11599_),
    .Y(_11980_));
 sg13g2_a21oi_1 _19660_ (.A1(net813),
    .A2(_11423_),
    .Y(_11981_),
    .B1(_11980_));
 sg13g2_nand2_1 _19661_ (.Y(_11982_),
    .A(net833),
    .B(_11981_));
 sg13g2_o21ai_1 _19662_ (.B1(_11982_),
    .Y(_11983_),
    .A1(_08418_),
    .A2(_00405_));
 sg13g2_nor2_1 _19663_ (.A(_11771_),
    .B(_11983_),
    .Y(_11984_));
 sg13g2_a21oi_1 _19664_ (.A1(net798),
    .A2(_00404_),
    .Y(_11985_),
    .B1(_11984_));
 sg13g2_nand2_1 _19665_ (.Y(_11986_),
    .A(net698),
    .B(_11985_));
 sg13g2_nand2_1 _19666_ (.Y(_11987_),
    .A(_11979_),
    .B(_11986_));
 sg13g2_buf_1 _19667_ (.A(_11987_),
    .X(_11988_));
 sg13g2_nand2_1 _19668_ (.Y(_11989_),
    .A(net282),
    .B(net457));
 sg13g2_xor2_1 _19669_ (.B(_09998_),
    .A(_09934_),
    .X(_11990_));
 sg13g2_mux2_1 _19670_ (.A0(_00412_),
    .A1(_11990_),
    .S(_11628_),
    .X(_11991_));
 sg13g2_mux2_1 _19671_ (.A0(_00018_),
    .A1(_11991_),
    .S(net726),
    .X(_11992_));
 sg13g2_nor2b_1 _19672_ (.A(_00413_),
    .B_N(net308),
    .Y(_11993_));
 sg13g2_nor2b_1 _19673_ (.A(_09902_),
    .B_N(_09837_),
    .Y(_11994_));
 sg13g2_nor3_1 _19674_ (.A(_09847_),
    .B(net308),
    .C(_11994_),
    .Y(_11995_));
 sg13g2_nor3_1 _19675_ (.A(net631),
    .B(_11993_),
    .C(_11995_),
    .Y(_11996_));
 sg13g2_a21oi_1 _19676_ (.A1(_11866_),
    .A2(_11992_),
    .Y(_11997_),
    .B1(_11996_));
 sg13g2_buf_1 _19677_ (.A(_11997_),
    .X(_11998_));
 sg13g2_buf_1 _19678_ (.A(_11998_),
    .X(_11999_));
 sg13g2_nor2_1 _19679_ (.A(_09933_),
    .B(_09934_),
    .Y(_12000_));
 sg13g2_nand2_1 _19680_ (.Y(_12001_),
    .A(_11967_),
    .B(_12000_));
 sg13g2_xnor2_1 _19681_ (.Y(_12002_),
    .A(_09932_),
    .B(_12001_));
 sg13g2_mux2_1 _19682_ (.A0(_00407_),
    .A1(_12002_),
    .S(net314),
    .X(_12003_));
 sg13g2_mux2_1 _19683_ (.A0(_00406_),
    .A1(_12003_),
    .S(net726),
    .X(_12004_));
 sg13g2_nor2b_1 _19684_ (.A(_00408_),
    .B_N(net308),
    .Y(_12005_));
 sg13g2_nor2_1 _19685_ (.A(_09836_),
    .B(_09837_),
    .Y(_12006_));
 sg13g2_nand2_1 _19686_ (.Y(_12007_),
    .A(_11972_),
    .B(_12006_));
 sg13g2_xnor2_1 _19687_ (.Y(_12008_),
    .A(_09835_),
    .B(_12007_));
 sg13g2_nor2_1 _19688_ (.A(net308),
    .B(_12008_),
    .Y(_12009_));
 sg13g2_nor3_1 _19689_ (.A(net631),
    .B(_12005_),
    .C(_12009_),
    .Y(_12010_));
 sg13g2_a21oi_1 _19690_ (.A1(net570),
    .A2(_12004_),
    .Y(_12011_),
    .B1(_12010_));
 sg13g2_buf_1 _19691_ (.A(_12011_),
    .X(_12012_));
 sg13g2_buf_2 _19692_ (.A(\rbzero.wall_tracer.stepDistX[-11] ),
    .X(_12013_));
 sg13g2_nand2_1 _19693_ (.Y(_12014_),
    .A(_08781_),
    .B(net699));
 sg13g2_nand2b_1 _19694_ (.Y(_12015_),
    .B(_09115_),
    .A_N(net699));
 sg13g2_nand3_1 _19695_ (.B(_12014_),
    .C(_12015_),
    .A(_08420_),
    .Y(_12016_));
 sg13g2_o21ai_1 _19696_ (.B1(_12016_),
    .Y(_12017_),
    .A1(net728),
    .A2(\rbzero.wall_tracer.size_full[-11] ));
 sg13g2_buf_2 _19697_ (.A(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_12018_));
 sg13g2_nand2_1 _19698_ (.Y(_12019_),
    .A(net726),
    .B(_12018_));
 sg13g2_o21ai_1 _19699_ (.B1(_12019_),
    .Y(_12020_),
    .A1(net684),
    .A2(_12017_));
 sg13g2_mux2_1 _19700_ (.A0(_12013_),
    .A1(_12020_),
    .S(net570),
    .X(_12021_));
 sg13g2_buf_2 _19701_ (.A(_12021_),
    .X(_12022_));
 sg13g2_buf_1 _19702_ (.A(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_12023_));
 sg13g2_nand2_1 _19703_ (.Y(_12024_),
    .A(net725),
    .B(_12023_));
 sg13g2_nand2_1 _19704_ (.Y(_12025_),
    .A(_08784_),
    .B(net699));
 sg13g2_nand2b_1 _19705_ (.Y(_12026_),
    .B(_09118_),
    .A_N(net699));
 sg13g2_nand3_1 _19706_ (.B(_12025_),
    .C(_12026_),
    .A(net800),
    .Y(_12027_));
 sg13g2_o21ai_1 _19707_ (.B1(_12027_),
    .Y(_12028_),
    .A1(_08419_),
    .A2(\rbzero.wall_tracer.size_full[-10] ));
 sg13g2_buf_1 _19708_ (.A(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_12029_));
 sg13g2_nand2_1 _19709_ (.Y(_12030_),
    .A(net798),
    .B(_12029_));
 sg13g2_o21ai_1 _19710_ (.B1(_12030_),
    .Y(_12031_),
    .A1(_08441_),
    .A2(_12028_));
 sg13g2_nand2_1 _19711_ (.Y(_12032_),
    .A(net631),
    .B(_12031_));
 sg13g2_nand2_1 _19712_ (.Y(_12033_),
    .A(_12024_),
    .B(_12032_));
 sg13g2_buf_1 _19713_ (.A(_12033_),
    .X(_12034_));
 sg13g2_nand4_1 _19714_ (.B(net281),
    .C(_12022_),
    .A(net266),
    .Y(_12035_),
    .D(net468));
 sg13g2_a22oi_1 _19715_ (.Y(_12036_),
    .B1(net468),
    .B2(net266),
    .A2(_12022_),
    .A1(net281));
 sg13g2_a21oi_1 _19716_ (.A1(_11989_),
    .A2(_12035_),
    .Y(_12037_),
    .B1(_12036_));
 sg13g2_o21ai_1 _19717_ (.B1(_11964_),
    .Y(_12038_),
    .A1(_11943_),
    .A2(_11944_));
 sg13g2_o21ai_1 _19718_ (.B1(_12038_),
    .Y(_12039_),
    .A1(_11965_),
    .A2(_12037_));
 sg13g2_buf_1 _19719_ (.A(_12039_),
    .X(_12040_));
 sg13g2_nand2_1 _19720_ (.Y(_12041_),
    .A(_11887_),
    .B(_11937_));
 sg13g2_a221oi_1 _19721_ (.B2(_11835_),
    .C1(_11874_),
    .B1(_11829_),
    .A1(net569),
    .Y(_12042_),
    .A2(_11870_));
 sg13g2_buf_1 _19722_ (.A(_12042_),
    .X(_12043_));
 sg13g2_a221oi_1 _19723_ (.B2(_11911_),
    .C1(_11933_),
    .B1(_11904_),
    .A1(net569),
    .Y(_12044_),
    .A2(_11927_));
 sg13g2_buf_1 _19724_ (.A(_12044_),
    .X(_12045_));
 sg13g2_xor2_1 _19725_ (.B(_12045_),
    .A(_12043_),
    .X(_12046_));
 sg13g2_xnor2_1 _19726_ (.Y(_12047_),
    .A(_12041_),
    .B(_12046_));
 sg13g2_nand2_1 _19727_ (.Y(_12048_),
    .A(net458),
    .B(net282));
 sg13g2_a221oi_1 _19728_ (.B2(_11986_),
    .C1(_11996_),
    .B1(_11979_),
    .A1(_11866_),
    .Y(_12049_),
    .A2(_11992_));
 sg13g2_buf_1 _19729_ (.A(_12049_),
    .X(_12050_));
 sg13g2_a21oi_1 _19730_ (.A1(_12011_),
    .A2(_12033_),
    .Y(_12051_),
    .B1(_12050_));
 sg13g2_nand3_1 _19731_ (.B(_12033_),
    .C(_12050_),
    .A(_12011_),
    .Y(_12052_));
 sg13g2_o21ai_1 _19732_ (.B1(_12052_),
    .Y(_12053_),
    .A1(_12048_),
    .A2(_12051_));
 sg13g2_buf_1 _19733_ (.A(_12053_),
    .X(_12054_));
 sg13g2_nand2_1 _19734_ (.Y(_12055_),
    .A(_11946_),
    .B(_11960_));
 sg13g2_a221oi_1 _19735_ (.B2(_11885_),
    .C1(_11874_),
    .B1(_11878_),
    .A1(net569),
    .Y(_12056_),
    .A2(_11870_));
 sg13g2_a21oi_1 _19736_ (.A1(_11937_),
    .A2(net407),
    .Y(_12057_),
    .B1(_12056_));
 sg13g2_nand3_1 _19737_ (.B(_11937_),
    .C(net407),
    .A(_12056_),
    .Y(_12058_));
 sg13g2_o21ai_1 _19738_ (.B1(_12058_),
    .Y(_12059_),
    .A1(_12055_),
    .A2(_12057_));
 sg13g2_buf_1 _19739_ (.A(_12059_),
    .X(_12060_));
 sg13g2_xor2_1 _19740_ (.B(_12060_),
    .A(_12054_),
    .X(_12061_));
 sg13g2_xnor2_1 _19741_ (.Y(_12062_),
    .A(_12047_),
    .B(_12061_));
 sg13g2_nand2_1 _19742_ (.Y(_12063_),
    .A(_12040_),
    .B(_12062_));
 sg13g2_nor2_1 _19743_ (.A(_12040_),
    .B(_12062_),
    .Y(_12064_));
 sg13g2_a21oi_1 _19744_ (.A1(_11865_),
    .A2(_12063_),
    .Y(_12065_),
    .B1(_12064_));
 sg13g2_buf_1 _19745_ (.A(_11876_),
    .X(_12066_));
 sg13g2_nand2_1 _19746_ (.Y(_12067_),
    .A(net265),
    .B(_11793_));
 sg13g2_and2_1 _19747_ (.A(_11878_),
    .B(_11885_),
    .X(_12068_));
 sg13g2_buf_1 _19748_ (.A(_12068_),
    .X(_12069_));
 sg13g2_a21o_1 _19749_ (.A2(_11927_),
    .A1(net570),
    .B1(_11933_),
    .X(_12070_));
 sg13g2_buf_2 _19750_ (.A(_12070_),
    .X(_12071_));
 sg13g2_nor2_1 _19751_ (.A(_12069_),
    .B(_12071_),
    .Y(_12072_));
 sg13g2_nand2_1 _19752_ (.Y(_12073_),
    .A(_11937_),
    .B(_11836_));
 sg13g2_xor2_1 _19753_ (.B(_12073_),
    .A(_12072_),
    .X(_12074_));
 sg13g2_xnor2_1 _19754_ (.Y(_12075_),
    .A(_12067_),
    .B(_12074_));
 sg13g2_nand2_1 _19755_ (.Y(_12076_),
    .A(_11946_),
    .B(net282));
 sg13g2_nand4_1 _19756_ (.B(_11998_),
    .C(net457),
    .A(_11958_),
    .Y(_12077_),
    .D(net281));
 sg13g2_a22oi_1 _19757_ (.Y(_12078_),
    .B1(net457),
    .B2(net281),
    .A2(_11998_),
    .A1(_11958_));
 sg13g2_a21oi_2 _19758_ (.B1(_12078_),
    .Y(_12079_),
    .A2(_12077_),
    .A1(_12076_));
 sg13g2_nand2_1 _19759_ (.Y(_12080_),
    .A(_12043_),
    .B(_12045_));
 sg13g2_nor2_1 _19760_ (.A(_12043_),
    .B(_12045_),
    .Y(_12081_));
 sg13g2_a21oi_2 _19761_ (.B1(_12081_),
    .Y(_12082_),
    .A2(_12080_),
    .A1(_12041_));
 sg13g2_xnor2_1 _19762_ (.Y(_12083_),
    .A(_12079_),
    .B(_12082_));
 sg13g2_xnor2_1 _19763_ (.Y(_12084_),
    .A(_12075_),
    .B(_12083_));
 sg13g2_nor2_1 _19764_ (.A(_12054_),
    .B(_12060_),
    .Y(_12085_));
 sg13g2_a21oi_1 _19765_ (.A1(_12054_),
    .A2(_12060_),
    .Y(_12086_),
    .B1(_12047_));
 sg13g2_nor2_1 _19766_ (.A(_11811_),
    .B(_11826_),
    .Y(_12087_));
 sg13g2_a21oi_1 _19767_ (.A1(net283),
    .A2(_11793_),
    .Y(_12088_),
    .B1(_12087_));
 sg13g2_a21o_1 _19768_ (.A2(_11826_),
    .A1(_11811_),
    .B1(_12088_),
    .X(_12089_));
 sg13g2_buf_1 _19769_ (.A(_12089_),
    .X(_12090_));
 sg13g2_a221oi_1 _19770_ (.B2(_11823_),
    .C1(_11778_),
    .B1(_11816_),
    .A1(net570),
    .Y(_12091_),
    .A2(_11773_));
 sg13g2_nand4_1 _19771_ (.B(_11767_),
    .C(_11796_),
    .A(_11783_),
    .Y(_12092_),
    .D(_11857_));
 sg13g2_buf_1 _19772_ (.A(_12092_),
    .X(_12093_));
 sg13g2_nand2_1 _19773_ (.Y(_12094_),
    .A(_11815_),
    .B(_11810_));
 sg13g2_xnor2_1 _19774_ (.Y(_12095_),
    .A(_12093_),
    .B(_12094_));
 sg13g2_xnor2_1 _19775_ (.Y(_12096_),
    .A(_12091_),
    .B(_12095_));
 sg13g2_xnor2_1 _19776_ (.Y(_12097_),
    .A(_09343_),
    .B(_09786_));
 sg13g2_xnor2_1 _19777_ (.Y(_12098_),
    .A(_11615_),
    .B(_12097_));
 sg13g2_xor2_1 _19778_ (.B(_09747_),
    .A(_09023_),
    .X(_12099_));
 sg13g2_xnor2_1 _19779_ (.Y(_12100_),
    .A(_11390_),
    .B(_12099_));
 sg13g2_nand2_1 _19780_ (.Y(_12101_),
    .A(_11711_),
    .B(_12100_));
 sg13g2_o21ai_1 _19781_ (.B1(_12101_),
    .Y(_12102_),
    .A1(net699),
    .A2(_12098_));
 sg13g2_xor2_1 _19782_ (.B(_11853_),
    .A(_00453_),
    .X(_12103_));
 sg13g2_nor2_1 _19783_ (.A(net800),
    .B(_12103_),
    .Y(_12104_));
 sg13g2_a21oi_1 _19784_ (.A1(net728),
    .A2(_12102_),
    .Y(_12105_),
    .B1(_12104_));
 sg13g2_nand2b_1 _19785_ (.Y(_12106_),
    .B(_08440_),
    .A_N(_00452_));
 sg13g2_o21ai_1 _19786_ (.B1(_12106_),
    .Y(_12107_),
    .A1(net726),
    .A2(_12105_));
 sg13g2_nand2_1 _19787_ (.Y(_12108_),
    .A(net631),
    .B(_12107_));
 sg13g2_o21ai_1 _19788_ (.B1(_12108_),
    .Y(_12109_),
    .A1(_11768_),
    .A2(_00451_));
 sg13g2_buf_1 _19789_ (.A(_12109_),
    .X(_12110_));
 sg13g2_nand2_1 _19790_ (.Y(_12111_),
    .A(net524),
    .B(_12110_));
 sg13g2_xor2_1 _19791_ (.B(_12111_),
    .A(_12096_),
    .X(_12112_));
 sg13g2_xnor2_1 _19792_ (.Y(_12113_),
    .A(_12090_),
    .B(_12112_));
 sg13g2_or3_1 _19793_ (.A(_12085_),
    .B(_12086_),
    .C(_12113_),
    .X(_12114_));
 sg13g2_o21ai_1 _19794_ (.B1(_12113_),
    .Y(_12115_),
    .A1(_12085_),
    .A2(_12086_));
 sg13g2_nand3_1 _19795_ (.B(_12114_),
    .C(_12115_),
    .A(_12084_),
    .Y(_12116_));
 sg13g2_buf_1 _19796_ (.A(_12116_),
    .X(_12117_));
 sg13g2_a21o_1 _19797_ (.A2(_12115_),
    .A1(_12114_),
    .B1(_12084_),
    .X(_12118_));
 sg13g2_buf_1 _19798_ (.A(_12118_),
    .X(_12119_));
 sg13g2_buf_1 _19799_ (.A(net468),
    .X(_12120_));
 sg13g2_nand2_1 _19800_ (.Y(_12121_),
    .A(net281),
    .B(net456));
 sg13g2_xnor2_1 _19801_ (.Y(_12122_),
    .A(_12050_),
    .B(_12048_));
 sg13g2_xnor2_1 _19802_ (.Y(_12123_),
    .A(_12121_),
    .B(_12122_));
 sg13g2_buf_1 _19803_ (.A(net458),
    .X(_12124_));
 sg13g2_nand2_1 _19804_ (.Y(_12125_),
    .A(net447),
    .B(net266));
 sg13g2_nand2_1 _19805_ (.Y(_12126_),
    .A(net457),
    .B(net281));
 sg13g2_xnor2_1 _19806_ (.Y(_12127_),
    .A(_12076_),
    .B(_12126_));
 sg13g2_xnor2_1 _19807_ (.Y(_12128_),
    .A(_12125_),
    .B(_12127_));
 sg13g2_buf_1 _19808_ (.A(_11783_),
    .X(_12129_));
 sg13g2_a21oi_1 _19809_ (.A1(_09947_),
    .A2(_11629_),
    .Y(_12130_),
    .B1(net697));
 sg13g2_a21o_1 _19810_ (.A2(_00399_),
    .A1(net697),
    .B1(_12130_),
    .X(_12131_));
 sg13g2_nand3b_1 _19811_ (.B(_09850_),
    .C(net725),
    .Y(_12132_),
    .A_N(_11440_));
 sg13g2_o21ai_1 _19812_ (.B1(_12132_),
    .Y(_12133_),
    .A1(net725),
    .A2(_12131_));
 sg13g2_buf_1 _19813_ (.A(_12133_),
    .X(_12134_));
 sg13g2_buf_1 _19814_ (.A(_12134_),
    .X(_12135_));
 sg13g2_and2_1 _19815_ (.A(_12024_),
    .B(_12032_),
    .X(_12136_));
 sg13g2_buf_1 _19816_ (.A(_12136_),
    .X(_12137_));
 sg13g2_buf_1 _19817_ (.A(_12137_),
    .X(_12138_));
 sg13g2_xnor2_1 _19818_ (.Y(_12139_),
    .A(net264),
    .B(net455));
 sg13g2_xnor2_1 _19819_ (.Y(_12140_),
    .A(_12128_),
    .B(_12139_));
 sg13g2_nand2b_1 _19820_ (.Y(_12141_),
    .B(net725),
    .A_N(_12013_));
 sg13g2_o21ai_1 _19821_ (.B1(_12141_),
    .Y(_12142_),
    .A1(net725),
    .A2(_12020_));
 sg13g2_buf_1 _19822_ (.A(_12142_),
    .X(_12143_));
 sg13g2_buf_1 _19823_ (.A(_12143_),
    .X(_12144_));
 sg13g2_xnor2_1 _19824_ (.Y(_12145_),
    .A(_09834_),
    .B(_09849_));
 sg13g2_mux2_1 _19825_ (.A0(_12145_),
    .A1(_00402_),
    .S(net302),
    .X(_12146_));
 sg13g2_nand2_1 _19826_ (.Y(_12147_),
    .A(net697),
    .B(_00400_));
 sg13g2_xnor2_1 _19827_ (.Y(_12148_),
    .A(_09931_),
    .B(_09946_));
 sg13g2_mux2_1 _19828_ (.A0(_00401_),
    .A1(_12148_),
    .S(net314),
    .X(_12149_));
 sg13g2_nand2_1 _19829_ (.Y(_12150_),
    .A(net684),
    .B(_12149_));
 sg13g2_a21oi_1 _19830_ (.A1(_12147_),
    .A2(_12150_),
    .Y(_12151_),
    .B1(net725));
 sg13g2_a21o_1 _19831_ (.A2(_12146_),
    .A1(net683),
    .B1(_12151_),
    .X(_12152_));
 sg13g2_buf_2 _19832_ (.A(_12152_),
    .X(_12153_));
 sg13g2_nor2_1 _19833_ (.A(net467),
    .B(_12153_),
    .Y(_12154_));
 sg13g2_nand3_1 _19834_ (.B(_12140_),
    .C(_12154_),
    .A(_12123_),
    .Y(_12155_));
 sg13g2_a21o_1 _19835_ (.A2(_12119_),
    .A1(_12117_),
    .B1(_12155_),
    .X(_12156_));
 sg13g2_nand3_1 _19836_ (.B(_12119_),
    .C(_12155_),
    .A(_12117_),
    .Y(_12157_));
 sg13g2_buf_1 _19837_ (.A(_12157_),
    .X(_12158_));
 sg13g2_nand3_1 _19838_ (.B(_12156_),
    .C(_12158_),
    .A(_12065_),
    .Y(_12159_));
 sg13g2_a21o_1 _19839_ (.A2(_12158_),
    .A1(_12156_),
    .B1(_12065_),
    .X(_12160_));
 sg13g2_nand2_1 _19840_ (.Y(_12161_),
    .A(net282),
    .B(net407));
 sg13g2_nand2_1 _19841_ (.Y(_12162_),
    .A(net458),
    .B(net281));
 sg13g2_nand2_1 _19842_ (.Y(_12163_),
    .A(_11998_),
    .B(_11946_));
 sg13g2_xnor2_1 _19843_ (.Y(_12164_),
    .A(_12162_),
    .B(_12163_));
 sg13g2_xnor2_1 _19844_ (.Y(_12165_),
    .A(_12161_),
    .B(_12164_));
 sg13g2_buf_1 _19845_ (.A(net457),
    .X(_12166_));
 sg13g2_nand2_2 _19846_ (.Y(_12167_),
    .A(_12134_),
    .B(net468));
 sg13g2_and2_1 _19847_ (.A(_08538_),
    .B(net630),
    .X(_12168_));
 sg13g2_buf_1 _19848_ (.A(_12168_),
    .X(_12169_));
 sg13g2_nor2_1 _19849_ (.A(_12143_),
    .B(net523),
    .Y(_12170_));
 sg13g2_a21oi_1 _19850_ (.A1(net683),
    .A2(_12146_),
    .Y(_12171_),
    .B1(_12151_));
 sg13g2_buf_1 _19851_ (.A(_12171_),
    .X(_12172_));
 sg13g2_a22oi_1 _19852_ (.Y(_12173_),
    .B1(_12170_),
    .B2(net280),
    .A2(_12167_),
    .A1(net467));
 sg13g2_and2_1 _19853_ (.A(_11979_),
    .B(_11986_),
    .X(_12174_));
 sg13g2_buf_1 _19854_ (.A(_12174_),
    .X(_12175_));
 sg13g2_nor2_1 _19855_ (.A(_12175_),
    .B(_12153_),
    .Y(_12176_));
 sg13g2_buf_1 _19856_ (.A(_12022_),
    .X(_12177_));
 sg13g2_nand2_1 _19857_ (.Y(_12178_),
    .A(_12022_),
    .B(net523));
 sg13g2_o21ai_1 _19858_ (.B1(_12178_),
    .Y(_12179_),
    .A1(net466),
    .A2(_12167_));
 sg13g2_xnor2_1 _19859_ (.Y(_12180_),
    .A(_12167_),
    .B(_12178_));
 sg13g2_a22oi_1 _19860_ (.Y(_12181_),
    .B1(_12180_),
    .B2(_12153_),
    .A2(_12179_),
    .A1(_12176_));
 sg13g2_o21ai_1 _19861_ (.B1(_12181_),
    .Y(_12182_),
    .A1(net446),
    .A2(_12173_));
 sg13g2_xor2_1 _19862_ (.B(_12182_),
    .A(_12165_),
    .X(_12183_));
 sg13g2_nand2_1 _19863_ (.Y(_12184_),
    .A(net466),
    .B(net264));
 sg13g2_nand2_1 _19864_ (.Y(_12185_),
    .A(net280),
    .B(net456));
 sg13g2_xnor2_1 _19865_ (.Y(_12186_),
    .A(_12184_),
    .B(_12185_));
 sg13g2_nor2_1 _19866_ (.A(_12128_),
    .B(_12186_),
    .Y(_12187_));
 sg13g2_xnor2_1 _19867_ (.Y(_12188_),
    .A(_12183_),
    .B(_12187_));
 sg13g2_a21oi_1 _19868_ (.A1(_12159_),
    .A2(_12160_),
    .Y(_12189_),
    .B1(_12188_));
 sg13g2_nand3_1 _19869_ (.B(_12160_),
    .C(_12188_),
    .A(_12159_),
    .Y(_12190_));
 sg13g2_nand2b_1 _19870_ (.Y(_12191_),
    .B(_12190_),
    .A_N(_12189_));
 sg13g2_xor2_1 _19871_ (.B(_12062_),
    .A(_11865_),
    .X(_12192_));
 sg13g2_xnor2_1 _19872_ (.Y(_12193_),
    .A(_12040_),
    .B(_12192_));
 sg13g2_a221oi_1 _19873_ (.B2(net569),
    .C1(_11778_),
    .B1(_11773_),
    .A1(_11878_),
    .Y(_12194_),
    .A2(_11885_));
 sg13g2_buf_1 _19874_ (.A(_12194_),
    .X(_12195_));
 sg13g2_and2_1 _19875_ (.A(_11829_),
    .B(_11835_),
    .X(_12196_));
 sg13g2_buf_1 _19876_ (.A(_12196_),
    .X(_12197_));
 sg13g2_a21o_1 _19877_ (.A2(_11812_),
    .A1(_11767_),
    .B1(_11813_),
    .X(_12198_));
 sg13g2_buf_1 _19878_ (.A(_12198_),
    .X(_12199_));
 sg13g2_nor2_1 _19879_ (.A(_12197_),
    .B(_12199_),
    .Y(_12200_));
 sg13g2_nand2_1 _19880_ (.Y(_12201_),
    .A(_11796_),
    .B(net630));
 sg13g2_buf_1 _19881_ (.A(_12201_),
    .X(_12202_));
 sg13g2_a21oi_1 _19882_ (.A1(_11782_),
    .A2(_11791_),
    .Y(_12203_),
    .B1(_12202_));
 sg13g2_o21ai_1 _19883_ (.B1(_12203_),
    .Y(_12204_),
    .A1(_12195_),
    .A2(_12200_));
 sg13g2_nand2_1 _19884_ (.Y(_12205_),
    .A(_12195_),
    .B(_12200_));
 sg13g2_nand2_1 _19885_ (.Y(_12206_),
    .A(_12204_),
    .B(_12205_));
 sg13g2_xnor2_1 _19886_ (.Y(_12207_),
    .A(_11840_),
    .B(_11842_));
 sg13g2_xnor2_1 _19887_ (.Y(_12208_),
    .A(_11838_),
    .B(_12207_));
 sg13g2_buf_1 _19888_ (.A(_11810_),
    .X(_12209_));
 sg13g2_nand2_1 _19889_ (.Y(_12210_),
    .A(net306),
    .B(net524));
 sg13g2_xnor2_1 _19890_ (.Y(_12211_),
    .A(_12208_),
    .B(_12210_));
 sg13g2_xnor2_1 _19891_ (.Y(_12212_),
    .A(_12206_),
    .B(_12211_));
 sg13g2_nor2_1 _19892_ (.A(_11943_),
    .B(_11944_),
    .Y(_12213_));
 sg13g2_xor2_1 _19893_ (.B(_12037_),
    .A(_11964_),
    .X(_12214_));
 sg13g2_xnor2_1 _19894_ (.Y(_12215_),
    .A(_12213_),
    .B(_12214_));
 sg13g2_nand2_1 _19895_ (.Y(_12216_),
    .A(_12212_),
    .B(_12215_));
 sg13g2_buf_1 _19896_ (.A(_11946_),
    .X(_12217_));
 sg13g2_nand2_1 _19897_ (.Y(_12218_),
    .A(net406),
    .B(net265));
 sg13g2_a221oi_1 _19898_ (.B2(net569),
    .C1(_11933_),
    .B1(_11927_),
    .A1(_11979_),
    .Y(_12219_),
    .A2(_11986_));
 sg13g2_buf_1 _19899_ (.A(_12219_),
    .X(_12220_));
 sg13g2_nand3_1 _19900_ (.B(net267),
    .C(_12220_),
    .A(net447),
    .Y(_12221_));
 sg13g2_a21oi_1 _19901_ (.A1(net447),
    .A2(net267),
    .Y(_12222_),
    .B1(_12220_));
 sg13g2_a21oi_1 _19902_ (.A1(_12218_),
    .A2(_12221_),
    .Y(_12223_),
    .B1(_12222_));
 sg13g2_nand2_1 _19903_ (.Y(_12224_),
    .A(net447),
    .B(_11960_));
 sg13g2_a21o_1 _19904_ (.A2(_11870_),
    .A1(net569),
    .B1(_11874_),
    .X(_12225_));
 sg13g2_buf_1 _19905_ (.A(_12225_),
    .X(_12226_));
 sg13g2_nor2_1 _19906_ (.A(net279),
    .B(_11913_),
    .Y(_12227_));
 sg13g2_xnor2_1 _19907_ (.Y(_12228_),
    .A(_12224_),
    .B(_12227_));
 sg13g2_xnor2_1 _19908_ (.Y(_12229_),
    .A(_11947_),
    .B(_12228_));
 sg13g2_and4_1 _19909_ (.A(net266),
    .B(net282),
    .C(_12022_),
    .D(net468),
    .X(_12230_));
 sg13g2_a21o_1 _19910_ (.A2(_12229_),
    .A1(_12223_),
    .B1(_12230_),
    .X(_12231_));
 sg13g2_o21ai_1 _19911_ (.B1(_12231_),
    .Y(_12232_),
    .A1(_12223_),
    .A2(_12229_));
 sg13g2_nor2_1 _19912_ (.A(_12212_),
    .B(_12215_),
    .Y(_12233_));
 sg13g2_a21oi_1 _19913_ (.A1(_12216_),
    .A2(_12232_),
    .Y(_12234_),
    .B1(_12233_));
 sg13g2_xor2_1 _19914_ (.B(_12234_),
    .A(_12193_),
    .X(_12235_));
 sg13g2_nor2_1 _19915_ (.A(net683),
    .B(_12131_),
    .Y(_12236_));
 sg13g2_nor2b_1 _19916_ (.A(_12236_),
    .B_N(_12132_),
    .Y(_12237_));
 sg13g2_buf_1 _19917_ (.A(_12237_),
    .X(_12238_));
 sg13g2_buf_1 _19918_ (.A(_12177_),
    .X(_12239_));
 sg13g2_nand3_1 _19919_ (.B(net455),
    .C(_12122_),
    .A(net454),
    .Y(_12240_));
 sg13g2_o21ai_1 _19920_ (.B1(_12240_),
    .Y(_12241_),
    .A1(net455),
    .A2(_12123_));
 sg13g2_xor2_1 _19921_ (.B(_12122_),
    .A(_12121_),
    .X(_12242_));
 sg13g2_o21ai_1 _19922_ (.B1(net454),
    .Y(_12243_),
    .A1(_12238_),
    .A2(_12242_));
 sg13g2_buf_1 _19923_ (.A(net456),
    .X(_12244_));
 sg13g2_a22oi_1 _19924_ (.Y(_12245_),
    .B1(_12243_),
    .B2(net445),
    .A2(_12241_),
    .A1(_12238_));
 sg13g2_o21ai_1 _19925_ (.B1(net280),
    .Y(_12246_),
    .A1(net445),
    .A2(_12122_));
 sg13g2_nand2b_1 _19926_ (.Y(_12247_),
    .B(_12246_),
    .A_N(_12184_));
 sg13g2_o21ai_1 _19927_ (.B1(_12247_),
    .Y(_12248_),
    .A1(_12153_),
    .A2(_12245_));
 sg13g2_xnor2_1 _19928_ (.Y(_12249_),
    .A(_12128_),
    .B(_12248_));
 sg13g2_nand2b_1 _19929_ (.Y(_12250_),
    .B(_12249_),
    .A_N(_12235_));
 sg13g2_nand2b_1 _19930_ (.Y(_12251_),
    .B(_12234_),
    .A_N(_12193_));
 sg13g2_a21o_1 _19931_ (.A2(_11828_),
    .A1(_11845_),
    .B1(_11863_),
    .X(_12252_));
 sg13g2_o21ai_1 _19932_ (.B1(_12252_),
    .Y(_12253_),
    .A1(_11845_),
    .A2(_11828_));
 sg13g2_xnor2_1 _19933_ (.Y(_12254_),
    .A(_12251_),
    .B(_12253_));
 sg13g2_xor2_1 _19934_ (.B(_12254_),
    .A(_12250_),
    .X(_12255_));
 sg13g2_xnor2_1 _19935_ (.Y(_12256_),
    .A(_12191_),
    .B(_12255_));
 sg13g2_xor2_1 _19936_ (.B(_12223_),
    .A(_12230_),
    .X(_12257_));
 sg13g2_xnor2_1 _19937_ (.Y(_12258_),
    .A(_12229_),
    .B(_12257_));
 sg13g2_nand2_1 _19938_ (.Y(_12259_),
    .A(_11836_),
    .B(_11800_));
 sg13g2_nand2_1 _19939_ (.Y(_12260_),
    .A(_11887_),
    .B(_11815_));
 sg13g2_nand2_1 _19940_ (.Y(_12261_),
    .A(_12259_),
    .B(_12260_));
 sg13g2_buf_1 _19941_ (.A(net569),
    .X(_12262_));
 sg13g2_a221oi_1 _19942_ (.B2(net522),
    .C1(_11778_),
    .B1(_11773_),
    .A1(_11904_),
    .Y(_12263_),
    .A2(_11911_));
 sg13g2_nor2_1 _19943_ (.A(_12259_),
    .B(_12260_),
    .Y(_12264_));
 sg13g2_a21oi_2 _19944_ (.B1(_12264_),
    .Y(_12265_),
    .A2(_12263_),
    .A1(_12261_));
 sg13g2_xor2_1 _19945_ (.B(_12200_),
    .A(_12203_),
    .X(_12266_));
 sg13g2_xnor2_1 _19946_ (.Y(_12267_),
    .A(_12195_),
    .B(_12266_));
 sg13g2_nand2_1 _19947_ (.Y(_12268_),
    .A(_11825_),
    .B(net524));
 sg13g2_xor2_1 _19948_ (.B(_12268_),
    .A(_12267_),
    .X(_12269_));
 sg13g2_xor2_1 _19949_ (.B(_12269_),
    .A(_12265_),
    .X(_12270_));
 sg13g2_nor2_1 _19950_ (.A(_12258_),
    .B(_12270_),
    .Y(_12271_));
 sg13g2_nand2_1 _19951_ (.Y(_12272_),
    .A(net458),
    .B(net267));
 sg13g2_a221oi_1 _19952_ (.B2(net522),
    .C1(_11874_),
    .B1(_11870_),
    .A1(_11915_),
    .Y(_12273_),
    .A2(_11923_));
 sg13g2_xnor2_1 _19953_ (.Y(_12274_),
    .A(_12273_),
    .B(_12220_));
 sg13g2_xnor2_1 _19954_ (.Y(_12275_),
    .A(_12272_),
    .B(_12274_));
 sg13g2_nand2_1 _19955_ (.Y(_12276_),
    .A(net457),
    .B(_11938_));
 sg13g2_a221oi_1 _19956_ (.B2(net570),
    .C1(_11933_),
    .B1(_11927_),
    .A1(_12024_),
    .Y(_12277_),
    .A2(_12032_));
 sg13g2_buf_1 _19957_ (.A(_12277_),
    .X(_12278_));
 sg13g2_a21oi_1 _19958_ (.A1(net458),
    .A2(_11876_),
    .Y(_12279_),
    .B1(_12278_));
 sg13g2_nand3_1 _19959_ (.B(net265),
    .C(_12278_),
    .A(net447),
    .Y(_12280_));
 sg13g2_o21ai_1 _19960_ (.B1(_12280_),
    .Y(_12281_),
    .A1(_12276_),
    .A2(_12279_));
 sg13g2_nor2b_1 _19961_ (.A(_12275_),
    .B_N(_12281_),
    .Y(_12282_));
 sg13g2_nand2_1 _19962_ (.Y(_12283_),
    .A(_12258_),
    .B(_12270_));
 sg13g2_o21ai_1 _19963_ (.B1(_12283_),
    .Y(_12284_),
    .A1(_12271_),
    .A2(_12282_));
 sg13g2_xor2_1 _19964_ (.B(_12215_),
    .A(_12212_),
    .X(_12285_));
 sg13g2_xnor2_1 _19965_ (.Y(_12286_),
    .A(_12232_),
    .B(_12285_));
 sg13g2_nand2b_1 _19966_ (.Y(_12287_),
    .B(_12286_),
    .A_N(_12284_));
 sg13g2_nor2_1 _19967_ (.A(_12208_),
    .B(_12210_),
    .Y(_12288_));
 sg13g2_nand2_1 _19968_ (.Y(_12289_),
    .A(_12208_),
    .B(_12210_));
 sg13g2_o21ai_1 _19969_ (.B1(_12289_),
    .Y(_12290_),
    .A1(_12206_),
    .A2(_12288_));
 sg13g2_nor2_1 _19970_ (.A(_12287_),
    .B(_12290_),
    .Y(_12291_));
 sg13g2_xor2_1 _19971_ (.B(_12286_),
    .A(_12284_),
    .X(_12292_));
 sg13g2_xnor2_1 _19972_ (.Y(_12293_),
    .A(_12242_),
    .B(_12154_));
 sg13g2_nor2b_1 _19973_ (.A(_12292_),
    .B_N(_12293_),
    .Y(_12294_));
 sg13g2_xnor2_1 _19974_ (.Y(_12295_),
    .A(_12249_),
    .B(_12235_));
 sg13g2_nor2_1 _19975_ (.A(_12294_),
    .B(_12295_),
    .Y(_12296_));
 sg13g2_xnor2_1 _19976_ (.Y(_12297_),
    .A(_12287_),
    .B(_12290_));
 sg13g2_nand2_1 _19977_ (.Y(_12298_),
    .A(_12294_),
    .B(_12295_));
 sg13g2_o21ai_1 _19978_ (.B1(_12298_),
    .Y(_12299_),
    .A1(_12296_),
    .A2(_12297_));
 sg13g2_nor2_1 _19979_ (.A(_12291_),
    .B(_12299_),
    .Y(_12300_));
 sg13g2_xor2_1 _19980_ (.B(_12300_),
    .A(_12256_),
    .X(_12301_));
 sg13g2_xnor2_1 _19981_ (.Y(_12302_),
    .A(_12294_),
    .B(_12297_));
 sg13g2_xnor2_1 _19982_ (.Y(_12303_),
    .A(_12295_),
    .B(_12302_));
 sg13g2_a21o_1 _19983_ (.A2(_12267_),
    .A1(_12265_),
    .B1(_12268_),
    .X(_12304_));
 sg13g2_o21ai_1 _19984_ (.B1(_12304_),
    .Y(_12305_),
    .A1(_12265_),
    .A2(_12267_));
 sg13g2_xnor2_1 _19985_ (.Y(_12306_),
    .A(_12270_),
    .B(_12282_));
 sg13g2_xor2_1 _19986_ (.B(_12306_),
    .A(_12258_),
    .X(_12307_));
 sg13g2_nand2_1 _19987_ (.Y(_12308_),
    .A(_11939_),
    .B(_11815_));
 sg13g2_nand2_1 _19988_ (.Y(_12309_),
    .A(_11887_),
    .B(_11800_));
 sg13g2_nand2_1 _19989_ (.Y(_12310_),
    .A(_12308_),
    .B(_12309_));
 sg13g2_a221oi_1 _19990_ (.B2(_11928_),
    .C1(_11778_),
    .B1(_11773_),
    .A1(_11915_),
    .Y(_12311_),
    .A2(_11923_));
 sg13g2_nor2_1 _19991_ (.A(_12308_),
    .B(_12309_),
    .Y(_12312_));
 sg13g2_a21oi_2 _19992_ (.B1(_12312_),
    .Y(_12313_),
    .A2(_12311_),
    .A1(_12310_));
 sg13g2_xnor2_1 _19993_ (.Y(_12314_),
    .A(_12259_),
    .B(_12260_));
 sg13g2_xor2_1 _19994_ (.B(_12314_),
    .A(_12263_),
    .X(_12315_));
 sg13g2_nand2_1 _19995_ (.Y(_12316_),
    .A(_11793_),
    .B(net524));
 sg13g2_xor2_1 _19996_ (.B(_12316_),
    .A(_12315_),
    .X(_12317_));
 sg13g2_xnor2_1 _19997_ (.Y(_12318_),
    .A(_12313_),
    .B(_12317_));
 sg13g2_xnor2_1 _19998_ (.Y(_12319_),
    .A(_12275_),
    .B(_12281_));
 sg13g2_nand2_1 _19999_ (.Y(_12320_),
    .A(_12318_),
    .B(_12319_));
 sg13g2_nand2_1 _20000_ (.Y(_12321_),
    .A(net458),
    .B(_11876_));
 sg13g2_o21ai_1 _20001_ (.B1(_12278_),
    .Y(_12322_),
    .A1(_12175_),
    .A2(_11902_));
 sg13g2_nand3b_1 _20002_ (.B(net457),
    .C(_11937_),
    .Y(_12323_),
    .A_N(_12278_));
 sg13g2_nand3_1 _20003_ (.B(_12322_),
    .C(_12323_),
    .A(_12321_),
    .Y(_12324_));
 sg13g2_a21o_1 _20004_ (.A2(_12323_),
    .A1(_12322_),
    .B1(_12321_),
    .X(_12325_));
 sg13g2_nand2_1 _20005_ (.Y(_12326_),
    .A(net457),
    .B(_11876_));
 sg13g2_a22oi_1 _20006_ (.Y(_12327_),
    .B1(net267),
    .B2(net468),
    .A2(_11960_),
    .A1(_12022_));
 sg13g2_nand4_1 _20007_ (.B(net468),
    .C(_11960_),
    .A(_12022_),
    .Y(_12328_),
    .D(net267));
 sg13g2_o21ai_1 _20008_ (.B1(_12328_),
    .Y(_12329_),
    .A1(_12326_),
    .A2(_12327_));
 sg13g2_nand3_1 _20009_ (.B(_12325_),
    .C(_12329_),
    .A(_12324_),
    .Y(_12330_));
 sg13g2_buf_1 _20010_ (.A(_12330_),
    .X(_12331_));
 sg13g2_nor2_1 _20011_ (.A(_12318_),
    .B(_12319_),
    .Y(_12332_));
 sg13g2_a21o_1 _20012_ (.A2(_12331_),
    .A1(_12320_),
    .B1(_12332_),
    .X(_12333_));
 sg13g2_nor2_1 _20013_ (.A(_12307_),
    .B(_12333_),
    .Y(_12334_));
 sg13g2_buf_1 _20014_ (.A(net266),
    .X(_12335_));
 sg13g2_nand2_1 _20015_ (.Y(_12336_),
    .A(net240),
    .B(net456));
 sg13g2_buf_1 _20016_ (.A(_12012_),
    .X(_12337_));
 sg13g2_nand2_1 _20017_ (.Y(_12338_),
    .A(net263),
    .B(net454));
 sg13g2_xnor2_1 _20018_ (.Y(_12339_),
    .A(_12336_),
    .B(_12338_));
 sg13g2_xnor2_1 _20019_ (.Y(_12340_),
    .A(_11989_),
    .B(_12339_));
 sg13g2_xor2_1 _20020_ (.B(_12333_),
    .A(_12307_),
    .X(_12341_));
 sg13g2_nor2b_1 _20021_ (.A(_12340_),
    .B_N(_12341_),
    .Y(_12342_));
 sg13g2_xnor2_1 _20022_ (.Y(_12343_),
    .A(_12305_),
    .B(_12334_));
 sg13g2_nand2b_1 _20023_ (.Y(_12344_),
    .B(_12343_),
    .A_N(_12342_));
 sg13g2_xnor2_1 _20024_ (.Y(_12345_),
    .A(_12292_),
    .B(_12293_));
 sg13g2_nor2b_1 _20025_ (.A(_12343_),
    .B_N(_12342_),
    .Y(_12346_));
 sg13g2_a221oi_1 _20026_ (.B2(_12345_),
    .C1(_12346_),
    .B1(_12344_),
    .A1(_12305_),
    .Y(_12347_),
    .A2(_12334_));
 sg13g2_xor2_1 _20027_ (.B(_12347_),
    .A(_12303_),
    .X(_12348_));
 sg13g2_a221oi_1 _20028_ (.B2(_11928_),
    .C1(_11778_),
    .B1(_11773_),
    .A1(_12024_),
    .Y(_12349_),
    .A2(_12032_));
 sg13g2_buf_1 _20029_ (.A(_12349_),
    .X(_12350_));
 sg13g2_a21oi_1 _20030_ (.A1(_11949_),
    .A2(_11956_),
    .Y(_12351_),
    .B1(_12202_));
 sg13g2_nand2_1 _20031_ (.Y(_12352_),
    .A(_11988_),
    .B(_11815_));
 sg13g2_nand2_1 _20032_ (.Y(_12353_),
    .A(_12350_),
    .B(_12351_));
 sg13g2_nand2_1 _20033_ (.Y(_12354_),
    .A(_12352_),
    .B(_12353_));
 sg13g2_o21ai_1 _20034_ (.B1(_12354_),
    .Y(_12355_),
    .A1(_12350_),
    .A2(_12351_));
 sg13g2_buf_1 _20035_ (.A(_12355_),
    .X(_12356_));
 sg13g2_nand2_1 _20036_ (.Y(_12357_),
    .A(net446),
    .B(net283));
 sg13g2_nand2_1 _20037_ (.Y(_12358_),
    .A(_11946_),
    .B(_11841_));
 sg13g2_nand2_1 _20038_ (.Y(_12359_),
    .A(net447),
    .B(net571));
 sg13g2_xnor2_1 _20039_ (.Y(_12360_),
    .A(_12358_),
    .B(_12359_));
 sg13g2_xnor2_1 _20040_ (.Y(_12361_),
    .A(_12357_),
    .B(_12360_));
 sg13g2_buf_1 _20041_ (.A(net407),
    .X(_12362_));
 sg13g2_buf_1 _20042_ (.A(_11848_),
    .X(_12363_));
 sg13g2_nand2_1 _20043_ (.Y(_12364_),
    .A(net363),
    .B(net505));
 sg13g2_o21ai_1 _20044_ (.B1(_12364_),
    .Y(_12365_),
    .A1(_12356_),
    .A2(_12361_));
 sg13g2_nand2_1 _20045_ (.Y(_12366_),
    .A(_12356_),
    .B(_12361_));
 sg13g2_nand2_1 _20046_ (.Y(_12367_),
    .A(_12365_),
    .B(_12366_));
 sg13g2_nand2_2 _20047_ (.Y(_12368_),
    .A(_11988_),
    .B(_11841_));
 sg13g2_nand2_2 _20048_ (.Y(_12369_),
    .A(net468),
    .B(net571));
 sg13g2_a21oi_1 _20049_ (.A1(_12368_),
    .A2(_12369_),
    .Y(_12370_),
    .B1(_12143_));
 sg13g2_nor2_1 _20050_ (.A(_12368_),
    .B(_12369_),
    .Y(_12371_));
 sg13g2_a21oi_2 _20051_ (.B1(_12371_),
    .Y(_12372_),
    .A2(_12370_),
    .A1(net283));
 sg13g2_xnor2_1 _20052_ (.Y(_12373_),
    .A(_12352_),
    .B(_12351_));
 sg13g2_xnor2_1 _20053_ (.Y(_12374_),
    .A(_12350_),
    .B(_12373_));
 sg13g2_nand2_1 _20054_ (.Y(_12375_),
    .A(_11946_),
    .B(net524));
 sg13g2_a21o_1 _20055_ (.A2(_12374_),
    .A1(_12372_),
    .B1(_12375_),
    .X(_12376_));
 sg13g2_o21ai_1 _20056_ (.B1(_12376_),
    .Y(_12377_),
    .A1(_12372_),
    .A2(_12374_));
 sg13g2_xnor2_1 _20057_ (.Y(_12378_),
    .A(_12361_),
    .B(_12364_));
 sg13g2_xnor2_1 _20058_ (.Y(_12379_),
    .A(_12356_),
    .B(_12378_));
 sg13g2_xor2_1 _20059_ (.B(_12375_),
    .A(_12374_),
    .X(_12380_));
 sg13g2_xor2_1 _20060_ (.B(_12380_),
    .A(_12372_),
    .X(_12381_));
 sg13g2_buf_1 _20061_ (.A(_12381_),
    .X(_12382_));
 sg13g2_buf_1 _20062_ (.A(net267),
    .X(_12383_));
 sg13g2_nor4_1 _20063_ (.A(net467),
    .B(net456),
    .C(net279),
    .D(net239),
    .Y(_12384_));
 sg13g2_nand2b_1 _20064_ (.Y(_12385_),
    .B(_12384_),
    .A_N(_12382_));
 sg13g2_nand4_1 _20065_ (.B(net455),
    .C(net239),
    .A(net454),
    .Y(_12386_),
    .D(_12382_));
 sg13g2_nand3_1 _20066_ (.B(net265),
    .C(net239),
    .A(net456),
    .Y(_12387_));
 sg13g2_buf_1 _20067_ (.A(_11902_),
    .X(_12388_));
 sg13g2_nand3_1 _20068_ (.B(net265),
    .C(net262),
    .A(net456),
    .Y(_12389_));
 sg13g2_mux2_1 _20069_ (.A0(_12387_),
    .A1(_12389_),
    .S(_12382_),
    .X(_12390_));
 sg13g2_buf_1 _20070_ (.A(net265),
    .X(_12391_));
 sg13g2_nor2_1 _20071_ (.A(_12022_),
    .B(_12137_),
    .Y(_12392_));
 sg13g2_nor2_1 _20072_ (.A(net238),
    .B(net262),
    .Y(_12393_));
 sg13g2_a22oi_1 _20073_ (.Y(_12394_),
    .B1(_12393_),
    .B2(net454),
    .A2(_12392_),
    .A1(net238));
 sg13g2_and4_1 _20074_ (.A(_12385_),
    .B(_12386_),
    .C(_12390_),
    .D(_12394_),
    .X(_12395_));
 sg13g2_xor2_1 _20075_ (.B(_12395_),
    .A(_12379_),
    .X(_12396_));
 sg13g2_nand2_1 _20076_ (.Y(_12397_),
    .A(_12377_),
    .B(_12396_));
 sg13g2_buf_1 _20077_ (.A(_12175_),
    .X(_12398_));
 sg13g2_o21ai_1 _20078_ (.B1(net444),
    .Y(_12399_),
    .A1(net467),
    .A2(net571));
 sg13g2_nand3_1 _20079_ (.B(net506),
    .C(_12399_),
    .A(_12120_),
    .Y(_12400_));
 sg13g2_o21ai_1 _20080_ (.B1(_12400_),
    .Y(_12401_),
    .A1(net467),
    .A2(_12352_));
 sg13g2_xnor2_1 _20081_ (.Y(_12402_),
    .A(_12368_),
    .B(_12369_));
 sg13g2_buf_1 _20082_ (.A(_12202_),
    .X(_12403_));
 sg13g2_nor2_1 _20083_ (.A(net467),
    .B(net504),
    .Y(_12404_));
 sg13g2_a22oi_1 _20084_ (.Y(_12405_),
    .B1(_12404_),
    .B2(net444),
    .A2(_12369_),
    .A1(net504));
 sg13g2_o21ai_1 _20085_ (.B1(_12368_),
    .Y(_12406_),
    .A1(net506),
    .A2(_12369_));
 sg13g2_nand3_1 _20086_ (.B(net268),
    .C(_12406_),
    .A(net466),
    .Y(_12407_));
 sg13g2_o21ai_1 _20087_ (.B1(_12407_),
    .Y(_12408_),
    .A1(net268),
    .A2(_12405_));
 sg13g2_a21oi_1 _20088_ (.A1(net467),
    .A2(_12402_),
    .Y(_12409_),
    .B1(_12408_));
 sg13g2_buf_1 _20089_ (.A(_12124_),
    .X(_12410_));
 sg13g2_o21ai_1 _20090_ (.B1(net405),
    .Y(_12411_),
    .A1(_12401_),
    .A2(_12409_));
 sg13g2_nand2_1 _20091_ (.Y(_12412_),
    .A(_12401_),
    .B(_12409_));
 sg13g2_nand2_1 _20092_ (.Y(_12413_),
    .A(_12411_),
    .B(_12412_));
 sg13g2_nand2_1 _20093_ (.Y(_12414_),
    .A(_11846_),
    .B(net630));
 sg13g2_buf_1 _20094_ (.A(_12414_),
    .X(_12415_));
 sg13g2_nand2_1 _20095_ (.Y(_12416_),
    .A(_12177_),
    .B(net238));
 sg13g2_xnor2_1 _20096_ (.Y(_12417_),
    .A(_12382_),
    .B(_12416_));
 sg13g2_nor2_1 _20097_ (.A(net521),
    .B(_12417_),
    .Y(_12418_));
 sg13g2_a21o_1 _20098_ (.A2(_11773_),
    .A1(net522),
    .B1(_11778_),
    .X(_12419_));
 sg13g2_buf_1 _20099_ (.A(_12419_),
    .X(_12420_));
 sg13g2_nand2_1 _20100_ (.Y(_12421_),
    .A(net444),
    .B(_12420_));
 sg13g2_nand3_1 _20101_ (.B(net505),
    .C(_12401_),
    .A(net405),
    .Y(_12422_));
 sg13g2_buf_1 _20102_ (.A(_12239_),
    .X(_12423_));
 sg13g2_buf_1 _20103_ (.A(net571),
    .X(_12424_));
 sg13g2_nand4_1 _20104_ (.B(net445),
    .C(net520),
    .A(net443),
    .Y(_12425_),
    .D(net506));
 sg13g2_a221oi_1 _20105_ (.B2(_12417_),
    .C1(_12425_),
    .B1(_12422_),
    .A1(_12357_),
    .Y(_12426_),
    .A2(_12421_));
 sg13g2_a21o_1 _20106_ (.A2(_12418_),
    .A1(_12413_),
    .B1(_12426_),
    .X(_12427_));
 sg13g2_o21ai_1 _20107_ (.B1(_12427_),
    .Y(_12428_),
    .A1(_12377_),
    .A2(_12396_));
 sg13g2_nand3_1 _20108_ (.B(_12397_),
    .C(_12428_),
    .A(_12367_),
    .Y(_12429_));
 sg13g2_nand2_1 _20109_ (.Y(_12430_),
    .A(net466),
    .B(_12034_));
 sg13g2_xnor2_1 _20110_ (.Y(_12431_),
    .A(net446),
    .B(_12071_));
 sg13g2_nor4_2 _20111_ (.A(net279),
    .B(_11902_),
    .C(_12430_),
    .Y(_12432_),
    .D(_12431_));
 sg13g2_a221oi_1 _20112_ (.B2(net522),
    .C1(_11778_),
    .B1(_11773_),
    .A1(_11949_),
    .Y(_12433_),
    .A2(_11956_));
 sg13g2_nand2_1 _20113_ (.Y(_12434_),
    .A(_11946_),
    .B(net571));
 sg13g2_nand2_1 _20114_ (.Y(_12435_),
    .A(_11939_),
    .B(net506));
 sg13g2_nand2_1 _20115_ (.Y(_12436_),
    .A(_12434_),
    .B(_12435_));
 sg13g2_nor2_1 _20116_ (.A(_12434_),
    .B(_12435_),
    .Y(_12437_));
 sg13g2_a21oi_2 _20117_ (.B1(_12437_),
    .Y(_12438_),
    .A2(_12436_),
    .A1(_12433_));
 sg13g2_nor2_1 _20118_ (.A(_12197_),
    .B(_12414_),
    .Y(_12439_));
 sg13g2_xor2_1 _20119_ (.B(_12309_),
    .A(_12308_),
    .X(_12440_));
 sg13g2_xnor2_1 _20120_ (.Y(_12441_),
    .A(_12311_),
    .B(_12440_));
 sg13g2_xnor2_1 _20121_ (.Y(_12442_),
    .A(_12439_),
    .B(_12441_));
 sg13g2_xor2_1 _20122_ (.B(_12442_),
    .A(_12438_),
    .X(_12443_));
 sg13g2_a21o_1 _20123_ (.A2(_12325_),
    .A1(_12324_),
    .B1(_12329_),
    .X(_12444_));
 sg13g2_buf_1 _20124_ (.A(_12444_),
    .X(_12445_));
 sg13g2_nand3_1 _20125_ (.B(_12443_),
    .C(_12445_),
    .A(_12331_),
    .Y(_12446_));
 sg13g2_a21o_1 _20126_ (.A2(_12445_),
    .A1(_12331_),
    .B1(_12443_),
    .X(_12447_));
 sg13g2_nand3_1 _20127_ (.B(_12446_),
    .C(_12447_),
    .A(_12432_),
    .Y(_12448_));
 sg13g2_buf_1 _20128_ (.A(_12448_),
    .X(_12449_));
 sg13g2_a21o_1 _20129_ (.A2(_12447_),
    .A1(_12446_),
    .B1(_12432_),
    .X(_12450_));
 sg13g2_buf_1 _20130_ (.A(_12450_),
    .X(_12451_));
 sg13g2_buf_1 _20131_ (.A(net282),
    .X(_12452_));
 sg13g2_nand2_1 _20132_ (.Y(_12453_),
    .A(net261),
    .B(net466));
 sg13g2_inv_1 _20133_ (.Y(_12454_),
    .A(_12453_));
 sg13g2_a21oi_1 _20134_ (.A1(_12034_),
    .A2(net239),
    .Y(_12455_),
    .B1(net466));
 sg13g2_buf_1 _20135_ (.A(_11960_),
    .X(_12456_));
 sg13g2_nor3_1 _20136_ (.A(_12143_),
    .B(net279),
    .C(net260),
    .Y(_12457_));
 sg13g2_o21ai_1 _20137_ (.B1(net444),
    .Y(_12458_),
    .A1(_12455_),
    .A2(_12457_));
 sg13g2_a22oi_1 _20138_ (.Y(_12459_),
    .B1(net239),
    .B2(_12392_),
    .A2(net260),
    .A1(net466));
 sg13g2_or2_1 _20139_ (.X(_12460_),
    .B(_12459_),
    .A(_12326_));
 sg13g2_nor4_1 _20140_ (.A(_12143_),
    .B(net455),
    .C(_12071_),
    .D(_11902_),
    .Y(_12461_));
 sg13g2_o21ai_1 _20141_ (.B1(net279),
    .Y(_12462_),
    .A1(_12327_),
    .A2(_12461_));
 sg13g2_nand3_1 _20142_ (.B(_12460_),
    .C(_12462_),
    .A(_12458_),
    .Y(_12463_));
 sg13g2_nand4_1 _20143_ (.B(net446),
    .C(_11780_),
    .A(net447),
    .Y(_12464_),
    .D(net571));
 sg13g2_a22oi_1 _20144_ (.Y(_12465_),
    .B1(_11839_),
    .B2(net447),
    .A2(_11780_),
    .A1(net446));
 sg13g2_a21o_1 _20145_ (.A2(_12464_),
    .A1(_12358_),
    .B1(_12465_),
    .X(_12466_));
 sg13g2_buf_1 _20146_ (.A(_12466_),
    .X(_12467_));
 sg13g2_nand2_1 _20147_ (.Y(_12468_),
    .A(_11887_),
    .B(net524));
 sg13g2_xor2_1 _20148_ (.B(_12435_),
    .A(_12434_),
    .X(_12469_));
 sg13g2_xnor2_1 _20149_ (.Y(_12470_),
    .A(_12433_),
    .B(_12469_));
 sg13g2_xnor2_1 _20150_ (.Y(_12471_),
    .A(_12468_),
    .B(_12470_));
 sg13g2_xnor2_1 _20151_ (.Y(_12472_),
    .A(_12467_),
    .B(_12471_));
 sg13g2_nor2_1 _20152_ (.A(_12463_),
    .B(_12472_),
    .Y(_12473_));
 sg13g2_xnor2_1 _20153_ (.Y(_12474_),
    .A(_12454_),
    .B(_12473_));
 sg13g2_nand3_1 _20154_ (.B(_12451_),
    .C(_12474_),
    .A(_12449_),
    .Y(_12475_));
 sg13g2_buf_1 _20155_ (.A(_12475_),
    .X(_12476_));
 sg13g2_a21o_1 _20156_ (.A2(_12451_),
    .A1(_12449_),
    .B1(_12474_),
    .X(_12477_));
 sg13g2_buf_1 _20157_ (.A(_12477_),
    .X(_12478_));
 sg13g2_and2_1 _20158_ (.A(_12476_),
    .B(_12478_),
    .X(_12479_));
 sg13g2_o21ai_1 _20159_ (.B1(_12468_),
    .Y(_12480_),
    .A1(_12467_),
    .A2(_12470_));
 sg13g2_nand2_1 _20160_ (.Y(_12481_),
    .A(_12467_),
    .B(_12470_));
 sg13g2_and2_1 _20161_ (.A(_12480_),
    .B(_12481_),
    .X(_12482_));
 sg13g2_xnor2_1 _20162_ (.Y(_12483_),
    .A(_12463_),
    .B(_12472_));
 sg13g2_nand2_1 _20163_ (.Y(_12484_),
    .A(net454),
    .B(net239));
 sg13g2_nor2_1 _20164_ (.A(_12138_),
    .B(net279),
    .Y(_12485_));
 sg13g2_xnor2_1 _20165_ (.Y(_12486_),
    .A(_12484_),
    .B(_12485_));
 sg13g2_nand2b_1 _20166_ (.Y(_12487_),
    .B(_12486_),
    .A_N(_12379_));
 sg13g2_nor2_1 _20167_ (.A(_12483_),
    .B(_12487_),
    .Y(_12488_));
 sg13g2_xnor2_1 _20168_ (.Y(_12489_),
    .A(_12482_),
    .B(_12488_));
 sg13g2_xnor2_1 _20169_ (.Y(_12490_),
    .A(_12479_),
    .B(_12489_));
 sg13g2_xor2_1 _20170_ (.B(_12487_),
    .A(_12483_),
    .X(_12491_));
 sg13g2_xnor2_1 _20171_ (.Y(_12492_),
    .A(_12138_),
    .B(net262));
 sg13g2_xnor2_1 _20172_ (.Y(_12493_),
    .A(_12379_),
    .B(_12492_));
 sg13g2_nor3_1 _20173_ (.A(_12382_),
    .B(_12416_),
    .C(_12493_),
    .Y(_12494_));
 sg13g2_or2_1 _20174_ (.X(_12495_),
    .B(_12494_),
    .A(_12491_));
 sg13g2_nand3_1 _20175_ (.B(_12490_),
    .C(_12495_),
    .A(_12429_),
    .Y(_12496_));
 sg13g2_inv_1 _20176_ (.Y(_12497_),
    .A(_12482_));
 sg13g2_nand3_1 _20177_ (.B(_12476_),
    .C(_12478_),
    .A(_12488_),
    .Y(_12498_));
 sg13g2_a21oi_1 _20178_ (.A1(_12476_),
    .A2(_12478_),
    .Y(_12499_),
    .B1(_12488_));
 sg13g2_a21oi_1 _20179_ (.A1(_12497_),
    .A2(_12498_),
    .Y(_12500_),
    .B1(_12499_));
 sg13g2_xnor2_1 _20180_ (.Y(_12501_),
    .A(_12438_),
    .B(_12442_));
 sg13g2_nor2_1 _20181_ (.A(_12432_),
    .B(_12501_),
    .Y(_12502_));
 sg13g2_a22oi_1 _20182_ (.Y(_12503_),
    .B1(_12445_),
    .B2(_12331_),
    .A2(_12501_),
    .A1(_12432_));
 sg13g2_nand2_1 _20183_ (.Y(_12504_),
    .A(_11977_),
    .B(net456));
 sg13g2_nand2_1 _20184_ (.Y(_12505_),
    .A(net266),
    .B(net466));
 sg13g2_xor2_1 _20185_ (.B(_12505_),
    .A(_12504_),
    .X(_12506_));
 sg13g2_o21ai_1 _20186_ (.B1(_12506_),
    .Y(_12507_),
    .A1(_12502_),
    .A2(_12503_));
 sg13g2_or3_1 _20187_ (.A(_12502_),
    .B(_12503_),
    .C(_12506_),
    .X(_12508_));
 sg13g2_xor2_1 _20188_ (.B(_12331_),
    .A(_12319_),
    .X(_12509_));
 sg13g2_xnor2_1 _20189_ (.Y(_12510_),
    .A(_12318_),
    .B(_12509_));
 sg13g2_a21o_1 _20190_ (.A2(_12508_),
    .A1(_12507_),
    .B1(_12510_),
    .X(_12511_));
 sg13g2_buf_1 _20191_ (.A(_12511_),
    .X(_12512_));
 sg13g2_nand3_1 _20192_ (.B(_12507_),
    .C(_12508_),
    .A(_12510_),
    .Y(_12513_));
 sg13g2_nor2_1 _20193_ (.A(_12438_),
    .B(_12441_),
    .Y(_12514_));
 sg13g2_nor2_1 _20194_ (.A(_12439_),
    .B(_12514_),
    .Y(_12515_));
 sg13g2_a21oi_1 _20195_ (.A1(_12438_),
    .A2(_12441_),
    .Y(_12516_),
    .B1(_12515_));
 sg13g2_inv_1 _20196_ (.Y(_12517_),
    .A(_12516_));
 sg13g2_a21oi_1 _20197_ (.A1(_12512_),
    .A2(_12513_),
    .Y(_12518_),
    .B1(_12517_));
 sg13g2_and3_1 _20198_ (.X(_12519_),
    .A(_12512_),
    .B(_12513_),
    .C(_12517_));
 sg13g2_inv_1 _20199_ (.Y(_12520_),
    .A(_12473_));
 sg13g2_nand3_1 _20200_ (.B(_12451_),
    .C(_12520_),
    .A(_12449_),
    .Y(_12521_));
 sg13g2_a21oi_1 _20201_ (.A1(_12449_),
    .A2(_12451_),
    .Y(_12522_),
    .B1(_12520_));
 sg13g2_a21oi_2 _20202_ (.B1(_12522_),
    .Y(_12523_),
    .A2(_12521_),
    .A1(_12454_));
 sg13g2_o21ai_1 _20203_ (.B1(_12523_),
    .Y(_12524_),
    .A1(_12518_),
    .A2(_12519_));
 sg13g2_or3_1 _20204_ (.A(_12523_),
    .B(_12518_),
    .C(_12519_),
    .X(_12525_));
 sg13g2_nand3_1 _20205_ (.B(_12524_),
    .C(_12525_),
    .A(_12500_),
    .Y(_12526_));
 sg13g2_and2_1 _20206_ (.A(_12491_),
    .B(_12494_),
    .X(_12527_));
 sg13g2_a21oi_1 _20207_ (.A1(_12397_),
    .A2(_12428_),
    .Y(_12528_),
    .B1(_12367_));
 sg13g2_nand2_1 _20208_ (.Y(_12529_),
    .A(_12527_),
    .B(_12528_));
 sg13g2_o21ai_1 _20209_ (.B1(_12490_),
    .Y(_12530_),
    .A1(_12527_),
    .A2(_12528_));
 sg13g2_nand4_1 _20210_ (.B(_12526_),
    .C(_12529_),
    .A(_12496_),
    .Y(_12531_),
    .D(_12530_));
 sg13g2_a21o_1 _20211_ (.A2(_12525_),
    .A1(_12524_),
    .B1(_12500_),
    .X(_12532_));
 sg13g2_and2_1 _20212_ (.A(_12512_),
    .B(_12513_),
    .X(_12533_));
 sg13g2_nor2_1 _20213_ (.A(_12523_),
    .B(_12533_),
    .Y(_12534_));
 sg13g2_a21oi_1 _20214_ (.A1(_12523_),
    .A2(_12533_),
    .Y(_12535_),
    .B1(_12517_));
 sg13g2_nor2_1 _20215_ (.A(_12534_),
    .B(_12535_),
    .Y(_12536_));
 sg13g2_xnor2_1 _20216_ (.Y(_12537_),
    .A(_12340_),
    .B(_12341_));
 sg13g2_or2_1 _20217_ (.X(_12538_),
    .B(_12503_),
    .A(_12502_));
 sg13g2_nor2_1 _20218_ (.A(_12506_),
    .B(_12510_),
    .Y(_12539_));
 sg13g2_nand2_1 _20219_ (.Y(_12540_),
    .A(_12506_),
    .B(_12510_));
 sg13g2_o21ai_1 _20220_ (.B1(_12540_),
    .Y(_12541_),
    .A1(_12538_),
    .A2(_12539_));
 sg13g2_a21o_1 _20221_ (.A2(_12315_),
    .A1(_12313_),
    .B1(_12316_),
    .X(_12542_));
 sg13g2_o21ai_1 _20222_ (.B1(_12542_),
    .Y(_12543_),
    .A1(_12313_),
    .A2(_12315_));
 sg13g2_buf_1 _20223_ (.A(_12543_),
    .X(_12544_));
 sg13g2_xor2_1 _20224_ (.B(_12544_),
    .A(_12541_),
    .X(_12545_));
 sg13g2_xnor2_1 _20225_ (.Y(_12546_),
    .A(_12537_),
    .B(_12545_));
 sg13g2_nor2_1 _20226_ (.A(_12536_),
    .B(_12546_),
    .Y(_12547_));
 sg13g2_a21oi_1 _20227_ (.A1(_12531_),
    .A2(_12532_),
    .Y(_12548_),
    .B1(_12547_));
 sg13g2_xor2_1 _20228_ (.B(_12343_),
    .A(_12342_),
    .X(_12549_));
 sg13g2_xnor2_1 _20229_ (.Y(_12550_),
    .A(_12345_),
    .B(_12549_));
 sg13g2_nand2_1 _20230_ (.Y(_12551_),
    .A(_12537_),
    .B(_12544_));
 sg13g2_o21ai_1 _20231_ (.B1(_12541_),
    .Y(_12552_),
    .A1(_12537_),
    .A2(_12544_));
 sg13g2_nand2_1 _20232_ (.Y(_12553_),
    .A(_12551_),
    .B(_12552_));
 sg13g2_a22oi_1 _20233_ (.Y(_12554_),
    .B1(_12546_),
    .B2(_12536_),
    .A2(_12553_),
    .A1(_12550_));
 sg13g2_o21ai_1 _20234_ (.B1(_12554_),
    .Y(_12555_),
    .A1(_12550_),
    .A2(_12553_));
 sg13g2_nand2_1 _20235_ (.Y(_12556_),
    .A(_12550_),
    .B(_12553_));
 sg13g2_o21ai_1 _20236_ (.B1(_12556_),
    .Y(_12557_),
    .A1(_12548_),
    .A2(_12555_));
 sg13g2_buf_1 _20237_ (.A(_12557_),
    .X(_12558_));
 sg13g2_nor2_1 _20238_ (.A(_12303_),
    .B(_12347_),
    .Y(_12559_));
 sg13g2_a21oi_1 _20239_ (.A1(_12348_),
    .A2(_12558_),
    .Y(_12560_),
    .B1(_12559_));
 sg13g2_a21o_1 _20240_ (.A2(_12191_),
    .A1(_12250_),
    .B1(_12254_),
    .X(_12561_));
 sg13g2_o21ai_1 _20241_ (.B1(_12561_),
    .Y(_12562_),
    .A1(_12250_),
    .A2(_12191_));
 sg13g2_nor2_1 _20242_ (.A(_12251_),
    .B(_12253_),
    .Y(_12563_));
 sg13g2_nand2_1 _20243_ (.Y(_12564_),
    .A(_12084_),
    .B(_12113_));
 sg13g2_or2_1 _20244_ (.X(_12565_),
    .B(_12086_),
    .A(_12085_));
 sg13g2_o21ai_1 _20245_ (.B1(_12565_),
    .Y(_12566_),
    .A1(_12084_),
    .A2(_12113_));
 sg13g2_and2_1 _20246_ (.A(_12564_),
    .B(_12566_),
    .X(_12567_));
 sg13g2_buf_1 _20247_ (.A(_12567_),
    .X(_12568_));
 sg13g2_nand2_1 _20248_ (.Y(_12569_),
    .A(_12183_),
    .B(_12187_));
 sg13g2_nand2_1 _20249_ (.Y(_12570_),
    .A(net265),
    .B(_11825_));
 sg13g2_nand2_1 _20250_ (.Y(_12571_),
    .A(_11938_),
    .B(_11793_));
 sg13g2_nand2_1 _20251_ (.Y(_12572_),
    .A(net260),
    .B(net333));
 sg13g2_xnor2_1 _20252_ (.Y(_12573_),
    .A(_12571_),
    .B(_12572_));
 sg13g2_xnor2_1 _20253_ (.Y(_12574_),
    .A(_12570_),
    .B(_12573_));
 sg13g2_and2_1 _20254_ (.A(_12161_),
    .B(_12163_),
    .X(_12575_));
 sg13g2_or2_1 _20255_ (.X(_12576_),
    .B(_12163_),
    .A(_12161_));
 sg13g2_o21ai_1 _20256_ (.B1(_12576_),
    .Y(_12577_),
    .A1(_12162_),
    .A2(_12575_));
 sg13g2_buf_1 _20257_ (.A(_12577_),
    .X(_12578_));
 sg13g2_nand2b_1 _20258_ (.Y(_12579_),
    .B(_12072_),
    .A_N(_12067_));
 sg13g2_a21oi_1 _20259_ (.A1(net265),
    .A2(_11793_),
    .Y(_12580_),
    .B1(_12072_));
 sg13g2_a21oi_1 _20260_ (.A1(_12073_),
    .A2(_12579_),
    .Y(_12581_),
    .B1(_12580_));
 sg13g2_xnor2_1 _20261_ (.Y(_12582_),
    .A(_12578_),
    .B(_12581_));
 sg13g2_xor2_1 _20262_ (.B(_12582_),
    .A(_12574_),
    .X(_12583_));
 sg13g2_nand2_1 _20263_ (.Y(_12584_),
    .A(_12079_),
    .B(_12082_));
 sg13g2_nor2_1 _20264_ (.A(_12079_),
    .B(_12082_),
    .Y(_12585_));
 sg13g2_a21o_1 _20265_ (.A2(_12584_),
    .A1(_12075_),
    .B1(_12585_),
    .X(_12586_));
 sg13g2_nand2_1 _20266_ (.Y(_12587_),
    .A(net283),
    .B(_11810_));
 sg13g2_and2_1 _20267_ (.A(_11800_),
    .B(_12110_),
    .X(_12588_));
 sg13g2_buf_1 _20268_ (.A(_12588_),
    .X(_12589_));
 sg13g2_and2_1 _20269_ (.A(net571),
    .B(_11862_),
    .X(_12590_));
 sg13g2_buf_1 _20270_ (.A(_12590_),
    .X(_12591_));
 sg13g2_xor2_1 _20271_ (.B(_12591_),
    .A(_12589_),
    .X(_12592_));
 sg13g2_xnor2_1 _20272_ (.Y(_12593_),
    .A(_12587_),
    .B(_12592_));
 sg13g2_nor2_1 _20273_ (.A(_12093_),
    .B(_12094_),
    .Y(_12594_));
 sg13g2_nor2_1 _20274_ (.A(_12091_),
    .B(_12594_),
    .Y(_12595_));
 sg13g2_a21oi_2 _20275_ (.B1(_12595_),
    .Y(_12596_),
    .A2(_12094_),
    .A1(_12093_));
 sg13g2_nor4_1 _20276_ (.A(_09343_),
    .B(_11606_),
    .C(_11610_),
    .D(_11614_),
    .Y(_12597_));
 sg13g2_or2_1 _20277_ (.X(_12598_),
    .B(_12597_),
    .A(_11616_));
 sg13g2_xor2_1 _20278_ (.B(_12598_),
    .A(_09357_),
    .X(_12599_));
 sg13g2_nand3b_1 _20279_ (.B(_09747_),
    .C(_11390_),
    .Y(_12600_),
    .A_N(_09023_));
 sg13g2_o21ai_1 _20280_ (.B1(_12600_),
    .Y(_12601_),
    .A1(_11390_),
    .A2(_11434_));
 sg13g2_xor2_1 _20281_ (.B(_12601_),
    .A(_09037_),
    .X(_12602_));
 sg13g2_mux2_1 _20282_ (.A0(_12599_),
    .A1(_12602_),
    .S(_11712_),
    .X(_12603_));
 sg13g2_o21ai_1 _20283_ (.B1(_00453_),
    .Y(_12604_),
    .A1(_11760_),
    .A2(_11853_));
 sg13g2_xor2_1 _20284_ (.B(_12604_),
    .A(_11727_),
    .X(_12605_));
 sg13g2_nor2_1 _20285_ (.A(net728),
    .B(_12605_),
    .Y(_12606_));
 sg13g2_a21oi_1 _20286_ (.A1(net728),
    .A2(_12603_),
    .Y(_12607_),
    .B1(_12606_));
 sg13g2_mux2_1 _20287_ (.A0(_00455_),
    .A1(_12607_),
    .S(net697),
    .X(_12608_));
 sg13g2_nand2b_1 _20288_ (.Y(_12609_),
    .B(_08445_),
    .A_N(_00454_));
 sg13g2_o21ai_1 _20289_ (.B1(_12609_),
    .Y(_12610_),
    .A1(_08445_),
    .A2(_12608_));
 sg13g2_buf_1 _20290_ (.A(_12610_),
    .X(_12611_));
 sg13g2_nand2_1 _20291_ (.Y(_12612_),
    .A(net524),
    .B(_12611_));
 sg13g2_xor2_1 _20292_ (.B(_12612_),
    .A(_12596_),
    .X(_12613_));
 sg13g2_xnor2_1 _20293_ (.Y(_12614_),
    .A(_12593_),
    .B(_12613_));
 sg13g2_xor2_1 _20294_ (.B(_12614_),
    .A(_12586_),
    .X(_12615_));
 sg13g2_xnor2_1 _20295_ (.Y(_12616_),
    .A(_12583_),
    .B(_12615_));
 sg13g2_xor2_1 _20296_ (.B(_12616_),
    .A(_12569_),
    .X(_12617_));
 sg13g2_xnor2_1 _20297_ (.Y(_12618_),
    .A(_12568_),
    .B(_12617_));
 sg13g2_xnor2_1 _20298_ (.Y(_12619_),
    .A(net444),
    .B(net523));
 sg13g2_nor3_1 _20299_ (.A(_12238_),
    .B(_12430_),
    .C(_12619_),
    .Y(_12620_));
 sg13g2_nor2_1 _20300_ (.A(_12165_),
    .B(_12182_),
    .Y(_12621_));
 sg13g2_a21oi_1 _20301_ (.A1(net280),
    .A2(_12620_),
    .Y(_12622_),
    .B1(_12621_));
 sg13g2_nand2_1 _20302_ (.Y(_12623_),
    .A(net282),
    .B(_11887_));
 sg13g2_nand2_1 _20303_ (.Y(_12624_),
    .A(net266),
    .B(net407));
 sg13g2_nand2_1 _20304_ (.Y(_12625_),
    .A(net406),
    .B(net281));
 sg13g2_xnor2_1 _20305_ (.Y(_12626_),
    .A(_12624_),
    .B(_12625_));
 sg13g2_xnor2_1 _20306_ (.Y(_12627_),
    .A(_12623_),
    .B(_12626_));
 sg13g2_nand2_1 _20307_ (.Y(_12628_),
    .A(net405),
    .B(net280));
 sg13g2_nand2_1 _20308_ (.Y(_12629_),
    .A(_08538_),
    .B(net630));
 sg13g2_buf_2 _20309_ (.A(_12629_),
    .X(_12630_));
 sg13g2_nor2_1 _20310_ (.A(net455),
    .B(_12630_),
    .Y(_12631_));
 sg13g2_nand2_1 _20311_ (.Y(_12632_),
    .A(net446),
    .B(_12134_));
 sg13g2_xor2_1 _20312_ (.B(_12632_),
    .A(_12631_),
    .X(_12633_));
 sg13g2_xnor2_1 _20313_ (.Y(_12634_),
    .A(_12628_),
    .B(_12633_));
 sg13g2_nand2_1 _20314_ (.Y(_12635_),
    .A(_12167_),
    .B(_12178_));
 sg13g2_nor2_1 _20315_ (.A(_12167_),
    .B(_12178_),
    .Y(_12636_));
 sg13g2_a21oi_1 _20316_ (.A1(_12176_),
    .A2(_12635_),
    .Y(_12637_),
    .B1(_12636_));
 sg13g2_xnor2_1 _20317_ (.Y(_12638_),
    .A(_12634_),
    .B(_12637_));
 sg13g2_xnor2_1 _20318_ (.Y(_12639_),
    .A(_12627_),
    .B(_12638_));
 sg13g2_xnor2_1 _20319_ (.Y(_12640_),
    .A(_12622_),
    .B(_12639_));
 sg13g2_and2_1 _20320_ (.A(_08537_),
    .B(net630),
    .X(_12641_));
 sg13g2_buf_2 _20321_ (.A(_12641_),
    .X(_12642_));
 sg13g2_nand2_2 _20322_ (.Y(_12643_),
    .A(net443),
    .B(_12642_));
 sg13g2_xor2_1 _20323_ (.B(_12643_),
    .A(_12640_),
    .X(_12644_));
 sg13g2_xor2_1 _20324_ (.B(_12644_),
    .A(_12618_),
    .X(_12645_));
 sg13g2_a21o_1 _20325_ (.A2(_12063_),
    .A1(_11865_),
    .B1(_12064_),
    .X(_12646_));
 sg13g2_a21oi_1 _20326_ (.A1(_12117_),
    .A2(_12119_),
    .Y(_12647_),
    .B1(_12155_));
 sg13g2_o21ai_1 _20327_ (.B1(_12158_),
    .Y(_12648_),
    .A1(_12646_),
    .A2(_12647_));
 sg13g2_nor2b_1 _20328_ (.A(_12096_),
    .B_N(_12090_),
    .Y(_12649_));
 sg13g2_nand2b_1 _20329_ (.Y(_12650_),
    .B(_12096_),
    .A_N(_12090_));
 sg13g2_o21ai_1 _20330_ (.B1(_12650_),
    .Y(_12651_),
    .A1(_12111_),
    .A2(_12649_));
 sg13g2_xnor2_1 _20331_ (.Y(_12652_),
    .A(_12648_),
    .B(_12651_));
 sg13g2_xnor2_1 _20332_ (.Y(_12653_),
    .A(_12189_),
    .B(_12652_));
 sg13g2_xnor2_1 _20333_ (.Y(_12654_),
    .A(_12645_),
    .B(_12653_));
 sg13g2_xor2_1 _20334_ (.B(_12654_),
    .A(_12563_),
    .X(_12655_));
 sg13g2_xnor2_1 _20335_ (.Y(_12656_),
    .A(_12562_),
    .B(_12655_));
 sg13g2_o21ai_1 _20336_ (.B1(_12656_),
    .Y(_12657_),
    .A1(_12301_),
    .A2(_12560_));
 sg13g2_or2_1 _20337_ (.X(_12658_),
    .B(_12301_),
    .A(_12656_));
 sg13g2_nor2b_1 _20338_ (.A(_12300_),
    .B_N(_12256_),
    .Y(_12659_));
 sg13g2_inv_1 _20339_ (.Y(_12660_),
    .A(_12659_));
 sg13g2_o21ai_1 _20340_ (.B1(_12660_),
    .Y(_12661_),
    .A1(_12560_),
    .A2(_12658_));
 sg13g2_and2_1 _20341_ (.A(_12657_),
    .B(_12661_),
    .X(_12662_));
 sg13g2_buf_1 _20342_ (.A(_12662_),
    .X(_12663_));
 sg13g2_a21o_1 _20343_ (.A2(_12645_),
    .A1(_12652_),
    .B1(_12189_),
    .X(_12664_));
 sg13g2_o21ai_1 _20344_ (.B1(_12664_),
    .Y(_12665_),
    .A1(_12652_),
    .A2(_12645_));
 sg13g2_buf_1 _20345_ (.A(_12665_),
    .X(_12666_));
 sg13g2_nor2b_1 _20346_ (.A(_12648_),
    .B_N(_12651_),
    .Y(_12667_));
 sg13g2_nand2_1 _20347_ (.Y(_12668_),
    .A(_12066_),
    .B(net306));
 sg13g2_nand2_1 _20348_ (.Y(_12669_),
    .A(_12383_),
    .B(_11825_));
 sg13g2_nand2_1 _20349_ (.Y(_12670_),
    .A(net260),
    .B(net307));
 sg13g2_xnor2_1 _20350_ (.Y(_12671_),
    .A(_12669_),
    .B(_12670_));
 sg13g2_xnor2_1 _20351_ (.Y(_12672_),
    .A(_12668_),
    .B(_12671_));
 sg13g2_and2_1 _20352_ (.A(_12623_),
    .B(_12624_),
    .X(_12673_));
 sg13g2_or2_1 _20353_ (.X(_12674_),
    .B(_12624_),
    .A(_12623_));
 sg13g2_o21ai_1 _20354_ (.B1(_12674_),
    .Y(_12675_),
    .A1(_12625_),
    .A2(_12673_));
 sg13g2_buf_1 _20355_ (.A(_12675_),
    .X(_12676_));
 sg13g2_and2_1 _20356_ (.A(_12570_),
    .B(_12572_),
    .X(_12677_));
 sg13g2_or2_1 _20357_ (.X(_12678_),
    .B(_12572_),
    .A(_12570_));
 sg13g2_o21ai_1 _20358_ (.B1(_12678_),
    .Y(_12679_),
    .A1(_12571_),
    .A2(_12677_));
 sg13g2_buf_1 _20359_ (.A(_12679_),
    .X(_12680_));
 sg13g2_xnor2_1 _20360_ (.Y(_12681_),
    .A(_12676_),
    .B(_12680_));
 sg13g2_xnor2_1 _20361_ (.Y(_12682_),
    .A(_12672_),
    .B(_12681_));
 sg13g2_nand2_1 _20362_ (.Y(_12683_),
    .A(_12578_),
    .B(_12581_));
 sg13g2_nor2_1 _20363_ (.A(_12578_),
    .B(_12581_),
    .Y(_12684_));
 sg13g2_a21oi_1 _20364_ (.A1(_12574_),
    .A2(_12683_),
    .Y(_12685_),
    .B1(_12684_));
 sg13g2_nand2_1 _20365_ (.Y(_12686_),
    .A(net506),
    .B(_12611_));
 sg13g2_nand2_1 _20366_ (.Y(_12687_),
    .A(net283),
    .B(_11862_));
 sg13g2_nand2_1 _20367_ (.Y(_12688_),
    .A(_11839_),
    .B(_12110_));
 sg13g2_xnor2_1 _20368_ (.Y(_12689_),
    .A(_12687_),
    .B(_12688_));
 sg13g2_xnor2_1 _20369_ (.Y(_12690_),
    .A(_12686_),
    .B(_12689_));
 sg13g2_a21oi_1 _20370_ (.A1(_09786_),
    .A2(_11615_),
    .Y(_12691_),
    .B1(_09357_));
 sg13g2_o21ai_1 _20371_ (.B1(_09357_),
    .Y(_12692_),
    .A1(_09786_),
    .A2(_11615_));
 sg13g2_o21ai_1 _20372_ (.B1(_12692_),
    .Y(_12693_),
    .A1(_09343_),
    .A2(_12691_));
 sg13g2_o21ai_1 _20373_ (.B1(_09037_),
    .Y(_12694_),
    .A1(_09747_),
    .A2(_11390_));
 sg13g2_a21oi_1 _20374_ (.A1(_09747_),
    .A2(_11390_),
    .Y(_12695_),
    .B1(_09037_));
 sg13g2_a21oi_1 _20375_ (.A1(_09023_),
    .A2(_12694_),
    .Y(_12696_),
    .B1(_12695_));
 sg13g2_nand2b_1 _20376_ (.Y(_12697_),
    .B(net699),
    .A_N(_12696_));
 sg13g2_o21ai_1 _20377_ (.B1(_12697_),
    .Y(_12698_),
    .A1(_11712_),
    .A2(_12693_));
 sg13g2_a21o_1 _20378_ (.A2(_12698_),
    .A1(net728),
    .B1(net684),
    .X(_12699_));
 sg13g2_buf_1 _20379_ (.A(_12699_),
    .X(_12700_));
 sg13g2_buf_1 _20380_ (.A(\rbzero.wall_tracer.size_full[3] ),
    .X(_12701_));
 sg13g2_nor3_2 _20381_ (.A(_11760_),
    .B(_11727_),
    .C(_11854_),
    .Y(_12702_));
 sg13g2_xor2_1 _20382_ (.B(_12702_),
    .A(_12701_),
    .X(_12703_));
 sg13g2_nor2_1 _20383_ (.A(net728),
    .B(_12703_),
    .Y(_12704_));
 sg13g2_nand2b_1 _20384_ (.Y(_12705_),
    .B(net684),
    .A_N(_00457_));
 sg13g2_o21ai_1 _20385_ (.B1(_12705_),
    .Y(_12706_),
    .A1(_12700_),
    .A2(_12704_));
 sg13g2_nand2_1 _20386_ (.Y(_12707_),
    .A(net683),
    .B(_00456_));
 sg13g2_o21ai_1 _20387_ (.B1(_12707_),
    .Y(_12708_),
    .A1(net683),
    .A2(_12706_));
 sg13g2_buf_1 _20388_ (.A(_12708_),
    .X(_12709_));
 sg13g2_nor2_1 _20389_ (.A(net521),
    .B(net278),
    .Y(_12710_));
 sg13g2_nor2_1 _20390_ (.A(_12589_),
    .B(_12591_),
    .Y(_12711_));
 sg13g2_a22oi_1 _20391_ (.Y(_12712_),
    .B1(_12589_),
    .B2(_12591_),
    .A2(_11810_),
    .A1(net283));
 sg13g2_or2_1 _20392_ (.X(_12713_),
    .B(_12712_),
    .A(_12711_));
 sg13g2_buf_1 _20393_ (.A(_12713_),
    .X(_12714_));
 sg13g2_xor2_1 _20394_ (.B(_12714_),
    .A(_12710_),
    .X(_12715_));
 sg13g2_xnor2_1 _20395_ (.Y(_12716_),
    .A(_12690_),
    .B(_12715_));
 sg13g2_xnor2_1 _20396_ (.Y(_12717_),
    .A(_12685_),
    .B(_12716_));
 sg13g2_xnor2_1 _20397_ (.Y(_12718_),
    .A(_12682_),
    .B(_12717_));
 sg13g2_nor2_1 _20398_ (.A(_12622_),
    .B(_12639_),
    .Y(_12719_));
 sg13g2_nor2_1 _20399_ (.A(_12583_),
    .B(_12614_),
    .Y(_12720_));
 sg13g2_nand2_1 _20400_ (.Y(_12721_),
    .A(_12583_),
    .B(_12614_));
 sg13g2_o21ai_1 _20401_ (.B1(_12721_),
    .Y(_12722_),
    .A1(_12586_),
    .A2(_12720_));
 sg13g2_buf_1 _20402_ (.A(_12722_),
    .X(_12723_));
 sg13g2_xor2_1 _20403_ (.B(_12723_),
    .A(_12719_),
    .X(_12724_));
 sg13g2_xnor2_1 _20404_ (.Y(_12725_),
    .A(_12718_),
    .B(_12724_));
 sg13g2_nor2_1 _20405_ (.A(_12640_),
    .B(_12643_),
    .Y(_12726_));
 sg13g2_buf_1 _20406_ (.A(net630),
    .X(_12727_));
 sg13g2_nand2_1 _20407_ (.Y(_12728_),
    .A(_08536_),
    .B(net567));
 sg13g2_buf_2 _20408_ (.A(_12728_),
    .X(_12729_));
 sg13g2_nor2_1 _20409_ (.A(net467),
    .B(_12729_),
    .Y(_12730_));
 sg13g2_nand2_1 _20410_ (.Y(_12731_),
    .A(_08537_),
    .B(net567));
 sg13g2_buf_1 _20411_ (.A(_12731_),
    .X(_12732_));
 sg13g2_nor2_1 _20412_ (.A(net455),
    .B(net503),
    .Y(_12733_));
 sg13g2_xnor2_1 _20413_ (.Y(_12734_),
    .A(_12730_),
    .B(_12733_));
 sg13g2_nand2_1 _20414_ (.Y(_12735_),
    .A(_12634_),
    .B(_12627_));
 sg13g2_o21ai_1 _20415_ (.B1(_12637_),
    .Y(_12736_),
    .A1(_12634_),
    .A2(_12627_));
 sg13g2_nand2_1 _20416_ (.Y(_12737_),
    .A(_12735_),
    .B(_12736_));
 sg13g2_nand2_1 _20417_ (.Y(_12738_),
    .A(net282),
    .B(net333));
 sg13g2_buf_1 _20418_ (.A(_11887_),
    .X(_12739_));
 sg13g2_nand2_1 _20419_ (.Y(_12740_),
    .A(net266),
    .B(net332));
 sg13g2_nand2_1 _20420_ (.Y(_12741_),
    .A(_12012_),
    .B(_11940_));
 sg13g2_xnor2_1 _20421_ (.Y(_12742_),
    .A(_12740_),
    .B(_12741_));
 sg13g2_xnor2_1 _20422_ (.Y(_12743_),
    .A(_12738_),
    .B(_12742_));
 sg13g2_nand3_1 _20423_ (.B(_12171_),
    .C(_12631_),
    .A(net405),
    .Y(_12744_));
 sg13g2_a21oi_1 _20424_ (.A1(net405),
    .A2(net280),
    .Y(_12745_),
    .B1(_12631_));
 sg13g2_a21o_1 _20425_ (.A2(_12744_),
    .A1(_12632_),
    .B1(_12745_),
    .X(_12746_));
 sg13g2_buf_1 _20426_ (.A(_12746_),
    .X(_12747_));
 sg13g2_nand2_1 _20427_ (.Y(_12748_),
    .A(net406),
    .B(net280));
 sg13g2_nand2_1 _20428_ (.Y(_12749_),
    .A(net446),
    .B(net523));
 sg13g2_nand2_1 _20429_ (.Y(_12750_),
    .A(_12124_),
    .B(net264));
 sg13g2_xor2_1 _20430_ (.B(_12750_),
    .A(_12749_),
    .X(_12751_));
 sg13g2_xnor2_1 _20431_ (.Y(_12752_),
    .A(_12748_),
    .B(_12751_));
 sg13g2_xor2_1 _20432_ (.B(_12752_),
    .A(_12747_),
    .X(_12753_));
 sg13g2_xnor2_1 _20433_ (.Y(_12754_),
    .A(_12743_),
    .B(_12753_));
 sg13g2_xnor2_1 _20434_ (.Y(_12755_),
    .A(_12737_),
    .B(_12754_));
 sg13g2_xnor2_1 _20435_ (.Y(_12756_),
    .A(_12734_),
    .B(_12755_));
 sg13g2_xor2_1 _20436_ (.B(_12756_),
    .A(_12726_),
    .X(_12757_));
 sg13g2_xnor2_1 _20437_ (.Y(_12758_),
    .A(_12725_),
    .B(_12757_));
 sg13g2_nand2_1 _20438_ (.Y(_12759_),
    .A(_12568_),
    .B(_12616_));
 sg13g2_nor2_1 _20439_ (.A(_12568_),
    .B(_12616_),
    .Y(_12760_));
 sg13g2_a21oi_1 _20440_ (.A1(_12569_),
    .A2(_12759_),
    .Y(_12761_),
    .B1(_12760_));
 sg13g2_buf_1 _20441_ (.A(_12611_),
    .X(_12762_));
 sg13g2_a22oi_1 _20442_ (.Y(_12763_),
    .B1(net277),
    .B2(net505),
    .A2(_12593_),
    .A1(_12596_));
 sg13g2_inv_1 _20443_ (.Y(_12764_),
    .A(_12763_));
 sg13g2_o21ai_1 _20444_ (.B1(_12764_),
    .Y(_12765_),
    .A1(_12596_),
    .A2(_12593_));
 sg13g2_xor2_1 _20445_ (.B(_12765_),
    .A(_12761_),
    .X(_12766_));
 sg13g2_nand2_1 _20446_ (.Y(_12767_),
    .A(_12618_),
    .B(_12644_));
 sg13g2_xor2_1 _20447_ (.B(_12767_),
    .A(_12766_),
    .X(_12768_));
 sg13g2_xnor2_1 _20448_ (.Y(_12769_),
    .A(_12758_),
    .B(_12768_));
 sg13g2_xor2_1 _20449_ (.B(_12769_),
    .A(_12667_),
    .X(_12770_));
 sg13g2_xnor2_1 _20450_ (.Y(_12771_),
    .A(_12666_),
    .B(_12770_));
 sg13g2_o21ai_1 _20451_ (.B1(_12654_),
    .Y(_12772_),
    .A1(_12563_),
    .A2(_12562_));
 sg13g2_nor2b_1 _20452_ (.A(_12771_),
    .B_N(_12772_),
    .Y(_12773_));
 sg13g2_nand2b_1 _20453_ (.Y(_12774_),
    .B(_12771_),
    .A_N(_12772_));
 sg13g2_inv_1 _20454_ (.Y(_12775_),
    .A(_12774_));
 sg13g2_nor2_1 _20455_ (.A(_12773_),
    .B(_12775_),
    .Y(_12776_));
 sg13g2_xor2_1 _20456_ (.B(_12776_),
    .A(_12663_),
    .X(_12777_));
 sg13g2_nand2_1 _20457_ (.Y(_12778_),
    .A(net450),
    .B(_12777_));
 sg13g2_nand2_1 _20458_ (.Y(_12779_),
    .A(\rbzero.traced_texVinit[0] ),
    .B(net448));
 sg13g2_a21oi_1 _20459_ (.A1(_12778_),
    .A2(_12779_),
    .Y(_01510_),
    .B1(net572));
 sg13g2_buf_1 _20460_ (.A(_08675_),
    .X(_12780_));
 sg13g2_nor2_1 _20461_ (.A(\rbzero.traced_texVinit[1] ),
    .B(_11714_),
    .Y(_12781_));
 sg13g2_a21oi_1 _20462_ (.A1(_12663_),
    .A2(_12776_),
    .Y(_12782_),
    .B1(_12775_));
 sg13g2_nand2b_1 _20463_ (.Y(_12783_),
    .B(_12666_),
    .A_N(_12769_));
 sg13g2_nor2b_1 _20464_ (.A(_12666_),
    .B_N(_12769_),
    .Y(_12784_));
 sg13g2_a21oi_2 _20465_ (.B1(_12784_),
    .Y(_12785_),
    .A2(_12783_),
    .A1(_12667_));
 sg13g2_nand2_1 _20466_ (.Y(_12786_),
    .A(_12725_),
    .B(_12756_));
 sg13g2_nor2_1 _20467_ (.A(_12725_),
    .B(_12756_),
    .Y(_12787_));
 sg13g2_a21oi_1 _20468_ (.A1(_12726_),
    .A2(_12786_),
    .Y(_12788_),
    .B1(_12787_));
 sg13g2_nand2_1 _20469_ (.Y(_12789_),
    .A(_12686_),
    .B(_12688_));
 sg13g2_o21ai_1 _20470_ (.B1(_12687_),
    .Y(_12790_),
    .A1(_12686_),
    .A2(_12688_));
 sg13g2_nand2_1 _20471_ (.Y(_12791_),
    .A(_12789_),
    .B(_12790_));
 sg13g2_nand2_1 _20472_ (.Y(_12792_),
    .A(net520),
    .B(_12611_));
 sg13g2_nand2_1 _20473_ (.Y(_12793_),
    .A(net268),
    .B(_12110_));
 sg13g2_nor2_1 _20474_ (.A(_12202_),
    .B(net278),
    .Y(_12794_));
 sg13g2_xnor2_1 _20475_ (.Y(_12795_),
    .A(_12793_),
    .B(_12794_));
 sg13g2_xnor2_1 _20476_ (.Y(_12796_),
    .A(_12792_),
    .B(_12795_));
 sg13g2_buf_1 _20477_ (.A(\rbzero.wall_tracer.size_full[4] ),
    .X(_12797_));
 sg13g2_nand2b_1 _20478_ (.Y(_12798_),
    .B(_12702_),
    .A_N(_12701_));
 sg13g2_xnor2_1 _20479_ (.Y(_12799_),
    .A(_12797_),
    .B(_12798_));
 sg13g2_inv_2 _20480_ (.Y(_12800_),
    .A(_12700_));
 sg13g2_o21ai_1 _20481_ (.B1(_12800_),
    .Y(_12801_),
    .A1(_08420_),
    .A2(_12799_));
 sg13g2_nand2b_1 _20482_ (.Y(_12802_),
    .B(net684),
    .A_N(_00459_));
 sg13g2_a21o_1 _20483_ (.A2(_12802_),
    .A1(_12801_),
    .B1(net683),
    .X(_12803_));
 sg13g2_o21ai_1 _20484_ (.B1(_12803_),
    .Y(_12804_),
    .A1(net522),
    .A2(_00458_));
 sg13g2_buf_1 _20485_ (.A(_12804_),
    .X(_12805_));
 sg13g2_and2_1 _20486_ (.A(net505),
    .B(_12805_),
    .X(_12806_));
 sg13g2_xnor2_1 _20487_ (.Y(_12807_),
    .A(_12796_),
    .B(_12806_));
 sg13g2_xnor2_1 _20488_ (.Y(_12808_),
    .A(_12791_),
    .B(_12807_));
 sg13g2_nor2_1 _20489_ (.A(_12676_),
    .B(_12680_),
    .Y(_12809_));
 sg13g2_nor2_1 _20490_ (.A(_12672_),
    .B(_12809_),
    .Y(_12810_));
 sg13g2_a21oi_2 _20491_ (.B1(_12810_),
    .Y(_12811_),
    .A2(_12680_),
    .A1(_12676_));
 sg13g2_nand2_1 _20492_ (.Y(_12812_),
    .A(_12066_),
    .B(_11862_));
 sg13g2_buf_1 _20493_ (.A(_11825_),
    .X(_12813_));
 sg13g2_nand2_1 _20494_ (.Y(_12814_),
    .A(net260),
    .B(net293));
 sg13g2_nand2_1 _20495_ (.Y(_12815_),
    .A(_12383_),
    .B(net306));
 sg13g2_xnor2_1 _20496_ (.Y(_12816_),
    .A(_12814_),
    .B(_12815_));
 sg13g2_xnor2_1 _20497_ (.Y(_12817_),
    .A(_12812_),
    .B(_12816_));
 sg13g2_and2_1 _20498_ (.A(_12740_),
    .B(_12741_),
    .X(_12818_));
 sg13g2_or2_1 _20499_ (.X(_12819_),
    .B(_12741_),
    .A(_12740_));
 sg13g2_o21ai_1 _20500_ (.B1(_12819_),
    .Y(_12820_),
    .A1(_12738_),
    .A2(_12818_));
 sg13g2_buf_1 _20501_ (.A(_12820_),
    .X(_12821_));
 sg13g2_or2_1 _20502_ (.X(_12822_),
    .B(_12670_),
    .A(_12668_));
 sg13g2_and2_1 _20503_ (.A(_12668_),
    .B(_12670_),
    .X(_12823_));
 sg13g2_a21oi_2 _20504_ (.B1(_12823_),
    .Y(_12824_),
    .A2(_12822_),
    .A1(_12669_));
 sg13g2_xnor2_1 _20505_ (.Y(_12825_),
    .A(_12821_),
    .B(_12824_));
 sg13g2_xnor2_1 _20506_ (.Y(_12826_),
    .A(_12817_),
    .B(_12825_));
 sg13g2_xor2_1 _20507_ (.B(_12826_),
    .A(_12811_),
    .X(_12827_));
 sg13g2_xnor2_1 _20508_ (.Y(_12828_),
    .A(_12808_),
    .B(_12827_));
 sg13g2_nand2_1 _20509_ (.Y(_12829_),
    .A(_12682_),
    .B(_12716_));
 sg13g2_nor2_1 _20510_ (.A(_12682_),
    .B(_12716_),
    .Y(_12830_));
 sg13g2_a21o_1 _20511_ (.A2(_12829_),
    .A1(_12685_),
    .B1(_12830_),
    .X(_12831_));
 sg13g2_buf_1 _20512_ (.A(_12831_),
    .X(_12832_));
 sg13g2_or2_1 _20513_ (.X(_12833_),
    .B(_12754_),
    .A(_12737_));
 sg13g2_xor2_1 _20514_ (.B(_12833_),
    .A(_12832_),
    .X(_12834_));
 sg13g2_xnor2_1 _20515_ (.Y(_12835_),
    .A(_12828_),
    .B(_12834_));
 sg13g2_and2_1 _20516_ (.A(_08536_),
    .B(_11798_),
    .X(_12836_));
 sg13g2_buf_1 _20517_ (.A(_12836_),
    .X(_12837_));
 sg13g2_nand2_1 _20518_ (.Y(_12838_),
    .A(_12120_),
    .B(net519));
 sg13g2_buf_2 _20519_ (.A(_12838_),
    .X(_12839_));
 sg13g2_and2_1 _20520_ (.A(_08535_),
    .B(_11798_),
    .X(_12840_));
 sg13g2_buf_1 _20521_ (.A(_12840_),
    .X(_12841_));
 sg13g2_nand2_1 _20522_ (.Y(_12842_),
    .A(net454),
    .B(net518));
 sg13g2_xor2_1 _20523_ (.B(_12842_),
    .A(_12839_),
    .X(_12843_));
 sg13g2_nand3_1 _20524_ (.B(_12642_),
    .C(net518),
    .A(_12239_),
    .Y(_12844_));
 sg13g2_o21ai_1 _20525_ (.B1(_12844_),
    .Y(_12845_),
    .A1(net443),
    .A2(_12839_));
 sg13g2_o21ai_1 _20526_ (.B1(_12842_),
    .Y(_12846_),
    .A1(net454),
    .A2(_12839_));
 sg13g2_nor3_1 _20527_ (.A(net444),
    .B(net503),
    .C(_12846_),
    .Y(_12847_));
 sg13g2_a221oi_1 _20528_ (.B2(net444),
    .C1(_12847_),
    .B1(_12845_),
    .A1(net503),
    .Y(_12848_),
    .A2(_12843_));
 sg13g2_nand2_1 _20529_ (.Y(_12849_),
    .A(_12747_),
    .B(_12743_));
 sg13g2_nor2_1 _20530_ (.A(_12747_),
    .B(_12743_),
    .Y(_12850_));
 sg13g2_a21oi_1 _20531_ (.A1(_12752_),
    .A2(_12849_),
    .Y(_12851_),
    .B1(_12850_));
 sg13g2_nand2_1 _20532_ (.Y(_12852_),
    .A(net261),
    .B(net307));
 sg13g2_nand2_1 _20533_ (.Y(_12853_),
    .A(_11999_),
    .B(_11837_));
 sg13g2_nand2_1 _20534_ (.Y(_12854_),
    .A(net263),
    .B(net332));
 sg13g2_xnor2_1 _20535_ (.Y(_12855_),
    .A(_12853_),
    .B(_12854_));
 sg13g2_xnor2_1 _20536_ (.Y(_12856_),
    .A(_12852_),
    .B(_12855_));
 sg13g2_nand2_1 _20537_ (.Y(_12857_),
    .A(_12172_),
    .B(_11940_));
 sg13g2_a21oi_2 _20538_ (.B1(_12630_),
    .Y(_12858_),
    .A2(_11956_),
    .A1(_11949_));
 sg13g2_nand2_1 _20539_ (.Y(_12859_),
    .A(net406),
    .B(_12134_));
 sg13g2_xor2_1 _20540_ (.B(_12859_),
    .A(_12858_),
    .X(_12860_));
 sg13g2_xnor2_1 _20541_ (.Y(_12861_),
    .A(_12857_),
    .B(_12860_));
 sg13g2_or2_1 _20542_ (.X(_12862_),
    .B(_12750_),
    .A(_12749_));
 sg13g2_and2_1 _20543_ (.A(_12749_),
    .B(_12750_),
    .X(_12863_));
 sg13g2_a21oi_1 _20544_ (.A1(_12748_),
    .A2(_12862_),
    .Y(_12864_),
    .B1(_12863_));
 sg13g2_xor2_1 _20545_ (.B(_12864_),
    .A(_12861_),
    .X(_12865_));
 sg13g2_xnor2_1 _20546_ (.Y(_12866_),
    .A(_12856_),
    .B(_12865_));
 sg13g2_xnor2_1 _20547_ (.Y(_12867_),
    .A(_12851_),
    .B(_12866_));
 sg13g2_xnor2_1 _20548_ (.Y(_12868_),
    .A(_12848_),
    .B(_12867_));
 sg13g2_nor2_1 _20549_ (.A(_12734_),
    .B(_12755_),
    .Y(_12869_));
 sg13g2_nor2b_1 _20550_ (.A(_12868_),
    .B_N(_12869_),
    .Y(_12870_));
 sg13g2_nand2b_1 _20551_ (.Y(_12871_),
    .B(_12868_),
    .A_N(_12869_));
 sg13g2_nand2b_1 _20552_ (.Y(_12872_),
    .B(_12871_),
    .A_N(_12870_));
 sg13g2_xnor2_1 _20553_ (.Y(_12873_),
    .A(_12835_),
    .B(_12872_));
 sg13g2_nand2_1 _20554_ (.Y(_12874_),
    .A(_12723_),
    .B(_12718_));
 sg13g2_o21ai_1 _20555_ (.B1(_12719_),
    .Y(_12875_),
    .A1(_12723_),
    .A2(_12718_));
 sg13g2_nand2_1 _20556_ (.Y(_12876_),
    .A(_12874_),
    .B(_12875_));
 sg13g2_nand2_1 _20557_ (.Y(_12877_),
    .A(_12690_),
    .B(_12714_));
 sg13g2_nor2_1 _20558_ (.A(_12690_),
    .B(_12714_),
    .Y(_12878_));
 sg13g2_a21oi_1 _20559_ (.A1(_12710_),
    .A2(_12877_),
    .Y(_12879_),
    .B1(_12878_));
 sg13g2_xnor2_1 _20560_ (.Y(_12880_),
    .A(_12876_),
    .B(_12879_));
 sg13g2_xor2_1 _20561_ (.B(_12880_),
    .A(_12873_),
    .X(_12881_));
 sg13g2_xnor2_1 _20562_ (.Y(_12882_),
    .A(_12788_),
    .B(_12881_));
 sg13g2_nor2b_1 _20563_ (.A(_12765_),
    .B_N(_12761_),
    .Y(_12883_));
 sg13g2_or2_1 _20564_ (.X(_12884_),
    .B(_12767_),
    .A(_12766_));
 sg13g2_and2_1 _20565_ (.A(_12766_),
    .B(_12767_),
    .X(_12885_));
 sg13g2_a21o_1 _20566_ (.A2(_12884_),
    .A1(_12758_),
    .B1(_12885_),
    .X(_12886_));
 sg13g2_xnor2_1 _20567_ (.Y(_12887_),
    .A(_12883_),
    .B(_12886_));
 sg13g2_xnor2_1 _20568_ (.Y(_12888_),
    .A(_12882_),
    .B(_12887_));
 sg13g2_xor2_1 _20569_ (.B(_12888_),
    .A(_12785_),
    .X(_12889_));
 sg13g2_xnor2_1 _20570_ (.Y(_12890_),
    .A(_12782_),
    .B(_12889_));
 sg13g2_nor2_1 _20571_ (.A(net464),
    .B(_12890_),
    .Y(_12891_));
 sg13g2_nor3_1 _20572_ (.A(net629),
    .B(_12781_),
    .C(_12891_),
    .Y(_01511_));
 sg13g2_nand2_1 _20573_ (.Y(_12892_),
    .A(_12785_),
    .B(_12888_));
 sg13g2_nor2b_1 _20574_ (.A(_12773_),
    .B_N(_12892_),
    .Y(_12893_));
 sg13g2_nor2_1 _20575_ (.A(_12785_),
    .B(_12888_),
    .Y(_12894_));
 sg13g2_a221oi_1 _20576_ (.B2(_12663_),
    .C1(_12894_),
    .B1(_12893_),
    .A1(_12775_),
    .Y(_12895_),
    .A2(_12892_));
 sg13g2_buf_1 _20577_ (.A(_12895_),
    .X(_12896_));
 sg13g2_nand2_1 _20578_ (.Y(_12897_),
    .A(_12883_),
    .B(_12882_));
 sg13g2_nor2_1 _20579_ (.A(_12883_),
    .B(_12882_),
    .Y(_12898_));
 sg13g2_a21oi_2 _20580_ (.B1(_12898_),
    .Y(_12899_),
    .A2(_12897_),
    .A1(_12886_));
 sg13g2_inv_1 _20581_ (.Y(_12900_),
    .A(_12899_));
 sg13g2_nand2_1 _20582_ (.Y(_12901_),
    .A(_12793_),
    .B(_12792_));
 sg13g2_nand2_1 _20583_ (.Y(_12902_),
    .A(_12794_),
    .B(_12901_));
 sg13g2_o21ai_1 _20584_ (.B1(_12902_),
    .Y(_12903_),
    .A1(_12793_),
    .A2(_12792_));
 sg13g2_buf_1 _20585_ (.A(_12903_),
    .X(_12904_));
 sg13g2_buf_1 _20586_ (.A(_12805_),
    .X(_12905_));
 sg13g2_nand2_1 _20587_ (.Y(_12906_),
    .A(net506),
    .B(net211));
 sg13g2_nand2_1 _20588_ (.Y(_12907_),
    .A(net268),
    .B(net277));
 sg13g2_nor2_1 _20589_ (.A(net568),
    .B(net278),
    .Y(_12908_));
 sg13g2_xnor2_1 _20590_ (.Y(_12909_),
    .A(_12907_),
    .B(_12908_));
 sg13g2_xnor2_1 _20591_ (.Y(_12910_),
    .A(_12906_),
    .B(_12909_));
 sg13g2_buf_1 _20592_ (.A(\rbzero.wall_tracer.size_full[5] ),
    .X(_12911_));
 sg13g2_or2_1 _20593_ (.X(_12912_),
    .B(_12798_),
    .A(_12797_));
 sg13g2_xnor2_1 _20594_ (.Y(_12913_),
    .A(_12911_),
    .B(_12912_));
 sg13g2_o21ai_1 _20595_ (.B1(_12800_),
    .Y(_12914_),
    .A1(net685),
    .A2(_12913_));
 sg13g2_nand2b_1 _20596_ (.Y(_12915_),
    .B(_08442_),
    .A_N(_00461_));
 sg13g2_a21o_1 _20597_ (.A2(_12915_),
    .A1(_12914_),
    .B1(net683),
    .X(_12916_));
 sg13g2_o21ai_1 _20598_ (.B1(_12916_),
    .Y(_12917_),
    .A1(net522),
    .A2(_00460_));
 sg13g2_buf_1 _20599_ (.A(_12917_),
    .X(_12918_));
 sg13g2_nand2_1 _20600_ (.Y(_12919_),
    .A(net505),
    .B(_12918_));
 sg13g2_xor2_1 _20601_ (.B(_12919_),
    .A(_12910_),
    .X(_12920_));
 sg13g2_xnor2_1 _20602_ (.Y(_12921_),
    .A(_12904_),
    .B(_12920_));
 sg13g2_nor2_1 _20603_ (.A(_12821_),
    .B(_12824_),
    .Y(_12922_));
 sg13g2_nor2_1 _20604_ (.A(_12817_),
    .B(_12922_),
    .Y(_12923_));
 sg13g2_a21oi_2 _20605_ (.B1(_12923_),
    .Y(_12924_),
    .A2(_12824_),
    .A1(_12821_));
 sg13g2_buf_1 _20606_ (.A(_12110_),
    .X(_12925_));
 sg13g2_nand2_1 _20607_ (.Y(_12926_),
    .A(net238),
    .B(net276));
 sg13g2_nand2_1 _20608_ (.Y(_12927_),
    .A(net260),
    .B(net306));
 sg13g2_buf_1 _20609_ (.A(_11862_),
    .X(_12928_));
 sg13g2_nand2_1 _20610_ (.Y(_12929_),
    .A(net239),
    .B(net292));
 sg13g2_xor2_1 _20611_ (.B(_12929_),
    .A(_12927_),
    .X(_12930_));
 sg13g2_xor2_1 _20612_ (.B(_12930_),
    .A(_12926_),
    .X(_12931_));
 sg13g2_nor2_1 _20613_ (.A(_12853_),
    .B(_12854_),
    .Y(_12932_));
 sg13g2_a21oi_1 _20614_ (.A1(_12853_),
    .A2(_12854_),
    .Y(_12933_),
    .B1(_12852_));
 sg13g2_or2_1 _20615_ (.X(_12934_),
    .B(_12933_),
    .A(_12932_));
 sg13g2_buf_1 _20616_ (.A(_12934_),
    .X(_12935_));
 sg13g2_a21o_1 _20617_ (.A2(_12814_),
    .A1(_12812_),
    .B1(_12815_),
    .X(_12936_));
 sg13g2_o21ai_1 _20618_ (.B1(_12936_),
    .Y(_12937_),
    .A1(_12812_),
    .A2(_12814_));
 sg13g2_buf_1 _20619_ (.A(_12937_),
    .X(_12938_));
 sg13g2_xnor2_1 _20620_ (.Y(_12939_),
    .A(_12935_),
    .B(_12938_));
 sg13g2_xnor2_1 _20621_ (.Y(_12940_),
    .A(_12931_),
    .B(_12939_));
 sg13g2_xor2_1 _20622_ (.B(_12940_),
    .A(_12924_),
    .X(_12941_));
 sg13g2_xnor2_1 _20623_ (.Y(_12942_),
    .A(_12921_),
    .B(_12941_));
 sg13g2_nand2_1 _20624_ (.Y(_12943_),
    .A(_12811_),
    .B(_12826_));
 sg13g2_o21ai_1 _20625_ (.B1(_12808_),
    .Y(_12944_),
    .A1(_12811_),
    .A2(_12826_));
 sg13g2_nand2_1 _20626_ (.Y(_12945_),
    .A(_12943_),
    .B(_12944_));
 sg13g2_or2_1 _20627_ (.X(_12946_),
    .B(_12866_),
    .A(_12851_));
 sg13g2_buf_1 _20628_ (.A(_12946_),
    .X(_12947_));
 sg13g2_xnor2_1 _20629_ (.Y(_12948_),
    .A(_12945_),
    .B(_12947_));
 sg13g2_xnor2_1 _20630_ (.Y(_12949_),
    .A(_12942_),
    .B(_12948_));
 sg13g2_nor2_1 _20631_ (.A(_12848_),
    .B(_12867_),
    .Y(_12950_));
 sg13g2_nand2_1 _20632_ (.Y(_12951_),
    .A(_12861_),
    .B(_12856_));
 sg13g2_nor2_1 _20633_ (.A(_12861_),
    .B(_12856_),
    .Y(_12952_));
 sg13g2_a21oi_1 _20634_ (.A1(_12864_),
    .A2(_12951_),
    .Y(_12953_),
    .B1(_12952_));
 sg13g2_nand2_1 _20635_ (.Y(_12954_),
    .A(net261),
    .B(net293));
 sg13g2_nand2_1 _20636_ (.Y(_12955_),
    .A(net263),
    .B(net333));
 sg13g2_nand2_1 _20637_ (.Y(_12956_),
    .A(net240),
    .B(net307));
 sg13g2_xnor2_1 _20638_ (.Y(_12957_),
    .A(_12955_),
    .B(_12956_));
 sg13g2_xnor2_1 _20639_ (.Y(_12958_),
    .A(_12954_),
    .B(_12957_));
 sg13g2_buf_1 _20640_ (.A(_12172_),
    .X(_12959_));
 sg13g2_nand3_1 _20641_ (.B(net363),
    .C(_12858_),
    .A(net259),
    .Y(_12960_));
 sg13g2_a21oi_1 _20642_ (.A1(net259),
    .A2(net363),
    .Y(_12961_),
    .B1(_12858_));
 sg13g2_a21oi_1 _20643_ (.A1(_12859_),
    .A2(_12960_),
    .Y(_12962_),
    .B1(_12961_));
 sg13g2_nand2_1 _20644_ (.Y(_12963_),
    .A(net259),
    .B(net332));
 sg13g2_nand2_1 _20645_ (.Y(_12964_),
    .A(net406),
    .B(net523));
 sg13g2_nand2_1 _20646_ (.Y(_12965_),
    .A(net264),
    .B(net363));
 sg13g2_xnor2_1 _20647_ (.Y(_12966_),
    .A(_12964_),
    .B(_12965_));
 sg13g2_xnor2_1 _20648_ (.Y(_12967_),
    .A(_12963_),
    .B(_12966_));
 sg13g2_xor2_1 _20649_ (.B(_12967_),
    .A(_12962_),
    .X(_12968_));
 sg13g2_xnor2_1 _20650_ (.Y(_12969_),
    .A(_12958_),
    .B(_12968_));
 sg13g2_xnor2_1 _20651_ (.Y(_12970_),
    .A(net444),
    .B(net518));
 sg13g2_nor3_2 _20652_ (.A(_12643_),
    .B(_12839_),
    .C(_12970_),
    .Y(_12971_));
 sg13g2_xor2_1 _20653_ (.B(_12971_),
    .A(_12969_),
    .X(_12972_));
 sg13g2_xnor2_1 _20654_ (.Y(_12973_),
    .A(_12953_),
    .B(_12972_));
 sg13g2_buf_1 _20655_ (.A(net446),
    .X(_12974_));
 sg13g2_nor2_1 _20656_ (.A(_12839_),
    .B(_12842_),
    .Y(_12975_));
 sg13g2_a21oi_1 _20657_ (.A1(net404),
    .A2(_12642_),
    .Y(_12976_),
    .B1(_12975_));
 sg13g2_a21o_1 _20658_ (.A2(_12842_),
    .A1(_12839_),
    .B1(_12976_),
    .X(_12977_));
 sg13g2_a21oi_2 _20659_ (.B1(net503),
    .Y(_12978_),
    .A2(_11956_),
    .A1(_11949_));
 sg13g2_nand2_2 _20660_ (.Y(_12979_),
    .A(_08535_),
    .B(net567));
 sg13g2_nor2_1 _20661_ (.A(net455),
    .B(_12979_),
    .Y(_12980_));
 sg13g2_nor2_1 _20662_ (.A(_12398_),
    .B(_12729_),
    .Y(_12981_));
 sg13g2_xnor2_1 _20663_ (.Y(_12982_),
    .A(_12980_),
    .B(_12981_));
 sg13g2_xnor2_1 _20664_ (.Y(_12983_),
    .A(_12978_),
    .B(_12982_));
 sg13g2_xor2_1 _20665_ (.B(_12983_),
    .A(_12977_),
    .X(_12984_));
 sg13g2_and2_1 _20666_ (.A(_08547_),
    .B(_12727_),
    .X(_12985_));
 sg13g2_buf_1 _20667_ (.A(_12985_),
    .X(_12986_));
 sg13g2_buf_1 _20668_ (.A(_12986_),
    .X(_12987_));
 sg13g2_nand2_1 _20669_ (.Y(_12988_),
    .A(net443),
    .B(net482));
 sg13g2_xor2_1 _20670_ (.B(_12988_),
    .A(_12984_),
    .X(_12989_));
 sg13g2_xor2_1 _20671_ (.B(_12989_),
    .A(_12973_),
    .X(_12990_));
 sg13g2_xor2_1 _20672_ (.B(_12990_),
    .A(_12950_),
    .X(_12991_));
 sg13g2_xnor2_1 _20673_ (.Y(_12992_),
    .A(_12949_),
    .B(_12991_));
 sg13g2_nand2_1 _20674_ (.Y(_12993_),
    .A(_12832_),
    .B(_12828_));
 sg13g2_nor2_1 _20675_ (.A(_12832_),
    .B(_12828_),
    .Y(_12994_));
 sg13g2_a21oi_1 _20676_ (.A1(_12833_),
    .A2(_12993_),
    .Y(_12995_),
    .B1(_12994_));
 sg13g2_nand2b_1 _20677_ (.Y(_12996_),
    .B(_12791_),
    .A_N(_12796_));
 sg13g2_nor2b_1 _20678_ (.A(_12791_),
    .B_N(_12796_),
    .Y(_12997_));
 sg13g2_a21oi_1 _20679_ (.A1(_12806_),
    .A2(_12996_),
    .Y(_12998_),
    .B1(_12997_));
 sg13g2_xnor2_1 _20680_ (.Y(_12999_),
    .A(_12995_),
    .B(_12998_));
 sg13g2_a21o_1 _20681_ (.A2(_12871_),
    .A1(_12835_),
    .B1(_12870_),
    .X(_13000_));
 sg13g2_buf_1 _20682_ (.A(_13000_),
    .X(_13001_));
 sg13g2_xnor2_1 _20683_ (.Y(_13002_),
    .A(_12999_),
    .B(_13001_));
 sg13g2_xnor2_1 _20684_ (.Y(_13003_),
    .A(_12992_),
    .B(_13002_));
 sg13g2_nand2b_1 _20685_ (.Y(_13004_),
    .B(_12876_),
    .A_N(_12879_));
 sg13g2_buf_1 _20686_ (.A(_13004_),
    .X(_13005_));
 sg13g2_nor2_1 _20687_ (.A(_12873_),
    .B(_12880_),
    .Y(_13006_));
 sg13g2_nor2_1 _20688_ (.A(_12788_),
    .B(_13006_),
    .Y(_13007_));
 sg13g2_a21oi_2 _20689_ (.B1(_13007_),
    .Y(_13008_),
    .A2(_12880_),
    .A1(_12873_));
 sg13g2_xnor2_1 _20690_ (.Y(_13009_),
    .A(_13005_),
    .B(_13008_));
 sg13g2_xnor2_1 _20691_ (.Y(_13010_),
    .A(_13003_),
    .B(_13009_));
 sg13g2_xnor2_1 _20692_ (.Y(_13011_),
    .A(_12900_),
    .B(_13010_));
 sg13g2_xnor2_1 _20693_ (.Y(_13012_),
    .A(_12896_),
    .B(_13011_));
 sg13g2_buf_2 _20694_ (.A(_13012_),
    .X(_13013_));
 sg13g2_nor2_1 _20695_ (.A(net464),
    .B(_13013_),
    .Y(_13014_));
 sg13g2_a21oi_1 _20696_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(net452),
    .Y(_13015_),
    .B1(_13014_));
 sg13g2_nor2_1 _20697_ (.A(net634),
    .B(_13015_),
    .Y(_01512_));
 sg13g2_nor2_1 _20698_ (.A(_12999_),
    .B(_13001_),
    .Y(_13016_));
 sg13g2_nor2_1 _20699_ (.A(_12992_),
    .B(_13016_),
    .Y(_13017_));
 sg13g2_a21oi_1 _20700_ (.A1(_12999_),
    .A2(_13001_),
    .Y(_13018_),
    .B1(_13017_));
 sg13g2_nor2b_1 _20701_ (.A(_12998_),
    .B_N(_12995_),
    .Y(_13019_));
 sg13g2_nand2_1 _20702_ (.Y(_13020_),
    .A(_12949_),
    .B(_12990_));
 sg13g2_nor2_1 _20703_ (.A(_12949_),
    .B(_12990_),
    .Y(_13021_));
 sg13g2_a21oi_1 _20704_ (.A1(_12950_),
    .A2(_13020_),
    .Y(_13022_),
    .B1(_13021_));
 sg13g2_buf_1 _20705_ (.A(net506),
    .X(_13023_));
 sg13g2_and2_1 _20706_ (.A(net481),
    .B(_12918_),
    .X(_13024_));
 sg13g2_nor2_1 _20707_ (.A(_12420_),
    .B(net278),
    .Y(_13025_));
 sg13g2_nand2_1 _20708_ (.Y(_13026_),
    .A(net520),
    .B(net211));
 sg13g2_xnor2_1 _20709_ (.Y(_13027_),
    .A(_13025_),
    .B(_13026_));
 sg13g2_xnor2_1 _20710_ (.Y(_13028_),
    .A(_13024_),
    .B(_13027_));
 sg13g2_nand3_1 _20711_ (.B(net211),
    .C(_12908_),
    .A(net481),
    .Y(_13029_));
 sg13g2_a21oi_1 _20712_ (.A1(net481),
    .A2(net211),
    .Y(_13030_),
    .B1(_12908_));
 sg13g2_a21o_1 _20713_ (.A2(_13029_),
    .A1(_12907_),
    .B1(_13030_),
    .X(_13031_));
 sg13g2_buf_1 _20714_ (.A(_13031_),
    .X(_13032_));
 sg13g2_buf_1 _20715_ (.A(\rbzero.wall_tracer.size_full[6] ),
    .X(_13033_));
 sg13g2_or2_1 _20716_ (.X(_13034_),
    .B(_12797_),
    .A(_12701_));
 sg13g2_nor4_2 _20717_ (.A(_11727_),
    .B(_12911_),
    .C(_12604_),
    .Y(_13035_),
    .D(_13034_));
 sg13g2_xor2_1 _20718_ (.B(_13035_),
    .A(_13033_),
    .X(_13036_));
 sg13g2_o21ai_1 _20719_ (.B1(_12800_),
    .Y(_13037_),
    .A1(net685),
    .A2(_13036_));
 sg13g2_o21ai_1 _20720_ (.B1(_13037_),
    .Y(_13038_),
    .A1(net697),
    .A2(_00463_));
 sg13g2_nand2_1 _20721_ (.Y(_13039_),
    .A(_08446_),
    .B(_00462_));
 sg13g2_o21ai_1 _20722_ (.B1(_13039_),
    .Y(_13040_),
    .A1(_08446_),
    .A2(_13038_));
 sg13g2_buf_1 _20723_ (.A(_13040_),
    .X(_13041_));
 sg13g2_nor2_1 _20724_ (.A(net521),
    .B(_13041_),
    .Y(_13042_));
 sg13g2_xnor2_1 _20725_ (.Y(_13043_),
    .A(_13032_),
    .B(_13042_));
 sg13g2_xnor2_1 _20726_ (.Y(_13044_),
    .A(_13028_),
    .B(_13043_));
 sg13g2_nor2_1 _20727_ (.A(_12935_),
    .B(_12938_),
    .Y(_13045_));
 sg13g2_nor2_1 _20728_ (.A(_12931_),
    .B(_13045_),
    .Y(_13046_));
 sg13g2_a21oi_1 _20729_ (.A1(_12935_),
    .A2(_12938_),
    .Y(_13047_),
    .B1(_13046_));
 sg13g2_nand2_1 _20730_ (.Y(_13048_),
    .A(net238),
    .B(net277));
 sg13g2_buf_1 _20731_ (.A(net239),
    .X(_13049_));
 sg13g2_nand2_1 _20732_ (.Y(_13050_),
    .A(net210),
    .B(net276));
 sg13g2_nand2_1 _20733_ (.Y(_13051_),
    .A(net260),
    .B(net292));
 sg13g2_xnor2_1 _20734_ (.Y(_13052_),
    .A(_13050_),
    .B(_13051_));
 sg13g2_xnor2_1 _20735_ (.Y(_13053_),
    .A(_13048_),
    .B(_13052_));
 sg13g2_a21oi_1 _20736_ (.A1(_12954_),
    .A2(_12955_),
    .Y(_13054_),
    .B1(_12956_));
 sg13g2_nor2_1 _20737_ (.A(_12954_),
    .B(_12955_),
    .Y(_13055_));
 sg13g2_nor2_1 _20738_ (.A(_13054_),
    .B(_13055_),
    .Y(_13056_));
 sg13g2_o21ai_1 _20739_ (.B1(_12929_),
    .Y(_13057_),
    .A1(_12926_),
    .A2(_12927_));
 sg13g2_nand2_1 _20740_ (.Y(_13058_),
    .A(_12926_),
    .B(_12927_));
 sg13g2_nand2_1 _20741_ (.Y(_13059_),
    .A(_13057_),
    .B(_13058_));
 sg13g2_xnor2_1 _20742_ (.Y(_13060_),
    .A(_13056_),
    .B(_13059_));
 sg13g2_xnor2_1 _20743_ (.Y(_13061_),
    .A(_13053_),
    .B(_13060_));
 sg13g2_nor2_1 _20744_ (.A(_13047_),
    .B(_13061_),
    .Y(_13062_));
 sg13g2_nand2_1 _20745_ (.Y(_13063_),
    .A(_13047_),
    .B(_13061_));
 sg13g2_nand2b_1 _20746_ (.Y(_13064_),
    .B(_13063_),
    .A_N(_13062_));
 sg13g2_xnor2_1 _20747_ (.Y(_13065_),
    .A(_13044_),
    .B(_13064_));
 sg13g2_nand2_1 _20748_ (.Y(_13066_),
    .A(_12924_),
    .B(_12940_));
 sg13g2_nor2_1 _20749_ (.A(_12924_),
    .B(_12940_),
    .Y(_13067_));
 sg13g2_a21oi_1 _20750_ (.A1(_12921_),
    .A2(_13066_),
    .Y(_13068_),
    .B1(_13067_));
 sg13g2_nand2b_1 _20751_ (.Y(_13069_),
    .B(_12971_),
    .A_N(_12969_));
 sg13g2_nor2b_1 _20752_ (.A(_12971_),
    .B_N(_12969_),
    .Y(_13070_));
 sg13g2_a21oi_1 _20753_ (.A1(_12953_),
    .A2(_13069_),
    .Y(_13071_),
    .B1(_13070_));
 sg13g2_xnor2_1 _20754_ (.Y(_13072_),
    .A(_13068_),
    .B(_13071_));
 sg13g2_xnor2_1 _20755_ (.Y(_13073_),
    .A(_13065_),
    .B(_13072_));
 sg13g2_nand2b_1 _20756_ (.Y(_13074_),
    .B(_12989_),
    .A_N(_12973_));
 sg13g2_nand2_1 _20757_ (.Y(_13075_),
    .A(_12958_),
    .B(_12967_));
 sg13g2_nor2_1 _20758_ (.A(_12958_),
    .B(_12967_),
    .Y(_13076_));
 sg13g2_a21oi_2 _20759_ (.B1(_13076_),
    .Y(_13077_),
    .A2(_13075_),
    .A1(_12962_));
 sg13g2_nand2b_1 _20760_ (.Y(_13078_),
    .B(_12983_),
    .A_N(_12977_));
 sg13g2_o21ai_1 _20761_ (.B1(_12964_),
    .Y(_13079_),
    .A1(_12963_),
    .A2(_12965_));
 sg13g2_nand2_1 _20762_ (.Y(_13080_),
    .A(_12963_),
    .B(_12965_));
 sg13g2_and2_1 _20763_ (.A(_13079_),
    .B(_13080_),
    .X(_13081_));
 sg13g2_nand2_1 _20764_ (.Y(_13082_),
    .A(net261),
    .B(net306));
 sg13g2_nand2_1 _20765_ (.Y(_13083_),
    .A(_11999_),
    .B(net293));
 sg13g2_nand2_1 _20766_ (.Y(_13084_),
    .A(net263),
    .B(net307));
 sg13g2_xnor2_1 _20767_ (.Y(_13085_),
    .A(_13083_),
    .B(_13084_));
 sg13g2_xnor2_1 _20768_ (.Y(_13086_),
    .A(_13082_),
    .B(_13085_));
 sg13g2_nand2_1 _20769_ (.Y(_13087_),
    .A(net280),
    .B(net333));
 sg13g2_nor2_1 _20770_ (.A(_11913_),
    .B(_12630_),
    .Y(_13088_));
 sg13g2_nand2_1 _20771_ (.Y(_13089_),
    .A(net264),
    .B(net332));
 sg13g2_xor2_1 _20772_ (.B(_13089_),
    .A(_13088_),
    .X(_13090_));
 sg13g2_xnor2_1 _20773_ (.Y(_13091_),
    .A(_13087_),
    .B(_13090_));
 sg13g2_xor2_1 _20774_ (.B(_13091_),
    .A(_13086_),
    .X(_13092_));
 sg13g2_xnor2_1 _20775_ (.Y(_13093_),
    .A(_13081_),
    .B(_13092_));
 sg13g2_xnor2_1 _20776_ (.Y(_13094_),
    .A(_13078_),
    .B(_13093_));
 sg13g2_xnor2_1 _20777_ (.Y(_13095_),
    .A(_13077_),
    .B(_13094_));
 sg13g2_nor2_1 _20778_ (.A(_12984_),
    .B(_12988_),
    .Y(_13096_));
 sg13g2_and2_1 _20779_ (.A(_08546_),
    .B(_12727_),
    .X(_13097_));
 sg13g2_buf_1 _20780_ (.A(_13097_),
    .X(_13098_));
 sg13g2_nand2_1 _20781_ (.Y(_13099_),
    .A(net443),
    .B(_13098_));
 sg13g2_nand2_1 _20782_ (.Y(_13100_),
    .A(net445),
    .B(_12986_));
 sg13g2_xnor2_1 _20783_ (.Y(_13101_),
    .A(_13099_),
    .B(_13100_));
 sg13g2_o21ai_1 _20784_ (.B1(_12981_),
    .Y(_13102_),
    .A1(_12978_),
    .A2(_12980_));
 sg13g2_nand2_1 _20785_ (.Y(_13103_),
    .A(_12978_),
    .B(_12980_));
 sg13g2_nand2_1 _20786_ (.Y(_13104_),
    .A(net406),
    .B(_12642_));
 sg13g2_nand2_1 _20787_ (.Y(_13105_),
    .A(_12166_),
    .B(net518));
 sg13g2_nand2_1 _20788_ (.Y(_13106_),
    .A(net405),
    .B(net519));
 sg13g2_xnor2_1 _20789_ (.Y(_13107_),
    .A(_13105_),
    .B(_13106_));
 sg13g2_xnor2_1 _20790_ (.Y(_13108_),
    .A(_13104_),
    .B(_13107_));
 sg13g2_a21oi_2 _20791_ (.B1(_13108_),
    .Y(_13109_),
    .A2(_13103_),
    .A1(_13102_));
 sg13g2_nand3_1 _20792_ (.B(_13103_),
    .C(_13108_),
    .A(_13102_),
    .Y(_13110_));
 sg13g2_nor2b_1 _20793_ (.A(_13109_),
    .B_N(_13110_),
    .Y(_13111_));
 sg13g2_xnor2_1 _20794_ (.Y(_13112_),
    .A(_13101_),
    .B(_13111_));
 sg13g2_xnor2_1 _20795_ (.Y(_13113_),
    .A(_13096_),
    .B(_13112_));
 sg13g2_xnor2_1 _20796_ (.Y(_13114_),
    .A(_13095_),
    .B(_13113_));
 sg13g2_xor2_1 _20797_ (.B(_13114_),
    .A(_13074_),
    .X(_13115_));
 sg13g2_xnor2_1 _20798_ (.Y(_13116_),
    .A(_13073_),
    .B(_13115_));
 sg13g2_a21o_1 _20799_ (.A2(_12947_),
    .A1(_12942_),
    .B1(_12945_),
    .X(_13117_));
 sg13g2_o21ai_1 _20800_ (.B1(_13117_),
    .Y(_13118_),
    .A1(_12942_),
    .A2(_12947_));
 sg13g2_nor2_1 _20801_ (.A(_12904_),
    .B(_12910_),
    .Y(_13119_));
 sg13g2_nand2_1 _20802_ (.Y(_13120_),
    .A(_12904_),
    .B(_12910_));
 sg13g2_o21ai_1 _20803_ (.B1(_13120_),
    .Y(_13121_),
    .A1(_12919_),
    .A2(_13119_));
 sg13g2_xor2_1 _20804_ (.B(_13121_),
    .A(_13118_),
    .X(_13122_));
 sg13g2_xnor2_1 _20805_ (.Y(_13123_),
    .A(_13116_),
    .B(_13122_));
 sg13g2_xnor2_1 _20806_ (.Y(_13124_),
    .A(_13022_),
    .B(_13123_));
 sg13g2_xnor2_1 _20807_ (.Y(_13125_),
    .A(_13019_),
    .B(_13124_));
 sg13g2_xnor2_1 _20808_ (.Y(_13126_),
    .A(_13018_),
    .B(_13125_));
 sg13g2_buf_1 _20809_ (.A(_13126_),
    .X(_13127_));
 sg13g2_nor2_1 _20810_ (.A(_13008_),
    .B(_13003_),
    .Y(_13128_));
 sg13g2_nand2_2 _20811_ (.Y(_13129_),
    .A(_13008_),
    .B(_13003_));
 sg13g2_o21ai_1 _20812_ (.B1(_13129_),
    .Y(_13130_),
    .A1(_12899_),
    .A2(_13128_));
 sg13g2_nand2_1 _20813_ (.Y(_13131_),
    .A(_12899_),
    .B(_13128_));
 sg13g2_o21ai_1 _20814_ (.B1(_13131_),
    .Y(_13132_),
    .A1(_12896_),
    .A2(_13130_));
 sg13g2_nor2_1 _20815_ (.A(_13005_),
    .B(_13132_),
    .Y(_13133_));
 sg13g2_nor2_1 _20816_ (.A(_12899_),
    .B(_13129_),
    .Y(_13134_));
 sg13g2_a21oi_1 _20817_ (.A1(_12896_),
    .A2(_13130_),
    .Y(_13135_),
    .B1(_13134_));
 sg13g2_and2_1 _20818_ (.A(_13005_),
    .B(_13135_),
    .X(_13136_));
 sg13g2_and2_1 _20819_ (.A(_12896_),
    .B(_12900_),
    .X(_13137_));
 sg13g2_buf_1 _20820_ (.A(_13137_),
    .X(_13138_));
 sg13g2_nand2b_1 _20821_ (.Y(_13139_),
    .B(_13138_),
    .A_N(_13129_));
 sg13g2_o21ai_1 _20822_ (.B1(_13139_),
    .Y(_13140_),
    .A1(_13133_),
    .A2(_13136_));
 sg13g2_xnor2_1 _20823_ (.Y(_13141_),
    .A(_13127_),
    .B(_13140_));
 sg13g2_buf_2 _20824_ (.A(_13141_),
    .X(_13142_));
 sg13g2_nand2_1 _20825_ (.Y(_13143_),
    .A(_11715_),
    .B(_13142_));
 sg13g2_buf_2 _20826_ (.A(\rbzero.traced_texVinit[3] ),
    .X(_13144_));
 sg13g2_nand2_1 _20827_ (.Y(_13145_),
    .A(_13144_),
    .B(net448));
 sg13g2_a21oi_1 _20828_ (.A1(_13143_),
    .A2(_13145_),
    .Y(_01513_),
    .B1(net572));
 sg13g2_buf_1 _20829_ (.A(\rbzero.traced_texVinit[4] ),
    .X(_13146_));
 sg13g2_nor2_1 _20830_ (.A(_13146_),
    .B(_11714_),
    .Y(_13147_));
 sg13g2_nand2_1 _20831_ (.Y(_13148_),
    .A(_13127_),
    .B(_13129_));
 sg13g2_nand2b_1 _20832_ (.Y(_13149_),
    .B(_12899_),
    .A_N(_12896_));
 sg13g2_a21o_1 _20833_ (.A2(_13149_),
    .A1(_13005_),
    .B1(_13138_),
    .X(_13150_));
 sg13g2_nand2b_1 _20834_ (.Y(_13151_),
    .B(_13127_),
    .A_N(_13138_));
 sg13g2_nor2b_1 _20835_ (.A(_13127_),
    .B_N(_13149_),
    .Y(_13152_));
 sg13g2_a21o_1 _20836_ (.A2(_13151_),
    .A1(_13005_),
    .B1(_13152_),
    .X(_13153_));
 sg13g2_inv_1 _20837_ (.Y(_13154_),
    .A(_13128_));
 sg13g2_nor2_1 _20838_ (.A(_13127_),
    .B(_13129_),
    .Y(_13155_));
 sg13g2_a221oi_1 _20839_ (.B2(_13154_),
    .C1(_13155_),
    .B1(_13153_),
    .A1(_13148_),
    .Y(_13156_),
    .A2(_13150_));
 sg13g2_nor2_1 _20840_ (.A(_13056_),
    .B(_13059_),
    .Y(_13157_));
 sg13g2_a21oi_1 _20841_ (.A1(_13056_),
    .A2(_13059_),
    .Y(_13158_),
    .B1(_13053_));
 sg13g2_nor2_1 _20842_ (.A(_13157_),
    .B(_13158_),
    .Y(_13159_));
 sg13g2_buf_1 _20843_ (.A(net260),
    .X(_13160_));
 sg13g2_nand2_1 _20844_ (.Y(_13161_),
    .A(net237),
    .B(net276));
 sg13g2_nand2_1 _20845_ (.Y(_13162_),
    .A(net210),
    .B(net277));
 sg13g2_nor2_1 _20846_ (.A(net279),
    .B(net278),
    .Y(_13163_));
 sg13g2_xor2_1 _20847_ (.B(_13163_),
    .A(_13162_),
    .X(_13164_));
 sg13g2_xnor2_1 _20848_ (.Y(_13165_),
    .A(_13161_),
    .B(_13164_));
 sg13g2_a21o_1 _20849_ (.A2(_13083_),
    .A1(_13082_),
    .B1(_13084_),
    .X(_13166_));
 sg13g2_o21ai_1 _20850_ (.B1(_13166_),
    .Y(_13167_),
    .A1(_13082_),
    .A2(_13083_));
 sg13g2_xor2_1 _20851_ (.B(_13167_),
    .A(_13165_),
    .X(_13168_));
 sg13g2_a21o_1 _20852_ (.A2(_13050_),
    .A1(_13048_),
    .B1(_13051_),
    .X(_13169_));
 sg13g2_o21ai_1 _20853_ (.B1(_13169_),
    .Y(_13170_),
    .A1(_13048_),
    .A2(_13050_));
 sg13g2_xnor2_1 _20854_ (.Y(_13171_),
    .A(_13168_),
    .B(_13170_));
 sg13g2_nor2_1 _20855_ (.A(net504),
    .B(_13041_),
    .Y(_13172_));
 sg13g2_nand2_1 _20856_ (.Y(_13173_),
    .A(_11781_),
    .B(net211));
 sg13g2_buf_1 _20857_ (.A(_12918_),
    .X(_13174_));
 sg13g2_nand2_1 _20858_ (.Y(_13175_),
    .A(net520),
    .B(net209));
 sg13g2_xnor2_1 _20859_ (.Y(_13176_),
    .A(_13173_),
    .B(_13175_));
 sg13g2_xnor2_1 _20860_ (.Y(_13177_),
    .A(_13172_),
    .B(_13176_));
 sg13g2_nand2b_1 _20861_ (.Y(_13178_),
    .B(_13026_),
    .A_N(_13025_));
 sg13g2_buf_1 _20862_ (.A(_12709_),
    .X(_13179_));
 sg13g2_nor3_1 _20863_ (.A(_12420_),
    .B(_13179_),
    .C(_13026_),
    .Y(_13180_));
 sg13g2_a21oi_2 _20864_ (.B1(_13180_),
    .Y(_13181_),
    .A2(_13178_),
    .A1(_13024_));
 sg13g2_buf_1 _20865_ (.A(\rbzero.wall_tracer.size_full[7] ),
    .X(_13182_));
 sg13g2_nor3_1 _20866_ (.A(_12911_),
    .B(_13033_),
    .C(_13034_),
    .Y(_13183_));
 sg13g2_nand2_1 _20867_ (.Y(_13184_),
    .A(_12702_),
    .B(_13183_));
 sg13g2_xnor2_1 _20868_ (.Y(_13185_),
    .A(_13182_),
    .B(_13184_));
 sg13g2_o21ai_1 _20869_ (.B1(_12800_),
    .Y(_13186_),
    .A1(net685),
    .A2(_13185_));
 sg13g2_o21ai_1 _20870_ (.B1(_13186_),
    .Y(_13187_),
    .A1(net697),
    .A2(_00465_));
 sg13g2_nand2_1 _20871_ (.Y(_13188_),
    .A(net611),
    .B(_00464_));
 sg13g2_o21ai_1 _20872_ (.B1(_13188_),
    .Y(_13189_),
    .A1(net611),
    .A2(_13187_));
 sg13g2_buf_1 _20873_ (.A(_13189_),
    .X(_13190_));
 sg13g2_buf_1 _20874_ (.A(_13190_),
    .X(_13191_));
 sg13g2_nor2_1 _20875_ (.A(_12415_),
    .B(net208),
    .Y(_13192_));
 sg13g2_xor2_1 _20876_ (.B(_13192_),
    .A(_13181_),
    .X(_13193_));
 sg13g2_xnor2_1 _20877_ (.Y(_13194_),
    .A(_13177_),
    .B(_13193_));
 sg13g2_nor2_1 _20878_ (.A(_13171_),
    .B(_13194_),
    .Y(_13195_));
 sg13g2_nand2_1 _20879_ (.Y(_13196_),
    .A(_13171_),
    .B(_13194_));
 sg13g2_nor2b_1 _20880_ (.A(_13195_),
    .B_N(_13196_),
    .Y(_13197_));
 sg13g2_xnor2_1 _20881_ (.Y(_13198_),
    .A(_13159_),
    .B(_13197_));
 sg13g2_a21oi_1 _20882_ (.A1(_13044_),
    .A2(_13063_),
    .Y(_13199_),
    .B1(_13062_));
 sg13g2_a21o_1 _20883_ (.A2(_13093_),
    .A1(_13077_),
    .B1(_13078_),
    .X(_13200_));
 sg13g2_o21ai_1 _20884_ (.B1(_13200_),
    .Y(_13201_),
    .A1(_13077_),
    .A2(_13093_));
 sg13g2_buf_1 _20885_ (.A(_13201_),
    .X(_13202_));
 sg13g2_xor2_1 _20886_ (.B(_13202_),
    .A(_13199_),
    .X(_13203_));
 sg13g2_xnor2_1 _20887_ (.Y(_13204_),
    .A(_13198_),
    .B(_13203_));
 sg13g2_inv_1 _20888_ (.Y(_13205_),
    .A(_13095_));
 sg13g2_nor2_1 _20889_ (.A(_13205_),
    .B(_13112_),
    .Y(_13206_));
 sg13g2_a21oi_1 _20890_ (.A1(_13205_),
    .A2(_13112_),
    .Y(_13207_),
    .B1(_13096_));
 sg13g2_nand2_1 _20891_ (.Y(_13208_),
    .A(_13086_),
    .B(_13091_));
 sg13g2_nor2_1 _20892_ (.A(_13086_),
    .B(_13091_),
    .Y(_13209_));
 sg13g2_a21oi_2 _20893_ (.B1(_13209_),
    .Y(_13210_),
    .A2(_13208_),
    .A1(_13081_));
 sg13g2_nand2_1 _20894_ (.Y(_13211_),
    .A(net261),
    .B(net292));
 sg13g2_nand2_1 _20895_ (.Y(_13212_),
    .A(net240),
    .B(net306));
 sg13g2_nand2_1 _20896_ (.Y(_13213_),
    .A(net263),
    .B(net293));
 sg13g2_xnor2_1 _20897_ (.Y(_13214_),
    .A(_13212_),
    .B(_13213_));
 sg13g2_xnor2_1 _20898_ (.Y(_13215_),
    .A(_13211_),
    .B(_13214_));
 sg13g2_buf_1 _20899_ (.A(net333),
    .X(_13216_));
 sg13g2_nand3_1 _20900_ (.B(net319),
    .C(_13088_),
    .A(net259),
    .Y(_13217_));
 sg13g2_a21oi_1 _20901_ (.A1(net259),
    .A2(net319),
    .Y(_13218_),
    .B1(_13088_));
 sg13g2_a21o_1 _20902_ (.A2(_13217_),
    .A1(_13089_),
    .B1(_13218_),
    .X(_13219_));
 sg13g2_buf_1 _20903_ (.A(_13219_),
    .X(_13220_));
 sg13g2_buf_1 _20904_ (.A(net307),
    .X(_13221_));
 sg13g2_nand2_1 _20905_ (.Y(_13222_),
    .A(_12959_),
    .B(net301));
 sg13g2_nor2_1 _20906_ (.A(_12069_),
    .B(_12630_),
    .Y(_13223_));
 sg13g2_nand2_1 _20907_ (.Y(_13224_),
    .A(net264),
    .B(net333));
 sg13g2_xnor2_1 _20908_ (.Y(_13225_),
    .A(_13223_),
    .B(_13224_));
 sg13g2_xnor2_1 _20909_ (.Y(_13226_),
    .A(_13222_),
    .B(_13225_));
 sg13g2_xor2_1 _20910_ (.B(_13226_),
    .A(_13220_),
    .X(_13227_));
 sg13g2_xnor2_1 _20911_ (.Y(_13228_),
    .A(_13215_),
    .B(_13227_));
 sg13g2_xor2_1 _20912_ (.B(_13228_),
    .A(_13109_),
    .X(_13229_));
 sg13g2_xnor2_1 _20913_ (.Y(_13230_),
    .A(_13210_),
    .B(_13229_));
 sg13g2_nor2b_1 _20914_ (.A(_13101_),
    .B_N(_13111_),
    .Y(_13231_));
 sg13g2_nor2_1 _20915_ (.A(_11913_),
    .B(net503),
    .Y(_13232_));
 sg13g2_a21oi_2 _20916_ (.B1(_12979_),
    .Y(_13233_),
    .A2(_11956_),
    .A1(_11949_));
 sg13g2_nand2_1 _20917_ (.Y(_13234_),
    .A(_12217_),
    .B(net519));
 sg13g2_xor2_1 _20918_ (.B(_13234_),
    .A(_13233_),
    .X(_13235_));
 sg13g2_xnor2_1 _20919_ (.Y(_13236_),
    .A(_13232_),
    .B(_13235_));
 sg13g2_a21o_1 _20920_ (.A2(_13104_),
    .A1(_13105_),
    .B1(_13106_),
    .X(_13237_));
 sg13g2_o21ai_1 _20921_ (.B1(_13237_),
    .Y(_13238_),
    .A1(_13105_),
    .A2(_13104_));
 sg13g2_buf_1 _20922_ (.A(_13238_),
    .X(_13239_));
 sg13g2_nand2_1 _20923_ (.Y(_13240_),
    .A(_12244_),
    .B(_13098_));
 sg13g2_or2_1 _20924_ (.X(_13241_),
    .B(_13240_),
    .A(_12988_));
 sg13g2_xor2_1 _20925_ (.B(_13241_),
    .A(_13239_),
    .X(_13242_));
 sg13g2_xnor2_1 _20926_ (.Y(_13243_),
    .A(_13236_),
    .B(_13242_));
 sg13g2_nand2_1 _20927_ (.Y(_13244_),
    .A(_12974_),
    .B(net482));
 sg13g2_and2_1 _20928_ (.A(_08545_),
    .B(net567),
    .X(_13245_));
 sg13g2_buf_1 _20929_ (.A(_13245_),
    .X(_13246_));
 sg13g2_nand2_1 _20930_ (.Y(_13247_),
    .A(_12423_),
    .B(net502));
 sg13g2_xor2_1 _20931_ (.B(_13247_),
    .A(_13240_),
    .X(_13248_));
 sg13g2_xnor2_1 _20932_ (.Y(_13249_),
    .A(_13244_),
    .B(_13248_));
 sg13g2_xor2_1 _20933_ (.B(_13249_),
    .A(_13243_),
    .X(_13250_));
 sg13g2_xnor2_1 _20934_ (.Y(_13251_),
    .A(_13231_),
    .B(_13250_));
 sg13g2_xnor2_1 _20935_ (.Y(_13252_),
    .A(_13230_),
    .B(_13251_));
 sg13g2_o21ai_1 _20936_ (.B1(_13252_),
    .Y(_13253_),
    .A1(_13206_),
    .A2(_13207_));
 sg13g2_or3_1 _20937_ (.A(_13252_),
    .B(_13206_),
    .C(_13207_),
    .X(_13254_));
 sg13g2_nand2_1 _20938_ (.Y(_13255_),
    .A(_13253_),
    .B(_13254_));
 sg13g2_xor2_1 _20939_ (.B(_13255_),
    .A(_13204_),
    .X(_13256_));
 sg13g2_nand2_1 _20940_ (.Y(_13257_),
    .A(_13073_),
    .B(_13114_));
 sg13g2_o21ai_1 _20941_ (.B1(_13074_),
    .Y(_13258_),
    .A1(_13073_),
    .A2(_13114_));
 sg13g2_nand2_1 _20942_ (.Y(_13259_),
    .A(_13257_),
    .B(_13258_));
 sg13g2_nand2_1 _20943_ (.Y(_13260_),
    .A(_13065_),
    .B(_13071_));
 sg13g2_nor2_1 _20944_ (.A(_13065_),
    .B(_13071_),
    .Y(_13261_));
 sg13g2_a21oi_1 _20945_ (.A1(_13068_),
    .A2(_13260_),
    .Y(_13262_),
    .B1(_13261_));
 sg13g2_nand2_1 _20946_ (.Y(_13263_),
    .A(_13032_),
    .B(_13028_));
 sg13g2_nor2_1 _20947_ (.A(_13032_),
    .B(_13028_),
    .Y(_13264_));
 sg13g2_a21oi_1 _20948_ (.A1(_13042_),
    .A2(_13263_),
    .Y(_13265_),
    .B1(_13264_));
 sg13g2_xor2_1 _20949_ (.B(_13265_),
    .A(_13262_),
    .X(_13266_));
 sg13g2_xor2_1 _20950_ (.B(_13266_),
    .A(_13259_),
    .X(_13267_));
 sg13g2_xnor2_1 _20951_ (.Y(_13268_),
    .A(_13256_),
    .B(_13267_));
 sg13g2_nand2_1 _20952_ (.Y(_13269_),
    .A(_13118_),
    .B(_13121_));
 sg13g2_nand2_1 _20953_ (.Y(_13270_),
    .A(_13116_),
    .B(_13122_));
 sg13g2_nor2_1 _20954_ (.A(_13116_),
    .B(_13122_),
    .Y(_13271_));
 sg13g2_a21oi_1 _20955_ (.A1(_13022_),
    .A2(_13270_),
    .Y(_13272_),
    .B1(_13271_));
 sg13g2_xnor2_1 _20956_ (.Y(_13273_),
    .A(_13269_),
    .B(_13272_));
 sg13g2_xnor2_1 _20957_ (.Y(_13274_),
    .A(_13268_),
    .B(_13273_));
 sg13g2_nand2_1 _20958_ (.Y(_13275_),
    .A(_13018_),
    .B(_13124_));
 sg13g2_nor2_1 _20959_ (.A(_13018_),
    .B(_13124_),
    .Y(_13276_));
 sg13g2_a21oi_1 _20960_ (.A1(_13019_),
    .A2(_13275_),
    .Y(_13277_),
    .B1(_13276_));
 sg13g2_or2_1 _20961_ (.X(_13278_),
    .B(_13277_),
    .A(_13274_));
 sg13g2_nand2_1 _20962_ (.Y(_13279_),
    .A(_13274_),
    .B(_13277_));
 sg13g2_nand2_1 _20963_ (.Y(_13280_),
    .A(_13278_),
    .B(_13279_));
 sg13g2_xnor2_1 _20964_ (.Y(_13281_),
    .A(_13156_),
    .B(_13280_));
 sg13g2_buf_2 _20965_ (.A(_13281_),
    .X(_13282_));
 sg13g2_nor2_1 _20966_ (.A(net464),
    .B(_13282_),
    .Y(_13283_));
 sg13g2_nor3_1 _20967_ (.A(net629),
    .B(_13147_),
    .C(_13283_),
    .Y(_01514_));
 sg13g2_buf_1 _20968_ (.A(\rbzero.traced_texVinit[5] ),
    .X(_13284_));
 sg13g2_inv_1 _20969_ (.Y(_13285_),
    .A(_13278_));
 sg13g2_a21o_1 _20970_ (.A2(_13279_),
    .A1(_13156_),
    .B1(_13285_),
    .X(_13286_));
 sg13g2_buf_1 _20971_ (.A(_13286_),
    .X(_13287_));
 sg13g2_nand2_1 _20972_ (.Y(_13288_),
    .A(_13272_),
    .B(_13268_));
 sg13g2_nand2_1 _20973_ (.Y(_13289_),
    .A(_13269_),
    .B(_13288_));
 sg13g2_o21ai_1 _20974_ (.B1(_13289_),
    .Y(_13290_),
    .A1(_13272_),
    .A2(_13268_));
 sg13g2_buf_1 _20975_ (.A(_13290_),
    .X(_13291_));
 sg13g2_a21oi_1 _20976_ (.A1(_13256_),
    .A2(_13266_),
    .Y(_13292_),
    .B1(_13259_));
 sg13g2_nor2_1 _20977_ (.A(_13256_),
    .B(_13266_),
    .Y(_13293_));
 sg13g2_nor2_1 _20978_ (.A(_13292_),
    .B(_13293_),
    .Y(_13294_));
 sg13g2_nor2b_1 _20979_ (.A(_13265_),
    .B_N(_13262_),
    .Y(_13295_));
 sg13g2_o21ai_1 _20980_ (.B1(_13196_),
    .Y(_13296_),
    .A1(_13159_),
    .A2(_13195_));
 sg13g2_nand2b_1 _20981_ (.Y(_13297_),
    .B(_13165_),
    .A_N(_13167_));
 sg13g2_nor2b_1 _20982_ (.A(_13165_),
    .B_N(_13167_),
    .Y(_13298_));
 sg13g2_a21oi_1 _20983_ (.A1(_13297_),
    .A2(_13170_),
    .Y(_13299_),
    .B1(_13298_));
 sg13g2_nand2b_1 _20984_ (.Y(_13300_),
    .B(_13163_),
    .A_N(_13161_));
 sg13g2_a21oi_1 _20985_ (.A1(net237),
    .A2(net276),
    .Y(_13301_),
    .B1(_13163_));
 sg13g2_a21oi_1 _20986_ (.A1(_13162_),
    .A2(_13300_),
    .Y(_13302_),
    .B1(_13301_));
 sg13g2_nand2_1 _20987_ (.Y(_13303_),
    .A(net238),
    .B(net211));
 sg13g2_nand2_1 _20988_ (.Y(_13304_),
    .A(_12456_),
    .B(net277));
 sg13g2_nor2_1 _20989_ (.A(net262),
    .B(net278),
    .Y(_13305_));
 sg13g2_xor2_1 _20990_ (.B(_13305_),
    .A(_13304_),
    .X(_13306_));
 sg13g2_xnor2_1 _20991_ (.Y(_13307_),
    .A(_13303_),
    .B(_13306_));
 sg13g2_a21o_1 _20992_ (.A2(_13212_),
    .A1(_13211_),
    .B1(_13213_),
    .X(_13308_));
 sg13g2_o21ai_1 _20993_ (.B1(_13308_),
    .Y(_13309_),
    .A1(_13211_),
    .A2(_13212_));
 sg13g2_xnor2_1 _20994_ (.Y(_13310_),
    .A(_13307_),
    .B(_13309_));
 sg13g2_xnor2_1 _20995_ (.Y(_13311_),
    .A(_13302_),
    .B(_13310_));
 sg13g2_nand2_1 _20996_ (.Y(_13312_),
    .A(net268),
    .B(net209));
 sg13g2_nor2_1 _20997_ (.A(net504),
    .B(_13190_),
    .Y(_13313_));
 sg13g2_nor2_1 _20998_ (.A(net568),
    .B(_13041_),
    .Y(_13314_));
 sg13g2_xor2_1 _20999_ (.B(_13314_),
    .A(_13313_),
    .X(_13315_));
 sg13g2_xnor2_1 _21000_ (.Y(_13316_),
    .A(_13312_),
    .B(_13315_));
 sg13g2_nand3_1 _21001_ (.B(net209),
    .C(_13172_),
    .A(_12424_),
    .Y(_13317_));
 sg13g2_a21oi_1 _21002_ (.A1(_12424_),
    .A2(net209),
    .Y(_13318_),
    .B1(_13172_));
 sg13g2_a21oi_2 _21003_ (.B1(_13318_),
    .Y(_13319_),
    .A2(_13317_),
    .A1(_13173_));
 sg13g2_buf_1 _21004_ (.A(\rbzero.wall_tracer.size_full[8] ),
    .X(_13320_));
 sg13g2_or2_1 _21005_ (.X(_13321_),
    .B(_13184_),
    .A(_13182_));
 sg13g2_xnor2_1 _21006_ (.Y(_13322_),
    .A(_13320_),
    .B(_13321_));
 sg13g2_o21ai_1 _21007_ (.B1(_12800_),
    .Y(_13323_),
    .A1(net685),
    .A2(_13322_));
 sg13g2_o21ai_1 _21008_ (.B1(_13323_),
    .Y(_13324_),
    .A1(_12129_),
    .A2(_00467_));
 sg13g2_nand2_1 _21009_ (.Y(_13325_),
    .A(net522),
    .B(_13324_));
 sg13g2_o21ai_1 _21010_ (.B1(_13325_),
    .Y(_13326_),
    .A1(net522),
    .A2(_00466_));
 sg13g2_buf_1 _21011_ (.A(_13326_),
    .X(_13327_));
 sg13g2_nand2_1 _21012_ (.Y(_13328_),
    .A(_12363_),
    .B(_13327_));
 sg13g2_xor2_1 _21013_ (.B(_13328_),
    .A(_13319_),
    .X(_13329_));
 sg13g2_xnor2_1 _21014_ (.Y(_13330_),
    .A(_13316_),
    .B(_13329_));
 sg13g2_xor2_1 _21015_ (.B(_13330_),
    .A(_13311_),
    .X(_13331_));
 sg13g2_xnor2_1 _21016_ (.Y(_13332_),
    .A(_13299_),
    .B(_13331_));
 sg13g2_nor2_1 _21017_ (.A(_13210_),
    .B(_13228_),
    .Y(_13333_));
 sg13g2_nand2_1 _21018_ (.Y(_13334_),
    .A(_13210_),
    .B(_13228_));
 sg13g2_o21ai_1 _21019_ (.B1(_13334_),
    .Y(_13335_),
    .A1(_13109_),
    .A2(_13333_));
 sg13g2_buf_1 _21020_ (.A(_13335_),
    .X(_13336_));
 sg13g2_xor2_1 _21021_ (.B(_13336_),
    .A(_13332_),
    .X(_13337_));
 sg13g2_xnor2_1 _21022_ (.Y(_13338_),
    .A(_13296_),
    .B(_13337_));
 sg13g2_nand2_1 _21023_ (.Y(_13339_),
    .A(_13220_),
    .B(_13215_));
 sg13g2_nor2_1 _21024_ (.A(_13220_),
    .B(_13215_),
    .Y(_13340_));
 sg13g2_a21oi_1 _21025_ (.A1(_13226_),
    .A2(_13339_),
    .Y(_13341_),
    .B1(_13340_));
 sg13g2_nand2_1 _21026_ (.Y(_13342_),
    .A(net261),
    .B(net276));
 sg13g2_nand2_1 _21027_ (.Y(_13343_),
    .A(net263),
    .B(net306));
 sg13g2_nand2_1 _21028_ (.Y(_13344_),
    .A(net240),
    .B(net292));
 sg13g2_xnor2_1 _21029_ (.Y(_13345_),
    .A(_13343_),
    .B(_13344_));
 sg13g2_xnor2_1 _21030_ (.Y(_13346_),
    .A(_13342_),
    .B(_13345_));
 sg13g2_nand3_1 _21031_ (.B(net307),
    .C(_13223_),
    .A(net259),
    .Y(_13347_));
 sg13g2_a21oi_1 _21032_ (.A1(net259),
    .A2(net307),
    .Y(_13348_),
    .B1(_13223_));
 sg13g2_a21o_1 _21033_ (.A2(_13347_),
    .A1(_13224_),
    .B1(_13348_),
    .X(_13349_));
 sg13g2_buf_1 _21034_ (.A(_13349_),
    .X(_13350_));
 sg13g2_buf_1 _21035_ (.A(net259),
    .X(_13351_));
 sg13g2_nand2_1 _21036_ (.Y(_13352_),
    .A(net236),
    .B(net293));
 sg13g2_nand2_1 _21037_ (.Y(_13353_),
    .A(net319),
    .B(_12169_));
 sg13g2_nand2_1 _21038_ (.Y(_13354_),
    .A(_12135_),
    .B(_11794_));
 sg13g2_xor2_1 _21039_ (.B(_13354_),
    .A(_13353_),
    .X(_13355_));
 sg13g2_xnor2_1 _21040_ (.Y(_13356_),
    .A(_13352_),
    .B(_13355_));
 sg13g2_xor2_1 _21041_ (.B(_13356_),
    .A(_13350_),
    .X(_13357_));
 sg13g2_xnor2_1 _21042_ (.Y(_13358_),
    .A(_13346_),
    .B(_13357_));
 sg13g2_nor2_1 _21043_ (.A(_13236_),
    .B(_13239_),
    .Y(_13359_));
 sg13g2_nand2_1 _21044_ (.Y(_13360_),
    .A(_13236_),
    .B(_13239_));
 sg13g2_o21ai_1 _21045_ (.B1(_13360_),
    .Y(_13361_),
    .A1(_13241_),
    .A2(_13359_));
 sg13g2_buf_1 _21046_ (.A(_13361_),
    .X(_13362_));
 sg13g2_xor2_1 _21047_ (.B(_13362_),
    .A(_13358_),
    .X(_13363_));
 sg13g2_xnor2_1 _21048_ (.Y(_13364_),
    .A(_13341_),
    .B(_13363_));
 sg13g2_and2_1 _21049_ (.A(_13243_),
    .B(_13249_),
    .X(_13365_));
 sg13g2_nor2_1 _21050_ (.A(_12069_),
    .B(net503),
    .Y(_13366_));
 sg13g2_buf_1 _21051_ (.A(_12217_),
    .X(_13367_));
 sg13g2_buf_1 _21052_ (.A(net518),
    .X(_13368_));
 sg13g2_nand2_1 _21053_ (.Y(_13369_),
    .A(net362),
    .B(_13368_));
 sg13g2_nor2_1 _21054_ (.A(_11913_),
    .B(_12729_),
    .Y(_13370_));
 sg13g2_xor2_1 _21055_ (.B(_13370_),
    .A(_13369_),
    .X(_13371_));
 sg13g2_xnor2_1 _21056_ (.Y(_13372_),
    .A(_13366_),
    .B(_13371_));
 sg13g2_and2_1 _21057_ (.A(_13240_),
    .B(_13247_),
    .X(_13373_));
 sg13g2_or2_1 _21058_ (.X(_13374_),
    .B(_13247_),
    .A(_13240_));
 sg13g2_o21ai_1 _21059_ (.B1(_13374_),
    .Y(_13375_),
    .A1(_13244_),
    .A2(_13373_));
 sg13g2_buf_1 _21060_ (.A(_13375_),
    .X(_13376_));
 sg13g2_a22oi_1 _21061_ (.Y(_13377_),
    .B1(_13232_),
    .B2(_13233_),
    .A2(net519),
    .A1(_13367_));
 sg13g2_nor2_1 _21062_ (.A(_13232_),
    .B(_13233_),
    .Y(_13378_));
 sg13g2_nor2_1 _21063_ (.A(_13377_),
    .B(_13378_),
    .Y(_13379_));
 sg13g2_xnor2_1 _21064_ (.Y(_13380_),
    .A(_13376_),
    .B(_13379_));
 sg13g2_xnor2_1 _21065_ (.Y(_13381_),
    .A(_13372_),
    .B(_13380_));
 sg13g2_and2_1 _21066_ (.A(_08542_),
    .B(net567),
    .X(_13382_));
 sg13g2_buf_1 _21067_ (.A(_13382_),
    .X(_13383_));
 sg13g2_buf_1 _21068_ (.A(_13383_),
    .X(_13384_));
 sg13g2_nand2_1 _21069_ (.Y(_13385_),
    .A(_12423_),
    .B(net480));
 sg13g2_nand2_1 _21070_ (.Y(_13386_),
    .A(_08547_),
    .B(net567));
 sg13g2_buf_2 _21071_ (.A(_13386_),
    .X(_13387_));
 sg13g2_a21oi_2 _21072_ (.B1(_13387_),
    .Y(_13388_),
    .A2(_11956_),
    .A1(_11949_));
 sg13g2_and2_1 _21073_ (.A(_12244_),
    .B(net502),
    .X(_13389_));
 sg13g2_buf_1 _21074_ (.A(_13389_),
    .X(_13390_));
 sg13g2_buf_1 _21075_ (.A(_13098_),
    .X(_13391_));
 sg13g2_nand2_1 _21076_ (.Y(_13392_),
    .A(net404),
    .B(net479));
 sg13g2_xor2_1 _21077_ (.B(_13392_),
    .A(_13390_),
    .X(_13393_));
 sg13g2_xnor2_1 _21078_ (.Y(_13394_),
    .A(_13388_),
    .B(_13393_));
 sg13g2_xnor2_1 _21079_ (.Y(_13395_),
    .A(_13385_),
    .B(_13394_));
 sg13g2_xor2_1 _21080_ (.B(_13395_),
    .A(_13381_),
    .X(_13396_));
 sg13g2_xnor2_1 _21081_ (.Y(_13397_),
    .A(_13365_),
    .B(_13396_));
 sg13g2_xnor2_1 _21082_ (.Y(_13398_),
    .A(_13364_),
    .B(_13397_));
 sg13g2_inv_1 _21083_ (.Y(_13399_),
    .A(_13250_));
 sg13g2_nand2_1 _21084_ (.Y(_13400_),
    .A(_13230_),
    .B(_13399_));
 sg13g2_nor2_1 _21085_ (.A(_13230_),
    .B(_13399_),
    .Y(_13401_));
 sg13g2_a21oi_1 _21086_ (.A1(_13231_),
    .A2(_13400_),
    .Y(_13402_),
    .B1(_13401_));
 sg13g2_xnor2_1 _21087_ (.Y(_13403_),
    .A(_13398_),
    .B(_13402_));
 sg13g2_xnor2_1 _21088_ (.Y(_13404_),
    .A(_13338_),
    .B(_13403_));
 sg13g2_inv_1 _21089_ (.Y(_13405_),
    .A(_13254_));
 sg13g2_o21ai_1 _21090_ (.B1(_13253_),
    .Y(_13406_),
    .A1(_13204_),
    .A2(_13405_));
 sg13g2_buf_1 _21091_ (.A(_13406_),
    .X(_13407_));
 sg13g2_nand2_1 _21092_ (.Y(_13408_),
    .A(_13198_),
    .B(_13202_));
 sg13g2_nor2_1 _21093_ (.A(_13198_),
    .B(_13202_),
    .Y(_13409_));
 sg13g2_a21oi_1 _21094_ (.A1(_13199_),
    .A2(_13408_),
    .Y(_13410_),
    .B1(_13409_));
 sg13g2_nand2b_1 _21095_ (.Y(_13411_),
    .B(_13181_),
    .A_N(_13177_));
 sg13g2_nor2b_1 _21096_ (.A(_13181_),
    .B_N(_13177_),
    .Y(_13412_));
 sg13g2_a21oi_1 _21097_ (.A1(_13192_),
    .A2(_13411_),
    .Y(_13413_),
    .B1(_13412_));
 sg13g2_inv_1 _21098_ (.Y(_13414_),
    .A(_13413_));
 sg13g2_xnor2_1 _21099_ (.Y(_13415_),
    .A(_13410_),
    .B(_13414_));
 sg13g2_xnor2_1 _21100_ (.Y(_13416_),
    .A(_13407_),
    .B(_13415_));
 sg13g2_xnor2_1 _21101_ (.Y(_13417_),
    .A(_13404_),
    .B(_13416_));
 sg13g2_xnor2_1 _21102_ (.Y(_13418_),
    .A(_13295_),
    .B(_13417_));
 sg13g2_xnor2_1 _21103_ (.Y(_13419_),
    .A(_13294_),
    .B(_13418_));
 sg13g2_xnor2_1 _21104_ (.Y(_13420_),
    .A(_13291_),
    .B(_13419_));
 sg13g2_xnor2_1 _21105_ (.Y(_13421_),
    .A(_13287_),
    .B(_13420_));
 sg13g2_buf_2 _21106_ (.A(_13421_),
    .X(_13422_));
 sg13g2_nor2_1 _21107_ (.A(net464),
    .B(_13422_),
    .Y(_13423_));
 sg13g2_a21oi_1 _21108_ (.A1(_13284_),
    .A2(_08682_),
    .Y(_13424_),
    .B1(_13423_));
 sg13g2_nor2_1 _21109_ (.A(net634),
    .B(_13424_),
    .Y(_01515_));
 sg13g2_or2_1 _21110_ (.X(_13425_),
    .B(_13417_),
    .A(_13294_));
 sg13g2_nand2_1 _21111_ (.Y(_13426_),
    .A(_13294_),
    .B(_13417_));
 sg13g2_nand2_1 _21112_ (.Y(_13427_),
    .A(_13295_),
    .B(_13426_));
 sg13g2_a21o_1 _21113_ (.A2(_13415_),
    .A1(_13407_),
    .B1(_13404_),
    .X(_13428_));
 sg13g2_o21ai_1 _21114_ (.B1(_13428_),
    .Y(_13429_),
    .A1(_13407_),
    .A2(_13415_));
 sg13g2_buf_1 _21115_ (.A(_13429_),
    .X(_13430_));
 sg13g2_nand2_1 _21116_ (.Y(_13431_),
    .A(_13410_),
    .B(_13414_));
 sg13g2_nand2_1 _21117_ (.Y(_13432_),
    .A(_13350_),
    .B(_13346_));
 sg13g2_nor2_1 _21118_ (.A(_13350_),
    .B(_13346_),
    .Y(_13433_));
 sg13g2_a21oi_2 _21119_ (.B1(_13433_),
    .Y(_13434_),
    .A2(_13432_),
    .A1(_13356_));
 sg13g2_a21o_1 _21120_ (.A2(_13379_),
    .A1(_13376_),
    .B1(_13372_),
    .X(_13435_));
 sg13g2_o21ai_1 _21121_ (.B1(_13435_),
    .Y(_13436_),
    .A1(_13376_),
    .A2(_13379_));
 sg13g2_and2_1 _21122_ (.A(_13352_),
    .B(_13353_),
    .X(_13437_));
 sg13g2_or2_1 _21123_ (.X(_13438_),
    .B(_13353_),
    .A(_13352_));
 sg13g2_o21ai_1 _21124_ (.B1(_13438_),
    .Y(_13439_),
    .A1(_13354_),
    .A2(_13437_));
 sg13g2_buf_1 _21125_ (.A(_13439_),
    .X(_13440_));
 sg13g2_nand2_1 _21126_ (.Y(_13441_),
    .A(net261),
    .B(net277));
 sg13g2_nand2_1 _21127_ (.Y(_13442_),
    .A(net263),
    .B(net292));
 sg13g2_nand2_1 _21128_ (.Y(_13443_),
    .A(net240),
    .B(_12925_));
 sg13g2_xnor2_1 _21129_ (.Y(_13444_),
    .A(_13442_),
    .B(_13443_));
 sg13g2_xnor2_1 _21130_ (.Y(_13445_),
    .A(_13441_),
    .B(_13444_));
 sg13g2_nand2_1 _21131_ (.Y(_13446_),
    .A(_12959_),
    .B(net306));
 sg13g2_nand2_1 _21132_ (.Y(_13447_),
    .A(net301),
    .B(net523));
 sg13g2_nand2_1 _21133_ (.Y(_13448_),
    .A(net264),
    .B(_12813_));
 sg13g2_xor2_1 _21134_ (.B(_13448_),
    .A(_13447_),
    .X(_13449_));
 sg13g2_xnor2_1 _21135_ (.Y(_13450_),
    .A(_13446_),
    .B(_13449_));
 sg13g2_xnor2_1 _21136_ (.Y(_13451_),
    .A(_13445_),
    .B(_13450_));
 sg13g2_xnor2_1 _21137_ (.Y(_13452_),
    .A(_13440_),
    .B(_13451_));
 sg13g2_xor2_1 _21138_ (.B(_13452_),
    .A(_13436_),
    .X(_13453_));
 sg13g2_xnor2_1 _21139_ (.Y(_13454_),
    .A(_13434_),
    .B(_13453_));
 sg13g2_nand2_1 _21140_ (.Y(_13455_),
    .A(_13381_),
    .B(_13395_));
 sg13g2_nand2_1 _21141_ (.Y(_13456_),
    .A(net333),
    .B(_12642_));
 sg13g2_nand2_1 _21142_ (.Y(_13457_),
    .A(net363),
    .B(net518));
 sg13g2_nand2_1 _21143_ (.Y(_13458_),
    .A(net332),
    .B(net519));
 sg13g2_xor2_1 _21144_ (.B(_13458_),
    .A(_13457_),
    .X(_13459_));
 sg13g2_xnor2_1 _21145_ (.Y(_13460_),
    .A(_13456_),
    .B(_13459_));
 sg13g2_a22oi_1 _21146_ (.Y(_13461_),
    .B1(_13388_),
    .B2(_13390_),
    .A2(net479),
    .A1(net404));
 sg13g2_nor2_1 _21147_ (.A(_13388_),
    .B(_13390_),
    .Y(_13462_));
 sg13g2_nor2_1 _21148_ (.A(_13461_),
    .B(_13462_),
    .Y(_13463_));
 sg13g2_a22oi_1 _21149_ (.Y(_13464_),
    .B1(_13366_),
    .B2(_13370_),
    .A2(net518),
    .A1(_13367_));
 sg13g2_nor2_1 _21150_ (.A(_13366_),
    .B(_13370_),
    .Y(_13465_));
 sg13g2_nor2_1 _21151_ (.A(_13464_),
    .B(_13465_),
    .Y(_13466_));
 sg13g2_xnor2_1 _21152_ (.Y(_13467_),
    .A(_13463_),
    .B(_13466_));
 sg13g2_xnor2_1 _21153_ (.Y(_13468_),
    .A(_13460_),
    .B(_13467_));
 sg13g2_a21oi_2 _21154_ (.B1(_13387_),
    .Y(_13469_),
    .A2(_11923_),
    .A1(_11915_));
 sg13g2_nand2_1 _21155_ (.Y(_13470_),
    .A(net404),
    .B(net502));
 sg13g2_nand2_1 _21156_ (.Y(_13471_),
    .A(net405),
    .B(_13098_));
 sg13g2_xnor2_1 _21157_ (.Y(_13472_),
    .A(_13470_),
    .B(_13471_));
 sg13g2_xor2_1 _21158_ (.B(_13472_),
    .A(_13469_),
    .X(_13473_));
 sg13g2_and2_1 _21159_ (.A(_08543_),
    .B(net567),
    .X(_13474_));
 sg13g2_buf_2 _21160_ (.A(_13474_),
    .X(_13475_));
 sg13g2_nand2_1 _21161_ (.Y(_13476_),
    .A(net443),
    .B(_13475_));
 sg13g2_nand2_1 _21162_ (.Y(_13477_),
    .A(net445),
    .B(net480));
 sg13g2_xnor2_1 _21163_ (.Y(_13478_),
    .A(_13476_),
    .B(_13477_));
 sg13g2_xor2_1 _21164_ (.B(_13478_),
    .A(_13473_),
    .X(_13479_));
 sg13g2_nand2b_1 _21165_ (.Y(_13480_),
    .B(_13394_),
    .A_N(_13385_));
 sg13g2_xor2_1 _21166_ (.B(_13480_),
    .A(_13479_),
    .X(_13481_));
 sg13g2_xnor2_1 _21167_ (.Y(_13482_),
    .A(_13468_),
    .B(_13481_));
 sg13g2_xor2_1 _21168_ (.B(_13482_),
    .A(_13455_),
    .X(_13483_));
 sg13g2_xnor2_1 _21169_ (.Y(_13484_),
    .A(_13454_),
    .B(_13483_));
 sg13g2_nor2b_1 _21170_ (.A(_13307_),
    .B_N(_13309_),
    .Y(_13485_));
 sg13g2_nand2b_1 _21171_ (.Y(_13486_),
    .B(_13307_),
    .A_N(_13309_));
 sg13g2_o21ai_1 _21172_ (.B1(_13486_),
    .Y(_13487_),
    .A1(_13302_),
    .A2(_13485_));
 sg13g2_nor2_1 _21173_ (.A(_13303_),
    .B(_13304_),
    .Y(_13488_));
 sg13g2_nor2_1 _21174_ (.A(_13305_),
    .B(_13488_),
    .Y(_13489_));
 sg13g2_a21oi_1 _21175_ (.A1(_13303_),
    .A2(_13304_),
    .Y(_13490_),
    .B1(_13489_));
 sg13g2_nand2_1 _21176_ (.Y(_13491_),
    .A(net238),
    .B(net209));
 sg13g2_nor2_1 _21177_ (.A(_12071_),
    .B(net278),
    .Y(_13492_));
 sg13g2_nand2_1 _21178_ (.Y(_13493_),
    .A(net210),
    .B(_12905_));
 sg13g2_xor2_1 _21179_ (.B(_13493_),
    .A(_13492_),
    .X(_13494_));
 sg13g2_xnor2_1 _21180_ (.Y(_13495_),
    .A(_13491_),
    .B(_13494_));
 sg13g2_a21o_1 _21181_ (.A2(_13344_),
    .A1(_13342_),
    .B1(_13343_),
    .X(_13496_));
 sg13g2_o21ai_1 _21182_ (.B1(_13496_),
    .Y(_13497_),
    .A1(_13342_),
    .A2(_13344_));
 sg13g2_xnor2_1 _21183_ (.Y(_13498_),
    .A(_13495_),
    .B(_13497_));
 sg13g2_xnor2_1 _21184_ (.Y(_13499_),
    .A(_13490_),
    .B(_13498_));
 sg13g2_nand2_1 _21185_ (.Y(_13500_),
    .A(_13313_),
    .B(_13314_));
 sg13g2_nand2_1 _21186_ (.Y(_13501_),
    .A(_13312_),
    .B(_13500_));
 sg13g2_o21ai_1 _21187_ (.B1(_13501_),
    .Y(_13502_),
    .A1(_13313_),
    .A2(_13314_));
 sg13g2_buf_1 _21188_ (.A(_13502_),
    .X(_13503_));
 sg13g2_and2_1 _21189_ (.A(net481),
    .B(_13327_),
    .X(_13504_));
 sg13g2_buf_1 _21190_ (.A(_13504_),
    .X(_13505_));
 sg13g2_inv_1 _21191_ (.Y(_13506_),
    .A(_13041_));
 sg13g2_nand2_1 _21192_ (.Y(_13507_),
    .A(net268),
    .B(_13506_));
 sg13g2_nor2_1 _21193_ (.A(net568),
    .B(net208),
    .Y(_13508_));
 sg13g2_xnor2_1 _21194_ (.Y(_13509_),
    .A(_13507_),
    .B(_13508_));
 sg13g2_xnor2_1 _21195_ (.Y(_13510_),
    .A(_13505_),
    .B(_13509_));
 sg13g2_nor2_1 _21196_ (.A(_13320_),
    .B(_13321_),
    .Y(_13511_));
 sg13g2_xor2_1 _21197_ (.B(_13511_),
    .A(\rbzero.wall_tracer.size_full[9] ),
    .X(_13512_));
 sg13g2_o21ai_1 _21198_ (.B1(_12800_),
    .Y(_13513_),
    .A1(_08421_),
    .A2(_13512_));
 sg13g2_o21ai_1 _21199_ (.B1(_13513_),
    .Y(_13514_),
    .A1(net697),
    .A2(_00469_));
 sg13g2_nor2_1 _21200_ (.A(_12262_),
    .B(_00468_),
    .Y(_13515_));
 sg13g2_a21oi_1 _21201_ (.A1(_12262_),
    .A2(_13514_),
    .Y(_13516_),
    .B1(_13515_));
 sg13g2_buf_1 _21202_ (.A(_13516_),
    .X(_13517_));
 sg13g2_nor2_1 _21203_ (.A(net521),
    .B(_13517_),
    .Y(_13518_));
 sg13g2_xor2_1 _21204_ (.B(_13518_),
    .A(_13510_),
    .X(_13519_));
 sg13g2_xnor2_1 _21205_ (.Y(_13520_),
    .A(_13503_),
    .B(_13519_));
 sg13g2_xnor2_1 _21206_ (.Y(_13521_),
    .A(_13499_),
    .B(_13520_));
 sg13g2_xnor2_1 _21207_ (.Y(_13522_),
    .A(_13487_),
    .B(_13521_));
 sg13g2_inv_1 _21208_ (.Y(_13523_),
    .A(_13311_));
 sg13g2_inv_1 _21209_ (.Y(_13524_),
    .A(_13330_));
 sg13g2_a21oi_1 _21210_ (.A1(_13311_),
    .A2(_13524_),
    .Y(_13525_),
    .B1(_13299_));
 sg13g2_a21oi_1 _21211_ (.A1(_13523_),
    .A2(_13330_),
    .Y(_13526_),
    .B1(_13525_));
 sg13g2_nand2b_1 _21212_ (.Y(_13527_),
    .B(_13362_),
    .A_N(_13358_));
 sg13g2_nor2b_1 _21213_ (.A(_13362_),
    .B_N(_13358_),
    .Y(_13528_));
 sg13g2_a21o_1 _21214_ (.A2(_13527_),
    .A1(_13341_),
    .B1(_13528_),
    .X(_13529_));
 sg13g2_buf_1 _21215_ (.A(_13529_),
    .X(_13530_));
 sg13g2_xor2_1 _21216_ (.B(_13530_),
    .A(_13526_),
    .X(_13531_));
 sg13g2_xnor2_1 _21217_ (.Y(_13532_),
    .A(_13522_),
    .B(_13531_));
 sg13g2_nand2b_1 _21218_ (.Y(_13533_),
    .B(_13364_),
    .A_N(_13396_));
 sg13g2_nor2b_1 _21219_ (.A(_13364_),
    .B_N(_13396_),
    .Y(_13534_));
 sg13g2_a21oi_1 _21220_ (.A1(_13365_),
    .A2(_13533_),
    .Y(_13535_),
    .B1(_13534_));
 sg13g2_xnor2_1 _21221_ (.Y(_13536_),
    .A(_13532_),
    .B(_13535_));
 sg13g2_xnor2_1 _21222_ (.Y(_13537_),
    .A(_13484_),
    .B(_13536_));
 sg13g2_a21o_1 _21223_ (.A2(_13402_),
    .A1(_13398_),
    .B1(_13338_),
    .X(_13538_));
 sg13g2_o21ai_1 _21224_ (.B1(_13538_),
    .Y(_13539_),
    .A1(_13398_),
    .A2(_13402_));
 sg13g2_buf_1 _21225_ (.A(_13539_),
    .X(_13540_));
 sg13g2_nand2_1 _21226_ (.Y(_13541_),
    .A(_13332_),
    .B(_13336_));
 sg13g2_nor2_1 _21227_ (.A(_13332_),
    .B(_13336_),
    .Y(_13542_));
 sg13g2_a21oi_1 _21228_ (.A1(_13296_),
    .A2(_13541_),
    .Y(_13543_),
    .B1(_13542_));
 sg13g2_nor2_1 _21229_ (.A(_13319_),
    .B(_13316_),
    .Y(_13544_));
 sg13g2_nand2_1 _21230_ (.Y(_13545_),
    .A(_13319_),
    .B(_13316_));
 sg13g2_o21ai_1 _21231_ (.B1(_13545_),
    .Y(_13546_),
    .A1(_13328_),
    .A2(_13544_));
 sg13g2_xnor2_1 _21232_ (.Y(_13547_),
    .A(_13543_),
    .B(_13546_));
 sg13g2_xor2_1 _21233_ (.B(_13547_),
    .A(_13540_),
    .X(_13548_));
 sg13g2_xnor2_1 _21234_ (.Y(_13549_),
    .A(_13537_),
    .B(_13548_));
 sg13g2_xnor2_1 _21235_ (.Y(_13550_),
    .A(_13431_),
    .B(_13549_));
 sg13g2_xnor2_1 _21236_ (.Y(_13551_),
    .A(_13430_),
    .B(_13550_));
 sg13g2_a21oi_2 _21237_ (.B1(_13551_),
    .Y(_13552_),
    .A2(_13427_),
    .A1(_13425_));
 sg13g2_and3_1 _21238_ (.X(_13553_),
    .A(_13551_),
    .B(_13425_),
    .C(_13427_));
 sg13g2_nor2_1 _21239_ (.A(_13552_),
    .B(_13553_),
    .Y(_13554_));
 sg13g2_nand2_1 _21240_ (.Y(_13555_),
    .A(_13287_),
    .B(_13419_));
 sg13g2_nor2_1 _21241_ (.A(_13287_),
    .B(_13419_),
    .Y(_13556_));
 sg13g2_a21oi_1 _21242_ (.A1(_13291_),
    .A2(_13555_),
    .Y(_13557_),
    .B1(_13556_));
 sg13g2_xor2_1 _21243_ (.B(_13557_),
    .A(_13554_),
    .X(_13558_));
 sg13g2_buf_2 _21244_ (.A(_13558_),
    .X(_13559_));
 sg13g2_nand2_1 _21245_ (.Y(_13560_),
    .A(net450),
    .B(_13559_));
 sg13g2_buf_1 _21246_ (.A(\rbzero.traced_texVinit[6] ),
    .X(_13561_));
 sg13g2_nand2_1 _21247_ (.Y(_13562_),
    .A(_13561_),
    .B(_11743_));
 sg13g2_a21oi_1 _21248_ (.A1(_13560_),
    .A2(_13562_),
    .Y(_01516_),
    .B1(net572));
 sg13g2_o21ai_1 _21249_ (.B1(_13555_),
    .Y(_13563_),
    .A1(_13291_),
    .A2(_13556_));
 sg13g2_nor2b_1 _21250_ (.A(_13553_),
    .B_N(_13563_),
    .Y(_13564_));
 sg13g2_nor2_2 _21251_ (.A(_13552_),
    .B(_13564_),
    .Y(_13565_));
 sg13g2_nand2_1 _21252_ (.Y(_13566_),
    .A(_13430_),
    .B(_13549_));
 sg13g2_nand2_1 _21253_ (.Y(_13567_),
    .A(_13431_),
    .B(_13566_));
 sg13g2_o21ai_1 _21254_ (.B1(_13567_),
    .Y(_13568_),
    .A1(_13430_),
    .A2(_13549_));
 sg13g2_buf_1 _21255_ (.A(_13568_),
    .X(_13569_));
 sg13g2_nand2_1 _21256_ (.Y(_13570_),
    .A(_13540_),
    .B(_13547_));
 sg13g2_nor2_1 _21257_ (.A(_13540_),
    .B(_13547_),
    .Y(_13571_));
 sg13g2_a21oi_1 _21258_ (.A1(_13537_),
    .A2(_13570_),
    .Y(_13572_),
    .B1(_13571_));
 sg13g2_buf_2 _21259_ (.A(_13572_),
    .X(_13573_));
 sg13g2_nand2b_1 _21260_ (.Y(_13574_),
    .B(_13546_),
    .A_N(_13543_));
 sg13g2_buf_2 _21261_ (.A(_13574_),
    .X(_13575_));
 sg13g2_inv_1 _21262_ (.Y(_13576_),
    .A(_13484_));
 sg13g2_inv_1 _21263_ (.Y(_13577_),
    .A(_13535_));
 sg13g2_a21oi_1 _21264_ (.A1(_13484_),
    .A2(_13577_),
    .Y(_13578_),
    .B1(_13532_));
 sg13g2_a21oi_1 _21265_ (.A1(_13576_),
    .A2(_13535_),
    .Y(_13579_),
    .B1(_13578_));
 sg13g2_nand2_1 _21266_ (.Y(_13580_),
    .A(net240),
    .B(net277));
 sg13g2_nand2_1 _21267_ (.Y(_13581_),
    .A(net263),
    .B(net276));
 sg13g2_nor2b_1 _21268_ (.A(net278),
    .B_N(net261),
    .Y(_13582_));
 sg13g2_xor2_1 _21269_ (.B(_13582_),
    .A(_13581_),
    .X(_13583_));
 sg13g2_xnor2_1 _21270_ (.Y(_13584_),
    .A(_13580_),
    .B(_13583_));
 sg13g2_nand2_1 _21271_ (.Y(_13585_),
    .A(net236),
    .B(net292));
 sg13g2_nand2_1 _21272_ (.Y(_13586_),
    .A(_12813_),
    .B(net523));
 sg13g2_nand2_1 _21273_ (.Y(_13587_),
    .A(_12135_),
    .B(_12209_));
 sg13g2_xor2_1 _21274_ (.B(_13587_),
    .A(_13586_),
    .X(_13588_));
 sg13g2_xnor2_1 _21275_ (.Y(_13589_),
    .A(_13585_),
    .B(_13588_));
 sg13g2_a21o_1 _21276_ (.A2(_13448_),
    .A1(_13446_),
    .B1(_13447_),
    .X(_13590_));
 sg13g2_o21ai_1 _21277_ (.B1(_13590_),
    .Y(_13591_),
    .A1(_13446_),
    .A2(_13448_));
 sg13g2_nor2_1 _21278_ (.A(_13589_),
    .B(_13591_),
    .Y(_13592_));
 sg13g2_nand2_1 _21279_ (.Y(_13593_),
    .A(_13589_),
    .B(_13591_));
 sg13g2_nand2b_1 _21280_ (.Y(_13594_),
    .B(_13593_),
    .A_N(_13592_));
 sg13g2_xnor2_1 _21281_ (.Y(_13595_),
    .A(_13584_),
    .B(_13594_));
 sg13g2_nor2_1 _21282_ (.A(_13440_),
    .B(_13450_),
    .Y(_13596_));
 sg13g2_nand2_1 _21283_ (.Y(_13597_),
    .A(_13440_),
    .B(_13450_));
 sg13g2_o21ai_1 _21284_ (.B1(_13597_),
    .Y(_13598_),
    .A1(_13445_),
    .A2(_13596_));
 sg13g2_a21o_1 _21285_ (.A2(_13466_),
    .A1(_13463_),
    .B1(_13460_),
    .X(_13599_));
 sg13g2_o21ai_1 _21286_ (.B1(_13599_),
    .Y(_13600_),
    .A1(_13463_),
    .A2(_13466_));
 sg13g2_buf_1 _21287_ (.A(_13600_),
    .X(_13601_));
 sg13g2_xnor2_1 _21288_ (.Y(_13602_),
    .A(_13598_),
    .B(_13601_));
 sg13g2_xnor2_1 _21289_ (.Y(_13603_),
    .A(_13595_),
    .B(_13602_));
 sg13g2_nor2_1 _21290_ (.A(_13468_),
    .B(_13479_),
    .Y(_13604_));
 sg13g2_nand2_1 _21291_ (.Y(_13605_),
    .A(_13468_),
    .B(_13479_));
 sg13g2_o21ai_1 _21292_ (.B1(_13605_),
    .Y(_13606_),
    .A1(_13480_),
    .A2(_13604_));
 sg13g2_nand2_1 _21293_ (.Y(_13607_),
    .A(_11794_),
    .B(_12642_));
 sg13g2_nand2_1 _21294_ (.Y(_13608_),
    .A(net332),
    .B(_12841_));
 sg13g2_nand2_1 _21295_ (.Y(_13609_),
    .A(_11837_),
    .B(net519));
 sg13g2_xor2_1 _21296_ (.B(_13609_),
    .A(_13608_),
    .X(_13610_));
 sg13g2_xnor2_1 _21297_ (.Y(_13611_),
    .A(_13607_),
    .B(_13610_));
 sg13g2_nor2b_1 _21298_ (.A(_13469_),
    .B_N(_13470_),
    .Y(_13612_));
 sg13g2_nand3_1 _21299_ (.B(net502),
    .C(_13469_),
    .A(net404),
    .Y(_13613_));
 sg13g2_o21ai_1 _21300_ (.B1(_13613_),
    .Y(_13614_),
    .A1(_13471_),
    .A2(_13612_));
 sg13g2_buf_1 _21301_ (.A(_13614_),
    .X(_13615_));
 sg13g2_a21o_1 _21302_ (.A2(_13458_),
    .A1(_13457_),
    .B1(_13456_),
    .X(_13616_));
 sg13g2_o21ai_1 _21303_ (.B1(_13616_),
    .Y(_13617_),
    .A1(_13457_),
    .A2(_13458_));
 sg13g2_buf_1 _21304_ (.A(_13617_),
    .X(_13618_));
 sg13g2_xnor2_1 _21305_ (.Y(_13619_),
    .A(_13615_),
    .B(_13618_));
 sg13g2_xnor2_1 _21306_ (.Y(_13620_),
    .A(_13611_),
    .B(_13619_));
 sg13g2_nor2_1 _21307_ (.A(_13473_),
    .B(_13478_),
    .Y(_13621_));
 sg13g2_nor2_1 _21308_ (.A(_11913_),
    .B(_13387_),
    .Y(_13622_));
 sg13g2_and2_1 _21309_ (.A(net405),
    .B(net502),
    .X(_13623_));
 sg13g2_buf_1 _21310_ (.A(_13623_),
    .X(_13624_));
 sg13g2_nand2_1 _21311_ (.Y(_13625_),
    .A(net406),
    .B(_13098_));
 sg13g2_xor2_1 _21312_ (.B(_13625_),
    .A(_13624_),
    .X(_13626_));
 sg13g2_xnor2_1 _21313_ (.Y(_13627_),
    .A(_13622_),
    .B(_13626_));
 sg13g2_nand2_2 _21314_ (.Y(_13628_),
    .A(net445),
    .B(_13475_));
 sg13g2_nand3_1 _21315_ (.B(_08481_),
    .C(_00023_),
    .A(_12129_),
    .Y(_13629_));
 sg13g2_buf_1 _21316_ (.A(_13629_),
    .X(_13630_));
 sg13g2_xnor2_1 _21317_ (.Y(_13631_),
    .A(_13628_),
    .B(net566));
 sg13g2_nand2_1 _21318_ (.Y(_13632_),
    .A(_08542_),
    .B(net567));
 sg13g2_buf_2 _21319_ (.A(_13632_),
    .X(_13633_));
 sg13g2_nor2_2 _21320_ (.A(_12398_),
    .B(_13633_),
    .Y(_13634_));
 sg13g2_nand2_1 _21321_ (.Y(_13635_),
    .A(_13631_),
    .B(_13634_));
 sg13g2_and2_1 _21322_ (.A(net445),
    .B(_13475_),
    .X(_13636_));
 sg13g2_buf_1 _21323_ (.A(_13636_),
    .X(_13637_));
 sg13g2_nand3_1 _21324_ (.B(_13637_),
    .C(net566),
    .A(_13633_),
    .Y(_13638_));
 sg13g2_nor3_1 _21325_ (.A(_13383_),
    .B(_13637_),
    .C(net566),
    .Y(_13639_));
 sg13g2_nor2_1 _21326_ (.A(net404),
    .B(_13631_),
    .Y(_13640_));
 sg13g2_o21ai_1 _21327_ (.B1(_12144_),
    .Y(_13641_),
    .A1(_13639_),
    .A2(_13640_));
 sg13g2_nor2_1 _21328_ (.A(_13383_),
    .B(_13628_),
    .Y(_13642_));
 sg13g2_o21ai_1 _21329_ (.B1(net443),
    .Y(_13643_),
    .A1(_13634_),
    .A2(_13642_));
 sg13g2_nand4_1 _21330_ (.B(_13638_),
    .C(_13641_),
    .A(_13635_),
    .Y(_13644_),
    .D(_13643_));
 sg13g2_xor2_1 _21331_ (.B(_13644_),
    .A(_13627_),
    .X(_13645_));
 sg13g2_xnor2_1 _21332_ (.Y(_13646_),
    .A(_13621_),
    .B(_13645_));
 sg13g2_xnor2_1 _21333_ (.Y(_13647_),
    .A(_13620_),
    .B(_13646_));
 sg13g2_and2_1 _21334_ (.A(_13606_),
    .B(_13647_),
    .X(_13648_));
 sg13g2_nor2_1 _21335_ (.A(_13606_),
    .B(_13647_),
    .Y(_13649_));
 sg13g2_nor2_1 _21336_ (.A(_13648_),
    .B(_13649_),
    .Y(_13650_));
 sg13g2_xnor2_1 _21337_ (.Y(_13651_),
    .A(_13603_),
    .B(_13650_));
 sg13g2_a21oi_1 _21338_ (.A1(_13434_),
    .A2(_13452_),
    .Y(_13652_),
    .B1(_13436_));
 sg13g2_inv_1 _21339_ (.Y(_13653_),
    .A(_13652_));
 sg13g2_o21ai_1 _21340_ (.B1(_13653_),
    .Y(_13654_),
    .A1(_13434_),
    .A2(_13452_));
 sg13g2_nand2b_1 _21341_ (.Y(_13655_),
    .B(_13495_),
    .A_N(_13497_));
 sg13g2_nor2b_1 _21342_ (.A(_13495_),
    .B_N(_13497_),
    .Y(_13656_));
 sg13g2_a21o_1 _21343_ (.A2(_13655_),
    .A1(_13490_),
    .B1(_13656_),
    .X(_13657_));
 sg13g2_buf_1 _21344_ (.A(_13657_),
    .X(_13658_));
 sg13g2_nand2_1 _21345_ (.Y(_13659_),
    .A(_13505_),
    .B(_13508_));
 sg13g2_nand2_1 _21346_ (.Y(_13660_),
    .A(_13507_),
    .B(_13659_));
 sg13g2_o21ai_1 _21347_ (.B1(_13660_),
    .Y(_13661_),
    .A1(_13505_),
    .A2(_13508_));
 sg13g2_buf_1 _21348_ (.A(_13661_),
    .X(_13662_));
 sg13g2_nor2_2 _21349_ (.A(net504),
    .B(_13517_),
    .Y(_13663_));
 sg13g2_inv_1 _21350_ (.Y(_13664_),
    .A(_13190_));
 sg13g2_nand2_1 _21351_ (.Y(_13665_),
    .A(_11781_),
    .B(_13664_));
 sg13g2_nand2_1 _21352_ (.Y(_13666_),
    .A(net520),
    .B(_13327_));
 sg13g2_xnor2_1 _21353_ (.Y(_13667_),
    .A(_13665_),
    .B(_13666_));
 sg13g2_xnor2_1 _21354_ (.Y(_13668_),
    .A(_13663_),
    .B(_13667_));
 sg13g2_inv_1 _21355_ (.Y(_13669_),
    .A(_00471_));
 sg13g2_nor4_1 _21356_ (.A(_13033_),
    .B(_13182_),
    .C(_13320_),
    .D(\rbzero.wall_tracer.size_full[9] ),
    .Y(_13670_));
 sg13g2_nand2_1 _21357_ (.Y(_13671_),
    .A(_13035_),
    .B(_13670_));
 sg13g2_xor2_1 _21358_ (.B(_13671_),
    .A(\rbzero.wall_tracer.size_full[10] ),
    .X(_13672_));
 sg13g2_nand2b_1 _21359_ (.Y(_13673_),
    .B(_13672_),
    .A_N(_08421_));
 sg13g2_a221oi_1 _21360_ (.B2(_13673_),
    .C1(net611),
    .B1(_12800_),
    .A1(_08442_),
    .Y(_13674_),
    .A2(_13669_));
 sg13g2_a21o_1 _21361_ (.A2(_00470_),
    .A1(_08447_),
    .B1(_13674_),
    .X(_13675_));
 sg13g2_buf_1 _21362_ (.A(_13675_),
    .X(_13676_));
 sg13g2_nor2_1 _21363_ (.A(net521),
    .B(_13676_),
    .Y(_13677_));
 sg13g2_xnor2_1 _21364_ (.Y(_13678_),
    .A(_13668_),
    .B(_13677_));
 sg13g2_xnor2_1 _21365_ (.Y(_13679_),
    .A(_13662_),
    .B(_13678_));
 sg13g2_nor2_1 _21366_ (.A(_12226_),
    .B(_13041_),
    .Y(_13680_));
 sg13g2_nand2_1 _21367_ (.Y(_13681_),
    .A(_12456_),
    .B(net211));
 sg13g2_nand2_1 _21368_ (.Y(_13682_),
    .A(net210),
    .B(_13174_));
 sg13g2_xnor2_1 _21369_ (.Y(_13683_),
    .A(_13681_),
    .B(_13682_));
 sg13g2_xnor2_1 _21370_ (.Y(_13684_),
    .A(_13680_),
    .B(_13683_));
 sg13g2_nand3_1 _21371_ (.B(net209),
    .C(_13492_),
    .A(net238),
    .Y(_13685_));
 sg13g2_a21oi_1 _21372_ (.A1(_12391_),
    .A2(net209),
    .Y(_13686_),
    .B1(_13492_));
 sg13g2_a21oi_2 _21373_ (.B1(_13686_),
    .Y(_13687_),
    .A2(_13685_),
    .A1(_13493_));
 sg13g2_a21o_1 _21374_ (.A2(_13443_),
    .A1(_13441_),
    .B1(_13442_),
    .X(_13688_));
 sg13g2_o21ai_1 _21375_ (.B1(_13688_),
    .Y(_13689_),
    .A1(_13441_),
    .A2(_13443_));
 sg13g2_buf_1 _21376_ (.A(_13689_),
    .X(_13690_));
 sg13g2_xor2_1 _21377_ (.B(_13690_),
    .A(_13687_),
    .X(_13691_));
 sg13g2_xnor2_1 _21378_ (.Y(_13692_),
    .A(_13684_),
    .B(_13691_));
 sg13g2_xnor2_1 _21379_ (.Y(_13693_),
    .A(_13679_),
    .B(_13692_));
 sg13g2_xnor2_1 _21380_ (.Y(_13694_),
    .A(_13658_),
    .B(_13693_));
 sg13g2_inv_1 _21381_ (.Y(_13695_),
    .A(_13694_));
 sg13g2_a21oi_1 _21382_ (.A1(_13499_),
    .A2(_13520_),
    .Y(_13696_),
    .B1(_13487_));
 sg13g2_nor2_1 _21383_ (.A(_13499_),
    .B(_13520_),
    .Y(_13697_));
 sg13g2_nor2_1 _21384_ (.A(_13696_),
    .B(_13697_),
    .Y(_13698_));
 sg13g2_nor2_1 _21385_ (.A(_13695_),
    .B(_13698_),
    .Y(_13699_));
 sg13g2_nand2_1 _21386_ (.Y(_13700_),
    .A(_13695_),
    .B(_13698_));
 sg13g2_nand2b_1 _21387_ (.Y(_13701_),
    .B(_13700_),
    .A_N(_13699_));
 sg13g2_xnor2_1 _21388_ (.Y(_13702_),
    .A(_13654_),
    .B(_13701_));
 sg13g2_nand2_1 _21389_ (.Y(_13703_),
    .A(_13454_),
    .B(_13482_));
 sg13g2_nand2_1 _21390_ (.Y(_13704_),
    .A(_13455_),
    .B(_13703_));
 sg13g2_o21ai_1 _21391_ (.B1(_13704_),
    .Y(_13705_),
    .A1(_13454_),
    .A2(_13482_));
 sg13g2_buf_1 _21392_ (.A(_13705_),
    .X(_13706_));
 sg13g2_xnor2_1 _21393_ (.Y(_13707_),
    .A(_13702_),
    .B(_13706_));
 sg13g2_xnor2_1 _21394_ (.Y(_13708_),
    .A(_13651_),
    .B(_13707_));
 sg13g2_o21ai_1 _21395_ (.B1(_13526_),
    .Y(_13709_),
    .A1(_13522_),
    .A2(_13530_));
 sg13g2_nand2_1 _21396_ (.Y(_13710_),
    .A(_13522_),
    .B(_13530_));
 sg13g2_nand2_1 _21397_ (.Y(_13711_),
    .A(_13709_),
    .B(_13710_));
 sg13g2_buf_1 _21398_ (.A(net566),
    .X(_13712_));
 sg13g2_nor2_1 _21399_ (.A(_13503_),
    .B(_13510_),
    .Y(_13713_));
 sg13g2_nand2_1 _21400_ (.Y(_13714_),
    .A(_13503_),
    .B(_13510_));
 sg13g2_o21ai_1 _21401_ (.B1(_13714_),
    .Y(_13715_),
    .A1(_13518_),
    .A2(_13713_));
 sg13g2_buf_1 _21402_ (.A(_13715_),
    .X(_13716_));
 sg13g2_xnor2_1 _21403_ (.Y(_13717_),
    .A(net517),
    .B(_13716_));
 sg13g2_xnor2_1 _21404_ (.Y(_13718_),
    .A(_13711_),
    .B(_13717_));
 sg13g2_xnor2_1 _21405_ (.Y(_13719_),
    .A(_13708_),
    .B(_13718_));
 sg13g2_xnor2_1 _21406_ (.Y(_13720_),
    .A(_13579_),
    .B(_13719_));
 sg13g2_xnor2_1 _21407_ (.Y(_13721_),
    .A(_13575_),
    .B(_13720_));
 sg13g2_xnor2_1 _21408_ (.Y(_13722_),
    .A(_13573_),
    .B(_13721_));
 sg13g2_xnor2_1 _21409_ (.Y(_13723_),
    .A(_13569_),
    .B(_13722_));
 sg13g2_xnor2_1 _21410_ (.Y(_13724_),
    .A(_13565_),
    .B(_13723_));
 sg13g2_nand2_1 _21411_ (.Y(_13725_),
    .A(net450),
    .B(_13724_));
 sg13g2_buf_1 _21412_ (.A(\rbzero.traced_texVinit[7] ),
    .X(_13726_));
 sg13g2_nand2_1 _21413_ (.Y(_13727_),
    .A(_13726_),
    .B(_11743_));
 sg13g2_a21oi_1 _21414_ (.A1(_13725_),
    .A2(_13727_),
    .Y(_01517_),
    .B1(net572));
 sg13g2_inv_1 _21415_ (.Y(_13728_),
    .A(_13708_));
 sg13g2_inv_1 _21416_ (.Y(_13729_),
    .A(_13718_));
 sg13g2_a21oi_1 _21417_ (.A1(_13708_),
    .A2(_13729_),
    .Y(_13730_),
    .B1(_13579_));
 sg13g2_a21oi_2 _21418_ (.B1(_13730_),
    .Y(_13731_),
    .A2(_13718_),
    .A1(_13728_));
 sg13g2_a21o_1 _21419_ (.A2(_13716_),
    .A1(_13711_),
    .B1(net517),
    .X(_13732_));
 sg13g2_o21ai_1 _21420_ (.B1(_13732_),
    .Y(_13733_),
    .A1(_13711_),
    .A2(_13716_));
 sg13g2_nand2_1 _21421_ (.Y(_13734_),
    .A(_13651_),
    .B(_13706_));
 sg13g2_nor2_1 _21422_ (.A(_13651_),
    .B(_13706_),
    .Y(_13735_));
 sg13g2_a21oi_1 _21423_ (.A1(_13702_),
    .A2(_13734_),
    .Y(_13736_),
    .B1(_13735_));
 sg13g2_inv_1 _21424_ (.Y(_13737_),
    .A(_13692_));
 sg13g2_inv_1 _21425_ (.Y(_13738_),
    .A(_13658_));
 sg13g2_a21oi_1 _21426_ (.A1(_13738_),
    .A2(_13692_),
    .Y(_13739_),
    .B1(_13679_));
 sg13g2_a21oi_1 _21427_ (.A1(_13658_),
    .A2(_13737_),
    .Y(_13740_),
    .B1(_13739_));
 sg13g2_a21o_1 _21428_ (.A2(_13690_),
    .A1(_13687_),
    .B1(_13684_),
    .X(_13741_));
 sg13g2_o21ai_1 _21429_ (.B1(_13741_),
    .Y(_13742_),
    .A1(_13687_),
    .A2(_13690_));
 sg13g2_nand3_1 _21430_ (.B(_13327_),
    .C(_13663_),
    .A(net520),
    .Y(_13743_));
 sg13g2_nor2b_1 _21431_ (.A(_13663_),
    .B_N(_13666_),
    .Y(_13744_));
 sg13g2_a21o_1 _21432_ (.A2(_13743_),
    .A1(_13665_),
    .B1(_13744_),
    .X(_13745_));
 sg13g2_buf_1 _21433_ (.A(_13745_),
    .X(_13746_));
 sg13g2_nor2_1 _21434_ (.A(net568),
    .B(_13517_),
    .Y(_13747_));
 sg13g2_buf_1 _21435_ (.A(net268),
    .X(_13748_));
 sg13g2_nand2_1 _21436_ (.Y(_13749_),
    .A(_13748_),
    .B(_13327_));
 sg13g2_xnor2_1 _21437_ (.Y(_13750_),
    .A(_13747_),
    .B(_13749_));
 sg13g2_a21oi_1 _21438_ (.A1(_08447_),
    .A2(_00470_),
    .Y(_13751_),
    .B1(_13674_));
 sg13g2_xnor2_1 _21439_ (.Y(_13752_),
    .A(net504),
    .B(net505));
 sg13g2_nand2_1 _21440_ (.Y(_13753_),
    .A(_13751_),
    .B(_13752_));
 sg13g2_xnor2_1 _21441_ (.Y(_13754_),
    .A(_13750_),
    .B(_13753_));
 sg13g2_xnor2_1 _21442_ (.Y(_13755_),
    .A(_13746_),
    .B(_13754_));
 sg13g2_nand2_1 _21443_ (.Y(_13756_),
    .A(net237),
    .B(net209));
 sg13g2_nor2_1 _21444_ (.A(_12226_),
    .B(_13191_),
    .Y(_13757_));
 sg13g2_buf_1 _21445_ (.A(_13041_),
    .X(_13758_));
 sg13g2_nor2_1 _21446_ (.A(net262),
    .B(net207),
    .Y(_13759_));
 sg13g2_xor2_1 _21447_ (.B(_13759_),
    .A(_13757_),
    .X(_13760_));
 sg13g2_xnor2_1 _21448_ (.Y(_13761_),
    .A(_13756_),
    .B(_13760_));
 sg13g2_nand2_1 _21449_ (.Y(_13762_),
    .A(_13681_),
    .B(_13682_));
 sg13g2_nand2_1 _21450_ (.Y(_13763_),
    .A(_13680_),
    .B(_13762_));
 sg13g2_o21ai_1 _21451_ (.B1(_13763_),
    .Y(_13764_),
    .A1(_13681_),
    .A2(_13682_));
 sg13g2_buf_1 _21452_ (.A(_13764_),
    .X(_13765_));
 sg13g2_nor2_1 _21453_ (.A(_13581_),
    .B(_13580_),
    .Y(_13766_));
 sg13g2_nor2_1 _21454_ (.A(_13582_),
    .B(_13766_),
    .Y(_13767_));
 sg13g2_a21oi_2 _21455_ (.B1(_13767_),
    .Y(_13768_),
    .A2(_13580_),
    .A1(_13581_));
 sg13g2_xnor2_1 _21456_ (.Y(_13769_),
    .A(_13765_),
    .B(_13768_));
 sg13g2_xnor2_1 _21457_ (.Y(_13770_),
    .A(_13761_),
    .B(_13769_));
 sg13g2_nor2_1 _21458_ (.A(_13755_),
    .B(_13770_),
    .Y(_13771_));
 sg13g2_nand2_1 _21459_ (.Y(_13772_),
    .A(_13755_),
    .B(_13770_));
 sg13g2_nand2b_1 _21460_ (.Y(_13773_),
    .B(_13772_),
    .A_N(_13771_));
 sg13g2_xnor2_1 _21461_ (.Y(_13774_),
    .A(_13742_),
    .B(_13773_));
 sg13g2_nor2_1 _21462_ (.A(_13595_),
    .B(_13601_),
    .Y(_13775_));
 sg13g2_nand2_1 _21463_ (.Y(_13776_),
    .A(_13595_),
    .B(_13601_));
 sg13g2_o21ai_1 _21464_ (.B1(_13776_),
    .Y(_13777_),
    .A1(_13598_),
    .A2(_13775_));
 sg13g2_buf_1 _21465_ (.A(_13777_),
    .X(_13778_));
 sg13g2_xor2_1 _21466_ (.B(_13778_),
    .A(_13774_),
    .X(_13779_));
 sg13g2_xnor2_1 _21467_ (.Y(_13780_),
    .A(_13740_),
    .B(_13779_));
 sg13g2_nand2_1 _21468_ (.Y(_13781_),
    .A(_12452_),
    .B(_12905_));
 sg13g2_and2_1 _21469_ (.A(_12337_),
    .B(net277),
    .X(_13782_));
 sg13g2_buf_1 _21470_ (.A(_13782_),
    .X(_13783_));
 sg13g2_nor2b_1 _21471_ (.A(net258),
    .B_N(net240),
    .Y(_13784_));
 sg13g2_xnor2_1 _21472_ (.Y(_13785_),
    .A(_13783_),
    .B(_13784_));
 sg13g2_xnor2_1 _21473_ (.Y(_13786_),
    .A(_13781_),
    .B(_13785_));
 sg13g2_nand2_1 _21474_ (.Y(_13787_),
    .A(net236),
    .B(net276));
 sg13g2_buf_1 _21475_ (.A(_12209_),
    .X(_13788_));
 sg13g2_buf_1 _21476_ (.A(net523),
    .X(_13789_));
 sg13g2_and2_1 _21477_ (.A(net300),
    .B(net500),
    .X(_13790_));
 sg13g2_buf_1 _21478_ (.A(net264),
    .X(_13791_));
 sg13g2_nand2_1 _21479_ (.Y(_13792_),
    .A(net234),
    .B(net292));
 sg13g2_xnor2_1 _21480_ (.Y(_13793_),
    .A(_13790_),
    .B(_13792_));
 sg13g2_xnor2_1 _21481_ (.Y(_13794_),
    .A(_13787_),
    .B(_13793_));
 sg13g2_and2_1 _21482_ (.A(_13585_),
    .B(_13586_),
    .X(_13795_));
 sg13g2_or2_1 _21483_ (.X(_13796_),
    .B(_13586_),
    .A(_13585_));
 sg13g2_o21ai_1 _21484_ (.B1(_13796_),
    .Y(_13797_),
    .A1(_13587_),
    .A2(_13795_));
 sg13g2_buf_1 _21485_ (.A(_13797_),
    .X(_13798_));
 sg13g2_xnor2_1 _21486_ (.Y(_13799_),
    .A(_13794_),
    .B(_13798_));
 sg13g2_xnor2_1 _21487_ (.Y(_13800_),
    .A(_13786_),
    .B(_13799_));
 sg13g2_o21ai_1 _21488_ (.B1(_13593_),
    .Y(_13801_),
    .A1(_13584_),
    .A2(_13592_));
 sg13g2_a21o_1 _21489_ (.A2(_13618_),
    .A1(_13615_),
    .B1(_13611_),
    .X(_13802_));
 sg13g2_o21ai_1 _21490_ (.B1(_13802_),
    .Y(_13803_),
    .A1(_13615_),
    .A2(_13618_));
 sg13g2_buf_1 _21491_ (.A(_13803_),
    .X(_13804_));
 sg13g2_xnor2_1 _21492_ (.Y(_13805_),
    .A(_13801_),
    .B(_13804_));
 sg13g2_xnor2_1 _21493_ (.Y(_13806_),
    .A(_13800_),
    .B(_13805_));
 sg13g2_buf_1 _21494_ (.A(_12642_),
    .X(_13807_));
 sg13g2_nand2_1 _21495_ (.Y(_13808_),
    .A(net293),
    .B(_13807_));
 sg13g2_nand2_1 _21496_ (.Y(_13809_),
    .A(net319),
    .B(net518));
 sg13g2_nand2_1 _21497_ (.Y(_13810_),
    .A(net301),
    .B(net519));
 sg13g2_xor2_1 _21498_ (.B(_13810_),
    .A(_13809_),
    .X(_13811_));
 sg13g2_xnor2_1 _21499_ (.Y(_13812_),
    .A(_13808_),
    .B(_13811_));
 sg13g2_and2_1 _21500_ (.A(_13608_),
    .B(_13609_),
    .X(_13813_));
 sg13g2_or2_1 _21501_ (.X(_13814_),
    .B(_13609_),
    .A(_13608_));
 sg13g2_o21ai_1 _21502_ (.B1(_13814_),
    .Y(_13815_),
    .A1(_13607_),
    .A2(_13813_));
 sg13g2_buf_1 _21503_ (.A(_13815_),
    .X(_13816_));
 sg13g2_a22oi_1 _21504_ (.Y(_13817_),
    .B1(_13622_),
    .B2(_13624_),
    .A2(net479),
    .A1(net362));
 sg13g2_nor2_1 _21505_ (.A(_13622_),
    .B(_13624_),
    .Y(_13818_));
 sg13g2_nor2_1 _21506_ (.A(_13817_),
    .B(_13818_),
    .Y(_13819_));
 sg13g2_xnor2_1 _21507_ (.Y(_13820_),
    .A(_13816_),
    .B(_13819_));
 sg13g2_xnor2_1 _21508_ (.Y(_13821_),
    .A(_13812_),
    .B(_13820_));
 sg13g2_nor2_1 _21509_ (.A(_12069_),
    .B(_13387_),
    .Y(_13822_));
 sg13g2_nand2_1 _21510_ (.Y(_13823_),
    .A(net406),
    .B(net502));
 sg13g2_and2_1 _21511_ (.A(net363),
    .B(_13098_),
    .X(_13824_));
 sg13g2_buf_1 _21512_ (.A(_13824_),
    .X(_13825_));
 sg13g2_xor2_1 _21513_ (.B(_13825_),
    .A(_13823_),
    .X(_13826_));
 sg13g2_xnor2_1 _21514_ (.Y(_13827_),
    .A(_13822_),
    .B(_13826_));
 sg13g2_a21oi_2 _21515_ (.B1(_13633_),
    .Y(_13828_),
    .A2(_11956_),
    .A1(_11949_));
 sg13g2_nor2_1 _21516_ (.A(net445),
    .B(_13630_),
    .Y(_13829_));
 sg13g2_nand2_1 _21517_ (.Y(_13830_),
    .A(_12166_),
    .B(_13475_));
 sg13g2_xor2_1 _21518_ (.B(_13830_),
    .A(_13829_),
    .X(_13831_));
 sg13g2_xnor2_1 _21519_ (.Y(_13832_),
    .A(_13828_),
    .B(_13831_));
 sg13g2_nand2b_1 _21520_ (.Y(_13833_),
    .B(_12144_),
    .A_N(net566));
 sg13g2_nand2_1 _21521_ (.Y(_13834_),
    .A(_13628_),
    .B(_13833_));
 sg13g2_nor2_1 _21522_ (.A(_13628_),
    .B(_13833_),
    .Y(_13835_));
 sg13g2_a21oi_1 _21523_ (.A1(_13634_),
    .A2(_13834_),
    .Y(_13836_),
    .B1(_13835_));
 sg13g2_xnor2_1 _21524_ (.Y(_13837_),
    .A(_13832_),
    .B(_13836_));
 sg13g2_xnor2_1 _21525_ (.Y(_13838_),
    .A(_13827_),
    .B(_13837_));
 sg13g2_nand2_1 _21526_ (.Y(_13839_),
    .A(_13637_),
    .B(net566));
 sg13g2_o21ai_1 _21527_ (.B1(_13839_),
    .Y(_13840_),
    .A1(_13637_),
    .A2(_13833_));
 sg13g2_nand2b_1 _21528_ (.Y(_13841_),
    .B(_13840_),
    .A_N(_13634_));
 sg13g2_o21ai_1 _21529_ (.B1(net443),
    .Y(_13842_),
    .A1(_13637_),
    .A2(_13634_));
 sg13g2_nand3_1 _21530_ (.B(_13841_),
    .C(_13842_),
    .A(_13635_),
    .Y(_13843_));
 sg13g2_nor3_1 _21531_ (.A(net404),
    .B(_13385_),
    .C(_13628_),
    .Y(_13844_));
 sg13g2_a21oi_2 _21532_ (.B1(_13844_),
    .Y(_13845_),
    .A2(_13843_),
    .A1(_13627_));
 sg13g2_xor2_1 _21533_ (.B(_13845_),
    .A(_13838_),
    .X(_13846_));
 sg13g2_xnor2_1 _21534_ (.Y(_13847_),
    .A(_13821_),
    .B(_13846_));
 sg13g2_nand2_1 _21535_ (.Y(_13848_),
    .A(_13620_),
    .B(_13645_));
 sg13g2_o21ai_1 _21536_ (.B1(_13621_),
    .Y(_13849_),
    .A1(_13620_),
    .A2(_13645_));
 sg13g2_and3_1 _21537_ (.X(_13850_),
    .A(_13847_),
    .B(_13848_),
    .C(_13849_));
 sg13g2_a21oi_1 _21538_ (.A1(_13848_),
    .A2(_13849_),
    .Y(_13851_),
    .B1(_13847_));
 sg13g2_nor2_1 _21539_ (.A(_13850_),
    .B(_13851_),
    .Y(_13852_));
 sg13g2_xnor2_1 _21540_ (.Y(_13853_),
    .A(_13806_),
    .B(_13852_));
 sg13g2_inv_1 _21541_ (.Y(_13854_),
    .A(_13649_));
 sg13g2_o21ai_1 _21542_ (.B1(_13854_),
    .Y(_13855_),
    .A1(_13603_),
    .A2(_13648_));
 sg13g2_nor2_1 _21543_ (.A(_13853_),
    .B(_13855_),
    .Y(_13856_));
 sg13g2_nand2_1 _21544_ (.Y(_13857_),
    .A(_13853_),
    .B(_13855_));
 sg13g2_nand2b_1 _21545_ (.Y(_13858_),
    .B(_13857_),
    .A_N(_13856_));
 sg13g2_xnor2_1 _21546_ (.Y(_13859_),
    .A(_13780_),
    .B(_13858_));
 sg13g2_o21ai_1 _21547_ (.B1(_13700_),
    .Y(_13860_),
    .A1(_13654_),
    .A2(_13699_));
 sg13g2_nor2b_1 _21548_ (.A(_13662_),
    .B_N(_13668_),
    .Y(_13861_));
 sg13g2_nand2b_1 _21549_ (.Y(_13862_),
    .B(_13662_),
    .A_N(_13668_));
 sg13g2_o21ai_1 _21550_ (.B1(_13862_),
    .Y(_13863_),
    .A1(_13677_),
    .A2(_13861_));
 sg13g2_xor2_1 _21551_ (.B(_13863_),
    .A(_13860_),
    .X(_13864_));
 sg13g2_xor2_1 _21552_ (.B(_13864_),
    .A(_13859_),
    .X(_13865_));
 sg13g2_xnor2_1 _21553_ (.Y(_13866_),
    .A(_13736_),
    .B(_13865_));
 sg13g2_xor2_1 _21554_ (.B(_13866_),
    .A(_13733_),
    .X(_13867_));
 sg13g2_xnor2_1 _21555_ (.Y(_13868_),
    .A(_13731_),
    .B(_13867_));
 sg13g2_nor2_1 _21556_ (.A(_13569_),
    .B(_13720_),
    .Y(_13869_));
 sg13g2_nand2_1 _21557_ (.Y(_13870_),
    .A(_13573_),
    .B(_13869_));
 sg13g2_nand2_1 _21558_ (.Y(_13871_),
    .A(_13569_),
    .B(_13720_));
 sg13g2_or2_1 _21559_ (.X(_13872_),
    .B(_13871_),
    .A(_13573_));
 sg13g2_mux2_1 _21560_ (.A0(_13870_),
    .A1(_13872_),
    .S(_13565_),
    .X(_13873_));
 sg13g2_nand2b_1 _21561_ (.Y(_13874_),
    .B(_13575_),
    .A_N(_13872_));
 sg13g2_o21ai_1 _21562_ (.B1(_13871_),
    .Y(_13875_),
    .A1(_13573_),
    .A2(_13869_));
 sg13g2_nand3_1 _21563_ (.B(_13575_),
    .C(_13875_),
    .A(_13565_),
    .Y(_13876_));
 sg13g2_o21ai_1 _21564_ (.B1(_13870_),
    .Y(_13877_),
    .A1(_13565_),
    .A2(_13875_));
 sg13g2_nand2b_1 _21565_ (.Y(_13878_),
    .B(_13877_),
    .A_N(_13575_));
 sg13g2_nand4_1 _21566_ (.B(_13874_),
    .C(_13876_),
    .A(_13873_),
    .Y(_13879_),
    .D(_13878_));
 sg13g2_xor2_1 _21567_ (.B(_13879_),
    .A(_13868_),
    .X(_13880_));
 sg13g2_nand2_1 _21568_ (.Y(_13881_),
    .A(net450),
    .B(_13880_));
 sg13g2_buf_1 _21569_ (.A(\rbzero.traced_texVinit[8] ),
    .X(_13882_));
 sg13g2_buf_1 _21570_ (.A(net464),
    .X(_13883_));
 sg13g2_nand2_1 _21571_ (.Y(_13884_),
    .A(_13882_),
    .B(net442));
 sg13g2_a21oi_1 _21572_ (.A1(_13881_),
    .A2(_13884_),
    .Y(_01518_),
    .B1(net572));
 sg13g2_or2_1 _21573_ (.X(_13885_),
    .B(_13720_),
    .A(_13569_));
 sg13g2_inv_1 _21574_ (.Y(_13886_),
    .A(_13871_));
 sg13g2_a21oi_1 _21575_ (.A1(_13575_),
    .A2(_13885_),
    .Y(_13887_),
    .B1(_13886_));
 sg13g2_nand2b_1 _21576_ (.Y(_13888_),
    .B(_13871_),
    .A_N(_13868_));
 sg13g2_a22oi_1 _21577_ (.Y(_13889_),
    .B1(_13888_),
    .B2(_13575_),
    .A2(_13885_),
    .A1(_13868_));
 sg13g2_o21ai_1 _21578_ (.B1(_13889_),
    .Y(_13890_),
    .A1(_13573_),
    .A2(_13887_));
 sg13g2_nand2b_1 _21579_ (.Y(_13891_),
    .B(_13890_),
    .A_N(_13552_));
 sg13g2_or2_1 _21580_ (.X(_13892_),
    .B(_13889_),
    .A(_13573_));
 sg13g2_o21ai_1 _21581_ (.B1(_13892_),
    .Y(_13893_),
    .A1(_13564_),
    .A2(_13891_));
 sg13g2_inv_1 _21582_ (.Y(_13894_),
    .A(_13887_));
 sg13g2_nor3_1 _21583_ (.A(_13552_),
    .B(_13564_),
    .C(_13573_),
    .Y(_13895_));
 sg13g2_o21ai_1 _21584_ (.B1(_13868_),
    .Y(_13896_),
    .A1(_13894_),
    .A2(_13895_));
 sg13g2_nor2b_1 _21585_ (.A(_13893_),
    .B_N(_13896_),
    .Y(_13897_));
 sg13g2_nand2_1 _21586_ (.Y(_13898_),
    .A(_13859_),
    .B(_13864_));
 sg13g2_nor2_1 _21587_ (.A(_13859_),
    .B(_13864_),
    .Y(_13899_));
 sg13g2_a21oi_1 _21588_ (.A1(_13736_),
    .A2(_13898_),
    .Y(_13900_),
    .B1(_13899_));
 sg13g2_nor2_1 _21589_ (.A(_13860_),
    .B(_13863_),
    .Y(_13901_));
 sg13g2_a21oi_1 _21590_ (.A1(_13780_),
    .A2(_13857_),
    .Y(_13902_),
    .B1(_13856_));
 sg13g2_buf_1 _21591_ (.A(_13327_),
    .X(_13903_));
 sg13g2_buf_1 _21592_ (.A(_13517_),
    .X(_13904_));
 sg13g2_nor2_1 _21593_ (.A(net481),
    .B(net206),
    .Y(_13905_));
 sg13g2_nand2_1 _21594_ (.Y(_13906_),
    .A(_13751_),
    .B(_13905_));
 sg13g2_nand3_1 _21595_ (.B(net174),
    .C(net206),
    .A(net481),
    .Y(_13907_));
 sg13g2_o21ai_1 _21596_ (.B1(_13907_),
    .Y(_13908_),
    .A1(net174),
    .A2(_13906_));
 sg13g2_a22oi_1 _21597_ (.Y(_13909_),
    .B1(_13908_),
    .B2(net235),
    .A2(_13676_),
    .A1(net174));
 sg13g2_buf_1 _21598_ (.A(_13751_),
    .X(_13910_));
 sg13g2_nand3_1 _21599_ (.B(_13505_),
    .C(net257),
    .A(net235),
    .Y(_13911_));
 sg13g2_inv_1 _21600_ (.Y(_13912_),
    .A(_13904_));
 sg13g2_buf_1 _21601_ (.A(_13912_),
    .X(_13913_));
 sg13g2_a22oi_1 _21602_ (.Y(_13914_),
    .B1(net257),
    .B2(net520),
    .A2(net150),
    .A1(net235));
 sg13g2_and2_1 _21603_ (.A(net568),
    .B(_13327_),
    .X(_13915_));
 sg13g2_a21o_1 _21604_ (.A2(_13915_),
    .A1(net257),
    .B1(_12420_),
    .X(_13916_));
 sg13g2_a22oi_1 _21605_ (.Y(_13917_),
    .B1(_13916_),
    .B2(_13663_),
    .A2(_13914_),
    .A1(_13911_));
 sg13g2_o21ai_1 _21606_ (.B1(_13917_),
    .Y(_13918_),
    .A1(net568),
    .A2(_13909_));
 sg13g2_xor2_1 _21607_ (.B(_13918_),
    .A(_13753_),
    .X(_13919_));
 sg13g2_buf_1 _21608_ (.A(_12391_),
    .X(_13920_));
 sg13g2_nand2_1 _21609_ (.Y(_13921_),
    .A(net205),
    .B(net174));
 sg13g2_nand2_1 _21610_ (.Y(_13922_),
    .A(net210),
    .B(_13664_));
 sg13g2_nor2_1 _21611_ (.A(_12071_),
    .B(net207),
    .Y(_13923_));
 sg13g2_xnor2_1 _21612_ (.Y(_13924_),
    .A(_13922_),
    .B(_13923_));
 sg13g2_xor2_1 _21613_ (.B(_13924_),
    .A(_13921_),
    .X(_13925_));
 sg13g2_nor2_1 _21614_ (.A(_13783_),
    .B(_13784_),
    .Y(_13926_));
 sg13g2_nand2_1 _21615_ (.Y(_13927_),
    .A(_13783_),
    .B(_13784_));
 sg13g2_o21ai_1 _21616_ (.B1(_13927_),
    .Y(_13928_),
    .A1(_13781_),
    .A2(_13926_));
 sg13g2_buf_1 _21617_ (.A(_13928_),
    .X(_13929_));
 sg13g2_nor2_1 _21618_ (.A(_13757_),
    .B(_13759_),
    .Y(_13930_));
 sg13g2_nand2_1 _21619_ (.Y(_13931_),
    .A(_13757_),
    .B(_13759_));
 sg13g2_o21ai_1 _21620_ (.B1(_13931_),
    .Y(_13932_),
    .A1(_13756_),
    .A2(_13930_));
 sg13g2_xnor2_1 _21621_ (.Y(_13933_),
    .A(_13929_),
    .B(_13932_));
 sg13g2_xnor2_1 _21622_ (.Y(_13934_),
    .A(_13925_),
    .B(_13933_));
 sg13g2_nand2_1 _21623_ (.Y(_13935_),
    .A(_13765_),
    .B(_13768_));
 sg13g2_o21ai_1 _21624_ (.B1(_13761_),
    .Y(_13936_),
    .A1(_13765_),
    .A2(_13768_));
 sg13g2_nand2_1 _21625_ (.Y(_13937_),
    .A(_13935_),
    .B(_13936_));
 sg13g2_xnor2_1 _21626_ (.Y(_13938_),
    .A(_13934_),
    .B(_13937_));
 sg13g2_xnor2_1 _21627_ (.Y(_13939_),
    .A(_13919_),
    .B(_13938_));
 sg13g2_a21oi_1 _21628_ (.A1(_13742_),
    .A2(_13772_),
    .Y(_13940_),
    .B1(_13771_));
 sg13g2_nor2_1 _21629_ (.A(_13800_),
    .B(_13804_),
    .Y(_13941_));
 sg13g2_nand2_1 _21630_ (.Y(_13942_),
    .A(_13800_),
    .B(_13804_));
 sg13g2_o21ai_1 _21631_ (.B1(_13942_),
    .Y(_13943_),
    .A1(_13801_),
    .A2(_13941_));
 sg13g2_buf_1 _21632_ (.A(_13943_),
    .X(_13944_));
 sg13g2_xnor2_1 _21633_ (.Y(_13945_),
    .A(_13940_),
    .B(_13944_));
 sg13g2_xnor2_1 _21634_ (.Y(_13946_),
    .A(_13939_),
    .B(_13945_));
 sg13g2_buf_1 _21635_ (.A(_12452_),
    .X(_13947_));
 sg13g2_buf_1 _21636_ (.A(_13174_),
    .X(_13948_));
 sg13g2_nand2_1 _21637_ (.Y(_13949_),
    .A(net233),
    .B(net173));
 sg13g2_buf_1 _21638_ (.A(_12337_),
    .X(_13950_));
 sg13g2_inv_1 _21639_ (.Y(_13951_),
    .A(net258));
 sg13g2_and2_1 _21640_ (.A(net232),
    .B(_13951_),
    .X(_13952_));
 sg13g2_buf_1 _21641_ (.A(_13952_),
    .X(_13953_));
 sg13g2_buf_1 _21642_ (.A(net211),
    .X(_13954_));
 sg13g2_nand2_1 _21643_ (.Y(_13955_),
    .A(net240),
    .B(net172));
 sg13g2_xor2_1 _21644_ (.B(_13955_),
    .A(_13953_),
    .X(_13956_));
 sg13g2_xnor2_1 _21645_ (.Y(_13957_),
    .A(_13949_),
    .B(_13956_));
 sg13g2_nand2_1 _21646_ (.Y(_13958_),
    .A(_13351_),
    .B(_12762_));
 sg13g2_nand2_1 _21647_ (.Y(_13959_),
    .A(net234),
    .B(_12925_));
 sg13g2_and2_1 _21648_ (.A(net292),
    .B(net500),
    .X(_13960_));
 sg13g2_xnor2_1 _21649_ (.Y(_13961_),
    .A(_13959_),
    .B(_13960_));
 sg13g2_xnor2_1 _21650_ (.Y(_13962_),
    .A(_13958_),
    .B(_13961_));
 sg13g2_nand2_1 _21651_ (.Y(_13963_),
    .A(_13787_),
    .B(_13792_));
 sg13g2_nand2_1 _21652_ (.Y(_13964_),
    .A(_13790_),
    .B(_13963_));
 sg13g2_o21ai_1 _21653_ (.B1(_13964_),
    .Y(_13965_),
    .A1(_13787_),
    .A2(_13792_));
 sg13g2_buf_1 _21654_ (.A(_13965_),
    .X(_13966_));
 sg13g2_xnor2_1 _21655_ (.Y(_13967_),
    .A(_13962_),
    .B(_13966_));
 sg13g2_xnor2_1 _21656_ (.Y(_13968_),
    .A(_13957_),
    .B(_13967_));
 sg13g2_nand2_1 _21657_ (.Y(_13969_),
    .A(_13794_),
    .B(_13798_));
 sg13g2_nor2_1 _21658_ (.A(_13794_),
    .B(_13798_),
    .Y(_13970_));
 sg13g2_a21oi_1 _21659_ (.A1(_13786_),
    .A2(_13969_),
    .Y(_13971_),
    .B1(_13970_));
 sg13g2_a21o_1 _21660_ (.A2(_13819_),
    .A1(_13816_),
    .B1(_13812_),
    .X(_13972_));
 sg13g2_o21ai_1 _21661_ (.B1(_13972_),
    .Y(_13973_),
    .A1(_13816_),
    .A2(_13819_));
 sg13g2_buf_1 _21662_ (.A(_13973_),
    .X(_13974_));
 sg13g2_xnor2_1 _21663_ (.Y(_13975_),
    .A(_13971_),
    .B(_13974_));
 sg13g2_xnor2_1 _21664_ (.Y(_13976_),
    .A(_13968_),
    .B(_13975_));
 sg13g2_and2_1 _21665_ (.A(net300),
    .B(net499),
    .X(_13977_));
 sg13g2_buf_1 _21666_ (.A(_13977_),
    .X(_13978_));
 sg13g2_nand2_1 _21667_ (.Y(_13979_),
    .A(net301),
    .B(net501));
 sg13g2_nand2_1 _21668_ (.Y(_13980_),
    .A(net293),
    .B(net519));
 sg13g2_xnor2_1 _21669_ (.Y(_13981_),
    .A(_13979_),
    .B(_13980_));
 sg13g2_xnor2_1 _21670_ (.Y(_13982_),
    .A(_13978_),
    .B(_13981_));
 sg13g2_and2_1 _21671_ (.A(_13808_),
    .B(_13809_),
    .X(_13983_));
 sg13g2_or2_1 _21672_ (.X(_13984_),
    .B(_13809_),
    .A(_13808_));
 sg13g2_o21ai_1 _21673_ (.B1(_13984_),
    .Y(_13985_),
    .A1(_13810_),
    .A2(_13983_));
 sg13g2_buf_1 _21674_ (.A(_13985_),
    .X(_13986_));
 sg13g2_a22oi_1 _21675_ (.Y(_13987_),
    .B1(_13822_),
    .B2(_13825_),
    .A2(net502),
    .A1(net362));
 sg13g2_nor2_1 _21676_ (.A(_13822_),
    .B(_13825_),
    .Y(_13988_));
 sg13g2_nor2_1 _21677_ (.A(_13987_),
    .B(_13988_),
    .Y(_13989_));
 sg13g2_xnor2_1 _21678_ (.Y(_13990_),
    .A(_13986_),
    .B(_13989_));
 sg13g2_xnor2_1 _21679_ (.Y(_13991_),
    .A(_13982_),
    .B(_13990_));
 sg13g2_nor2_1 _21680_ (.A(_12197_),
    .B(_13387_),
    .Y(_13992_));
 sg13g2_nand2_1 _21681_ (.Y(_13993_),
    .A(net363),
    .B(net502));
 sg13g2_and2_1 _21682_ (.A(net332),
    .B(net479),
    .X(_13994_));
 sg13g2_buf_1 _21683_ (.A(_13994_),
    .X(_13995_));
 sg13g2_xor2_1 _21684_ (.B(_13995_),
    .A(_13993_),
    .X(_13996_));
 sg13g2_xnor2_1 _21685_ (.Y(_13997_),
    .A(_13992_),
    .B(_13996_));
 sg13g2_a22oi_1 _21686_ (.Y(_13998_),
    .B1(_13828_),
    .B2(_13829_),
    .A2(_13475_),
    .A1(_12974_));
 sg13g2_nor2_1 _21687_ (.A(_13828_),
    .B(_13829_),
    .Y(_13999_));
 sg13g2_nor2_1 _21688_ (.A(_13998_),
    .B(_13999_),
    .Y(_14000_));
 sg13g2_nand2_1 _21689_ (.Y(_14001_),
    .A(net362),
    .B(net480));
 sg13g2_nor2_1 _21690_ (.A(net404),
    .B(net566),
    .Y(_14002_));
 sg13g2_and2_1 _21691_ (.A(_12410_),
    .B(_13475_),
    .X(_14003_));
 sg13g2_buf_1 _21692_ (.A(_14003_),
    .X(_14004_));
 sg13g2_xor2_1 _21693_ (.B(_14004_),
    .A(_14002_),
    .X(_14005_));
 sg13g2_xnor2_1 _21694_ (.Y(_14006_),
    .A(_14001_),
    .B(_14005_));
 sg13g2_and2_1 _21695_ (.A(_14000_),
    .B(_14006_),
    .X(_14007_));
 sg13g2_or2_1 _21696_ (.X(_14008_),
    .B(_14006_),
    .A(_14000_));
 sg13g2_nor2b_1 _21697_ (.A(_14007_),
    .B_N(_14008_),
    .Y(_14009_));
 sg13g2_xnor2_1 _21698_ (.Y(_14010_),
    .A(_13997_),
    .B(_14009_));
 sg13g2_nand2b_1 _21699_ (.Y(_14011_),
    .B(_13836_),
    .A_N(_13832_));
 sg13g2_nor2b_1 _21700_ (.A(_13836_),
    .B_N(_13832_),
    .Y(_14012_));
 sg13g2_a21oi_1 _21701_ (.A1(_13827_),
    .A2(_14011_),
    .Y(_14013_),
    .B1(_14012_));
 sg13g2_xnor2_1 _21702_ (.Y(_14014_),
    .A(_14010_),
    .B(_14013_));
 sg13g2_xnor2_1 _21703_ (.Y(_14015_),
    .A(_13991_),
    .B(_14014_));
 sg13g2_nor2_1 _21704_ (.A(_13838_),
    .B(_13845_),
    .Y(_14016_));
 sg13g2_nand2_1 _21705_ (.Y(_14017_),
    .A(_13838_),
    .B(_13845_));
 sg13g2_o21ai_1 _21706_ (.B1(_14017_),
    .Y(_14018_),
    .A1(_13821_),
    .A2(_14016_));
 sg13g2_buf_1 _21707_ (.A(_14018_),
    .X(_14019_));
 sg13g2_xor2_1 _21708_ (.B(_14019_),
    .A(_14015_),
    .X(_14020_));
 sg13g2_xnor2_1 _21709_ (.Y(_14021_),
    .A(_13976_),
    .B(_14020_));
 sg13g2_nor2_1 _21710_ (.A(_13806_),
    .B(_13851_),
    .Y(_14022_));
 sg13g2_nor2_1 _21711_ (.A(_13850_),
    .B(_14022_),
    .Y(_14023_));
 sg13g2_xnor2_1 _21712_ (.Y(_14024_),
    .A(_14021_),
    .B(_14023_));
 sg13g2_xnor2_1 _21713_ (.Y(_14025_),
    .A(_13946_),
    .B(_14024_));
 sg13g2_nand2_1 _21714_ (.Y(_14026_),
    .A(_13774_),
    .B(_13778_));
 sg13g2_o21ai_1 _21715_ (.B1(_13740_),
    .Y(_14027_),
    .A1(_13774_),
    .A2(_13778_));
 sg13g2_nand2_1 _21716_ (.Y(_14028_),
    .A(net481),
    .B(net257));
 sg13g2_nand2_1 _21717_ (.Y(_14029_),
    .A(_13750_),
    .B(_14028_));
 sg13g2_nand2_1 _21718_ (.Y(_14030_),
    .A(net504),
    .B(_13750_));
 sg13g2_a21oi_1 _21719_ (.A1(_13746_),
    .A2(_14030_),
    .Y(_14031_),
    .B1(net521));
 sg13g2_or2_1 _21720_ (.X(_14032_),
    .B(_13750_),
    .A(net504));
 sg13g2_a21oi_1 _21721_ (.A1(net521),
    .A2(_13746_),
    .Y(_14033_),
    .B1(_14032_));
 sg13g2_o21ai_1 _21722_ (.B1(net257),
    .Y(_14034_),
    .A1(_14031_),
    .A2(_14033_));
 sg13g2_o21ai_1 _21723_ (.B1(_14034_),
    .Y(_14035_),
    .A1(_13746_),
    .A2(_14029_));
 sg13g2_nand3_1 _21724_ (.B(_14027_),
    .C(_14035_),
    .A(_14026_),
    .Y(_14036_));
 sg13g2_buf_1 _21725_ (.A(_14036_),
    .X(_14037_));
 sg13g2_a21o_1 _21726_ (.A2(_14027_),
    .A1(_14026_),
    .B1(_14035_),
    .X(_14038_));
 sg13g2_and2_1 _21727_ (.A(_14037_),
    .B(_14038_),
    .X(_14039_));
 sg13g2_nor2_1 _21728_ (.A(_14025_),
    .B(_14039_),
    .Y(_14040_));
 sg13g2_nand2_1 _21729_ (.Y(_14041_),
    .A(_14025_),
    .B(_14039_));
 sg13g2_nor2b_1 _21730_ (.A(_14040_),
    .B_N(_14041_),
    .Y(_14042_));
 sg13g2_xnor2_1 _21731_ (.Y(_14043_),
    .A(_13902_),
    .B(_14042_));
 sg13g2_xnor2_1 _21732_ (.Y(_14044_),
    .A(_13901_),
    .B(_14043_));
 sg13g2_xnor2_1 _21733_ (.Y(_14045_),
    .A(_13900_),
    .B(_14044_));
 sg13g2_o21ai_1 _21734_ (.B1(_13733_),
    .Y(_14046_),
    .A1(_13731_),
    .A2(_13866_));
 sg13g2_nand2_1 _21735_ (.Y(_14047_),
    .A(_13731_),
    .B(_13866_));
 sg13g2_nand2_1 _21736_ (.Y(_14048_),
    .A(_14046_),
    .B(_14047_));
 sg13g2_xor2_1 _21737_ (.B(_14048_),
    .A(_14045_),
    .X(_14049_));
 sg13g2_xnor2_1 _21738_ (.Y(_14050_),
    .A(_13897_),
    .B(_14049_));
 sg13g2_nor2_1 _21739_ (.A(_08681_),
    .B(_14050_),
    .Y(_14051_));
 sg13g2_a21oi_1 _21740_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(net452),
    .Y(_14052_),
    .B1(_14051_));
 sg13g2_nor2_1 _21741_ (.A(net634),
    .B(_14052_),
    .Y(_01519_));
 sg13g2_nor2_1 _21742_ (.A(_14045_),
    .B(_14048_),
    .Y(_14053_));
 sg13g2_nor2_1 _21743_ (.A(_13893_),
    .B(_14053_),
    .Y(_14054_));
 sg13g2_a22oi_1 _21744_ (.Y(_14055_),
    .B1(_14054_),
    .B2(_13896_),
    .A2(_14048_),
    .A1(_14045_));
 sg13g2_o21ai_1 _21745_ (.B1(_13900_),
    .Y(_14056_),
    .A1(_13901_),
    .A2(_14043_));
 sg13g2_nand2_1 _21746_ (.Y(_14057_),
    .A(_13901_),
    .B(_14043_));
 sg13g2_o21ai_1 _21747_ (.B1(_13946_),
    .Y(_14058_),
    .A1(_14021_),
    .A2(_14023_));
 sg13g2_inv_1 _21748_ (.Y(_14059_),
    .A(_14058_));
 sg13g2_a21oi_1 _21749_ (.A1(_14021_),
    .A2(_14023_),
    .Y(_14060_),
    .B1(_14059_));
 sg13g2_nand2_1 _21750_ (.Y(_14061_),
    .A(_13919_),
    .B(_13937_));
 sg13g2_nor2_1 _21751_ (.A(_13919_),
    .B(_13937_),
    .Y(_14062_));
 sg13g2_a21oi_1 _21752_ (.A1(_13934_),
    .A2(_14061_),
    .Y(_14063_),
    .B1(_14062_));
 sg13g2_nand2_1 _21753_ (.Y(_14064_),
    .A(net205),
    .B(net150));
 sg13g2_nor2_1 _21754_ (.A(_12071_),
    .B(net208),
    .Y(_14065_));
 sg13g2_inv_1 _21755_ (.Y(_14066_),
    .A(_14065_));
 sg13g2_nand2_1 _21756_ (.Y(_14067_),
    .A(net210),
    .B(net174));
 sg13g2_xnor2_1 _21757_ (.Y(_14068_),
    .A(_14066_),
    .B(_14067_));
 sg13g2_xnor2_1 _21758_ (.Y(_14069_),
    .A(_14064_),
    .B(_14068_));
 sg13g2_nor2b_1 _21759_ (.A(_13953_),
    .B_N(_13955_),
    .Y(_14070_));
 sg13g2_buf_1 _21760_ (.A(_12335_),
    .X(_14071_));
 sg13g2_nand3_1 _21761_ (.B(net172),
    .C(_13953_),
    .A(net204),
    .Y(_14072_));
 sg13g2_o21ai_1 _21762_ (.B1(_14072_),
    .Y(_14073_),
    .A1(_13949_),
    .A2(_14070_));
 sg13g2_buf_1 _21763_ (.A(_14073_),
    .X(_14074_));
 sg13g2_a21oi_1 _21764_ (.A1(net205),
    .A2(net174),
    .Y(_14075_),
    .B1(_13923_));
 sg13g2_nand3_1 _21765_ (.B(net174),
    .C(_13923_),
    .A(net205),
    .Y(_14076_));
 sg13g2_o21ai_1 _21766_ (.B1(_14076_),
    .Y(_14077_),
    .A1(_13922_),
    .A2(_14075_));
 sg13g2_buf_1 _21767_ (.A(_14077_),
    .X(_14078_));
 sg13g2_xnor2_1 _21768_ (.Y(_14079_),
    .A(_14074_),
    .B(_14078_));
 sg13g2_xnor2_1 _21769_ (.Y(_14080_),
    .A(_14069_),
    .B(_14079_));
 sg13g2_or2_1 _21770_ (.X(_14081_),
    .B(_13932_),
    .A(_13929_));
 sg13g2_nand2_1 _21771_ (.Y(_14082_),
    .A(_13929_),
    .B(_13932_));
 sg13g2_nand2_1 _21772_ (.Y(_14083_),
    .A(_13925_),
    .B(_14082_));
 sg13g2_nand2_1 _21773_ (.Y(_14084_),
    .A(net481),
    .B(net206));
 sg13g2_o21ai_1 _21774_ (.B1(_14084_),
    .Y(_14085_),
    .A1(net568),
    .A2(_13905_));
 sg13g2_nand2_1 _21775_ (.Y(_14086_),
    .A(net568),
    .B(_12403_));
 sg13g2_nor2_1 _21776_ (.A(net235),
    .B(_14086_),
    .Y(_14087_));
 sg13g2_a21oi_1 _21777_ (.A1(net235),
    .A2(_14085_),
    .Y(_14088_),
    .B1(_14087_));
 sg13g2_xnor2_1 _21778_ (.Y(_14089_),
    .A(_12415_),
    .B(_14088_));
 sg13g2_a22oi_1 _21779_ (.Y(_14090_),
    .B1(_14089_),
    .B2(net257),
    .A2(_14083_),
    .A1(_14081_));
 sg13g2_nand4_1 _21780_ (.B(_14081_),
    .C(_14083_),
    .A(net257),
    .Y(_14091_),
    .D(_14089_));
 sg13g2_nand2b_1 _21781_ (.Y(_14092_),
    .B(_14091_),
    .A_N(_14090_));
 sg13g2_xor2_1 _21782_ (.B(_14092_),
    .A(_14080_),
    .X(_14093_));
 sg13g2_inv_1 _21783_ (.Y(_14094_),
    .A(_14093_));
 sg13g2_nor2_1 _21784_ (.A(_13968_),
    .B(_13974_),
    .Y(_14095_));
 sg13g2_nand2_1 _21785_ (.Y(_14096_),
    .A(_13968_),
    .B(_13974_));
 sg13g2_o21ai_1 _21786_ (.B1(_14096_),
    .Y(_14097_),
    .A1(_13971_),
    .A2(_14095_));
 sg13g2_nor2_1 _21787_ (.A(_14094_),
    .B(_14097_),
    .Y(_14098_));
 sg13g2_nand2_1 _21788_ (.Y(_14099_),
    .A(_14094_),
    .B(_14097_));
 sg13g2_nor2b_1 _21789_ (.A(_14098_),
    .B_N(_14099_),
    .Y(_14100_));
 sg13g2_xnor2_1 _21790_ (.Y(_14101_),
    .A(_14063_),
    .B(_14100_));
 sg13g2_nand2_1 _21791_ (.Y(_14102_),
    .A(_13962_),
    .B(_13966_));
 sg13g2_nand2_1 _21792_ (.Y(_14103_),
    .A(_13957_),
    .B(_14102_));
 sg13g2_o21ai_1 _21793_ (.B1(_14103_),
    .Y(_14104_),
    .A1(_13962_),
    .A2(_13966_));
 sg13g2_buf_1 _21794_ (.A(net276),
    .X(_01810_));
 sg13g2_nand2_1 _21795_ (.Y(_01811_),
    .A(net256),
    .B(net500));
 sg13g2_buf_1 _21796_ (.A(_12762_),
    .X(_01812_));
 sg13g2_nand2_1 _21797_ (.Y(_01813_),
    .A(net234),
    .B(net255));
 sg13g2_nor2_1 _21798_ (.A(_12153_),
    .B(net258),
    .Y(_01814_));
 sg13g2_xnor2_1 _21799_ (.Y(_01815_),
    .A(_01813_),
    .B(_01814_));
 sg13g2_xnor2_1 _21800_ (.Y(_01816_),
    .A(_01811_),
    .B(_01815_));
 sg13g2_nor2_1 _21801_ (.A(_13958_),
    .B(_13959_),
    .Y(_01817_));
 sg13g2_nor2_1 _21802_ (.A(_13960_),
    .B(_01817_),
    .Y(_01818_));
 sg13g2_a21oi_1 _21803_ (.A1(_13958_),
    .A2(_13959_),
    .Y(_01819_),
    .B1(_01818_));
 sg13g2_nor2b_1 _21804_ (.A(net207),
    .B_N(net233),
    .Y(_01820_));
 sg13g2_nand2_1 _21805_ (.Y(_01821_),
    .A(net232),
    .B(net172));
 sg13g2_nand2_1 _21806_ (.Y(_01822_),
    .A(_12335_),
    .B(net173));
 sg13g2_xnor2_1 _21807_ (.Y(_01823_),
    .A(_01821_),
    .B(_01822_));
 sg13g2_xnor2_1 _21808_ (.Y(_01824_),
    .A(_01820_),
    .B(_01823_));
 sg13g2_xnor2_1 _21809_ (.Y(_01825_),
    .A(_01819_),
    .B(_01824_));
 sg13g2_xnor2_1 _21810_ (.Y(_01826_),
    .A(_01816_),
    .B(_01825_));
 sg13g2_o21ai_1 _21811_ (.B1(_13989_),
    .Y(_01827_),
    .A1(_13986_),
    .A2(_13982_));
 sg13g2_nand2_1 _21812_ (.Y(_01828_),
    .A(_13986_),
    .B(_13982_));
 sg13g2_nand2_1 _21813_ (.Y(_01829_),
    .A(_01827_),
    .B(_01828_));
 sg13g2_nor2_1 _21814_ (.A(_01826_),
    .B(_01829_),
    .Y(_01830_));
 sg13g2_nand2_1 _21815_ (.Y(_01831_),
    .A(_01826_),
    .B(_01829_));
 sg13g2_nand2b_1 _21816_ (.Y(_01832_),
    .B(_01831_),
    .A_N(_01830_));
 sg13g2_xnor2_1 _21817_ (.Y(_01833_),
    .A(_14104_),
    .B(_01832_));
 sg13g2_inv_1 _21818_ (.Y(_01834_),
    .A(_13991_));
 sg13g2_a21oi_1 _21819_ (.A1(_14010_),
    .A2(_14013_),
    .Y(_01835_),
    .B1(_01834_));
 sg13g2_nor2_1 _21820_ (.A(_14010_),
    .B(_14013_),
    .Y(_01836_));
 sg13g2_and2_1 _21821_ (.A(_12928_),
    .B(net499),
    .X(_01837_));
 sg13g2_buf_1 _21822_ (.A(_01837_),
    .X(_01838_));
 sg13g2_buf_1 _21823_ (.A(net293),
    .X(_01839_));
 sg13g2_nand2_1 _21824_ (.Y(_01840_),
    .A(net288),
    .B(net501));
 sg13g2_buf_1 _21825_ (.A(_12837_),
    .X(_01841_));
 sg13g2_and2_1 _21826_ (.A(net300),
    .B(net498),
    .X(_01842_));
 sg13g2_buf_1 _21827_ (.A(_01842_),
    .X(_01843_));
 sg13g2_xor2_1 _21828_ (.B(_01843_),
    .A(_01840_),
    .X(_01844_));
 sg13g2_xnor2_1 _21829_ (.Y(_01845_),
    .A(_01838_),
    .B(_01844_));
 sg13g2_buf_1 _21830_ (.A(_13246_),
    .X(_01846_));
 sg13g2_a22oi_1 _21831_ (.Y(_01847_),
    .B1(_13992_),
    .B2(_13995_),
    .A2(net478),
    .A1(net363));
 sg13g2_nor2_1 _21832_ (.A(_13992_),
    .B(_13995_),
    .Y(_01848_));
 sg13g2_nor2_1 _21833_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sg13g2_nor2b_1 _21834_ (.A(_13978_),
    .B_N(_13980_),
    .Y(_01850_));
 sg13g2_nand3_1 _21835_ (.B(net498),
    .C(_13978_),
    .A(net288),
    .Y(_01851_));
 sg13g2_o21ai_1 _21836_ (.B1(_01851_),
    .Y(_01852_),
    .A1(_13979_),
    .A2(_01850_));
 sg13g2_buf_1 _21837_ (.A(_01852_),
    .X(_01853_));
 sg13g2_xnor2_1 _21838_ (.Y(_01854_),
    .A(_01849_),
    .B(_01853_));
 sg13g2_xnor2_1 _21839_ (.Y(_01855_),
    .A(_01845_),
    .B(_01854_));
 sg13g2_a21oi_2 _21840_ (.B1(_13387_),
    .Y(_01856_),
    .A2(_11791_),
    .A1(_11782_));
 sg13g2_nand2_1 _21841_ (.Y(_01857_),
    .A(net332),
    .B(_13246_));
 sg13g2_nand2_1 _21842_ (.Y(_01858_),
    .A(net319),
    .B(net479));
 sg13g2_xnor2_1 _21843_ (.Y(_01859_),
    .A(_01857_),
    .B(_01858_));
 sg13g2_xnor2_1 _21844_ (.Y(_01860_),
    .A(_01856_),
    .B(_01859_));
 sg13g2_nor2_1 _21845_ (.A(_11913_),
    .B(_13633_),
    .Y(_01861_));
 sg13g2_nor2_1 _21846_ (.A(_12410_),
    .B(net566),
    .Y(_01862_));
 sg13g2_buf_1 _21847_ (.A(_13475_),
    .X(_01863_));
 sg13g2_nand2_1 _21848_ (.Y(_01864_),
    .A(net362),
    .B(net477));
 sg13g2_xor2_1 _21849_ (.B(_01864_),
    .A(_01862_),
    .X(_01865_));
 sg13g2_xnor2_1 _21850_ (.Y(_01866_),
    .A(_01861_),
    .B(_01865_));
 sg13g2_a22oi_1 _21851_ (.Y(_01867_),
    .B1(_14002_),
    .B2(_14004_),
    .A2(net480),
    .A1(net362));
 sg13g2_nor2_1 _21852_ (.A(_14002_),
    .B(_14004_),
    .Y(_01868_));
 sg13g2_nor2_1 _21853_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sg13g2_xnor2_1 _21854_ (.Y(_01870_),
    .A(_01866_),
    .B(_01869_));
 sg13g2_xnor2_1 _21855_ (.Y(_01871_),
    .A(_01860_),
    .B(_01870_));
 sg13g2_a21o_1 _21856_ (.A2(_14008_),
    .A1(_13997_),
    .B1(_14007_),
    .X(_01872_));
 sg13g2_buf_1 _21857_ (.A(_01872_),
    .X(_01873_));
 sg13g2_xnor2_1 _21858_ (.Y(_01874_),
    .A(_01871_),
    .B(_01873_));
 sg13g2_xnor2_1 _21859_ (.Y(_01875_),
    .A(_01855_),
    .B(_01874_));
 sg13g2_o21ai_1 _21860_ (.B1(_01875_),
    .Y(_01876_),
    .A1(_01835_),
    .A2(_01836_));
 sg13g2_or3_1 _21861_ (.A(_01875_),
    .B(_01835_),
    .C(_01836_),
    .X(_01877_));
 sg13g2_nand2_1 _21862_ (.Y(_01878_),
    .A(_01876_),
    .B(_01877_));
 sg13g2_xnor2_1 _21863_ (.Y(_01879_),
    .A(_01833_),
    .B(_01878_));
 sg13g2_inv_1 _21864_ (.Y(_01880_),
    .A(_14015_));
 sg13g2_nand2_1 _21865_ (.Y(_01881_),
    .A(_01880_),
    .B(_14019_));
 sg13g2_nor2_1 _21866_ (.A(_01880_),
    .B(_14019_),
    .Y(_01882_));
 sg13g2_a21oi_2 _21867_ (.B1(_01882_),
    .Y(_01883_),
    .A2(_01881_),
    .A1(_13976_));
 sg13g2_xor2_1 _21868_ (.B(_01883_),
    .A(_01879_),
    .X(_01884_));
 sg13g2_xnor2_1 _21869_ (.Y(_01885_),
    .A(_14101_),
    .B(_01884_));
 sg13g2_nor2_1 _21870_ (.A(_13939_),
    .B(_13944_),
    .Y(_01886_));
 sg13g2_nand2_1 _21871_ (.Y(_01887_),
    .A(_13939_),
    .B(_13944_));
 sg13g2_o21ai_1 _21872_ (.B1(_01887_),
    .Y(_01888_),
    .A1(_13940_),
    .A2(_01886_));
 sg13g2_a21oi_1 _21873_ (.A1(net206),
    .A2(_13915_),
    .Y(_01889_),
    .B1(_13747_));
 sg13g2_buf_1 _21874_ (.A(_13903_),
    .X(_01890_));
 sg13g2_buf_1 _21875_ (.A(_13676_),
    .X(_01891_));
 sg13g2_nand3_1 _21876_ (.B(net231),
    .C(_13747_),
    .A(_01890_),
    .Y(_01892_));
 sg13g2_o21ai_1 _21877_ (.B1(_01892_),
    .Y(_01893_),
    .A1(_14028_),
    .A2(_01889_));
 sg13g2_xnor2_1 _21878_ (.Y(_01894_),
    .A(_13023_),
    .B(_13918_));
 sg13g2_a22oi_1 _21879_ (.Y(_01895_),
    .B1(_01894_),
    .B2(_13677_),
    .A2(_01893_),
    .A1(net235));
 sg13g2_xor2_1 _21880_ (.B(_01895_),
    .A(_01888_),
    .X(_01896_));
 sg13g2_xor2_1 _21881_ (.B(_01896_),
    .A(_01885_),
    .X(_01897_));
 sg13g2_xnor2_1 _21882_ (.Y(_01898_),
    .A(_14060_),
    .B(_01897_));
 sg13g2_a21oi_1 _21883_ (.A1(_13902_),
    .A2(_14041_),
    .Y(_01899_),
    .B1(_14040_));
 sg13g2_xnor2_1 _21884_ (.Y(_01900_),
    .A(_14037_),
    .B(_01899_));
 sg13g2_xnor2_1 _21885_ (.Y(_01901_),
    .A(_01898_),
    .B(_01900_));
 sg13g2_and3_1 _21886_ (.X(_01902_),
    .A(_14056_),
    .B(_14057_),
    .C(_01901_));
 sg13g2_a21o_1 _21887_ (.A2(_14057_),
    .A1(_14056_),
    .B1(_01901_),
    .X(_01903_));
 sg13g2_nor2b_1 _21888_ (.A(_01902_),
    .B_N(_01903_),
    .Y(_01904_));
 sg13g2_xnor2_1 _21889_ (.Y(_01905_),
    .A(_14055_),
    .B(_01904_));
 sg13g2_nand2_1 _21890_ (.Y(_01906_),
    .A(net450),
    .B(_01905_));
 sg13g2_nand2_1 _21891_ (.Y(_01907_),
    .A(\rbzero.traced_texVinit[10] ),
    .B(net442));
 sg13g2_a21oi_1 _21892_ (.A1(_01906_),
    .A2(_01907_),
    .Y(_01520_),
    .B1(net572));
 sg13g2_nand2_1 _21893_ (.Y(_01908_),
    .A(_11846_),
    .B(net449));
 sg13g2_nand2_1 _21894_ (.Y(_01909_),
    .A(_09540_),
    .B(net442));
 sg13g2_a21oi_1 _21895_ (.A1(_01908_),
    .A2(_01909_),
    .Y(_01521_),
    .B1(net572));
 sg13g2_nand2_1 _21896_ (.Y(_01910_),
    .A(_08533_),
    .B(net449));
 sg13g2_nand2_1 _21897_ (.Y(_01911_),
    .A(_09583_),
    .B(net442));
 sg13g2_a21oi_1 _21898_ (.A1(_01910_),
    .A2(_01911_),
    .Y(_01522_),
    .B1(_11765_));
 sg13g2_buf_1 _21899_ (.A(_08808_),
    .X(_01912_));
 sg13g2_nand2_1 _21900_ (.Y(_01913_),
    .A(_08532_),
    .B(_01912_));
 sg13g2_nand2_1 _21901_ (.Y(_01914_),
    .A(_09591_),
    .B(net442));
 sg13g2_a21oi_1 _21902_ (.A1(_01913_),
    .A2(_01914_),
    .Y(_01523_),
    .B1(net572));
 sg13g2_nand2_1 _21903_ (.Y(_01915_),
    .A(_08538_),
    .B(net441));
 sg13g2_nand2_1 _21904_ (.Y(_01916_),
    .A(_09595_),
    .B(_13883_));
 sg13g2_buf_1 _21905_ (.A(_11764_),
    .X(_01917_));
 sg13g2_a21oi_1 _21906_ (.A1(_01915_),
    .A2(_01916_),
    .Y(_01524_),
    .B1(net565));
 sg13g2_nand2_1 _21907_ (.Y(_01918_),
    .A(_08537_),
    .B(net441));
 sg13g2_nand2_1 _21908_ (.Y(_01919_),
    .A(_09605_),
    .B(_13883_));
 sg13g2_a21oi_1 _21909_ (.A1(_01918_),
    .A2(_01919_),
    .Y(_01525_),
    .B1(net565));
 sg13g2_nand2_1 _21910_ (.Y(_01920_),
    .A(_08536_),
    .B(net441));
 sg13g2_nand2_1 _21911_ (.Y(_01921_),
    .A(_09612_),
    .B(net442));
 sg13g2_a21oi_1 _21912_ (.A1(_01920_),
    .A2(_01921_),
    .Y(_01526_),
    .B1(_01917_));
 sg13g2_nand2_1 _21913_ (.Y(_01922_),
    .A(_08535_),
    .B(_01912_));
 sg13g2_nand2_1 _21914_ (.Y(_01923_),
    .A(_09620_),
    .B(net442));
 sg13g2_a21oi_1 _21915_ (.A1(_01922_),
    .A2(_01923_),
    .Y(_01527_),
    .B1(_01917_));
 sg13g2_nand2_1 _21916_ (.Y(_01924_),
    .A(_08547_),
    .B(net441));
 sg13g2_nand2_1 _21917_ (.Y(_01925_),
    .A(_09628_),
    .B(net442));
 sg13g2_a21oi_1 _21918_ (.A1(_01924_),
    .A2(_01925_),
    .Y(_01528_),
    .B1(net565));
 sg13g2_nand2_1 _21919_ (.Y(_01926_),
    .A(_08546_),
    .B(net441));
 sg13g2_buf_1 _21920_ (.A(_08681_),
    .X(_01927_));
 sg13g2_nand2_1 _21921_ (.Y(_01928_),
    .A(_09632_),
    .B(net440));
 sg13g2_a21oi_1 _21922_ (.A1(_01926_),
    .A2(_01928_),
    .Y(_01529_),
    .B1(net565));
 sg13g2_nand2_1 _21923_ (.Y(_01929_),
    .A(_08545_),
    .B(net441));
 sg13g2_nand2_1 _21924_ (.Y(_01930_),
    .A(_09643_),
    .B(net440));
 sg13g2_a21oi_1 _21925_ (.A1(_01929_),
    .A2(_01930_),
    .Y(_01530_),
    .B1(net565));
 sg13g2_nand2_1 _21926_ (.Y(_01931_),
    .A(_08542_),
    .B(net441));
 sg13g2_nand2_1 _21927_ (.Y(_01932_),
    .A(_09647_),
    .B(_01927_));
 sg13g2_a21oi_1 _21928_ (.A1(_01931_),
    .A2(_01932_),
    .Y(_01531_),
    .B1(net565));
 sg13g2_nand2_1 _21929_ (.Y(_01933_),
    .A(_11796_),
    .B(net441));
 sg13g2_nand2_1 _21930_ (.Y(_01934_),
    .A(_09554_),
    .B(net440));
 sg13g2_a21oi_1 _21931_ (.A1(_01933_),
    .A2(_01934_),
    .Y(_01532_),
    .B1(net565));
 sg13g2_buf_1 _21932_ (.A(_08808_),
    .X(_01935_));
 sg13g2_nand2_1 _21933_ (.Y(_01936_),
    .A(_08543_),
    .B(net439));
 sg13g2_nand2_1 _21934_ (.Y(_01937_),
    .A(_09669_),
    .B(net440));
 sg13g2_a21oi_1 _21935_ (.A1(_01936_),
    .A2(_01937_),
    .Y(_01533_),
    .B1(net565));
 sg13g2_nand2_1 _21936_ (.Y(_01938_),
    .A(_08481_),
    .B(net439));
 sg13g2_nand2_1 _21937_ (.Y(_01939_),
    .A(\rbzero.traced_texa[10] ),
    .B(net440));
 sg13g2_buf_1 _21938_ (.A(_11764_),
    .X(_01940_));
 sg13g2_a21oi_1 _21939_ (.A1(_01938_),
    .A2(_01939_),
    .Y(_01534_),
    .B1(net564));
 sg13g2_nand2_1 _21940_ (.Y(_01941_),
    .A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_01935_));
 sg13g2_nand2_1 _21941_ (.Y(_01942_),
    .A(_09552_),
    .B(net440));
 sg13g2_a21oi_1 _21942_ (.A1(_01941_),
    .A2(_01942_),
    .Y(_01535_),
    .B1(net564));
 sg13g2_nand2_1 _21943_ (.Y(_01943_),
    .A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(net439));
 sg13g2_nand2_1 _21944_ (.Y(_01944_),
    .A(_09551_),
    .B(net440));
 sg13g2_a21oi_1 _21945_ (.A1(_01943_),
    .A2(_01944_),
    .Y(_01536_),
    .B1(net564));
 sg13g2_nand2_1 _21946_ (.Y(_01945_),
    .A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(net439));
 sg13g2_nand2_1 _21947_ (.Y(_01946_),
    .A(_09549_),
    .B(net440));
 sg13g2_a21oi_1 _21948_ (.A1(_01945_),
    .A2(_01946_),
    .Y(_01537_),
    .B1(net564));
 sg13g2_nand2_1 _21949_ (.Y(_01947_),
    .A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(net439));
 sg13g2_nand2_1 _21950_ (.Y(_01948_),
    .A(_09548_),
    .B(_01927_));
 sg13g2_a21oi_1 _21951_ (.A1(_01947_),
    .A2(_01948_),
    .Y(_01538_),
    .B1(net564));
 sg13g2_nand2_1 _21952_ (.Y(_01949_),
    .A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_01935_));
 sg13g2_buf_1 _21953_ (.A(_08981_),
    .X(_01950_));
 sg13g2_nand2_1 _21954_ (.Y(_01951_),
    .A(_09546_),
    .B(net438));
 sg13g2_a21oi_1 _21955_ (.A1(_01949_),
    .A2(_01951_),
    .Y(_01539_),
    .B1(net564));
 sg13g2_nand2_1 _21956_ (.Y(_01952_),
    .A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(net439));
 sg13g2_nand2_1 _21957_ (.Y(_01953_),
    .A(_09545_),
    .B(net438));
 sg13g2_a21oi_1 _21958_ (.A1(_01952_),
    .A2(_01953_),
    .Y(_01540_),
    .B1(net564));
 sg13g2_nand2_1 _21959_ (.Y(_01954_),
    .A(_08541_),
    .B(net439));
 sg13g2_nand2_1 _21960_ (.Y(_01955_),
    .A(_09543_),
    .B(_01950_));
 sg13g2_a21oi_1 _21961_ (.A1(_01954_),
    .A2(_01955_),
    .Y(_01541_),
    .B1(net564));
 sg13g2_nand2_1 _21962_ (.Y(_01956_),
    .A(_08540_),
    .B(net439));
 sg13g2_nand2_1 _21963_ (.Y(_01957_),
    .A(_09542_),
    .B(_01950_));
 sg13g2_a21oi_1 _21964_ (.A1(_01956_),
    .A2(_01957_),
    .Y(_01542_),
    .B1(_01940_));
 sg13g2_nand2_1 _21965_ (.Y(_01958_),
    .A(\rbzero.wall_tracer.texu[0] ),
    .B(net459));
 sg13g2_buf_1 _21966_ (.A(\rbzero.row_render.texu[0] ),
    .X(_01959_));
 sg13g2_nand2_1 _21967_ (.Y(_01960_),
    .A(_01959_),
    .B(net438));
 sg13g2_a21oi_1 _21968_ (.A1(_01958_),
    .A2(_01960_),
    .Y(_01543_),
    .B1(_01940_));
 sg13g2_nand2_1 _21969_ (.Y(_01961_),
    .A(\rbzero.wall_tracer.texu[1] ),
    .B(net459));
 sg13g2_nand2_1 _21970_ (.Y(_01962_),
    .A(\rbzero.row_render.texu[1] ),
    .B(net438));
 sg13g2_buf_1 _21971_ (.A(_11764_),
    .X(_01963_));
 sg13g2_a21oi_1 _21972_ (.A1(_01961_),
    .A2(_01962_),
    .Y(_01544_),
    .B1(net563));
 sg13g2_nand2_1 _21973_ (.Y(_01964_),
    .A(\rbzero.wall_tracer.texu[2] ),
    .B(net459));
 sg13g2_buf_1 _21974_ (.A(\rbzero.row_render.texu[2] ),
    .X(_01965_));
 sg13g2_nand2_1 _21975_ (.Y(_01966_),
    .A(_01965_),
    .B(net438));
 sg13g2_a21oi_1 _21976_ (.A1(_01964_),
    .A2(_01966_),
    .Y(_01545_),
    .B1(net563));
 sg13g2_nand2_1 _21977_ (.Y(_01967_),
    .A(\rbzero.wall_tracer.texu[3] ),
    .B(net459));
 sg13g2_nand2_1 _21978_ (.Y(_01968_),
    .A(\rbzero.row_render.texu[3] ),
    .B(net438));
 sg13g2_a21oi_1 _21979_ (.A1(_01967_),
    .A2(_01968_),
    .Y(_01546_),
    .B1(_01963_));
 sg13g2_nand2_1 _21980_ (.Y(_01969_),
    .A(\rbzero.wall_tracer.texu[4] ),
    .B(net459));
 sg13g2_nand2_1 _21981_ (.Y(_01970_),
    .A(\rbzero.row_render.texu[4] ),
    .B(net438));
 sg13g2_a21oi_1 _21982_ (.A1(_01969_),
    .A2(_01970_),
    .Y(_01547_),
    .B1(_01963_));
 sg13g2_nand2_1 _21983_ (.Y(_01971_),
    .A(\rbzero.wall_tracer.texu[0] ),
    .B(net547));
 sg13g2_nand2_1 _21984_ (.Y(_01972_),
    .A(\rbzero.texu_hot[0] ),
    .B(net525));
 sg13g2_a21oi_1 _21985_ (.A1(_01971_),
    .A2(_01972_),
    .Y(_01548_),
    .B1(net563));
 sg13g2_nand2_1 _21986_ (.Y(_01973_),
    .A(\rbzero.wall_tracer.texu[1] ),
    .B(net547));
 sg13g2_buf_1 _21987_ (.A(\rbzero.texu_hot[1] ),
    .X(_01974_));
 sg13g2_nand2_1 _21988_ (.Y(_01975_),
    .A(_01974_),
    .B(net525));
 sg13g2_a21oi_1 _21989_ (.A1(_01973_),
    .A2(_01975_),
    .Y(_01549_),
    .B1(net563));
 sg13g2_nand2_1 _21990_ (.Y(_01976_),
    .A(\rbzero.wall_tracer.texu[2] ),
    .B(net547));
 sg13g2_nand2_1 _21991_ (.Y(_01977_),
    .A(\rbzero.texu_hot[2] ),
    .B(net525));
 sg13g2_a21oi_1 _21992_ (.A1(_01976_),
    .A2(_01977_),
    .Y(_01550_),
    .B1(net563));
 sg13g2_nand2_1 _21993_ (.Y(_01978_),
    .A(\rbzero.wall_tracer.texu[3] ),
    .B(net547));
 sg13g2_buf_1 _21994_ (.A(\rbzero.texu_hot[3] ),
    .X(_01979_));
 sg13g2_nand2_1 _21995_ (.Y(_01980_),
    .A(_01979_),
    .B(net525));
 sg13g2_a21oi_1 _21996_ (.A1(_01978_),
    .A2(_01980_),
    .Y(_01551_),
    .B1(net563));
 sg13g2_nand2_1 _21997_ (.Y(_01981_),
    .A(\rbzero.wall_tracer.texu[4] ),
    .B(_08477_));
 sg13g2_nand2_1 _21998_ (.Y(_01982_),
    .A(\rbzero.texu_hot[4] ),
    .B(net525));
 sg13g2_a21oi_1 _21999_ (.A1(_01981_),
    .A2(_01982_),
    .Y(_01552_),
    .B1(net563));
 sg13g2_nand2_1 _22000_ (.Y(_01983_),
    .A(\rbzero.wall_tracer.texu[5] ),
    .B(net547));
 sg13g2_buf_1 _22001_ (.A(\rbzero.texu_hot[5] ),
    .X(_01984_));
 sg13g2_nand2_1 _22002_ (.Y(_01985_),
    .A(_01984_),
    .B(net525));
 sg13g2_a21oi_1 _22003_ (.A1(_01983_),
    .A2(_01985_),
    .Y(_01553_),
    .B1(net563));
 sg13g2_nand2_1 _22004_ (.Y(_01986_),
    .A(\rbzero.wall_tracer.wall[0] ),
    .B(net459));
 sg13g2_buf_1 _22005_ (.A(\rbzero.row_render.wall[0] ),
    .X(_01987_));
 sg13g2_nand2_1 _22006_ (.Y(_01988_),
    .A(net810),
    .B(net438));
 sg13g2_buf_1 _22007_ (.A(_11764_),
    .X(_01989_));
 sg13g2_a21oi_1 _22008_ (.A1(_01986_),
    .A2(_01988_),
    .Y(_01554_),
    .B1(net562));
 sg13g2_nand2_1 _22009_ (.Y(_01990_),
    .A(\rbzero.wall_tracer.wall[1] ),
    .B(net459));
 sg13g2_buf_1 _22010_ (.A(\rbzero.row_render.wall[1] ),
    .X(_01991_));
 sg13g2_nand2_1 _22011_ (.Y(_01992_),
    .A(net809),
    .B(net464));
 sg13g2_a21oi_1 _22012_ (.A1(_01990_),
    .A2(_01992_),
    .Y(_01555_),
    .B1(net562));
 sg13g2_nand2_1 _22013_ (.Y(_01993_),
    .A(\rbzero.wall_tracer.wall[0] ),
    .B(net547));
 sg13g2_buf_1 _22014_ (.A(\rbzero.wall_hot[0] ),
    .X(_01994_));
 sg13g2_buf_1 _22015_ (.A(_01994_),
    .X(_01995_));
 sg13g2_buf_1 _22016_ (.A(net739),
    .X(_01996_));
 sg13g2_buf_1 _22017_ (.A(_01996_),
    .X(_01997_));
 sg13g2_nand2_1 _22018_ (.Y(_01998_),
    .A(net628),
    .B(net525));
 sg13g2_a21oi_1 _22019_ (.A1(_01993_),
    .A2(_01998_),
    .Y(_01556_),
    .B1(net562));
 sg13g2_nand2_1 _22020_ (.Y(_01999_),
    .A(\rbzero.wall_tracer.wall[1] ),
    .B(net547));
 sg13g2_buf_4 _22021_ (.X(_02000_),
    .A(\rbzero.wall_hot[1] ));
 sg13g2_buf_1 _22022_ (.A(_02000_),
    .X(_02001_));
 sg13g2_buf_2 _22023_ (.A(_02001_),
    .X(_02002_));
 sg13g2_buf_1 _22024_ (.A(net695),
    .X(_02003_));
 sg13g2_nand2_1 _22025_ (.Y(_02004_),
    .A(_02003_),
    .B(net525));
 sg13g2_a21oi_1 _22026_ (.A1(_01999_),
    .A2(_02004_),
    .Y(_01557_),
    .B1(net562));
 sg13g2_buf_2 _22027_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[10] ),
    .X(_02005_));
 sg13g2_inv_1 _22028_ (.Y(_02006_),
    .A(_02005_));
 sg13g2_buf_1 _22029_ (.A(_02006_),
    .X(_02007_));
 sg13g2_buf_1 _22030_ (.A(net694),
    .X(_02008_));
 sg13g2_buf_2 _22031_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-2] ),
    .X(_02009_));
 sg13g2_inv_2 _22032_ (.Y(_02010_),
    .A(_02009_));
 sg13g2_nor2_1 _22033_ (.A(_02008_),
    .B(_02010_),
    .Y(_02011_));
 sg13g2_buf_2 _22034_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-3] ),
    .X(_02012_));
 sg13g2_buf_1 _22035_ (.A(_02012_),
    .X(_02013_));
 sg13g2_buf_8 _22036_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-10] ),
    .X(_02014_));
 sg13g2_buf_8 _22037_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-9] ),
    .X(_02015_));
 sg13g2_buf_2 _22038_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-8] ),
    .X(_02016_));
 sg13g2_nor4_1 _22039_ (.A(_02014_),
    .B(\rbzero.wall_tracer.rcp_fsm.operand[-11] ),
    .C(_02015_),
    .D(_02016_),
    .Y(_02017_));
 sg13g2_buf_1 _22040_ (.A(_02017_),
    .X(_02018_));
 sg13g2_buf_1 _22041_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-7] ),
    .X(_02019_));
 sg13g2_buf_1 _22042_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-6] ),
    .X(_02020_));
 sg13g2_buf_8 _22043_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-5] ),
    .X(_02021_));
 sg13g2_nor4_1 _22044_ (.A(_02019_),
    .B(_02020_),
    .C(_02021_),
    .D(\rbzero.wall_tracer.rcp_fsm.operand[-4] ),
    .Y(_02022_));
 sg13g2_buf_1 _22045_ (.A(_02022_),
    .X(_02023_));
 sg13g2_and2_1 _22046_ (.A(net693),
    .B(net692),
    .X(_02024_));
 sg13g2_buf_2 _22047_ (.A(_02024_),
    .X(_02025_));
 sg13g2_xnor2_1 _22048_ (.Y(_02026_),
    .A(net737),
    .B(_02025_));
 sg13g2_buf_1 _22049_ (.A(_02005_),
    .X(_02027_));
 sg13g2_buf_1 _22050_ (.A(net736),
    .X(_02028_));
 sg13g2_buf_1 _22051_ (.A(net691),
    .X(_02029_));
 sg13g2_nor2_1 _22052_ (.A(net625),
    .B(_02009_),
    .Y(_02030_));
 sg13g2_buf_8 _22053_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-4] ),
    .X(_02031_));
 sg13g2_inv_2 _22054_ (.Y(_02032_),
    .A(_02012_));
 sg13g2_nand2_1 _22055_ (.Y(_02033_),
    .A(net807),
    .B(_02032_));
 sg13g2_a22oi_1 _22056_ (.Y(_02034_),
    .B1(_02030_),
    .B2(_02033_),
    .A2(_02026_),
    .A1(_02011_));
 sg13g2_buf_1 _22057_ (.A(_02020_),
    .X(_02035_));
 sg13g2_or3_1 _22058_ (.A(_02019_),
    .B(_02035_),
    .C(net808),
    .X(_02036_));
 sg13g2_buf_2 _22059_ (.A(_00474_),
    .X(_02037_));
 sg13g2_nand2b_1 _22060_ (.Y(_02038_),
    .B(_02037_),
    .A_N(_02014_));
 sg13g2_nor4_1 _22061_ (.A(_02015_),
    .B(_02016_),
    .C(_02036_),
    .D(_02038_),
    .Y(_02039_));
 sg13g2_buf_2 _22062_ (.A(_02039_),
    .X(_02040_));
 sg13g2_o21ai_1 _22063_ (.B1(net807),
    .Y(_02041_),
    .A1(net626),
    .A2(_02040_));
 sg13g2_buf_1 _22064_ (.A(_02041_),
    .X(_02042_));
 sg13g2_or3_1 _22065_ (.A(net626),
    .B(net807),
    .C(_02040_),
    .X(_02043_));
 sg13g2_buf_1 _22066_ (.A(_02043_),
    .X(_02044_));
 sg13g2_nand2_1 _22067_ (.Y(_02045_),
    .A(_02005_),
    .B(net737));
 sg13g2_buf_1 _22068_ (.A(net693),
    .X(_02046_));
 sg13g2_nand4_1 _22069_ (.B(_02010_),
    .C(_02046_),
    .A(_02032_),
    .Y(_02047_),
    .D(net692));
 sg13g2_buf_1 _22070_ (.A(_02047_),
    .X(_02048_));
 sg13g2_o21ai_1 _22071_ (.B1(_02048_),
    .Y(_02049_),
    .A1(_02010_),
    .A2(_02045_));
 sg13g2_nand3_1 _22072_ (.B(_02044_),
    .C(_02049_),
    .A(_02042_),
    .Y(_02050_));
 sg13g2_buf_1 _22073_ (.A(_02050_),
    .X(_02051_));
 sg13g2_and3_1 _22074_ (.X(_02052_),
    .A(net736),
    .B(net807),
    .C(net737));
 sg13g2_nor3_1 _22075_ (.A(net807),
    .B(net693),
    .C(_02045_),
    .Y(_02053_));
 sg13g2_mux2_1 _22076_ (.A0(_02052_),
    .A1(_02053_),
    .S(_02040_),
    .X(_02054_));
 sg13g2_nor2_1 _22077_ (.A(_02015_),
    .B(_02016_),
    .Y(_02055_));
 sg13g2_buf_1 _22078_ (.A(_02055_),
    .X(_02056_));
 sg13g2_nor3_1 _22079_ (.A(_02019_),
    .B(_02020_),
    .C(net808),
    .Y(_02057_));
 sg13g2_buf_2 _22080_ (.A(_02057_),
    .X(_02058_));
 sg13g2_nor2b_1 _22081_ (.A(_02014_),
    .B_N(_02037_),
    .Y(_02059_));
 sg13g2_buf_2 _22082_ (.A(_02059_),
    .X(_02060_));
 sg13g2_nand4_1 _22083_ (.B(net693),
    .C(_02058_),
    .A(_02056_),
    .Y(_02061_),
    .D(_02060_));
 sg13g2_or2_1 _22084_ (.X(_02062_),
    .B(_02013_),
    .A(net807));
 sg13g2_a21oi_1 _22085_ (.A1(net736),
    .A2(_02061_),
    .Y(_02063_),
    .B1(_02062_));
 sg13g2_buf_1 _22086_ (.A(_02019_),
    .X(_02064_));
 sg13g2_nor2_1 _22087_ (.A(net734),
    .B(net735),
    .Y(_02065_));
 sg13g2_a21o_1 _22088_ (.A2(_02065_),
    .A1(net624),
    .B1(net694),
    .X(_02066_));
 sg13g2_xnor2_1 _22089_ (.Y(_02067_),
    .A(net808),
    .B(_02066_));
 sg13g2_o21ai_1 _22090_ (.B1(_02067_),
    .Y(_02068_),
    .A1(_02054_),
    .A2(_02063_));
 sg13g2_buf_1 _22091_ (.A(net625),
    .X(_02069_));
 sg13g2_a21oi_1 _22092_ (.A1(_02032_),
    .A2(_02068_),
    .Y(_02070_),
    .B1(_02069_));
 sg13g2_nor2_1 _22093_ (.A(_02032_),
    .B(_02025_),
    .Y(_02071_));
 sg13g2_nand3_1 _22094_ (.B(net693),
    .C(net692),
    .A(_02032_),
    .Y(_02072_));
 sg13g2_buf_2 _22095_ (.A(_02072_),
    .X(_02073_));
 sg13g2_nand2_1 _22096_ (.Y(_02074_),
    .A(_02011_),
    .B(_02073_));
 sg13g2_a21oi_1 _22097_ (.A1(_02071_),
    .A2(_02068_),
    .Y(_02075_),
    .B1(_02074_));
 sg13g2_a221oi_1 _22098_ (.B2(_02010_),
    .C1(_02075_),
    .B1(_02070_),
    .A1(_02034_),
    .Y(_02076_),
    .A2(_02051_));
 sg13g2_buf_1 _22099_ (.A(_02076_),
    .X(_02077_));
 sg13g2_nand3_1 _22100_ (.B(_02031_),
    .C(_02013_),
    .A(net625),
    .Y(_02078_));
 sg13g2_or3_1 _22101_ (.A(_02031_),
    .B(_02046_),
    .C(_02045_),
    .X(_02079_));
 sg13g2_mux2_1 _22102_ (.A0(_02078_),
    .A1(_02079_),
    .S(_02040_),
    .X(_02080_));
 sg13g2_a21o_1 _22103_ (.A2(_02061_),
    .A1(net625),
    .B1(_02062_),
    .X(_02081_));
 sg13g2_nor2_1 _22104_ (.A(_02006_),
    .B(_02009_),
    .Y(_02082_));
 sg13g2_a21oi_1 _22105_ (.A1(net625),
    .A2(_02073_),
    .Y(_02083_),
    .B1(_02010_));
 sg13g2_a221oi_1 _22106_ (.B2(_02073_),
    .C1(_02083_),
    .B1(_02082_),
    .A1(_02080_),
    .Y(_02084_),
    .A2(_02081_));
 sg13g2_o21ai_1 _22107_ (.B1(net736),
    .Y(_02085_),
    .A1(_02015_),
    .A2(_02038_));
 sg13g2_xor2_1 _22108_ (.B(_02085_),
    .A(_02016_),
    .X(_02086_));
 sg13g2_buf_2 _22109_ (.A(_02086_),
    .X(_02087_));
 sg13g2_buf_1 _22110_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-11] ),
    .X(_02088_));
 sg13g2_o21ai_1 _22111_ (.B1(_02027_),
    .Y(_02089_),
    .A1(_02014_),
    .A2(net806));
 sg13g2_xor2_1 _22112_ (.B(_02089_),
    .A(_02015_),
    .X(_02090_));
 sg13g2_xnor2_1 _22113_ (.Y(_02091_),
    .A(_02014_),
    .B(net806));
 sg13g2_nor2b_1 _22114_ (.A(net691),
    .B_N(_00472_),
    .Y(_02092_));
 sg13g2_a21oi_1 _22115_ (.A1(net625),
    .A2(_02091_),
    .Y(_02093_),
    .B1(_02092_));
 sg13g2_buf_1 _22116_ (.A(_02093_),
    .X(_02094_));
 sg13g2_nand2_1 _22117_ (.Y(_02095_),
    .A(_02090_),
    .B(_02094_));
 sg13g2_a21o_1 _22118_ (.A2(net624),
    .A1(_02037_),
    .B1(net694),
    .X(_02096_));
 sg13g2_inv_1 _22119_ (.Y(_02097_),
    .A(net735));
 sg13g2_inv_1 _22120_ (.Y(_02098_),
    .A(net808));
 sg13g2_nor3_1 _22121_ (.A(net694),
    .B(_02097_),
    .C(_02098_),
    .Y(_02099_));
 sg13g2_nor2_1 _22122_ (.A(_02037_),
    .B(net734),
    .Y(_02100_));
 sg13g2_mux2_1 _22123_ (.A0(net734),
    .A1(_02100_),
    .S(net624),
    .X(_02101_));
 sg13g2_a22oi_1 _22124_ (.Y(_02102_),
    .B1(_02099_),
    .B2(_02101_),
    .A2(_02096_),
    .A1(_02058_));
 sg13g2_buf_1 _22125_ (.A(_02102_),
    .X(_02103_));
 sg13g2_a21oi_1 _22126_ (.A1(_02087_),
    .A2(_02095_),
    .Y(_02104_),
    .B1(_02103_));
 sg13g2_a21oi_1 _22127_ (.A1(net690),
    .A2(_02060_),
    .Y(_02105_),
    .B1(net624));
 sg13g2_nor2_1 _22128_ (.A(net735),
    .B(_02098_),
    .Y(_02106_));
 sg13g2_o21ai_1 _22129_ (.B1(_02106_),
    .Y(_02107_),
    .A1(net734),
    .A2(_02105_));
 sg13g2_nand4_1 _22130_ (.B(net808),
    .C(net690),
    .A(net735),
    .Y(_02108_),
    .D(_02060_));
 sg13g2_nor2_1 _22131_ (.A(_02014_),
    .B(net806),
    .Y(_02109_));
 sg13g2_nor2_1 _22132_ (.A(net735),
    .B(net808),
    .Y(_02110_));
 sg13g2_nand4_1 _22133_ (.B(net690),
    .C(_02110_),
    .A(_02109_),
    .Y(_02111_),
    .D(_02038_));
 sg13g2_a21o_1 _22134_ (.A2(_02111_),
    .A1(_02108_),
    .B1(_02064_),
    .X(_02112_));
 sg13g2_a21oi_1 _22135_ (.A1(_02107_),
    .A2(_02112_),
    .Y(_02113_),
    .B1(net626));
 sg13g2_nor3_1 _22136_ (.A(net561),
    .B(_02097_),
    .C(net808),
    .Y(_02114_));
 sg13g2_or3_1 _22137_ (.A(_02104_),
    .B(_02113_),
    .C(_02114_),
    .X(_02115_));
 sg13g2_nor2_1 _22138_ (.A(net737),
    .B(_02010_),
    .Y(_02116_));
 sg13g2_nor2_1 _22139_ (.A(net736),
    .B(_02010_),
    .Y(_02117_));
 sg13g2_a221oi_1 _22140_ (.B2(_02073_),
    .C1(_02117_),
    .B1(_02082_),
    .A1(_02025_),
    .Y(_02118_),
    .A2(_02116_));
 sg13g2_buf_2 _22141_ (.A(_02118_),
    .X(_02119_));
 sg13g2_o21ai_1 _22142_ (.B1(_02119_),
    .Y(_02120_),
    .A1(_02054_),
    .A2(_02063_));
 sg13g2_buf_1 _22143_ (.A(_02120_),
    .X(_02121_));
 sg13g2_nand3b_1 _22144_ (.B(_02087_),
    .C(_02090_),
    .Y(_02122_),
    .A_N(_02103_));
 sg13g2_nor2_1 _22145_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sg13g2_nand2b_1 _22146_ (.Y(_02124_),
    .B(_02014_),
    .A_N(net806));
 sg13g2_nand2_1 _22147_ (.Y(_02125_),
    .A(net806),
    .B(_02094_));
 sg13g2_and2_1 _22148_ (.A(_02124_),
    .B(_02125_),
    .X(_02126_));
 sg13g2_nor3_1 _22149_ (.A(net691),
    .B(net735),
    .C(net808),
    .Y(_02127_));
 sg13g2_a21o_1 _22150_ (.A2(_02099_),
    .A1(net624),
    .B1(_02127_),
    .X(_02128_));
 sg13g2_nand2_1 _22151_ (.Y(_02129_),
    .A(net690),
    .B(_02060_));
 sg13g2_xnor2_1 _22152_ (.Y(_02130_),
    .A(net735),
    .B(_02129_));
 sg13g2_nor4_1 _22153_ (.A(net626),
    .B(net734),
    .C(_02098_),
    .D(net624),
    .Y(_02131_));
 sg13g2_a22oi_1 _22154_ (.Y(_02132_),
    .B1(_02130_),
    .B2(_02131_),
    .A2(_02128_),
    .A1(net734));
 sg13g2_xnor2_1 _22155_ (.Y(_02133_),
    .A(_02015_),
    .B(_02089_));
 sg13g2_buf_2 _22156_ (.A(_02133_),
    .X(_02134_));
 sg13g2_nand3b_1 _22157_ (.B(_02087_),
    .C(_02134_),
    .Y(_02135_),
    .A_N(_02103_));
 sg13g2_a21oi_1 _22158_ (.A1(_02132_),
    .A2(_02135_),
    .Y(_02136_),
    .B1(_02121_));
 sg13g2_a221oi_1 _22159_ (.B2(_02126_),
    .C1(_02136_),
    .B1(_02123_),
    .A1(_02084_),
    .Y(_02137_),
    .A2(_02115_));
 sg13g2_buf_1 _22160_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[3] ),
    .X(_02138_));
 sg13g2_buf_1 _22161_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[-1] ),
    .X(_02139_));
 sg13g2_buf_1 _22162_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[0] ),
    .X(_02140_));
 sg13g2_nor4_1 _22163_ (.A(_02012_),
    .B(_02009_),
    .C(net804),
    .D(net803),
    .Y(_02141_));
 sg13g2_buf_2 _22164_ (.A(_02141_),
    .X(_02142_));
 sg13g2_buf_2 _22165_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[1] ),
    .X(_02143_));
 sg13g2_buf_2 _22166_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[2] ),
    .X(_02144_));
 sg13g2_nor2_1 _22167_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sg13g2_and3_1 _22168_ (.X(_02146_),
    .A(net805),
    .B(_02142_),
    .C(_02145_));
 sg13g2_nor2_1 _22169_ (.A(_02006_),
    .B(net805),
    .Y(_02147_));
 sg13g2_nand4_1 _22170_ (.B(net692),
    .C(_02142_),
    .A(net693),
    .Y(_02148_),
    .D(_02145_));
 sg13g2_buf_2 _22171_ (.A(_02148_),
    .X(_02149_));
 sg13g2_nor2b_1 _22172_ (.A(net736),
    .B_N(net805),
    .Y(_02150_));
 sg13g2_a221oi_1 _22173_ (.B2(_02149_),
    .C1(_02150_),
    .B1(_02147_),
    .A1(_02025_),
    .Y(_02151_),
    .A2(_02146_));
 sg13g2_buf_2 _22174_ (.A(_02151_),
    .X(_02152_));
 sg13g2_nor4_2 _22175_ (.A(net807),
    .B(_02012_),
    .C(_02009_),
    .Y(_02153_),
    .D(net804));
 sg13g2_and3_1 _22176_ (.X(_02154_),
    .A(net690),
    .B(_02060_),
    .C(_02153_));
 sg13g2_buf_1 _22177_ (.A(_02154_),
    .X(_02155_));
 sg13g2_nor2_1 _22178_ (.A(net803),
    .B(_02143_),
    .Y(_02156_));
 sg13g2_and3_1 _22179_ (.X(_02157_),
    .A(_02144_),
    .B(_02058_),
    .C(_02156_));
 sg13g2_a22oi_1 _22180_ (.Y(_02158_),
    .B1(_02155_),
    .B2(_02157_),
    .A2(_02144_),
    .A1(net694));
 sg13g2_buf_1 _22181_ (.A(_02158_),
    .X(_02159_));
 sg13g2_nand3_1 _22182_ (.B(_02060_),
    .C(_02153_),
    .A(net690),
    .Y(_02160_));
 sg13g2_buf_1 _22183_ (.A(_02160_),
    .X(_02161_));
 sg13g2_nand2_1 _22184_ (.Y(_02162_),
    .A(_02058_),
    .B(_02156_));
 sg13g2_nor2_1 _22185_ (.A(_02007_),
    .B(_02144_),
    .Y(_02163_));
 sg13g2_o21ai_1 _22186_ (.B1(_02163_),
    .Y(_02164_),
    .A1(_02161_),
    .A2(_02162_));
 sg13g2_buf_1 _22187_ (.A(_02164_),
    .X(_02165_));
 sg13g2_nand3_1 _22188_ (.B(_02159_),
    .C(_02165_),
    .A(_02152_),
    .Y(_02166_));
 sg13g2_buf_1 _22189_ (.A(_02166_),
    .X(_02167_));
 sg13g2_nand2_1 _22190_ (.Y(_02168_),
    .A(net693),
    .B(net692));
 sg13g2_or2_1 _22191_ (.X(_02169_),
    .B(_02009_),
    .A(_02012_));
 sg13g2_buf_1 _22192_ (.A(_02169_),
    .X(_02170_));
 sg13g2_buf_1 _22193_ (.A(_02143_),
    .X(_02171_));
 sg13g2_and2_1 _22194_ (.A(_02005_),
    .B(net733),
    .X(_02172_));
 sg13g2_a21oi_1 _22195_ (.A1(net803),
    .A2(_02172_),
    .Y(_02173_),
    .B1(_02156_));
 sg13g2_nor4_1 _22196_ (.A(net804),
    .B(_02168_),
    .C(_02170_),
    .D(_02173_),
    .Y(_02174_));
 sg13g2_nand2_1 _22197_ (.Y(_02175_),
    .A(net804),
    .B(_02172_));
 sg13g2_inv_1 _22198_ (.Y(_02176_),
    .A(net804));
 sg13g2_nor2_1 _22199_ (.A(_02005_),
    .B(net733),
    .Y(_02177_));
 sg13g2_and3_1 _22200_ (.X(_02178_),
    .A(net736),
    .B(net804),
    .C(net733));
 sg13g2_a22oi_1 _22201_ (.Y(_02179_),
    .B1(_02178_),
    .B2(_02170_),
    .A2(_02177_),
    .A1(_02176_));
 sg13g2_o21ai_1 _22202_ (.B1(_02179_),
    .Y(_02180_),
    .A1(_02025_),
    .A2(_02175_));
 sg13g2_and2_1 _22203_ (.A(net803),
    .B(_02153_),
    .X(_02181_));
 sg13g2_nor2_1 _22204_ (.A(_02006_),
    .B(net803),
    .Y(_02182_));
 sg13g2_nand4_1 _22205_ (.B(_02058_),
    .C(_02060_),
    .A(net690),
    .Y(_02183_),
    .D(_02153_));
 sg13g2_buf_1 _22206_ (.A(_02183_),
    .X(_02184_));
 sg13g2_nor2b_1 _22207_ (.A(_02005_),
    .B_N(net803),
    .Y(_02185_));
 sg13g2_a221oi_1 _22208_ (.B2(_02184_),
    .C1(_02185_),
    .B1(_02182_),
    .A1(_02040_),
    .Y(_02186_),
    .A2(_02181_));
 sg13g2_buf_1 _22209_ (.A(_02186_),
    .X(_02187_));
 sg13g2_o21ai_1 _22210_ (.B1(net497),
    .Y(_02188_),
    .A1(_02174_),
    .A2(_02180_));
 sg13g2_buf_1 _22211_ (.A(_02188_),
    .X(_02189_));
 sg13g2_nor2_1 _22212_ (.A(_02167_),
    .B(_02189_),
    .Y(_02190_));
 sg13g2_buf_1 _22213_ (.A(_02190_),
    .X(_02191_));
 sg13g2_nor4_1 _22214_ (.A(net803),
    .B(net733),
    .C(_02144_),
    .D(net805),
    .Y(_02192_));
 sg13g2_nand2_1 _22215_ (.Y(_02193_),
    .A(_02058_),
    .B(_02192_));
 sg13g2_or2_1 _22216_ (.X(_02194_),
    .B(_02193_),
    .A(_02161_));
 sg13g2_buf_2 _22217_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[4] ),
    .X(_02195_));
 sg13g2_nor2_1 _22218_ (.A(net626),
    .B(_02195_),
    .Y(_02196_));
 sg13g2_buf_1 _22219_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[5] ),
    .X(_02197_));
 sg13g2_buf_1 _22220_ (.A(_02197_),
    .X(_02198_));
 sg13g2_buf_1 _22221_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[6] ),
    .X(_02199_));
 sg13g2_nor2_1 _22222_ (.A(net732),
    .B(net802),
    .Y(_02200_));
 sg13g2_and3_1 _22223_ (.X(_02201_),
    .A(net693),
    .B(net692),
    .C(_02142_));
 sg13g2_buf_1 _22224_ (.A(_02201_),
    .X(_02202_));
 sg13g2_nor4_2 _22225_ (.A(net805),
    .B(_02195_),
    .C(_02197_),
    .Y(_02203_),
    .D(net802));
 sg13g2_and2_1 _22226_ (.A(_02145_),
    .B(_02203_),
    .X(_02204_));
 sg13g2_buf_1 _22227_ (.A(_02204_),
    .X(_02205_));
 sg13g2_a22oi_1 _22228_ (.Y(_02206_),
    .B1(_02202_),
    .B2(_02205_),
    .A2(_02200_),
    .A1(net694));
 sg13g2_buf_1 _22229_ (.A(_02206_),
    .X(_02207_));
 sg13g2_nor4_1 _22230_ (.A(_02143_),
    .B(_02144_),
    .C(net805),
    .D(_02195_),
    .Y(_02208_));
 sg13g2_nand4_1 _22231_ (.B(net692),
    .C(_02142_),
    .A(_02018_),
    .Y(_02209_),
    .D(_02208_));
 sg13g2_buf_2 _22232_ (.A(_02209_),
    .X(_02210_));
 sg13g2_nand4_1 _22233_ (.B(net732),
    .C(net802),
    .A(_02027_),
    .Y(_02211_),
    .D(_02210_));
 sg13g2_buf_1 _22234_ (.A(_02211_),
    .X(_02212_));
 sg13g2_and4_1 _22235_ (.A(_02098_),
    .B(_02195_),
    .C(_02065_),
    .D(_02192_),
    .X(_02213_));
 sg13g2_nor2b_1 _22236_ (.A(net691),
    .B_N(_02195_),
    .Y(_02214_));
 sg13g2_a21o_1 _22237_ (.A2(_02213_),
    .A1(_02155_),
    .B1(_02214_),
    .X(_02215_));
 sg13g2_a221oi_1 _22238_ (.B2(_02212_),
    .C1(_02215_),
    .B1(_02207_),
    .A1(_02194_),
    .Y(_02216_),
    .A2(_02196_));
 sg13g2_buf_1 _22239_ (.A(_02216_),
    .X(_02217_));
 sg13g2_buf_1 _22240_ (.A(_02217_),
    .X(_02218_));
 sg13g2_buf_2 _22241_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[7] ),
    .X(_02219_));
 sg13g2_buf_1 _22242_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[8] ),
    .X(_02220_));
 sg13g2_or2_1 _22243_ (.X(_02221_),
    .B(_02220_),
    .A(_02219_));
 sg13g2_buf_1 _22244_ (.A(_02221_),
    .X(_02222_));
 sg13g2_nor2_1 _22245_ (.A(net691),
    .B(_02222_),
    .Y(_02223_));
 sg13g2_nand3_1 _22246_ (.B(_02219_),
    .C(_02220_),
    .A(_02028_),
    .Y(_02224_));
 sg13g2_a21oi_1 _22247_ (.A1(_02202_),
    .A2(_02205_),
    .Y(_02225_),
    .B1(_02224_));
 sg13g2_nor2_1 _22248_ (.A(_02223_),
    .B(_02225_),
    .Y(_02226_));
 sg13g2_nor2_1 _22249_ (.A(_02007_),
    .B(_02219_),
    .Y(_02227_));
 sg13g2_nand4_1 _22250_ (.B(_02202_),
    .C(_02205_),
    .A(_02220_),
    .Y(_02228_),
    .D(_02227_));
 sg13g2_nand2b_1 _22251_ (.Y(_02229_),
    .B(_02203_),
    .A_N(_02222_));
 sg13g2_or2_1 _22252_ (.X(_02230_),
    .B(_02229_),
    .A(_02149_));
 sg13g2_buf_2 _22253_ (.A(_02230_),
    .X(_02231_));
 sg13g2_nor3_1 _22254_ (.A(net803),
    .B(_02143_),
    .C(_02144_),
    .Y(_02232_));
 sg13g2_nand3b_1 _22255_ (.B(_02203_),
    .C(_02232_),
    .Y(_02233_),
    .A_N(_02219_));
 sg13g2_nor2_1 _22256_ (.A(_02184_),
    .B(_02233_),
    .Y(_02234_));
 sg13g2_mux2_1 _22257_ (.A0(_02228_),
    .A1(_02231_),
    .S(_02234_),
    .X(_02235_));
 sg13g2_buf_1 _22258_ (.A(\rbzero.wall_tracer.rcp_fsm.operand[9] ),
    .X(_02236_));
 sg13g2_or4_1 _22259_ (.A(net805),
    .B(_02195_),
    .C(_02197_),
    .D(net802),
    .X(_02237_));
 sg13g2_nand4_1 _22260_ (.B(_02060_),
    .C(_02153_),
    .A(net690),
    .Y(_02238_),
    .D(_02232_));
 sg13g2_nor4_1 _22261_ (.A(_00473_),
    .B(_02036_),
    .C(_02237_),
    .D(_02238_),
    .Y(_02239_));
 sg13g2_or3_1 _22262_ (.A(_02236_),
    .B(_02231_),
    .C(_02239_),
    .X(_02240_));
 sg13g2_inv_1 _22263_ (.Y(_02241_),
    .A(_02236_));
 sg13g2_nor2_1 _22264_ (.A(net694),
    .B(_02241_),
    .Y(_02242_));
 sg13g2_nor2_1 _22265_ (.A(net691),
    .B(_02236_),
    .Y(_02243_));
 sg13g2_nand2_1 _22266_ (.Y(_02244_),
    .A(_02058_),
    .B(_02203_));
 sg13g2_or4_1 _22267_ (.A(_00473_),
    .B(_02222_),
    .C(_02238_),
    .D(_02244_),
    .X(_02245_));
 sg13g2_a22oi_1 _22268_ (.Y(_02246_),
    .B1(_02243_),
    .B2(_02245_),
    .A2(_02242_),
    .A1(_02231_));
 sg13g2_a22oi_1 _22269_ (.Y(_02247_),
    .B1(_02240_),
    .B2(_02246_),
    .A2(_02235_),
    .A1(_02226_));
 sg13g2_buf_1 _22270_ (.A(_02247_),
    .X(_02248_));
 sg13g2_buf_8 _22271_ (.A(_02248_),
    .X(_02249_));
 sg13g2_nand3_1 _22272_ (.B(net465),
    .C(net453),
    .A(_02191_),
    .Y(_02250_));
 sg13g2_buf_2 _22273_ (.A(_02250_),
    .X(_02251_));
 sg13g2_a21oi_1 _22274_ (.A1(_02077_),
    .A2(_02137_),
    .Y(_02252_),
    .B1(_02251_));
 sg13g2_buf_1 _22275_ (.A(_02252_),
    .X(_02253_));
 sg13g2_buf_1 _22276_ (.A(_02253_),
    .X(_02254_));
 sg13g2_nand2_1 _22277_ (.Y(_02255_),
    .A(_02159_),
    .B(_02165_));
 sg13g2_or2_1 _22278_ (.X(_02256_),
    .B(_02189_),
    .A(_02255_));
 sg13g2_nand4_1 _22279_ (.B(net465),
    .C(net453),
    .A(_02152_),
    .Y(_02257_),
    .D(_02256_));
 sg13g2_buf_1 _22280_ (.A(_02257_),
    .X(_02258_));
 sg13g2_o21ai_1 _22281_ (.B1(_02258_),
    .Y(_02259_),
    .A1(_02251_),
    .A2(_02077_));
 sg13g2_buf_2 _22282_ (.A(_02259_),
    .X(_02260_));
 sg13g2_and3_1 _22283_ (.X(_02261_),
    .A(_02191_),
    .B(_02218_),
    .C(_02248_));
 sg13g2_buf_1 _22284_ (.A(_02261_),
    .X(_02262_));
 sg13g2_a22oi_1 _22285_ (.Y(_02263_),
    .B1(_02030_),
    .B2(net737),
    .A2(_02026_),
    .A1(_02011_));
 sg13g2_inv_1 _22286_ (.Y(_02264_),
    .A(_02263_));
 sg13g2_or2_1 _22287_ (.X(_02265_),
    .B(_02189_),
    .A(_02167_));
 sg13g2_xnor2_1 _22288_ (.Y(_02266_),
    .A(_02016_),
    .B(_02085_));
 sg13g2_nor2_1 _22289_ (.A(_02124_),
    .B(_02094_),
    .Y(_02267_));
 sg13g2_nor4_1 _22290_ (.A(_02103_),
    .B(_02266_),
    .C(_02134_),
    .D(_02267_),
    .Y(_02268_));
 sg13g2_a22oi_1 _22291_ (.Y(_02269_),
    .B1(_02084_),
    .B2(_02268_),
    .A2(_02051_),
    .A1(_02034_));
 sg13g2_o21ai_1 _22292_ (.B1(net465),
    .Y(_02270_),
    .A1(_02265_),
    .A2(_02269_));
 sg13g2_xnor2_1 _22293_ (.Y(_02271_),
    .A(_02098_),
    .B(_02066_));
 sg13g2_buf_2 _22294_ (.A(_02271_),
    .X(_02272_));
 sg13g2_or4_1 _22295_ (.A(_02255_),
    .B(_02189_),
    .C(_02272_),
    .D(_02121_),
    .X(_02273_));
 sg13g2_nor3_1 _22296_ (.A(_02236_),
    .B(_02231_),
    .C(_02239_),
    .Y(_02274_));
 sg13g2_nand2_1 _22297_ (.Y(_02275_),
    .A(net626),
    .B(_02241_));
 sg13g2_nor4_1 _22298_ (.A(_00473_),
    .B(_02222_),
    .C(_02238_),
    .D(_02244_),
    .Y(_02276_));
 sg13g2_o21ai_1 _22299_ (.B1(_02242_),
    .Y(_02277_),
    .A1(_02149_),
    .A2(_02229_));
 sg13g2_o21ai_1 _22300_ (.B1(_02277_),
    .Y(_02278_),
    .A1(_02275_),
    .A2(_02276_));
 sg13g2_o21ai_1 _22301_ (.B1(_02217_),
    .Y(_02279_),
    .A1(_02274_),
    .A2(_02278_));
 sg13g2_a221oi_1 _22302_ (.B2(_02152_),
    .C1(_02279_),
    .B1(_02273_),
    .A1(_02226_),
    .Y(_02280_),
    .A2(_02235_));
 sg13g2_buf_1 _22303_ (.A(_02280_),
    .X(_02281_));
 sg13g2_buf_8 _22304_ (.A(_02281_),
    .X(_02282_));
 sg13g2_a221oi_1 _22305_ (.B2(net453),
    .C1(net403),
    .B1(_02270_),
    .A1(_02262_),
    .Y(_02283_),
    .A2(_02264_));
 sg13g2_buf_2 _22306_ (.A(_02283_),
    .X(_02284_));
 sg13g2_nor2_1 _22307_ (.A(_02260_),
    .B(_02284_),
    .Y(_02285_));
 sg13g2_buf_2 _22308_ (.A(_02285_),
    .X(_02286_));
 sg13g2_nand2_1 _22309_ (.Y(_02287_),
    .A(_02069_),
    .B(_02231_));
 sg13g2_xnor2_1 _22310_ (.Y(_02288_),
    .A(_02241_),
    .B(_02287_));
 sg13g2_o21ai_1 _22311_ (.B1(net625),
    .Y(_02289_),
    .A1(_02149_),
    .A2(_02237_));
 sg13g2_xor2_1 _22312_ (.B(_02289_),
    .A(_02219_),
    .X(_02290_));
 sg13g2_xor2_1 _22313_ (.B(_02210_),
    .A(net732),
    .X(_02291_));
 sg13g2_inv_1 _22314_ (.Y(_02292_),
    .A(net802));
 sg13g2_nor2_1 _22315_ (.A(_02008_),
    .B(_02292_),
    .Y(_02293_));
 sg13g2_nor2_1 _22316_ (.A(_02029_),
    .B(net802),
    .Y(_02294_));
 sg13g2_a22oi_1 _22317_ (.Y(_02295_),
    .B1(_02294_),
    .B2(net732),
    .A2(_02293_),
    .A1(_02291_));
 sg13g2_o21ai_1 _22318_ (.B1(_02029_),
    .Y(_02296_),
    .A1(_02184_),
    .A2(_02233_));
 sg13g2_xnor2_1 _22319_ (.Y(_02297_),
    .A(_02220_),
    .B(_02296_));
 sg13g2_a21o_1 _22320_ (.A2(_02295_),
    .A1(_02290_),
    .B1(_02297_),
    .X(_02298_));
 sg13g2_a22oi_1 _22321_ (.Y(_02299_),
    .B1(_02288_),
    .B2(_02298_),
    .A2(_02276_),
    .A1(_02241_));
 sg13g2_a21o_1 _22322_ (.A2(_02091_),
    .A1(net625),
    .B1(_02092_),
    .X(_02300_));
 sg13g2_buf_1 _22323_ (.A(_02300_),
    .X(_02301_));
 sg13g2_and2_1 _22324_ (.A(net806),
    .B(_02301_),
    .X(_02302_));
 sg13g2_nor4_1 _22325_ (.A(_02167_),
    .B(_02189_),
    .C(_02121_),
    .D(_02122_),
    .Y(_02303_));
 sg13g2_and4_1 _22326_ (.A(net465),
    .B(net453),
    .C(_02302_),
    .D(_02303_),
    .X(_02304_));
 sg13g2_buf_1 _22327_ (.A(_02304_),
    .X(_02305_));
 sg13g2_nor2_1 _22328_ (.A(_02299_),
    .B(_02305_),
    .Y(_02306_));
 sg13g2_buf_8 _22329_ (.A(_02306_),
    .X(_02307_));
 sg13g2_and4_1 _22330_ (.A(_02191_),
    .B(net465),
    .C(net453),
    .D(_02136_),
    .X(_02308_));
 sg13g2_nand2_1 _22331_ (.Y(_02309_),
    .A(_02207_),
    .B(_02212_));
 sg13g2_a21oi_1 _22332_ (.A1(_02155_),
    .A2(_02213_),
    .Y(_02310_),
    .B1(_02214_));
 sg13g2_o21ai_1 _22333_ (.B1(_02196_),
    .Y(_02311_),
    .A1(_02161_),
    .A2(_02193_));
 sg13g2_buf_1 _22334_ (.A(_02311_),
    .X(_02312_));
 sg13g2_nand2_1 _22335_ (.Y(_02313_),
    .A(_02310_),
    .B(_02312_));
 sg13g2_nor2_1 _22336_ (.A(_02313_),
    .B(_02263_),
    .Y(_02314_));
 sg13g2_and4_1 _22337_ (.A(_02191_),
    .B(_02309_),
    .C(_02249_),
    .D(_02314_),
    .X(_02315_));
 sg13g2_nand2_1 _22338_ (.Y(_02316_),
    .A(_02028_),
    .B(_02149_));
 sg13g2_xnor2_1 _22339_ (.Y(_02317_),
    .A(_02138_),
    .B(_02316_));
 sg13g2_nor2_1 _22340_ (.A(_02317_),
    .B(_02255_),
    .Y(_02318_));
 sg13g2_nand2_1 _22341_ (.Y(_02319_),
    .A(net736),
    .B(net733));
 sg13g2_nor2_1 _22342_ (.A(net804),
    .B(_02319_),
    .Y(_02320_));
 sg13g2_nor3_1 _22343_ (.A(_02176_),
    .B(_02170_),
    .C(_02319_),
    .Y(_02321_));
 sg13g2_and2_1 _22344_ (.A(net804),
    .B(_02177_),
    .X(_02322_));
 sg13g2_a221oi_1 _22345_ (.B2(_02025_),
    .C1(_02322_),
    .B1(_02321_),
    .A1(_02048_),
    .Y(_02323_),
    .A2(_02320_));
 sg13g2_nand2b_1 _22346_ (.Y(_02324_),
    .B(net497),
    .A_N(_02323_));
 sg13g2_and2_1 _22347_ (.A(net733),
    .B(_02142_),
    .X(_02325_));
 sg13g2_nor2_1 _22348_ (.A(net694),
    .B(net733),
    .Y(_02326_));
 sg13g2_nand3_1 _22349_ (.B(_02023_),
    .C(_02142_),
    .A(_02018_),
    .Y(_02327_));
 sg13g2_nor2b_1 _22350_ (.A(net691),
    .B_N(_02171_),
    .Y(_02328_));
 sg13g2_a221oi_1 _22351_ (.B2(_02327_),
    .C1(_02328_),
    .B1(_02326_),
    .A1(_02025_),
    .Y(_02329_),
    .A2(_02325_));
 sg13g2_buf_2 _22352_ (.A(_02329_),
    .X(_02330_));
 sg13g2_nand2_1 _22353_ (.Y(_02331_),
    .A(_02324_),
    .B(_02330_));
 sg13g2_and4_1 _22354_ (.A(_02318_),
    .B(_02217_),
    .C(_02248_),
    .D(_02331_),
    .X(_02332_));
 sg13g2_buf_1 _22355_ (.A(_02332_),
    .X(_02333_));
 sg13g2_nor4_1 _22356_ (.A(_02308_),
    .B(_02281_),
    .C(_02315_),
    .D(_02333_),
    .Y(_02334_));
 sg13g2_buf_1 _22357_ (.A(_02334_),
    .X(_02335_));
 sg13g2_xor2_1 _22358_ (.B(_02015_),
    .A(net691),
    .X(_02336_));
 sg13g2_nor2_1 _22359_ (.A(_02109_),
    .B(_02336_),
    .Y(_02337_));
 sg13g2_a21o_1 _22360_ (.A2(_02337_),
    .A1(_02087_),
    .B1(_02103_),
    .X(_02338_));
 sg13g2_nand2_1 _22361_ (.Y(_02339_),
    .A(net737),
    .B(_02009_));
 sg13g2_a21o_1 _22362_ (.A2(net692),
    .A1(net624),
    .B1(net626),
    .X(_02340_));
 sg13g2_buf_1 _22363_ (.A(_02340_),
    .X(_02341_));
 sg13g2_mux2_1 _22364_ (.A0(_02339_),
    .A1(_02170_),
    .S(_02341_),
    .X(_02342_));
 sg13g2_a21o_1 _22365_ (.A2(_02044_),
    .A1(_02042_),
    .B1(_02342_),
    .X(_02343_));
 sg13g2_o21ai_1 _22366_ (.B1(_02343_),
    .Y(_02344_),
    .A1(_02121_),
    .A2(_02338_));
 sg13g2_nand4_1 _22367_ (.B(_02218_),
    .C(_02249_),
    .A(_02191_),
    .Y(_02345_),
    .D(_02344_));
 sg13g2_nor2b_1 _22368_ (.A(net403),
    .B_N(_02345_),
    .Y(_02346_));
 sg13g2_nand2b_1 _22369_ (.Y(_02347_),
    .B(_02330_),
    .A_N(net497));
 sg13g2_a221oi_1 _22370_ (.B2(_02347_),
    .C1(_02167_),
    .B1(_02324_),
    .A1(_02207_),
    .Y(_02348_),
    .A2(_02212_));
 sg13g2_a22oi_1 _22371_ (.Y(_02349_),
    .B1(_02207_),
    .B2(_02212_),
    .A2(_02312_),
    .A1(_02310_));
 sg13g2_a21o_1 _22372_ (.A2(_02235_),
    .A1(_02226_),
    .B1(_02349_),
    .X(_02350_));
 sg13g2_nand2_1 _22373_ (.Y(_02351_),
    .A(_02240_),
    .B(_02246_));
 sg13g2_o21ai_1 _22374_ (.B1(_02351_),
    .Y(_02352_),
    .A1(_02348_),
    .A2(_02350_));
 sg13g2_buf_2 _22375_ (.A(_02352_),
    .X(_02353_));
 sg13g2_a221oi_1 _22376_ (.B2(_02353_),
    .C1(_02260_),
    .B1(_02346_),
    .A1(_02307_),
    .Y(_02354_),
    .A2(_02335_));
 sg13g2_buf_1 _22377_ (.A(_02258_),
    .X(_02355_));
 sg13g2_nand3b_1 _22378_ (.B(_02345_),
    .C(_02353_),
    .Y(_02356_),
    .A_N(_02281_));
 sg13g2_buf_8 _22379_ (.A(_02356_),
    .X(_02357_));
 sg13g2_nor2_1 _22380_ (.A(net361),
    .B(_02357_),
    .Y(_02358_));
 sg13g2_buf_1 _22381_ (.A(_02358_),
    .X(_02359_));
 sg13g2_or2_1 _22382_ (.X(_02360_),
    .B(_02305_),
    .A(_02299_));
 sg13g2_buf_1 _22383_ (.A(_02360_),
    .X(_02361_));
 sg13g2_or4_1 _22384_ (.A(_02308_),
    .B(_02281_),
    .C(_02315_),
    .D(_02333_),
    .X(_02362_));
 sg13g2_buf_8 _22385_ (.A(_02362_),
    .X(_02363_));
 sg13g2_nor3_2 _22386_ (.A(net361),
    .B(net345),
    .C(_02363_),
    .Y(_02364_));
 sg13g2_or4_1 _22387_ (.A(_02286_),
    .B(_02354_),
    .C(net330),
    .D(_02364_),
    .X(_02365_));
 sg13g2_buf_1 _22388_ (.A(_02365_),
    .X(_02366_));
 sg13g2_buf_1 _22389_ (.A(_02366_),
    .X(_02367_));
 sg13g2_buf_8 _22390_ (.A(_02284_),
    .X(_02368_));
 sg13g2_o21ai_1 _22391_ (.B1(_02357_),
    .Y(_02369_),
    .A1(net345),
    .A2(_02363_));
 sg13g2_buf_2 _22392_ (.A(_02369_),
    .X(_02370_));
 sg13g2_a21oi_1 _22393_ (.A1(net329),
    .A2(_02370_),
    .Y(_02371_),
    .B1(net403));
 sg13g2_buf_2 _22394_ (.A(_02371_),
    .X(_02372_));
 sg13g2_buf_1 _22395_ (.A(_02372_),
    .X(_02373_));
 sg13g2_nand2_1 _22396_ (.Y(_02374_),
    .A(net346),
    .B(_02335_));
 sg13g2_buf_2 _22397_ (.A(_02374_),
    .X(_02375_));
 sg13g2_buf_8 _22398_ (.A(_02375_),
    .X(_02376_));
 sg13g2_buf_1 _22399_ (.A(net313),
    .X(_02377_));
 sg13g2_nor3_1 _22400_ (.A(_02134_),
    .B(_02124_),
    .C(_02094_),
    .Y(_02378_));
 sg13g2_nor4_1 _22401_ (.A(_02121_),
    .B(_02103_),
    .C(_02266_),
    .D(_02378_),
    .Y(_02379_));
 sg13g2_and4_1 _22402_ (.A(_02191_),
    .B(net465),
    .C(net453),
    .D(_02379_),
    .X(_02380_));
 sg13g2_buf_1 _22403_ (.A(_02380_),
    .X(_02381_));
 sg13g2_inv_1 _22404_ (.Y(_02382_),
    .A(_02381_));
 sg13g2_nor4_1 _22405_ (.A(_02286_),
    .B(_02354_),
    .C(_02359_),
    .D(_02364_),
    .Y(_02383_));
 sg13g2_buf_1 _22406_ (.A(_02383_),
    .X(_02384_));
 sg13g2_a21o_1 _22407_ (.A2(_02370_),
    .A1(net329),
    .B1(net403),
    .X(_02385_));
 sg13g2_buf_1 _22408_ (.A(_02385_),
    .X(_02386_));
 sg13g2_nor2_1 _22409_ (.A(_02361_),
    .B(_02363_),
    .Y(_02387_));
 sg13g2_buf_4 _22410_ (.X(_02388_),
    .A(_02387_));
 sg13g2_mux2_1 _22411_ (.A0(_02266_),
    .A1(_02094_),
    .S(_02357_),
    .X(_02389_));
 sg13g2_buf_8 _22412_ (.A(_02357_),
    .X(_02390_));
 sg13g2_nor2_1 _22413_ (.A(net626),
    .B(net624),
    .Y(_02391_));
 sg13g2_xnor2_1 _22414_ (.Y(_02392_),
    .A(net734),
    .B(_02391_));
 sg13g2_buf_1 _22415_ (.A(_02392_),
    .X(_02393_));
 sg13g2_nand2_1 _22416_ (.Y(_02394_),
    .A(net344),
    .B(_02393_));
 sg13g2_buf_1 _22417_ (.A(_02335_),
    .X(_02395_));
 sg13g2_or2_1 _22418_ (.X(_02396_),
    .B(_02350_),
    .A(_02348_));
 sg13g2_a221oi_1 _22419_ (.B2(_02351_),
    .C1(net403),
    .B1(_02396_),
    .A1(_02262_),
    .Y(_02397_),
    .A2(_02344_));
 sg13g2_buf_8 _22420_ (.A(_02397_),
    .X(_02398_));
 sg13g2_a22oi_1 _22421_ (.Y(_02399_),
    .B1(_02398_),
    .B2(_02090_),
    .A2(net343),
    .A1(net346));
 sg13g2_a22oi_1 _22422_ (.Y(_02400_),
    .B1(_02394_),
    .B2(_02399_),
    .A2(_02389_),
    .A1(_02388_));
 sg13g2_nand2_1 _22423_ (.Y(_02401_),
    .A(net806),
    .B(_02282_));
 sg13g2_o21ai_1 _22424_ (.B1(_02401_),
    .Y(_02402_),
    .A1(_02386_),
    .A2(_02400_));
 sg13g2_buf_2 _22425_ (.A(_02402_),
    .X(_02403_));
 sg13g2_nor2_1 _22426_ (.A(_02384_),
    .B(_02403_),
    .Y(_02404_));
 sg13g2_nor2_1 _22427_ (.A(_02382_),
    .B(_02404_),
    .Y(_02405_));
 sg13g2_buf_1 _22428_ (.A(_02405_),
    .X(_02406_));
 sg13g2_buf_1 _22429_ (.A(net254),
    .X(_02407_));
 sg13g2_nor2_1 _22430_ (.A(net305),
    .B(_02407_),
    .Y(_02408_));
 sg13g2_buf_2 _22431_ (.A(_02408_),
    .X(_02409_));
 sg13g2_nand2_1 _22432_ (.Y(_02410_),
    .A(net331),
    .B(_02383_));
 sg13g2_buf_8 _22433_ (.A(_02398_),
    .X(_02411_));
 sg13g2_mux4_1 _22434_ (.S0(_02375_),
    .A0(_02037_),
    .A1(_02087_),
    .A2(_02090_),
    .A3(_02301_),
    .S1(net328),
    .X(_02412_));
 sg13g2_buf_2 _22435_ (.A(_02412_),
    .X(_02413_));
 sg13g2_and2_1 _22436_ (.A(_02042_),
    .B(_02044_),
    .X(_02414_));
 sg13g2_buf_1 _22437_ (.A(_02414_),
    .X(_02415_));
 sg13g2_o21ai_1 _22438_ (.B1(net561),
    .Y(_02416_),
    .A1(net734),
    .A2(_02129_));
 sg13g2_xnor2_1 _22439_ (.Y(_02417_),
    .A(_02097_),
    .B(_02416_));
 sg13g2_mux4_1 _22440_ (.S0(_02388_),
    .A0(_02415_),
    .A1(_02393_),
    .A2(_02417_),
    .A3(_02272_),
    .S1(_02411_),
    .X(_02418_));
 sg13g2_mux2_1 _22441_ (.A0(_02413_),
    .A1(_02418_),
    .S(_02372_),
    .X(_02419_));
 sg13g2_nor2_1 _22442_ (.A(_02410_),
    .B(_02419_),
    .Y(_02420_));
 sg13g2_buf_1 _22443_ (.A(_02420_),
    .X(_02421_));
 sg13g2_buf_1 _22444_ (.A(_02286_),
    .X(_02422_));
 sg13g2_and2_1 _22445_ (.A(_02159_),
    .B(_02165_),
    .X(_02423_));
 sg13g2_buf_1 _22446_ (.A(_02423_),
    .X(_02424_));
 sg13g2_mux4_1 _22447_ (.S0(_02375_),
    .A0(_02152_),
    .A1(_02424_),
    .A2(_02330_),
    .A3(net497),
    .S1(_02390_),
    .X(_02425_));
 sg13g2_nand2_1 _22448_ (.Y(_02426_),
    .A(net312),
    .B(_02425_));
 sg13g2_o21ai_1 _22449_ (.B1(net561),
    .Y(_02427_),
    .A1(net732),
    .A2(_02210_));
 sg13g2_xnor2_1 _22450_ (.Y(_02428_),
    .A(net802),
    .B(_02427_));
 sg13g2_nand2_1 _22451_ (.Y(_02429_),
    .A(net561),
    .B(_02210_));
 sg13g2_xnor2_1 _22452_ (.Y(_02430_),
    .A(net732),
    .B(_02429_));
 sg13g2_xnor2_1 _22453_ (.Y(_02431_),
    .A(_02219_),
    .B(_02289_));
 sg13g2_buf_8 _22454_ (.A(_02388_),
    .X(_02432_));
 sg13g2_mux4_1 _22455_ (.S0(net328),
    .A0(_02313_),
    .A1(_02428_),
    .A2(_02430_),
    .A3(_02431_),
    .S1(_02432_),
    .X(_02433_));
 sg13g2_and4_1 _22456_ (.A(_02152_),
    .B(net465),
    .C(net453),
    .D(_02256_),
    .X(_02434_));
 sg13g2_buf_1 _22457_ (.A(_02434_),
    .X(_02435_));
 sg13g2_nor2_1 _22458_ (.A(_02435_),
    .B(_02286_),
    .Y(_02436_));
 sg13g2_buf_2 _22459_ (.A(_02436_),
    .X(_02437_));
 sg13g2_nand2b_1 _22460_ (.Y(_02438_),
    .B(_02437_),
    .A_N(_02433_));
 sg13g2_nand2_1 _22461_ (.Y(_02439_),
    .A(net561),
    .B(_02048_));
 sg13g2_xnor2_1 _22462_ (.Y(_02440_),
    .A(_02176_),
    .B(_02439_));
 sg13g2_buf_1 _22463_ (.A(_02440_),
    .X(_02441_));
 sg13g2_nand3_1 _22464_ (.B(net343),
    .C(_02441_),
    .A(net346),
    .Y(_02442_));
 sg13g2_o21ai_1 _22465_ (.B1(_02119_),
    .Y(_02443_),
    .A1(net345),
    .A2(_02363_));
 sg13g2_nand2_1 _22466_ (.Y(_02444_),
    .A(_02442_),
    .B(_02443_));
 sg13g2_nor2_2 _22467_ (.A(net361),
    .B(_02398_),
    .Y(_02445_));
 sg13g2_xnor2_1 _22468_ (.Y(_02446_),
    .A(_02032_),
    .B(_02341_));
 sg13g2_buf_1 _22469_ (.A(_02446_),
    .X(_02447_));
 sg13g2_mux2_1 _22470_ (.A0(_02415_),
    .A1(_02447_),
    .S(_02388_),
    .X(_02448_));
 sg13g2_a221oi_1 _22471_ (.B2(_02448_),
    .C1(_02253_),
    .B1(_02445_),
    .A1(net330),
    .Y(_02449_),
    .A2(_02444_));
 sg13g2_buf_1 _22472_ (.A(_02449_),
    .X(_02450_));
 sg13g2_and3_1 _22473_ (.X(_02451_),
    .A(_02426_),
    .B(_02438_),
    .C(_02450_));
 sg13g2_buf_1 _22474_ (.A(_02451_),
    .X(_02452_));
 sg13g2_nor2_1 _22475_ (.A(net287),
    .B(net286),
    .Y(_02453_));
 sg13g2_buf_2 _22476_ (.A(_02453_),
    .X(_02454_));
 sg13g2_buf_1 _22477_ (.A(_02454_),
    .X(_02455_));
 sg13g2_buf_1 _22478_ (.A(net229),
    .X(_02456_));
 sg13g2_buf_1 _22479_ (.A(net203),
    .X(_02457_));
 sg13g2_and2_1 _22480_ (.A(net361),
    .B(net329),
    .X(_02458_));
 sg13g2_buf_1 _22481_ (.A(_02458_),
    .X(_02459_));
 sg13g2_mux4_1 _22482_ (.S0(net344),
    .A0(net497),
    .A1(_02119_),
    .A2(_02441_),
    .A3(_02447_),
    .S1(net313),
    .X(_02460_));
 sg13g2_nand2_1 _22483_ (.Y(_02461_),
    .A(_02459_),
    .B(_02460_));
 sg13g2_nand2_1 _22484_ (.Y(_02462_),
    .A(_02042_),
    .B(_02044_));
 sg13g2_xnor2_1 _22485_ (.Y(_02463_),
    .A(net735),
    .B(_02416_));
 sg13g2_mux2_1 _22486_ (.A0(_02462_),
    .A1(_02463_),
    .S(_02357_),
    .X(_02464_));
 sg13g2_a22oi_1 _22487_ (.Y(_02465_),
    .B1(_02398_),
    .B2(_02272_),
    .A2(_02395_),
    .A1(net346));
 sg13g2_a22oi_1 _22488_ (.Y(_02466_),
    .B1(_02465_),
    .B2(_02394_),
    .A2(_02464_),
    .A1(_02388_));
 sg13g2_nand2_1 _22489_ (.Y(_02467_),
    .A(_02037_),
    .B(net344));
 sg13g2_a22oi_1 _22490_ (.Y(_02468_),
    .B1(_02399_),
    .B2(_02467_),
    .A2(_02389_),
    .A1(net311));
 sg13g2_buf_1 _22491_ (.A(_02435_),
    .X(_02469_));
 sg13g2_a221oi_1 _22492_ (.B2(net360),
    .C1(net331),
    .B1(_02468_),
    .A1(_02286_),
    .Y(_02470_),
    .A2(_02466_));
 sg13g2_buf_1 _22493_ (.A(_02470_),
    .X(_02471_));
 sg13g2_nand2_1 _22494_ (.Y(_02472_),
    .A(_02461_),
    .B(_02471_));
 sg13g2_and2_1 _22495_ (.A(_02310_),
    .B(_02312_),
    .X(_02473_));
 sg13g2_buf_1 _22496_ (.A(_02473_),
    .X(_02474_));
 sg13g2_xor2_1 _22497_ (.B(_02429_),
    .A(net732),
    .X(_02475_));
 sg13g2_mux4_1 _22498_ (.S0(_02388_),
    .A0(_02474_),
    .A1(_02475_),
    .A2(_02187_),
    .A3(_02330_),
    .S1(net329),
    .X(_02476_));
 sg13g2_nor2_1 _22499_ (.A(_02251_),
    .B(_02077_),
    .Y(_02477_));
 sg13g2_o21ai_1 _22500_ (.B1(net361),
    .Y(_02478_),
    .A1(_02477_),
    .A2(_02284_));
 sg13g2_buf_1 _22501_ (.A(_02478_),
    .X(_02479_));
 sg13g2_nor2_1 _22502_ (.A(net344),
    .B(net318),
    .Y(_02480_));
 sg13g2_nand2_1 _22503_ (.Y(_02481_),
    .A(net329),
    .B(net344));
 sg13g2_a21oi_1 _22504_ (.A1(_02442_),
    .A2(_02443_),
    .Y(_02482_),
    .B1(_02481_));
 sg13g2_nand2b_1 _22505_ (.Y(_02483_),
    .B(net344),
    .A_N(net329));
 sg13g2_nor2_1 _22506_ (.A(net318),
    .B(_02483_),
    .Y(_02484_));
 sg13g2_a221oi_1 _22507_ (.B2(net361),
    .C1(_02484_),
    .B1(_02482_),
    .A1(_02476_),
    .Y(_02485_),
    .A2(_02480_));
 sg13g2_buf_1 _22508_ (.A(_02485_),
    .X(_02486_));
 sg13g2_buf_1 _22509_ (.A(_02363_),
    .X(_02487_));
 sg13g2_o21ai_1 _22510_ (.B1(_02087_),
    .Y(_02488_),
    .A1(net345),
    .A2(net342));
 sg13g2_nand3_1 _22511_ (.B(net343),
    .C(_02393_),
    .A(net346),
    .Y(_02489_));
 sg13g2_nand2_1 _22512_ (.Y(_02490_),
    .A(_02435_),
    .B(_02353_));
 sg13g2_a21o_1 _22513_ (.A2(_02489_),
    .A1(_02488_),
    .B1(_02490_),
    .X(_02491_));
 sg13g2_buf_1 _22514_ (.A(net345),
    .X(_02492_));
 sg13g2_nor3_1 _22515_ (.A(_02134_),
    .B(net327),
    .C(net342),
    .Y(_02493_));
 sg13g2_buf_8 _22516_ (.A(_02307_),
    .X(_02494_));
 sg13g2_buf_1 _22517_ (.A(_02335_),
    .X(_02495_));
 sg13g2_a21oi_1 _22518_ (.A1(net326),
    .A2(net341),
    .Y(_02496_),
    .B1(_02094_));
 sg13g2_o21ai_1 _22519_ (.B1(_02445_),
    .Y(_02497_),
    .A1(_02493_),
    .A2(_02496_));
 sg13g2_mux2_1 _22520_ (.A0(_02272_),
    .A1(_02447_),
    .S(_02398_),
    .X(_02498_));
 sg13g2_buf_1 _22521_ (.A(_02498_),
    .X(_02499_));
 sg13g2_nor4_1 _22522_ (.A(_02260_),
    .B(_02284_),
    .C(net345),
    .D(_02363_),
    .Y(_02500_));
 sg13g2_a21oi_1 _22523_ (.A1(_02034_),
    .A2(_02051_),
    .Y(_02501_),
    .B1(_02075_));
 sg13g2_nand2_1 _22524_ (.Y(_02502_),
    .A(_02010_),
    .B(_02070_));
 sg13g2_nand2_1 _22525_ (.Y(_02503_),
    .A(_02501_),
    .B(_02502_));
 sg13g2_a221oi_1 _22526_ (.B2(net343),
    .C1(net329),
    .B1(net346),
    .A1(_02262_),
    .Y(_02504_),
    .A2(_02503_));
 sg13g2_mux2_1 _22527_ (.A0(_02415_),
    .A1(_02417_),
    .S(_02357_),
    .X(_02505_));
 sg13g2_a221oi_1 _22528_ (.B2(_02505_),
    .C1(_02253_),
    .B1(_02504_),
    .A1(_02499_),
    .Y(_02506_),
    .A2(_02500_));
 sg13g2_and3_1 _22529_ (.X(_02507_),
    .A(_02491_),
    .B(_02497_),
    .C(_02506_));
 sg13g2_buf_1 _22530_ (.A(_02507_),
    .X(_02508_));
 sg13g2_nor2_1 _22531_ (.A(net403),
    .B(_02368_),
    .Y(_02509_));
 sg13g2_nor4_1 _22532_ (.A(_02037_),
    .B(net345),
    .C(net342),
    .D(_02357_),
    .Y(_02510_));
 sg13g2_a221oi_1 _22533_ (.B2(_02353_),
    .C1(_02301_),
    .B1(_02346_),
    .A1(net346),
    .Y(_02511_),
    .A2(net343));
 sg13g2_a21o_1 _22534_ (.A2(_02510_),
    .A1(_02509_),
    .B1(_02511_),
    .X(_02512_));
 sg13g2_buf_1 _22535_ (.A(_02512_),
    .X(_02513_));
 sg13g2_nand2_1 _22536_ (.Y(_02514_),
    .A(_02262_),
    .B(_02503_));
 sg13g2_nor2_1 _22537_ (.A(_02514_),
    .B(_02282_),
    .Y(_02515_));
 sg13g2_and2_1 _22538_ (.A(_02513_),
    .B(_02515_),
    .X(_02516_));
 sg13g2_a21oi_1 _22539_ (.A1(_02486_),
    .A2(_02508_),
    .Y(_02517_),
    .B1(_02516_));
 sg13g2_buf_8 _22540_ (.A(net311),
    .X(_02518_));
 sg13g2_a22oi_1 _22541_ (.Y(_02519_),
    .B1(_02445_),
    .B2(_02090_),
    .A2(_02499_),
    .A1(_02286_));
 sg13g2_or2_1 _22542_ (.X(_02520_),
    .B(_02519_),
    .A(net303));
 sg13g2_buf_1 _22543_ (.A(_02520_),
    .X(_02521_));
 sg13g2_nand3_1 _22544_ (.B(net326),
    .C(net343),
    .A(_02424_),
    .Y(_02522_));
 sg13g2_o21ai_1 _22545_ (.B1(_02330_),
    .Y(_02523_),
    .A1(net327),
    .A2(net342));
 sg13g2_nand3_1 _22546_ (.B(_02368_),
    .C(_02398_),
    .A(net361),
    .Y(_02524_));
 sg13g2_a21o_1 _22547_ (.A2(_02523_),
    .A1(_02522_),
    .B1(_02524_),
    .X(_02525_));
 sg13g2_nand3_1 _22548_ (.B(net346),
    .C(_02395_),
    .A(net497),
    .Y(_02526_));
 sg13g2_o21ai_1 _22549_ (.B1(_02441_),
    .Y(_02527_),
    .A1(net345),
    .A2(_02487_));
 sg13g2_a21o_1 _22550_ (.A2(_02527_),
    .A1(_02526_),
    .B1(_02481_),
    .X(_02528_));
 sg13g2_nor3_1 _22551_ (.A(net327),
    .B(net342),
    .C(_02463_),
    .Y(_02529_));
 sg13g2_inv_1 _22552_ (.Y(_02530_),
    .A(_02393_));
 sg13g2_a21oi_1 _22553_ (.A1(net326),
    .A2(net343),
    .Y(_02531_),
    .B1(_02530_));
 sg13g2_o21ai_1 _22554_ (.B1(net330),
    .Y(_02532_),
    .A1(_02529_),
    .A2(_02531_));
 sg13g2_nor3_1 _22555_ (.A(_02266_),
    .B(net327),
    .C(net342),
    .Y(_02533_));
 sg13g2_mux2_1 _22556_ (.A0(_02415_),
    .A1(_02119_),
    .S(_02398_),
    .X(_02534_));
 sg13g2_a221oi_1 _22557_ (.B2(_02500_),
    .C1(_02253_),
    .B1(_02534_),
    .A1(_02445_),
    .Y(_02535_),
    .A2(_02533_));
 sg13g2_and4_1 _22558_ (.A(_02525_),
    .B(_02528_),
    .C(_02532_),
    .D(_02535_),
    .X(_02536_));
 sg13g2_buf_8 _22559_ (.A(_02536_),
    .X(_02537_));
 sg13g2_a21oi_1 _22560_ (.A1(net326),
    .A2(net343),
    .Y(_02538_),
    .B1(_02398_));
 sg13g2_and2_1 _22561_ (.A(_02088_),
    .B(net328),
    .X(_02539_));
 sg13g2_nor4_1 _22562_ (.A(_02301_),
    .B(net327),
    .C(net342),
    .D(net344),
    .Y(_02540_));
 sg13g2_a221oi_1 _22563_ (.B2(_02376_),
    .C1(_02540_),
    .B1(_02539_),
    .A1(_02134_),
    .Y(_02541_),
    .A2(_02538_));
 sg13g2_buf_1 _22564_ (.A(_02541_),
    .X(_02542_));
 sg13g2_nor2b_1 _22565_ (.A(_02542_),
    .B_N(_02515_),
    .Y(_02543_));
 sg13g2_a21oi_1 _22566_ (.A1(_02521_),
    .A2(_02537_),
    .Y(_02544_),
    .B1(_02543_));
 sg13g2_buf_2 _22567_ (.A(_02544_),
    .X(_02545_));
 sg13g2_o21ai_1 _22568_ (.B1(_02545_),
    .Y(_02546_),
    .A1(_02472_),
    .A2(_02517_));
 sg13g2_buf_1 _22569_ (.A(_02546_),
    .X(_02547_));
 sg13g2_buf_1 _22570_ (.A(_02547_),
    .X(_02548_));
 sg13g2_nand2_1 _22571_ (.Y(_02549_),
    .A(_02488_),
    .B(_02489_));
 sg13g2_mux4_1 _22572_ (.S0(net328),
    .A0(_02415_),
    .A1(_02119_),
    .A2(_02447_),
    .A3(_02441_),
    .S1(net311),
    .X(_02550_));
 sg13g2_a22oi_1 _22573_ (.Y(_02551_),
    .B1(_02550_),
    .B2(net312),
    .A2(_02445_),
    .A1(_02549_));
 sg13g2_mux2_1 _22574_ (.A0(_02272_),
    .A1(_02417_),
    .S(_02376_),
    .X(_02552_));
 sg13g2_a221oi_1 _22575_ (.B2(_02459_),
    .C1(_02477_),
    .B1(_02425_),
    .A1(net330),
    .Y(_02553_),
    .A2(_02552_));
 sg13g2_buf_1 _22576_ (.A(_02553_),
    .X(_02554_));
 sg13g2_a21o_1 _22577_ (.A2(_02137_),
    .A1(_02077_),
    .B1(_02251_),
    .X(_02555_));
 sg13g2_buf_1 _22578_ (.A(_02555_),
    .X(_02556_));
 sg13g2_buf_1 _22579_ (.A(_02556_),
    .X(_02557_));
 sg13g2_buf_8 _22580_ (.A(_02386_),
    .X(_02558_));
 sg13g2_nor4_1 _22581_ (.A(net325),
    .B(_02366_),
    .C(_02558_),
    .D(_02413_),
    .Y(_02559_));
 sg13g2_a21oi_1 _22582_ (.A1(_02551_),
    .A2(_02554_),
    .Y(_02560_),
    .B1(_02559_));
 sg13g2_buf_2 _22583_ (.A(_02560_),
    .X(_02561_));
 sg13g2_nor2_1 _22584_ (.A(_02317_),
    .B(_02492_),
    .Y(_02562_));
 sg13g2_a221oi_1 _22585_ (.B2(_02495_),
    .C1(_02481_),
    .B1(_02562_),
    .A1(_02424_),
    .Y(_02563_),
    .A2(net313));
 sg13g2_nor2_1 _22586_ (.A(_02492_),
    .B(_02430_),
    .Y(_02564_));
 sg13g2_buf_8 _22587_ (.A(net329),
    .X(_02565_));
 sg13g2_nand2_1 _22588_ (.Y(_02566_),
    .A(net317),
    .B(net328));
 sg13g2_a221oi_1 _22589_ (.B2(net341),
    .C1(_02566_),
    .B1(_02564_),
    .A1(_02474_),
    .Y(_02567_),
    .A2(net313));
 sg13g2_or3_1 _22590_ (.A(net318),
    .B(_02563_),
    .C(_02567_),
    .X(_02568_));
 sg13g2_buf_8 _22591_ (.A(net344),
    .X(_02569_));
 sg13g2_mux4_1 _22592_ (.S0(net324),
    .A0(net497),
    .A1(_02119_),
    .A2(_02330_),
    .A3(_02441_),
    .S1(net311),
    .X(_02570_));
 sg13g2_and2_1 _22593_ (.A(_02364_),
    .B(_02499_),
    .X(_02571_));
 sg13g2_a221oi_1 _22594_ (.B2(net312),
    .C1(_02571_),
    .B1(_02570_),
    .A1(_02333_),
    .Y(_02572_),
    .A2(_02505_));
 sg13g2_mux4_1 _22595_ (.S0(net311),
    .A0(_02266_),
    .A1(_02530_),
    .A2(_02463_),
    .A3(_02134_),
    .S1(net324),
    .X(_02573_));
 sg13g2_or2_1 _22596_ (.X(_02574_),
    .B(_02510_),
    .A(_02511_));
 sg13g2_mux2_1 _22597_ (.A0(_02573_),
    .A1(_02574_),
    .S(net297),
    .X(_02575_));
 sg13g2_nor2_1 _22598_ (.A(_02556_),
    .B(_02366_),
    .Y(_02576_));
 sg13g2_buf_1 _22599_ (.A(_02576_),
    .X(_02577_));
 sg13g2_a22oi_1 _22600_ (.Y(_02578_),
    .B1(_02575_),
    .B2(net291),
    .A2(_02572_),
    .A1(_02568_));
 sg13g2_buf_1 _22601_ (.A(_02578_),
    .X(_02579_));
 sg13g2_a221oi_1 _22602_ (.B2(_02286_),
    .C1(_02253_),
    .B1(_02460_),
    .A1(net360),
    .Y(_02580_),
    .A2(_02466_));
 sg13g2_buf_1 _22603_ (.A(_02580_),
    .X(_02581_));
 sg13g2_nand2_1 _22604_ (.Y(_02582_),
    .A(net561),
    .B(_02327_));
 sg13g2_xnor2_1 _22605_ (.Y(_02583_),
    .A(_02171_),
    .B(_02582_));
 sg13g2_mux4_1 _22606_ (.S0(_02388_),
    .A0(_02317_),
    .A1(_02313_),
    .A2(_02583_),
    .A3(_02255_),
    .S1(_02390_),
    .X(_02584_));
 sg13g2_a21o_1 _22607_ (.A2(_02584_),
    .A1(net317),
    .B1(net318),
    .X(_02585_));
 sg13g2_buf_1 _22608_ (.A(_02585_),
    .X(_02586_));
 sg13g2_a22oi_1 _22609_ (.Y(_02587_),
    .B1(_02581_),
    .B2(_02586_),
    .A2(_02577_),
    .A1(_02403_));
 sg13g2_buf_1 _22610_ (.A(_02587_),
    .X(_02588_));
 sg13g2_nor3_1 _22611_ (.A(_02561_),
    .B(_02579_),
    .C(_02588_),
    .Y(_02589_));
 sg13g2_buf_1 _22612_ (.A(_02589_),
    .X(_02590_));
 sg13g2_mux4_1 _22613_ (.S0(net311),
    .A0(_02272_),
    .A1(_02087_),
    .A2(_02393_),
    .A3(_02417_),
    .S1(_02411_),
    .X(_02591_));
 sg13g2_mux2_1 _22614_ (.A0(_02591_),
    .A1(_02542_),
    .S(net297),
    .X(_02592_));
 sg13g2_buf_1 _22615_ (.A(_02592_),
    .X(_02593_));
 sg13g2_nand2b_1 _22616_ (.Y(_02594_),
    .B(net291),
    .A_N(_02593_));
 sg13g2_and2_1 _22617_ (.A(net317),
    .B(net324),
    .X(_02595_));
 sg13g2_buf_1 _22618_ (.A(_02595_),
    .X(_02596_));
 sg13g2_mux2_1 _22619_ (.A0(_02317_),
    .A1(_02313_),
    .S(net303),
    .X(_02597_));
 sg13g2_nand3_1 _22620_ (.B(_02293_),
    .C(net326),
    .A(_02210_),
    .Y(_02598_));
 sg13g2_and2_1 _22621_ (.A(net561),
    .B(_02198_),
    .X(_02599_));
 sg13g2_nand4_1 _22622_ (.B(net326),
    .C(net341),
    .A(_02199_),
    .Y(_02600_),
    .D(_02599_));
 sg13g2_nand3_1 _22623_ (.B(net327),
    .C(_02599_),
    .A(_02210_),
    .Y(_02601_));
 sg13g2_and3_1 _22624_ (.X(_02602_),
    .A(_02598_),
    .B(_02600_),
    .C(_02601_));
 sg13g2_o21ai_1 _22625_ (.B1(_02198_),
    .Y(_02603_),
    .A1(net327),
    .A2(_02487_));
 sg13g2_nor3_1 _22626_ (.A(_02292_),
    .B(_02299_),
    .C(_02305_),
    .Y(_02604_));
 sg13g2_inv_1 _22627_ (.Y(_02605_),
    .A(_02427_));
 sg13g2_a21oi_1 _22628_ (.A1(net341),
    .A2(_02604_),
    .Y(_02606_),
    .B1(_02605_));
 sg13g2_a21oi_1 _22629_ (.A1(_02603_),
    .A2(_02606_),
    .Y(_02607_),
    .B1(_02566_));
 sg13g2_a221oi_1 _22630_ (.B2(_02607_),
    .C1(net318),
    .B1(_02602_),
    .A1(_02596_),
    .Y(_02608_),
    .A2(_02597_));
 sg13g2_mux2_1 _22631_ (.A0(_02499_),
    .A1(_02534_),
    .S(net303),
    .X(_02609_));
 sg13g2_mux4_1 _22632_ (.S0(net324),
    .A0(_02424_),
    .A1(net497),
    .A2(_02330_),
    .A3(_02441_),
    .S1(net313),
    .X(_02610_));
 sg13g2_a221oi_1 _22633_ (.B2(net312),
    .C1(net331),
    .B1(_02610_),
    .A1(net360),
    .Y(_02611_),
    .A2(_02609_));
 sg13g2_nand2b_1 _22634_ (.Y(_02612_),
    .B(_02611_),
    .A_N(_02608_));
 sg13g2_nand2_1 _22635_ (.Y(_02613_),
    .A(_02594_),
    .B(_02612_));
 sg13g2_buf_1 _22636_ (.A(_02613_),
    .X(_02614_));
 sg13g2_buf_1 _22637_ (.A(_02614_),
    .X(_02615_));
 sg13g2_buf_1 _22638_ (.A(net201),
    .X(_02616_));
 sg13g2_a21oi_1 _22639_ (.A1(net202),
    .A2(net228),
    .Y(_02617_),
    .B1(net170));
 sg13g2_xnor2_1 _22640_ (.Y(_02618_),
    .A(net171),
    .B(_02617_));
 sg13g2_buf_1 _22641_ (.A(_02618_),
    .X(_02619_));
 sg13g2_or2_1 _22642_ (.X(_02620_),
    .B(_02476_),
    .A(_02437_));
 sg13g2_a221oi_1 _22643_ (.B2(_02495_),
    .C1(_02483_),
    .B1(_02562_),
    .A1(_02424_),
    .Y(_02621_),
    .A2(net313));
 sg13g2_and3_1 _22644_ (.X(_02622_),
    .A(_02288_),
    .B(net326),
    .C(net341));
 sg13g2_a21oi_1 _22645_ (.A1(_02494_),
    .A2(net341),
    .Y(_02623_),
    .B1(_02297_));
 sg13g2_o21ai_1 _22646_ (.B1(net325),
    .Y(_02624_),
    .A1(_02622_),
    .A2(_02623_));
 sg13g2_and4_1 _22647_ (.A(net360),
    .B(_02442_),
    .C(_02443_),
    .D(_02596_),
    .X(_02625_));
 sg13g2_a21oi_1 _22648_ (.A1(_02494_),
    .A2(net341),
    .Y(_02626_),
    .B1(_02428_));
 sg13g2_a221oi_1 _22649_ (.B2(_02353_),
    .C1(_02626_),
    .B1(_02346_),
    .A1(_02290_),
    .Y(_02627_),
    .A2(net303));
 sg13g2_nor4_1 _22650_ (.A(_02621_),
    .B(_02624_),
    .C(_02625_),
    .D(_02627_),
    .Y(_02628_));
 sg13g2_a221oi_1 _22651_ (.B2(_02370_),
    .C1(net403),
    .B1(net317),
    .A1(_02355_),
    .Y(_02629_),
    .A2(_02514_));
 sg13g2_buf_2 _22652_ (.A(_02629_),
    .X(_02630_));
 sg13g2_xnor2_1 _22653_ (.Y(_02631_),
    .A(net737),
    .B(_02341_));
 sg13g2_mux2_1 _22654_ (.A0(_02067_),
    .A1(_02631_),
    .S(net328),
    .X(_02632_));
 sg13g2_a21o_1 _22655_ (.A2(_02082_),
    .A1(_02073_),
    .B1(_02083_),
    .X(_02633_));
 sg13g2_mux2_1 _22656_ (.A0(_02462_),
    .A1(_02633_),
    .S(net324),
    .X(_02634_));
 sg13g2_mux2_1 _22657_ (.A0(_02632_),
    .A1(_02634_),
    .S(net313),
    .X(_02635_));
 sg13g2_a221oi_1 _22658_ (.B2(_02381_),
    .C1(_02557_),
    .B1(_02513_),
    .A1(_02630_),
    .Y(_02636_),
    .A2(_02635_));
 sg13g2_nand3_1 _22659_ (.B(net297),
    .C(_02573_),
    .A(net304),
    .Y(_02637_));
 sg13g2_a22oi_1 _22660_ (.Y(_02638_),
    .B1(_02636_),
    .B2(_02637_),
    .A2(_02628_),
    .A1(_02620_));
 sg13g2_buf_2 _22661_ (.A(_02638_),
    .X(_02639_));
 sg13g2_buf_8 _22662_ (.A(_02639_),
    .X(_02640_));
 sg13g2_buf_1 _22663_ (.A(_02640_),
    .X(_02641_));
 sg13g2_or2_1 _22664_ (.X(_02642_),
    .B(net317),
    .A(_02260_));
 sg13g2_buf_1 _22665_ (.A(_02642_),
    .X(_02643_));
 sg13g2_nand2_1 _22666_ (.Y(_02644_),
    .A(_02526_),
    .B(_02527_));
 sg13g2_nand3_1 _22667_ (.B(net326),
    .C(net341),
    .A(_02119_),
    .Y(_02645_));
 sg13g2_o21ai_1 _22668_ (.B1(_02447_),
    .Y(_02646_),
    .A1(net327),
    .A2(net342));
 sg13g2_a221oi_1 _22669_ (.B2(_02646_),
    .C1(net361),
    .B1(_02645_),
    .A1(_02346_),
    .Y(_02647_),
    .A2(_02353_));
 sg13g2_a21oi_1 _22670_ (.A1(net330),
    .A2(_02644_),
    .Y(_02648_),
    .B1(_02647_));
 sg13g2_o21ai_1 _22671_ (.B1(_02648_),
    .Y(_02649_),
    .A1(_02643_),
    .A2(_02584_));
 sg13g2_or2_1 _22672_ (.X(_02650_),
    .B(_02419_),
    .A(_02410_));
 sg13g2_buf_1 _22673_ (.A(_02650_),
    .X(_02651_));
 sg13g2_nand3_1 _22674_ (.B(_02438_),
    .C(_02450_),
    .A(_02426_),
    .Y(_02652_));
 sg13g2_buf_1 _22675_ (.A(_02652_),
    .X(_02653_));
 sg13g2_nand2_1 _22676_ (.Y(_02654_),
    .A(net324),
    .B(_02447_));
 sg13g2_and2_1 _22677_ (.A(_02088_),
    .B(_02381_),
    .X(_02655_));
 sg13g2_a21o_1 _22678_ (.A2(_02655_),
    .A1(net317),
    .B1(_02556_),
    .X(_02656_));
 sg13g2_a221oi_1 _22679_ (.B2(_02654_),
    .C1(_02656_),
    .B1(_02465_),
    .A1(net311),
    .Y(_02657_),
    .A2(_02464_));
 sg13g2_a221oi_1 _22680_ (.B2(_02399_),
    .C1(_02656_),
    .B1(_02394_),
    .A1(net311),
    .Y(_02658_),
    .A2(_02389_));
 sg13g2_mux2_1 _22681_ (.A0(_02657_),
    .A1(_02658_),
    .S(net297),
    .X(_02659_));
 sg13g2_buf_1 _22682_ (.A(net328),
    .X(_02660_));
 sg13g2_mux2_1 _22683_ (.A0(_02297_),
    .A1(_02431_),
    .S(net313),
    .X(_02661_));
 sg13g2_a21oi_1 _22684_ (.A1(_02603_),
    .A2(_02606_),
    .Y(_02662_),
    .B1(net328));
 sg13g2_nand2b_1 _22685_ (.Y(_02663_),
    .B(_02557_),
    .A_N(net318));
 sg13g2_a221oi_1 _22686_ (.B2(_02662_),
    .C1(_02663_),
    .B1(_02602_),
    .A1(net316),
    .Y(_02664_),
    .A2(_02661_));
 sg13g2_or2_1 _22687_ (.X(_02665_),
    .B(_02664_),
    .A(_02659_));
 sg13g2_buf_2 _22688_ (.A(_02665_),
    .X(_02666_));
 sg13g2_a221oi_1 _22689_ (.B2(_02653_),
    .C1(_02666_),
    .B1(_02651_),
    .A1(net325),
    .Y(_02667_),
    .A2(_02649_));
 sg13g2_buf_2 _22690_ (.A(_02667_),
    .X(_02668_));
 sg13g2_buf_8 _22691_ (.A(_02668_),
    .X(_02669_));
 sg13g2_nand3_1 _22692_ (.B(net201),
    .C(net200),
    .A(net227),
    .Y(_02670_));
 sg13g2_buf_1 _22693_ (.A(_02670_),
    .X(_02671_));
 sg13g2_buf_1 _22694_ (.A(_02561_),
    .X(_02672_));
 sg13g2_buf_1 _22695_ (.A(_02579_),
    .X(_02673_));
 sg13g2_nor2_1 _22696_ (.A(net252),
    .B(net251),
    .Y(_02674_));
 sg13g2_buf_1 _22697_ (.A(_02588_),
    .X(_02675_));
 sg13g2_nor2b_1 _22698_ (.A(net250),
    .B_N(net253),
    .Y(_02676_));
 sg13g2_nand4_1 _22699_ (.B(_02674_),
    .C(net200),
    .A(net202),
    .Y(_02677_),
    .D(_02676_));
 sg13g2_buf_1 _22700_ (.A(_02677_),
    .X(_02678_));
 sg13g2_nand2_2 _22701_ (.Y(_02679_),
    .A(_02671_),
    .B(_02678_));
 sg13g2_buf_1 _22702_ (.A(_02617_),
    .X(_02680_));
 sg13g2_buf_1 _22703_ (.A(_02594_),
    .X(_02681_));
 sg13g2_buf_8 _22704_ (.A(_02612_),
    .X(_02682_));
 sg13g2_buf_8 _22705_ (.A(_02545_),
    .X(_02683_));
 sg13g2_buf_1 _22706_ (.A(net248),
    .X(_02684_));
 sg13g2_buf_8 _22707_ (.A(net226),
    .X(_02685_));
 sg13g2_buf_1 _22708_ (.A(net199),
    .X(_02686_));
 sg13g2_buf_1 _22709_ (.A(_02517_),
    .X(_02687_));
 sg13g2_buf_1 _22710_ (.A(net285),
    .X(_02688_));
 sg13g2_a221oi_1 _22711_ (.B2(_02471_),
    .C1(_02543_),
    .B1(_02461_),
    .A1(_02521_),
    .Y(_02689_),
    .A2(_02537_));
 sg13g2_a221oi_1 _22712_ (.B2(net274),
    .C1(_02689_),
    .B1(net169),
    .A1(net249),
    .Y(_02690_),
    .A2(net275));
 sg13g2_and2_1 _22713_ (.A(net228),
    .B(_02690_),
    .X(_02691_));
 sg13g2_buf_2 _22714_ (.A(_02691_),
    .X(_02692_));
 sg13g2_nor2_1 _22715_ (.A(net122),
    .B(_02692_),
    .Y(_02693_));
 sg13g2_buf_1 _22716_ (.A(_02693_),
    .X(_02694_));
 sg13g2_buf_1 _22717_ (.A(_02694_),
    .X(_02695_));
 sg13g2_mux4_1 _22718_ (.S0(_02432_),
    .A0(_02152_),
    .A1(_02474_),
    .A2(_02330_),
    .A3(_02424_),
    .S1(net324),
    .X(_02696_));
 sg13g2_a221oi_1 _22719_ (.B2(net312),
    .C1(_02647_),
    .B1(_02696_),
    .A1(net330),
    .Y(_02697_),
    .A2(_02644_));
 sg13g2_or2_1 _22720_ (.X(_02698_),
    .B(_02697_),
    .A(net331));
 sg13g2_buf_8 _22721_ (.A(_02698_),
    .X(_02699_));
 sg13g2_nor2_1 _22722_ (.A(_02659_),
    .B(_02664_),
    .Y(_02700_));
 sg13g2_buf_2 _22723_ (.A(_02700_),
    .X(_02701_));
 sg13g2_nand2_1 _22724_ (.Y(_02702_),
    .A(_02699_),
    .B(_02701_));
 sg13g2_buf_1 _22725_ (.A(_02702_),
    .X(_02703_));
 sg13g2_buf_8 _22726_ (.A(net225),
    .X(_02704_));
 sg13g2_buf_1 _22727_ (.A(net198),
    .X(_02705_));
 sg13g2_buf_1 _22728_ (.A(_02705_),
    .X(_02706_));
 sg13g2_nand2_1 _22729_ (.Y(_02707_),
    .A(_02620_),
    .B(_02628_));
 sg13g2_nand2_1 _22730_ (.Y(_02708_),
    .A(_02636_),
    .B(_02637_));
 sg13g2_nand2_1 _22731_ (.Y(_02709_),
    .A(_02707_),
    .B(_02708_));
 sg13g2_buf_2 _22732_ (.A(_02709_),
    .X(_02710_));
 sg13g2_buf_1 _22733_ (.A(_02710_),
    .X(_02711_));
 sg13g2_buf_1 _22734_ (.A(net224),
    .X(_02712_));
 sg13g2_nand2_2 _22735_ (.Y(_02713_),
    .A(net228),
    .B(_02690_));
 sg13g2_nor2_1 _22736_ (.A(net171),
    .B(net122),
    .Y(_02714_));
 sg13g2_o21ai_1 _22737_ (.B1(_02714_),
    .Y(_02715_),
    .A1(net197),
    .A2(_02713_));
 sg13g2_nor2_1 _22738_ (.A(_02410_),
    .B(_02593_),
    .Y(_02716_));
 sg13g2_nor2b_1 _22739_ (.A(_02608_),
    .B_N(_02611_),
    .Y(_02717_));
 sg13g2_buf_2 _22740_ (.A(_02717_),
    .X(_02718_));
 sg13g2_nor2_1 _22741_ (.A(_02716_),
    .B(_02718_),
    .Y(_02719_));
 sg13g2_buf_2 _22742_ (.A(_02719_),
    .X(_02720_));
 sg13g2_buf_8 _22743_ (.A(_02720_),
    .X(_02721_));
 sg13g2_buf_1 _22744_ (.A(net196),
    .X(_02722_));
 sg13g2_nand2_1 _22745_ (.Y(_02723_),
    .A(_02486_),
    .B(_02508_));
 sg13g2_a221oi_1 _22746_ (.B2(_02513_),
    .C1(_02543_),
    .B1(_02515_),
    .A1(_02521_),
    .Y(_02724_),
    .A2(_02537_));
 sg13g2_buf_1 _22747_ (.A(_02724_),
    .X(_02725_));
 sg13g2_a221oi_1 _22748_ (.B2(_02725_),
    .C1(_02561_),
    .B1(_02723_),
    .A1(_02545_),
    .Y(_02726_),
    .A2(_02472_));
 sg13g2_buf_8 _22749_ (.A(_02726_),
    .X(_02727_));
 sg13g2_buf_1 _22750_ (.A(net223),
    .X(_02728_));
 sg13g2_nor2_1 _22751_ (.A(net251),
    .B(net250),
    .Y(_02729_));
 sg13g2_buf_1 _22752_ (.A(_02729_),
    .X(_02730_));
 sg13g2_a21oi_1 _22753_ (.A1(net195),
    .A2(net194),
    .Y(_02731_),
    .B1(_02704_));
 sg13g2_or2_1 _22754_ (.X(_02732_),
    .B(_02731_),
    .A(net167));
 sg13g2_buf_1 _22755_ (.A(net227),
    .X(_02733_));
 sg13g2_buf_1 _22756_ (.A(net193),
    .X(_02734_));
 sg13g2_nor2_1 _22757_ (.A(_02734_),
    .B(net171),
    .Y(_02735_));
 sg13g2_a22oi_1 _22758_ (.Y(_02736_),
    .B1(_02732_),
    .B2(_02735_),
    .A2(_02715_),
    .A1(_02706_));
 sg13g2_buf_1 _22759_ (.A(_02736_),
    .X(_02737_));
 sg13g2_nor3_2 _22760_ (.A(net297),
    .B(_02382_),
    .C(_02413_),
    .Y(_02738_));
 sg13g2_nand2_1 _22761_ (.Y(_02739_),
    .A(_02738_),
    .B(net254));
 sg13g2_buf_1 _22762_ (.A(_02739_),
    .X(_02740_));
 sg13g2_o21ai_1 _22763_ (.B1(_02366_),
    .Y(_02741_),
    .A1(_02558_),
    .A2(_02542_));
 sg13g2_a21oi_1 _22764_ (.A1(net331),
    .A2(_02741_),
    .Y(_02742_),
    .B1(_02251_));
 sg13g2_buf_2 _22765_ (.A(_02742_),
    .X(_02743_));
 sg13g2_nor2_2 _22766_ (.A(net253),
    .B(_02743_),
    .Y(_02744_));
 sg13g2_buf_8 _22767_ (.A(net251),
    .X(_02745_));
 sg13g2_a21oi_2 _22768_ (.B1(net222),
    .Y(_02746_),
    .A2(net275),
    .A1(net249));
 sg13g2_nand3_1 _22769_ (.B(_02744_),
    .C(_02746_),
    .A(net171),
    .Y(_02747_));
 sg13g2_buf_1 _22770_ (.A(_02747_),
    .X(_02748_));
 sg13g2_buf_1 _22771_ (.A(_02669_),
    .X(_02749_));
 sg13g2_nand3_1 _22772_ (.B(net122),
    .C(net165),
    .A(net197),
    .Y(_02750_));
 sg13g2_a21oi_1 _22773_ (.A1(net249),
    .A2(net275),
    .Y(_02751_),
    .B1(_02640_));
 sg13g2_o21ai_1 _22774_ (.B1(net148),
    .Y(_02752_),
    .A1(net171),
    .A2(_02751_));
 sg13g2_nand2_1 _22775_ (.Y(_02753_),
    .A(net166),
    .B(_02457_));
 sg13g2_nand3_1 _22776_ (.B(_02752_),
    .C(_02753_),
    .A(_02750_),
    .Y(_02754_));
 sg13g2_buf_1 _22777_ (.A(_02651_),
    .X(_02755_));
 sg13g2_buf_8 _22778_ (.A(_02653_),
    .X(_02756_));
 sg13g2_nand2_1 _22779_ (.Y(_02757_),
    .A(net273),
    .B(net272));
 sg13g2_buf_2 _22780_ (.A(_02757_),
    .X(_02758_));
 sg13g2_buf_1 _22781_ (.A(_02758_),
    .X(_02759_));
 sg13g2_buf_1 _22782_ (.A(net191),
    .X(_02760_));
 sg13g2_buf_1 _22783_ (.A(net164),
    .X(_02761_));
 sg13g2_and2_1 _22784_ (.A(_02461_),
    .B(_02471_),
    .X(_02762_));
 sg13g2_buf_1 _22785_ (.A(_02762_),
    .X(_02763_));
 sg13g2_a21o_1 _22786_ (.A2(_02508_),
    .A1(_02486_),
    .B1(_02516_),
    .X(_02764_));
 sg13g2_buf_8 _22787_ (.A(_02764_),
    .X(_02765_));
 sg13g2_a21o_1 _22788_ (.A2(_02537_),
    .A1(_02521_),
    .B1(_02543_),
    .X(_02766_));
 sg13g2_buf_1 _22789_ (.A(_02766_),
    .X(_02767_));
 sg13g2_a21oi_1 _22790_ (.A1(_02763_),
    .A2(_02765_),
    .Y(_02768_),
    .B1(net271));
 sg13g2_buf_2 _22791_ (.A(_02768_),
    .X(_02769_));
 sg13g2_buf_1 _22792_ (.A(_02769_),
    .X(_02770_));
 sg13g2_or3_1 _22793_ (.A(_02561_),
    .B(net251),
    .C(_02588_),
    .X(_02771_));
 sg13g2_buf_2 _22794_ (.A(_02771_),
    .X(_02772_));
 sg13g2_o21ai_1 _22795_ (.B1(net196),
    .Y(_02773_),
    .A1(net190),
    .A2(net189));
 sg13g2_buf_8 _22796_ (.A(_02773_),
    .X(_02774_));
 sg13g2_nor2_1 _22797_ (.A(net147),
    .B(net146),
    .Y(_02775_));
 sg13g2_a21o_1 _22798_ (.A2(_02741_),
    .A1(net331),
    .B1(_02251_),
    .X(_02776_));
 sg13g2_buf_2 _22799_ (.A(_02776_),
    .X(_02777_));
 sg13g2_a22oi_1 _22800_ (.Y(_02778_),
    .B1(_02775_),
    .B2(_02777_),
    .A2(_02714_),
    .A1(net166));
 sg13g2_nor2_1 _22801_ (.A(net148),
    .B(_02778_),
    .Y(_02779_));
 sg13g2_nor2_2 _22802_ (.A(net331),
    .B(_02697_),
    .Y(_02780_));
 sg13g2_nor2_1 _22803_ (.A(_02780_),
    .B(_02666_),
    .Y(_02781_));
 sg13g2_buf_2 _22804_ (.A(_02781_),
    .X(_02782_));
 sg13g2_buf_1 _22805_ (.A(_02782_),
    .X(_02783_));
 sg13g2_nor2_1 _22806_ (.A(net197),
    .B(net146),
    .Y(_02784_));
 sg13g2_a21oi_1 _22807_ (.A1(net146),
    .A2(_02744_),
    .Y(_02785_),
    .B1(_02784_));
 sg13g2_nor3_1 _22808_ (.A(net188),
    .B(net171),
    .C(_02785_),
    .Y(_02786_));
 sg13g2_nor2_1 _22809_ (.A(net197),
    .B(net122),
    .Y(_02787_));
 sg13g2_a22oi_1 _22810_ (.Y(_02788_),
    .B1(_02787_),
    .B2(net148),
    .A2(_02744_),
    .A1(net122));
 sg13g2_nor2_1 _22811_ (.A(_02769_),
    .B(net189),
    .Y(_02789_));
 sg13g2_buf_1 _22812_ (.A(_02789_),
    .X(_02790_));
 sg13g2_a22oi_1 _22813_ (.Y(_02791_),
    .B1(_02681_),
    .B2(_02682_),
    .A2(net272),
    .A1(net273));
 sg13g2_buf_1 _22814_ (.A(_02791_),
    .X(_02792_));
 sg13g2_a21oi_1 _22815_ (.A1(net145),
    .A2(net187),
    .Y(_02793_),
    .B1(net254));
 sg13g2_o21ai_1 _22816_ (.B1(_02793_),
    .Y(_02794_),
    .A1(net147),
    .A2(_02788_));
 sg13g2_nor3_1 _22817_ (.A(_02779_),
    .B(_02786_),
    .C(_02794_),
    .Y(_02795_));
 sg13g2_a21oi_1 _22818_ (.A1(_02748_),
    .A2(_02754_),
    .Y(_02796_),
    .B1(_02795_));
 sg13g2_nor2_1 _22819_ (.A(_02748_),
    .B(_02754_),
    .Y(_02797_));
 sg13g2_nor2_1 _22820_ (.A(_02797_),
    .B(_02796_),
    .Y(_02798_));
 sg13g2_xnor2_1 _22821_ (.Y(_02799_),
    .A(_02761_),
    .B(_02680_));
 sg13g2_buf_1 _22822_ (.A(_02799_),
    .X(_02800_));
 sg13g2_nand2_1 _22823_ (.Y(_02801_),
    .A(net146),
    .B(_02749_));
 sg13g2_nand2_1 _22824_ (.Y(_02802_),
    .A(net148),
    .B(net203));
 sg13g2_nand2_1 _22825_ (.Y(_02803_),
    .A(_02801_),
    .B(_02802_));
 sg13g2_a22oi_1 _22826_ (.Y(_02804_),
    .B1(_02803_),
    .B2(_02712_),
    .A2(_02800_),
    .A1(net148));
 sg13g2_nor2_1 _22827_ (.A(net297),
    .B(_02413_),
    .Y(_02805_));
 sg13g2_nand2_1 _22828_ (.Y(_02806_),
    .A(_02381_),
    .B(_02805_));
 sg13g2_buf_2 _22829_ (.A(_02806_),
    .X(_02807_));
 sg13g2_o21ai_1 _22830_ (.B1(_02807_),
    .Y(_02808_),
    .A1(_02743_),
    .A2(_02804_));
 sg13g2_buf_1 _22831_ (.A(_02808_),
    .X(_02809_));
 sg13g2_mux2_1 _22832_ (.A0(_02796_),
    .A1(_02798_),
    .S(_02809_),
    .X(_02810_));
 sg13g2_a21oi_1 _22833_ (.A1(net192),
    .A2(_02810_),
    .Y(_02811_),
    .B1(_02797_));
 sg13g2_xnor2_1 _22834_ (.Y(_02812_),
    .A(_02737_),
    .B(_02811_));
 sg13g2_a21o_1 _22835_ (.A2(net83),
    .A1(_02679_),
    .B1(_02812_),
    .X(_02813_));
 sg13g2_o21ai_1 _22836_ (.B1(_02381_),
    .Y(_02814_),
    .A1(_02384_),
    .A2(_02403_));
 sg13g2_buf_1 _22837_ (.A(_02814_),
    .X(_02815_));
 sg13g2_nor2_1 _22838_ (.A(_02807_),
    .B(_02815_),
    .Y(_02816_));
 sg13g2_buf_2 _22839_ (.A(_02816_),
    .X(_02817_));
 sg13g2_nor2_1 _22840_ (.A(_02817_),
    .B(_02795_),
    .Y(_02818_));
 sg13g2_a221oi_1 _22841_ (.B2(net188),
    .C1(net197),
    .B1(_02694_),
    .A1(net273),
    .Y(_02819_),
    .A2(net272));
 sg13g2_o21ai_1 _22842_ (.B1(_02713_),
    .Y(_02820_),
    .A1(net148),
    .A2(net146));
 sg13g2_a21oi_1 _22843_ (.A1(net147),
    .A2(_02820_),
    .Y(_02821_),
    .B1(net166));
 sg13g2_o21ai_1 _22844_ (.B1(_02752_),
    .Y(_02822_),
    .A1(_02819_),
    .A2(_02821_));
 sg13g2_xnor2_1 _22845_ (.Y(_02823_),
    .A(_02748_),
    .B(_02822_));
 sg13g2_xnor2_1 _22846_ (.Y(_02824_),
    .A(_02818_),
    .B(_02823_));
 sg13g2_nand2_1 _22847_ (.Y(_02825_),
    .A(_02403_),
    .B(net291));
 sg13g2_nand2_1 _22848_ (.Y(_02826_),
    .A(_02581_),
    .B(_02586_));
 sg13g2_nand2_1 _22849_ (.Y(_02827_),
    .A(_02825_),
    .B(_02826_));
 sg13g2_buf_1 _22850_ (.A(_02827_),
    .X(_02828_));
 sg13g2_inv_2 _22851_ (.Y(_02829_),
    .A(net222));
 sg13g2_a21oi_1 _22852_ (.A1(_02828_),
    .A2(net223),
    .Y(_02830_),
    .B1(_02829_));
 sg13g2_nor2_1 _22853_ (.A(net145),
    .B(_02830_),
    .Y(_02831_));
 sg13g2_buf_2 _22854_ (.A(_02831_),
    .X(_02832_));
 sg13g2_nand2_1 _22855_ (.Y(_02833_),
    .A(_02807_),
    .B(_02815_));
 sg13g2_buf_1 _22856_ (.A(_02833_),
    .X(_02834_));
 sg13g2_nand2_1 _22857_ (.Y(_02835_),
    .A(net192),
    .B(_02834_));
 sg13g2_o21ai_1 _22858_ (.B1(_02835_),
    .Y(_02836_),
    .A1(_02743_),
    .A2(_02832_));
 sg13g2_buf_1 _22859_ (.A(_02836_),
    .X(_02837_));
 sg13g2_xnor2_1 _22860_ (.Y(_02838_),
    .A(_02828_),
    .B(net223));
 sg13g2_buf_2 _22861_ (.A(_02838_),
    .X(_02839_));
 sg13g2_a21oi_1 _22862_ (.A1(_02777_),
    .A2(_02839_),
    .Y(_02840_),
    .B1(_02738_));
 sg13g2_nor3_2 _22863_ (.A(net224),
    .B(_02832_),
    .C(_02840_),
    .Y(_02841_));
 sg13g2_inv_1 _22864_ (.Y(_02842_),
    .A(_02841_));
 sg13g2_a21oi_1 _22865_ (.A1(_02711_),
    .A2(net146),
    .Y(_02843_),
    .B1(_02692_));
 sg13g2_mux2_1 _22866_ (.A0(net146),
    .A1(_02843_),
    .S(_02783_),
    .X(_02844_));
 sg13g2_nor4_2 _22867_ (.A(_02780_),
    .B(_02666_),
    .C(net287),
    .Y(_02845_),
    .D(net286));
 sg13g2_nor2_1 _22868_ (.A(net224),
    .B(_02749_),
    .Y(_02846_));
 sg13g2_a22oi_1 _22869_ (.Y(_02847_),
    .B1(_02694_),
    .B2(_02846_),
    .A2(_02845_),
    .A1(net122));
 sg13g2_o21ai_1 _22870_ (.B1(_02847_),
    .Y(_02848_),
    .A1(net171),
    .A2(_02844_));
 sg13g2_buf_1 _22871_ (.A(_02848_),
    .X(_02849_));
 sg13g2_xnor2_1 _22872_ (.Y(_02850_),
    .A(_02842_),
    .B(_02849_));
 sg13g2_buf_1 _22873_ (.A(net170),
    .X(_02851_));
 sg13g2_nand2_1 _22874_ (.Y(_02852_),
    .A(net202),
    .B(_02590_));
 sg13g2_buf_1 _22875_ (.A(_02852_),
    .X(_02853_));
 sg13g2_nor4_1 _22876_ (.A(net166),
    .B(net148),
    .C(net190),
    .D(net189),
    .Y(_02854_));
 sg13g2_a21oi_1 _22877_ (.A1(net166),
    .A2(net143),
    .Y(_02855_),
    .B1(_02854_));
 sg13g2_buf_1 _22878_ (.A(_02745_),
    .X(_02856_));
 sg13g2_buf_1 _22879_ (.A(net186),
    .X(_02857_));
 sg13g2_or2_1 _22880_ (.X(_02858_),
    .B(_02857_),
    .A(net193));
 sg13g2_nand2_1 _22881_ (.Y(_02859_),
    .A(net144),
    .B(_02858_));
 sg13g2_buf_1 _22882_ (.A(net163),
    .X(_02860_));
 sg13g2_buf_1 _22883_ (.A(net142),
    .X(_02861_));
 sg13g2_nor2b_1 _22884_ (.A(net166),
    .B_N(net121),
    .Y(_02862_));
 sg13g2_and3_1 _22885_ (.X(_02863_),
    .A(net253),
    .B(_02681_),
    .C(_02682_));
 sg13g2_buf_1 _22886_ (.A(_02863_),
    .X(_02864_));
 sg13g2_a21o_1 _22887_ (.A2(_02862_),
    .A1(_02792_),
    .B1(_02864_),
    .X(_02865_));
 sg13g2_a22oi_1 _22888_ (.Y(_02866_),
    .B1(_02865_),
    .B2(net148),
    .A2(_02859_),
    .A1(net171));
 sg13g2_o21ai_1 _22889_ (.B1(_02866_),
    .Y(_02867_),
    .A1(net144),
    .A2(_02855_));
 sg13g2_buf_1 _22890_ (.A(_02867_),
    .X(_02868_));
 sg13g2_a21oi_1 _22891_ (.A1(net195),
    .A2(net165),
    .Y(_02869_),
    .B1(net144));
 sg13g2_or2_1 _22892_ (.X(_02870_),
    .B(net250),
    .A(net251));
 sg13g2_buf_2 _22893_ (.A(_02870_),
    .X(_02871_));
 sg13g2_nor2_1 _22894_ (.A(net166),
    .B(_02871_),
    .Y(_02872_));
 sg13g2_nand2_2 _22895_ (.Y(_02873_),
    .A(_02782_),
    .B(net191));
 sg13g2_a21oi_1 _22896_ (.A1(_02873_),
    .A2(_02802_),
    .Y(_02874_),
    .B1(net146));
 sg13g2_nor2_1 _22897_ (.A(_02692_),
    .B(_02874_),
    .Y(_02875_));
 sg13g2_a221oi_1 _22898_ (.B2(_02841_),
    .C1(_02679_),
    .B1(_02875_),
    .A1(_02869_),
    .Y(_02876_),
    .A2(_02872_));
 sg13g2_buf_1 _22899_ (.A(_02876_),
    .X(_02877_));
 sg13g2_nand2_1 _22900_ (.Y(_02878_),
    .A(_02868_),
    .B(_02877_));
 sg13g2_o21ai_1 _22901_ (.B1(net197),
    .Y(_02879_),
    .A1(_02680_),
    .A2(_02692_));
 sg13g2_nand2_1 _22902_ (.Y(_02880_),
    .A(net193),
    .B(net191));
 sg13g2_mux2_1 _22903_ (.A0(net147),
    .A1(_02880_),
    .S(_02713_),
    .X(_02881_));
 sg13g2_a21oi_1 _22904_ (.A1(_02879_),
    .A2(_02881_),
    .Y(_02882_),
    .B1(_02834_));
 sg13g2_o21ai_1 _22905_ (.B1(_02882_),
    .Y(_02883_),
    .A1(_02868_),
    .A2(_02877_));
 sg13g2_a22oi_1 _22906_ (.Y(_02884_),
    .B1(_02878_),
    .B2(_02883_),
    .A2(_02850_),
    .A1(_02837_));
 sg13g2_nand3_1 _22907_ (.B(_02882_),
    .C(_02877_),
    .A(_02868_),
    .Y(_02885_));
 sg13g2_nor2b_1 _22908_ (.A(_02884_),
    .B_N(_02885_),
    .Y(_02886_));
 sg13g2_xnor2_1 _22909_ (.Y(_02887_),
    .A(_02824_),
    .B(_02886_));
 sg13g2_nor3_1 _22910_ (.A(_02704_),
    .B(_02770_),
    .C(net189),
    .Y(_02888_));
 sg13g2_buf_1 _22911_ (.A(_02828_),
    .X(_02889_));
 sg13g2_nand3_1 _22912_ (.B(_02701_),
    .C(net186),
    .A(_02699_),
    .Y(_02890_));
 sg13g2_a21oi_1 _22913_ (.A1(net221),
    .A2(net195),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_buf_1 _22914_ (.A(_02472_),
    .X(_02892_));
 sg13g2_a21o_1 _22915_ (.A2(_02554_),
    .A1(_02551_),
    .B1(_02559_),
    .X(_02893_));
 sg13g2_buf_2 _22916_ (.A(_02893_),
    .X(_02894_));
 sg13g2_a221oi_1 _22917_ (.B2(_02725_),
    .C1(_02894_),
    .B1(_02723_),
    .A1(net248),
    .Y(_02895_),
    .A2(net270));
 sg13g2_buf_1 _22918_ (.A(_02895_),
    .X(_02896_));
 sg13g2_nand2_1 _22919_ (.Y(_02897_),
    .A(_02805_),
    .B(net291));
 sg13g2_nand2_1 _22920_ (.Y(_02898_),
    .A(_02551_),
    .B(_02554_));
 sg13g2_a221oi_1 _22921_ (.B2(_02898_),
    .C1(net271),
    .B1(_02897_),
    .A1(_02763_),
    .Y(_02899_),
    .A2(_02765_));
 sg13g2_buf_1 _22922_ (.A(_02899_),
    .X(_02900_));
 sg13g2_nor3_1 _22923_ (.A(_02743_),
    .B(_02896_),
    .C(_02900_),
    .Y(_02901_));
 sg13g2_nor3_1 _22924_ (.A(_02888_),
    .B(_02891_),
    .C(_02901_),
    .Y(_02902_));
 sg13g2_nand2_1 _22925_ (.Y(_02903_),
    .A(_02733_),
    .B(_02839_));
 sg13g2_and2_1 _22926_ (.A(_02672_),
    .B(net222),
    .X(_02904_));
 sg13g2_xnor2_1 _22927_ (.Y(_02905_),
    .A(net251),
    .B(net250));
 sg13g2_a22oi_1 _22928_ (.Y(_02906_),
    .B1(_02905_),
    .B2(_02728_),
    .A2(_02904_),
    .A1(net190));
 sg13g2_nand2b_1 _22929_ (.Y(_02907_),
    .B(net188),
    .A_N(_02906_));
 sg13g2_o21ai_1 _22930_ (.B1(_02907_),
    .Y(_02908_),
    .A1(_02902_),
    .A2(_02903_));
 sg13g2_a21oi_1 _22931_ (.A1(net145),
    .A2(_02802_),
    .Y(_02909_),
    .B1(_02851_));
 sg13g2_nand2_1 _22932_ (.Y(_02910_),
    .A(_02692_),
    .B(_02845_));
 sg13g2_nor2b_1 _22933_ (.A(_02909_),
    .B_N(_02910_),
    .Y(_02911_));
 sg13g2_a22oi_1 _22934_ (.Y(_02912_),
    .B1(_02908_),
    .B2(_02911_),
    .A2(net187),
    .A1(net143));
 sg13g2_buf_1 _22935_ (.A(_02672_),
    .X(_02913_));
 sg13g2_buf_1 _22936_ (.A(_02675_),
    .X(_02914_));
 sg13g2_nor2_1 _22937_ (.A(net220),
    .B(net219),
    .Y(_02915_));
 sg13g2_and3_1 _22938_ (.X(_02916_),
    .A(_02777_),
    .B(_02671_),
    .C(_02678_));
 sg13g2_buf_1 _22939_ (.A(_02916_),
    .X(_02917_));
 sg13g2_nand2b_1 _22940_ (.Y(_02918_),
    .B(net227),
    .A_N(net200));
 sg13g2_nor2_1 _22941_ (.A(net253),
    .B(net250),
    .Y(_02919_));
 sg13g2_nand4_1 _22942_ (.B(_02674_),
    .C(net200),
    .A(net202),
    .Y(_02920_),
    .D(_02919_));
 sg13g2_or2_1 _22943_ (.X(_02921_),
    .B(net222),
    .A(net252));
 sg13g2_o21ai_1 _22944_ (.B1(_02864_),
    .Y(_02922_),
    .A1(_02921_),
    .A2(net219));
 sg13g2_a22oi_1 _22945_ (.Y(_02923_),
    .B1(_02864_),
    .B2(net190),
    .A2(_02751_),
    .A1(net200));
 sg13g2_and4_1 _22946_ (.A(_02918_),
    .B(_02920_),
    .C(_02922_),
    .D(_02923_),
    .X(_02924_));
 sg13g2_buf_1 _22947_ (.A(_02924_),
    .X(_02925_));
 sg13g2_buf_1 _22948_ (.A(_02925_),
    .X(_02926_));
 sg13g2_nand4_1 _22949_ (.B(_02915_),
    .C(_02917_),
    .A(_02861_),
    .Y(_02927_),
    .D(net106));
 sg13g2_nor4_1 _22950_ (.A(_02706_),
    .B(_02456_),
    .C(_02851_),
    .D(net142),
    .Y(_02928_));
 sg13g2_and2_1 _22951_ (.A(_02828_),
    .B(net223),
    .X(_02929_));
 sg13g2_buf_2 _22952_ (.A(_02929_),
    .X(_02930_));
 sg13g2_a221oi_1 _22953_ (.B2(_02930_),
    .C1(net224),
    .B1(_02928_),
    .A1(net121),
    .Y(_02931_),
    .A2(_02873_));
 sg13g2_and2_1 _22954_ (.A(net142),
    .B(net165),
    .X(_02932_));
 sg13g2_buf_1 _22955_ (.A(_02889_),
    .X(_02933_));
 sg13g2_nor4_1 _22956_ (.A(net167),
    .B(_02860_),
    .C(net185),
    .D(net165),
    .Y(_02934_));
 sg13g2_a221oi_1 _22957_ (.B2(net165),
    .C1(net144),
    .B1(net195),
    .A1(_02825_),
    .Y(_02935_),
    .A2(_02826_));
 sg13g2_nor4_1 _22958_ (.A(_02734_),
    .B(_02932_),
    .C(_02934_),
    .D(_02935_),
    .Y(_02936_));
 sg13g2_nand2_1 _22959_ (.Y(_02937_),
    .A(_02721_),
    .B(net222));
 sg13g2_o21ai_1 _22960_ (.B1(_02937_),
    .Y(_02938_),
    .A1(_02931_),
    .A2(_02936_));
 sg13g2_a21oi_1 _22961_ (.A1(_02912_),
    .A2(_02927_),
    .Y(_02939_),
    .B1(_02938_));
 sg13g2_xnor2_1 _22962_ (.Y(_02940_),
    .A(_02868_),
    .B(_02882_));
 sg13g2_xnor2_1 _22963_ (.Y(_02941_),
    .A(_02877_),
    .B(_02940_));
 sg13g2_a21oi_1 _22964_ (.A1(_02837_),
    .A2(_02850_),
    .Y(_02942_),
    .B1(_02941_));
 sg13g2_and3_1 _22965_ (.X(_02943_),
    .A(_02837_),
    .B(_02850_),
    .C(_02941_));
 sg13g2_nor3_1 _22966_ (.A(_02939_),
    .B(_02942_),
    .C(_02943_),
    .Y(_02944_));
 sg13g2_o21ai_1 _22967_ (.B1(_02840_),
    .Y(_02945_),
    .A1(_02712_),
    .A2(_02832_));
 sg13g2_nand2b_1 _22968_ (.Y(_02946_),
    .B(_02945_),
    .A_N(_02841_));
 sg13g2_nand2_1 _22969_ (.Y(_02947_),
    .A(net147),
    .B(net143));
 sg13g2_nand3b_1 _22970_ (.B(_02910_),
    .C(_02947_),
    .Y(_02948_),
    .A_N(_02909_));
 sg13g2_xnor2_1 _22971_ (.Y(_02949_),
    .A(_02908_),
    .B(_02948_));
 sg13g2_nor2b_1 _22972_ (.A(_02946_),
    .B_N(_02949_),
    .Y(_02950_));
 sg13g2_nand2b_1 _22973_ (.Y(_02951_),
    .B(_02837_),
    .A_N(_02841_));
 sg13g2_mux2_1 _22974_ (.A0(_02951_),
    .A1(_02842_),
    .S(_02849_),
    .X(_02952_));
 sg13g2_nand2b_1 _22975_ (.Y(_02953_),
    .B(_02849_),
    .A_N(_02837_));
 sg13g2_xnor2_1 _22976_ (.Y(_02954_),
    .A(_02938_),
    .B(_02927_));
 sg13g2_xnor2_1 _22977_ (.Y(_02955_),
    .A(_02912_),
    .B(_02954_));
 sg13g2_nand3_1 _22978_ (.B(_02953_),
    .C(_02955_),
    .A(_02952_),
    .Y(_02956_));
 sg13g2_a21oi_1 _22979_ (.A1(_02952_),
    .A2(_02953_),
    .Y(_02957_),
    .B1(_02955_));
 sg13g2_a21oi_1 _22980_ (.A1(_02950_),
    .A2(_02956_),
    .Y(_02958_),
    .B1(_02957_));
 sg13g2_o21ai_1 _22981_ (.B1(_02939_),
    .Y(_02959_),
    .A1(_02942_),
    .A2(_02943_));
 sg13g2_o21ai_1 _22982_ (.B1(_02959_),
    .Y(_02960_),
    .A1(_02944_),
    .A2(_02958_));
 sg13g2_buf_1 _22983_ (.A(_02960_),
    .X(_02961_));
 sg13g2_nand2b_1 _22984_ (.Y(_02962_),
    .B(_02961_),
    .A_N(_02887_));
 sg13g2_and2_1 _22985_ (.A(_02878_),
    .B(_02883_),
    .X(_02963_));
 sg13g2_nor2_1 _22986_ (.A(_02868_),
    .B(_02877_),
    .Y(_02964_));
 sg13g2_a21o_1 _22987_ (.A2(_02881_),
    .A1(_02879_),
    .B1(_02834_),
    .X(_02965_));
 sg13g2_o21ai_1 _22988_ (.B1(_02965_),
    .Y(_02966_),
    .A1(_02824_),
    .A2(_02964_));
 sg13g2_nand2_1 _22989_ (.Y(_02967_),
    .A(_02824_),
    .B(_02878_));
 sg13g2_nand2_1 _22990_ (.Y(_02968_),
    .A(_02837_),
    .B(_02850_));
 sg13g2_a21oi_1 _22991_ (.A1(_02966_),
    .A2(_02967_),
    .Y(_02969_),
    .B1(_02968_));
 sg13g2_a21oi_1 _22992_ (.A1(_02824_),
    .A2(_02963_),
    .Y(_02970_),
    .B1(_02969_));
 sg13g2_nand2b_1 _22993_ (.Y(_02971_),
    .B(_02812_),
    .A_N(_02970_));
 sg13g2_nand2_1 _22994_ (.Y(_02972_),
    .A(_02962_),
    .B(_02971_));
 sg13g2_xor2_1 _22995_ (.B(_02961_),
    .A(_02887_),
    .X(_02973_));
 sg13g2_buf_1 _22996_ (.A(_02973_),
    .X(_02974_));
 sg13g2_and2_1 _22997_ (.A(_02952_),
    .B(_02953_),
    .X(_02975_));
 sg13g2_xnor2_1 _22998_ (.Y(_02976_),
    .A(_02950_),
    .B(_02955_));
 sg13g2_xnor2_1 _22999_ (.Y(_02977_),
    .A(_02975_),
    .B(_02976_));
 sg13g2_buf_2 _23000_ (.A(_02977_),
    .X(_02978_));
 sg13g2_and2_1 _23001_ (.A(net144),
    .B(net200),
    .X(_02979_));
 sg13g2_nor2_1 _23002_ (.A(net224),
    .B(_02860_),
    .Y(_02980_));
 sg13g2_buf_1 _23003_ (.A(net219),
    .X(_02981_));
 sg13g2_a22oi_1 _23004_ (.Y(_02982_),
    .B1(_02858_),
    .B2(_02981_),
    .A2(net165),
    .A1(net144));
 sg13g2_a221oi_1 _23005_ (.B2(_02980_),
    .C1(_02982_),
    .B1(_02979_),
    .A1(net224),
    .Y(_02983_),
    .A2(net185));
 sg13g2_buf_1 _23006_ (.A(_02983_),
    .X(_02984_));
 sg13g2_or2_1 _23007_ (.X(_02985_),
    .B(_02830_),
    .A(_02790_));
 sg13g2_buf_1 _23008_ (.A(_02985_),
    .X(_02986_));
 sg13g2_or2_1 _23009_ (.X(_02987_),
    .B(_02900_),
    .A(_02896_));
 sg13g2_buf_8 _23010_ (.A(_02987_),
    .X(_02988_));
 sg13g2_nor2_1 _23011_ (.A(_02988_),
    .B(_02880_),
    .Y(_02989_));
 sg13g2_xnor2_1 _23012_ (.Y(_02990_),
    .A(_02914_),
    .B(net223));
 sg13g2_buf_1 _23013_ (.A(_02990_),
    .X(_02991_));
 sg13g2_nor2_1 _23014_ (.A(net198),
    .B(_02991_),
    .Y(_02992_));
 sg13g2_nor2_1 _23015_ (.A(net229),
    .B(_02829_),
    .Y(_02993_));
 sg13g2_nor2_1 _23016_ (.A(_02455_),
    .B(net186),
    .Y(_02994_));
 sg13g2_mux2_1 _23017_ (.A0(_02993_),
    .A1(_02994_),
    .S(_02930_),
    .X(_02995_));
 sg13g2_nor4_1 _23018_ (.A(_02710_),
    .B(net168),
    .C(_02991_),
    .D(_02988_),
    .Y(_02996_));
 sg13g2_a221oi_1 _23019_ (.B2(_02995_),
    .C1(_02996_),
    .B1(_02992_),
    .A1(_02986_),
    .Y(_02997_),
    .A2(_02989_));
 sg13g2_and2_1 _23020_ (.A(_02438_),
    .B(_02450_),
    .X(_02998_));
 sg13g2_a221oi_1 _23021_ (.B2(_02998_),
    .C1(_02420_),
    .B1(_02426_),
    .A1(_02699_),
    .Y(_02999_),
    .A2(_02701_));
 sg13g2_buf_2 _23022_ (.A(_02999_),
    .X(_03000_));
 sg13g2_a21oi_1 _23023_ (.A1(net185),
    .A2(_03000_),
    .Y(_03001_),
    .B1(_02979_));
 sg13g2_or3_1 _23024_ (.A(net121),
    .B(net145),
    .C(_03001_),
    .X(_03002_));
 sg13g2_nand2_1 _23025_ (.Y(_03003_),
    .A(_02783_),
    .B(_02933_));
 sg13g2_o21ai_1 _23026_ (.B1(_03003_),
    .Y(_03004_),
    .A1(_02861_),
    .A2(net145));
 sg13g2_nand3_1 _23027_ (.B(_02616_),
    .C(net221),
    .A(net229),
    .Y(_03005_));
 sg13g2_a21oi_1 _23028_ (.A1(_02857_),
    .A2(_03005_),
    .Y(_03006_),
    .B1(net188));
 sg13g2_a21oi_1 _23029_ (.A1(_02714_),
    .A2(_03004_),
    .Y(_03007_),
    .B1(_03006_));
 sg13g2_a21oi_1 _23030_ (.A1(_02997_),
    .A2(_03002_),
    .Y(_03008_),
    .B1(_03007_));
 sg13g2_buf_1 _23031_ (.A(_02894_),
    .X(_03009_));
 sg13g2_buf_1 _23032_ (.A(net247),
    .X(_03010_));
 sg13g2_xnor2_1 _23033_ (.Y(_03011_),
    .A(net218),
    .B(net121));
 sg13g2_and2_1 _23034_ (.A(_02919_),
    .B(_03011_),
    .X(_03012_));
 sg13g2_nand2_1 _23035_ (.Y(_03013_),
    .A(_02801_),
    .B(_03012_));
 sg13g2_nand2_1 _23036_ (.Y(_03014_),
    .A(net271),
    .B(_02894_));
 sg13g2_nor4_2 _23037_ (.A(net166),
    .B(_02933_),
    .C(_02743_),
    .Y(_03015_),
    .D(_03014_));
 sg13g2_a21oi_1 _23038_ (.A1(_03008_),
    .A2(_03013_),
    .Y(_03016_),
    .B1(_03015_));
 sg13g2_nor2_1 _23039_ (.A(_02984_),
    .B(_03016_),
    .Y(_03017_));
 sg13g2_inv_1 _23040_ (.Y(_03018_),
    .A(_03017_));
 sg13g2_xor2_1 _23041_ (.B(_02949_),
    .A(_02946_),
    .X(_03019_));
 sg13g2_o21ai_1 _23042_ (.B1(_03015_),
    .Y(_03020_),
    .A1(net122),
    .A2(_02873_));
 sg13g2_mux2_1 _23043_ (.A0(_03015_),
    .A1(_03020_),
    .S(_02984_),
    .X(_03021_));
 sg13g2_nor2_1 _23044_ (.A(_02617_),
    .B(_02873_),
    .Y(_03022_));
 sg13g2_buf_2 _23045_ (.A(_03022_),
    .X(_03023_));
 sg13g2_nand2b_1 _23046_ (.Y(_03024_),
    .B(_03023_),
    .A_N(_02984_));
 sg13g2_o21ai_1 _23047_ (.B1(_03024_),
    .Y(_03025_),
    .A1(_03012_),
    .A2(_03021_));
 sg13g2_xnor2_1 _23048_ (.Y(_03026_),
    .A(_03008_),
    .B(_03025_));
 sg13g2_nand2_1 _23049_ (.Y(_03027_),
    .A(_03019_),
    .B(_03026_));
 sg13g2_nor2_1 _23050_ (.A(_02888_),
    .B(_02891_),
    .Y(_03028_));
 sg13g2_xnor2_1 _23051_ (.Y(_03029_),
    .A(_03028_),
    .B(_02901_));
 sg13g2_xnor2_1 _23052_ (.Y(_03030_),
    .A(_02903_),
    .B(_03029_));
 sg13g2_a22oi_1 _23053_ (.Y(_03031_),
    .B1(net195),
    .B2(net194),
    .A2(net186),
    .A1(_02616_));
 sg13g2_nor3_1 _23054_ (.A(net168),
    .B(_02981_),
    .C(_03031_),
    .Y(_03032_));
 sg13g2_o21ai_1 _23055_ (.B1(net168),
    .Y(_03033_),
    .A1(net195),
    .A2(_02871_));
 sg13g2_nand2_1 _23056_ (.Y(_03034_),
    .A(_02456_),
    .B(_03033_));
 sg13g2_o21ai_1 _23057_ (.B1(_03034_),
    .Y(_03035_),
    .A1(_03006_),
    .A2(_03032_));
 sg13g2_xor2_1 _23058_ (.B(_03035_),
    .A(_02997_),
    .X(_03036_));
 sg13g2_o21ai_1 _23059_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_02406_),
    .A2(_03030_));
 sg13g2_buf_1 _23060_ (.A(_02763_),
    .X(_03038_));
 sg13g2_nand2_1 _23061_ (.Y(_03039_),
    .A(net246),
    .B(_02765_));
 sg13g2_buf_1 _23062_ (.A(_03039_),
    .X(_03040_));
 sg13g2_buf_8 _23063_ (.A(_02765_),
    .X(_03041_));
 sg13g2_nor2_1 _23064_ (.A(net246),
    .B(net269),
    .Y(_03042_));
 sg13g2_buf_2 _23065_ (.A(_03042_),
    .X(_03043_));
 sg13g2_a22oi_1 _23066_ (.Y(_03044_),
    .B1(_02777_),
    .B2(_03043_),
    .A2(_03009_),
    .A1(net183));
 sg13g2_nand3_1 _23067_ (.B(net246),
    .C(net269),
    .A(_02684_),
    .Y(_03045_));
 sg13g2_o21ai_1 _23068_ (.B1(_03045_),
    .Y(_03046_),
    .A1(net169),
    .A2(_03044_));
 sg13g2_nand2_1 _23069_ (.Y(_03047_),
    .A(_02733_),
    .B(_03046_));
 sg13g2_buf_1 _23070_ (.A(net270),
    .X(_03048_));
 sg13g2_buf_1 _23071_ (.A(net245),
    .X(_03049_));
 sg13g2_nor3_1 _23072_ (.A(net199),
    .B(net217),
    .C(_02688_),
    .Y(_03050_));
 sg13g2_buf_2 _23073_ (.A(_03050_),
    .X(_03051_));
 sg13g2_nor2_1 _23074_ (.A(net190),
    .B(_03051_),
    .Y(_03052_));
 sg13g2_o21ai_1 _23075_ (.B1(_03052_),
    .Y(_03053_),
    .A1(net224),
    .A2(_02913_));
 sg13g2_nand3_1 _23076_ (.B(net270),
    .C(net285),
    .A(net271),
    .Y(_03054_));
 sg13g2_buf_1 _23077_ (.A(_03054_),
    .X(_03055_));
 sg13g2_and3_1 _23078_ (.X(_03056_),
    .A(_03045_),
    .B(_03053_),
    .C(_03055_));
 sg13g2_xor2_1 _23079_ (.B(_02992_),
    .A(_02995_),
    .X(_03057_));
 sg13g2_mux2_1 _23080_ (.A0(_03047_),
    .A1(_03056_),
    .S(_03057_),
    .X(_03058_));
 sg13g2_nor3_1 _23081_ (.A(_02406_),
    .B(_03030_),
    .C(_03036_),
    .Y(_03059_));
 sg13g2_a21oi_1 _23082_ (.A1(_03037_),
    .A2(_03058_),
    .Y(_03060_),
    .B1(_03059_));
 sg13g2_nor2_1 _23083_ (.A(_03019_),
    .B(_03026_),
    .Y(_03061_));
 sg13g2_a21oi_1 _23084_ (.A1(_03027_),
    .A2(_03060_),
    .Y(_03062_),
    .B1(_03061_));
 sg13g2_buf_2 _23085_ (.A(_03062_),
    .X(_03063_));
 sg13g2_nand2_1 _23086_ (.Y(_03064_),
    .A(_03018_),
    .B(_03063_));
 sg13g2_nor2_1 _23087_ (.A(_03018_),
    .B(_03063_),
    .Y(_03065_));
 sg13g2_a21oi_1 _23088_ (.A1(_02978_),
    .A2(_03064_),
    .Y(_03066_),
    .B1(_03065_));
 sg13g2_buf_1 _23089_ (.A(net169),
    .X(_03067_));
 sg13g2_buf_1 _23090_ (.A(net274),
    .X(_03068_));
 sg13g2_buf_1 _23091_ (.A(net244),
    .X(_03069_));
 sg13g2_buf_1 _23092_ (.A(_02917_),
    .X(_03070_));
 sg13g2_nand2_1 _23093_ (.Y(_03071_),
    .A(net96),
    .B(net106));
 sg13g2_nor4_1 _23094_ (.A(_03067_),
    .B(_03069_),
    .C(_03010_),
    .D(_03071_),
    .Y(_03072_));
 sg13g2_buf_1 _23095_ (.A(net184),
    .X(_03073_));
 sg13g2_buf_1 _23096_ (.A(net220),
    .X(_03074_));
 sg13g2_nor2_1 _23097_ (.A(net182),
    .B(_02679_),
    .Y(_03075_));
 sg13g2_nor2_1 _23098_ (.A(net253),
    .B(net248),
    .Y(_03076_));
 sg13g2_nand2_1 _23099_ (.Y(_03077_),
    .A(_02801_),
    .B(_03076_));
 sg13g2_nand2_1 _23100_ (.Y(_03078_),
    .A(_03075_),
    .B(_03077_));
 sg13g2_buf_1 _23101_ (.A(net271),
    .X(_03079_));
 sg13g2_buf_1 _23102_ (.A(net243),
    .X(_03080_));
 sg13g2_buf_1 _23103_ (.A(net215),
    .X(_03081_));
 sg13g2_nand4_1 _23104_ (.B(_02920_),
    .C(_02922_),
    .A(_02918_),
    .Y(_03082_),
    .D(_02923_));
 sg13g2_buf_1 _23105_ (.A(_03082_),
    .X(_03083_));
 sg13g2_nor3_1 _23106_ (.A(net181),
    .B(_03073_),
    .C(net120),
    .Y(_03084_));
 sg13g2_nor2_1 _23107_ (.A(net106),
    .B(_03075_),
    .Y(_03085_));
 sg13g2_a221oi_1 _23108_ (.B2(_03075_),
    .C1(_03085_),
    .B1(_03084_),
    .A1(_03073_),
    .Y(_03086_),
    .A2(_03078_));
 sg13g2_nand3b_1 _23109_ (.B(_02746_),
    .C(net229),
    .Y(_03087_),
    .A_N(_02727_));
 sg13g2_nand3_1 _23110_ (.B(_02727_),
    .C(net187),
    .A(net221),
    .Y(_03088_));
 sg13g2_nor4_2 _23111_ (.A(_02421_),
    .B(_02452_),
    .C(_02716_),
    .Y(_03089_),
    .D(_02718_));
 sg13g2_nand2_1 _23112_ (.Y(_03090_),
    .A(net221),
    .B(_03089_));
 sg13g2_nor2b_2 _23113_ (.A(net222),
    .B_N(_02675_),
    .Y(_03091_));
 sg13g2_nor2b_1 _23114_ (.A(net219),
    .B_N(net222),
    .Y(_03092_));
 sg13g2_a22oi_1 _23115_ (.Y(_03093_),
    .B1(_03092_),
    .B2(net187),
    .A2(_03091_),
    .A1(_02615_));
 sg13g2_and4_1 _23116_ (.A(_03087_),
    .B(_03088_),
    .C(_03090_),
    .D(_03093_),
    .X(_03094_));
 sg13g2_a221oi_1 _23117_ (.B2(_02826_),
    .C1(net251),
    .B1(_02825_),
    .A1(_02755_),
    .Y(_03095_),
    .A2(_02756_));
 sg13g2_nor3_1 _23118_ (.A(_02703_),
    .B(net187),
    .C(_03095_),
    .Y(_03096_));
 sg13g2_nor4_1 _23119_ (.A(_02782_),
    .B(_02454_),
    .C(_02769_),
    .D(_02871_),
    .Y(_03097_));
 sg13g2_nor3_1 _23120_ (.A(net225),
    .B(_02548_),
    .C(net187),
    .Y(_03098_));
 sg13g2_a21o_1 _23121_ (.A2(net187),
    .A1(net225),
    .B1(net252),
    .X(_03099_));
 sg13g2_nor4_2 _23122_ (.A(_03096_),
    .B(_03097_),
    .C(_03098_),
    .Y(_03100_),
    .D(_03099_));
 sg13g2_nand2b_1 _23123_ (.Y(_03101_),
    .B(_03100_),
    .A_N(_03094_));
 sg13g2_xnor2_1 _23124_ (.Y(_03102_),
    .A(net167),
    .B(net195));
 sg13g2_nand2_1 _23125_ (.Y(_03103_),
    .A(_03102_),
    .B(_03095_));
 sg13g2_nand2_1 _23126_ (.Y(_03104_),
    .A(_03101_),
    .B(_03103_));
 sg13g2_nor2_1 _23127_ (.A(_02873_),
    .B(_02988_),
    .Y(_03105_));
 sg13g2_and2_1 _23128_ (.A(net222),
    .B(_02914_),
    .X(_03106_));
 sg13g2_nand2b_1 _23129_ (.Y(_03107_),
    .B(_03106_),
    .A_N(_02728_));
 sg13g2_nand2_1 _23130_ (.Y(_03108_),
    .A(_02853_),
    .B(_03107_));
 sg13g2_nor3_1 _23131_ (.A(_02705_),
    .B(net167),
    .C(_02906_),
    .Y(_03109_));
 sg13g2_a221oi_1 _23132_ (.B2(_02792_),
    .C1(_03109_),
    .B1(_03108_),
    .A1(_02839_),
    .Y(_03110_),
    .A2(_03105_));
 sg13g2_nor2_1 _23133_ (.A(net196),
    .B(_02871_),
    .Y(_03111_));
 sg13g2_a21oi_1 _23134_ (.A1(net196),
    .A2(_02856_),
    .Y(_03112_),
    .B1(_02760_));
 sg13g2_o21ai_1 _23135_ (.B1(_02731_),
    .Y(_03113_),
    .A1(_03111_),
    .A2(_03112_));
 sg13g2_mux2_1 _23136_ (.A0(_02856_),
    .A1(net221),
    .S(_02721_),
    .X(_03114_));
 sg13g2_o21ai_1 _23137_ (.B1(_02889_),
    .Y(_03115_),
    .A1(net188),
    .A2(net203));
 sg13g2_a22oi_1 _23138_ (.Y(_03116_),
    .B1(_03114_),
    .B2(_03115_),
    .A2(_03091_),
    .A1(net203));
 sg13g2_nand2_1 _23139_ (.Y(_03117_),
    .A(net168),
    .B(net221));
 sg13g2_a21o_1 _23140_ (.A2(_02937_),
    .A1(net143),
    .B1(_03117_),
    .X(_03118_));
 sg13g2_nand3_1 _23141_ (.B(_03116_),
    .C(_03118_),
    .A(_03113_),
    .Y(_03119_));
 sg13g2_xnor2_1 _23142_ (.Y(_03120_),
    .A(_03110_),
    .B(_03119_));
 sg13g2_nor2b_1 _23143_ (.A(_03110_),
    .B_N(_03119_),
    .Y(_03121_));
 sg13g2_a21oi_1 _23144_ (.A1(_03104_),
    .A2(_03120_),
    .Y(_03122_),
    .B1(_03121_));
 sg13g2_nor2_1 _23145_ (.A(_03074_),
    .B(net185),
    .Y(_03123_));
 sg13g2_nor2_1 _23146_ (.A(net247),
    .B(net184),
    .Y(_03124_));
 sg13g2_a221oi_1 _23147_ (.B2(_03124_),
    .C1(net181),
    .B1(net106),
    .A1(_02744_),
    .Y(_03125_),
    .A2(_03123_));
 sg13g2_nand3_1 _23148_ (.B(_02671_),
    .C(_02678_),
    .A(_02777_),
    .Y(_03126_));
 sg13g2_buf_1 _23149_ (.A(_03126_),
    .X(_03127_));
 sg13g2_buf_1 _23150_ (.A(_03127_),
    .X(_03128_));
 sg13g2_buf_1 _23151_ (.A(net269),
    .X(_03129_));
 sg13g2_nand3_1 _23152_ (.B(net220),
    .C(net184),
    .A(net242),
    .Y(_03130_));
 sg13g2_nand2b_1 _23153_ (.Y(_03131_),
    .B(_02688_),
    .A_N(net219));
 sg13g2_o21ai_1 _23154_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net95),
    .A2(_03130_));
 sg13g2_a21oi_1 _23155_ (.A1(net106),
    .A2(_03132_),
    .Y(_03133_),
    .B1(_03067_));
 sg13g2_nor2_1 _23156_ (.A(net169),
    .B(net184),
    .Y(_03134_));
 sg13g2_nand2b_1 _23157_ (.Y(_03135_),
    .B(_02925_),
    .A_N(_03134_));
 sg13g2_a22oi_1 _23158_ (.Y(_03136_),
    .B1(_03135_),
    .B2(net218),
    .A2(net95),
    .A1(net185));
 sg13g2_o21ai_1 _23159_ (.B1(_03136_),
    .Y(_03137_),
    .A1(_03125_),
    .A2(_03133_));
 sg13g2_nor2b_1 _23160_ (.A(_03122_),
    .B_N(_03137_),
    .Y(_03138_));
 sg13g2_a21oi_2 _23161_ (.B1(_03138_),
    .Y(_03139_),
    .A2(_03086_),
    .A1(_03072_));
 sg13g2_xor2_1 _23162_ (.B(_03026_),
    .A(_03019_),
    .X(_03140_));
 sg13g2_xnor2_1 _23163_ (.Y(_03141_),
    .A(_03060_),
    .B(_03140_));
 sg13g2_nor2_1 _23164_ (.A(_03139_),
    .B(_03141_),
    .Y(_03142_));
 sg13g2_nand2_1 _23165_ (.Y(_03143_),
    .A(_02710_),
    .B(_03041_));
 sg13g2_and2_1 _23166_ (.A(_02639_),
    .B(net285),
    .X(_03144_));
 sg13g2_buf_1 _23167_ (.A(_03144_),
    .X(_03145_));
 sg13g2_nand2_1 _23168_ (.Y(_03146_),
    .A(net198),
    .B(_03145_));
 sg13g2_nand3_1 _23169_ (.B(_03143_),
    .C(_03146_),
    .A(_03038_),
    .Y(_03147_));
 sg13g2_nand2_1 _23170_ (.Y(_03148_),
    .A(_02641_),
    .B(net269));
 sg13g2_a21oi_1 _23171_ (.A1(net217),
    .A2(_03148_),
    .Y(_03149_),
    .B1(net199));
 sg13g2_nand2_1 _23172_ (.Y(_03150_),
    .A(net270),
    .B(_02517_));
 sg13g2_buf_2 _23173_ (.A(_03150_),
    .X(_03151_));
 sg13g2_nand2_1 _23174_ (.Y(_03152_),
    .A(_02710_),
    .B(_03038_));
 sg13g2_a21oi_1 _23175_ (.A1(_03151_),
    .A2(_03152_),
    .Y(_03153_),
    .B1(net198));
 sg13g2_nand2_1 _23176_ (.Y(_03154_),
    .A(_02685_),
    .B(_02777_));
 sg13g2_nor2_1 _23177_ (.A(net270),
    .B(net285),
    .Y(_03155_));
 sg13g2_buf_2 _23178_ (.A(_03155_),
    .X(_03156_));
 sg13g2_o21ai_1 _23179_ (.B1(_03156_),
    .Y(_03157_),
    .A1(net227),
    .A2(net198));
 sg13g2_nor2_1 _23180_ (.A(net243),
    .B(_02743_),
    .Y(_03158_));
 sg13g2_o21ai_1 _23181_ (.B1(_03043_),
    .Y(_03159_),
    .A1(_02744_),
    .A2(_03158_));
 sg13g2_o21ai_1 _23182_ (.B1(_03159_),
    .Y(_03160_),
    .A1(_03154_),
    .A2(_03157_));
 sg13g2_a221oi_1 _23183_ (.B2(net215),
    .C1(_03160_),
    .B1(_03153_),
    .A1(_03147_),
    .Y(_03161_),
    .A2(_03149_));
 sg13g2_o21ai_1 _23184_ (.B1(net170),
    .Y(_03162_),
    .A1(_02790_),
    .A2(_02830_));
 sg13g2_and4_1 _23185_ (.A(net225),
    .B(net191),
    .C(_02828_),
    .D(net223),
    .X(_03163_));
 sg13g2_nor3_1 _23186_ (.A(_02780_),
    .B(_02666_),
    .C(_02894_),
    .Y(_03164_));
 sg13g2_o21ai_1 _23187_ (.B1(net250),
    .Y(_03165_),
    .A1(net287),
    .A2(net286));
 sg13g2_a221oi_1 _23188_ (.B2(_02769_),
    .C1(_03165_),
    .B1(_03164_),
    .A1(net225),
    .Y(_03166_),
    .A2(net223));
 sg13g2_and3_1 _23189_ (.X(_03167_),
    .A(_02769_),
    .B(_03165_),
    .C(_03164_));
 sg13g2_nor4_1 _23190_ (.A(net198),
    .B(net191),
    .C(_02769_),
    .D(net252),
    .Y(_03168_));
 sg13g2_nor4_1 _23191_ (.A(_03163_),
    .B(_03166_),
    .C(_03167_),
    .D(_03168_),
    .Y(_03169_));
 sg13g2_xnor2_1 _23192_ (.Y(_03170_),
    .A(_03162_),
    .B(_03169_));
 sg13g2_buf_1 _23193_ (.A(net246),
    .X(_03171_));
 sg13g2_nor2_1 _23194_ (.A(net188),
    .B(_03129_),
    .Y(_03172_));
 sg13g2_nand2_1 _23195_ (.Y(_03173_),
    .A(net193),
    .B(net215));
 sg13g2_nor2_1 _23196_ (.A(_02639_),
    .B(net285),
    .Y(_03174_));
 sg13g2_buf_1 _23197_ (.A(_03174_),
    .X(_03175_));
 sg13g2_nand3_1 _23198_ (.B(net169),
    .C(_03175_),
    .A(net188),
    .Y(_03176_));
 sg13g2_o21ai_1 _23199_ (.B1(_03176_),
    .Y(_03177_),
    .A1(_03172_),
    .A2(_03173_));
 sg13g2_nand2_1 _23200_ (.Y(_03178_),
    .A(_03171_),
    .B(_03177_));
 sg13g2_o21ai_1 _23201_ (.B1(_03178_),
    .Y(_03179_),
    .A1(_03161_),
    .A2(_03170_));
 sg13g2_nor2_1 _23202_ (.A(_02683_),
    .B(net270),
    .Y(_03180_));
 sg13g2_nand2_1 _23203_ (.Y(_03181_),
    .A(_03048_),
    .B(_03041_));
 sg13g2_nor2_1 _23204_ (.A(net220),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_a21oi_1 _23205_ (.A1(net183),
    .A2(_03055_),
    .Y(_03183_),
    .B1(net247));
 sg13g2_nor3_1 _23206_ (.A(net199),
    .B(net245),
    .C(net269),
    .Y(_03184_));
 sg13g2_and2_1 _23207_ (.A(net247),
    .B(_03184_),
    .X(_03185_));
 sg13g2_or3_1 _23208_ (.A(_03182_),
    .B(_03183_),
    .C(_03185_),
    .X(_03186_));
 sg13g2_nor2_1 _23209_ (.A(_02738_),
    .B(net193),
    .Y(_03187_));
 sg13g2_a22oi_1 _23210_ (.Y(_03188_),
    .B1(_03187_),
    .B2(net183),
    .A2(net247),
    .A1(net244));
 sg13g2_nor2_1 _23211_ (.A(net215),
    .B(_03188_),
    .Y(_03189_));
 sg13g2_a221oi_1 _23212_ (.B2(net193),
    .C1(_03189_),
    .B1(_03186_),
    .A1(_03180_),
    .Y(_03190_),
    .A2(_03175_));
 sg13g2_xnor2_1 _23213_ (.Y(_03191_),
    .A(_03057_),
    .B(_03190_));
 sg13g2_xnor2_1 _23214_ (.Y(_03192_),
    .A(_03104_),
    .B(_03120_));
 sg13g2_nand2_1 _23215_ (.Y(_03193_),
    .A(_03191_),
    .B(_03192_));
 sg13g2_nor2_1 _23216_ (.A(_03191_),
    .B(_03192_),
    .Y(_03194_));
 sg13g2_a21oi_1 _23217_ (.A1(_03179_),
    .A2(_03193_),
    .Y(_03195_),
    .B1(_03194_));
 sg13g2_nor2_1 _23218_ (.A(net254),
    .B(_03030_),
    .Y(_03196_));
 sg13g2_xor2_1 _23219_ (.B(_03058_),
    .A(_03036_),
    .X(_03197_));
 sg13g2_xnor2_1 _23220_ (.Y(_03198_),
    .A(_03196_),
    .B(_03197_));
 sg13g2_xor2_1 _23221_ (.B(_03137_),
    .A(_03122_),
    .X(_03199_));
 sg13g2_and2_1 _23222_ (.A(_03198_),
    .B(_03199_),
    .X(_03200_));
 sg13g2_or2_1 _23223_ (.X(_03201_),
    .B(_03199_),
    .A(_03198_));
 sg13g2_o21ai_1 _23224_ (.B1(_03201_),
    .Y(_03202_),
    .A1(_03195_),
    .A2(_03200_));
 sg13g2_nand2_1 _23225_ (.Y(_03203_),
    .A(_03139_),
    .B(_03141_));
 sg13g2_o21ai_1 _23226_ (.B1(_03203_),
    .Y(_03204_),
    .A1(_03142_),
    .A2(_03202_));
 sg13g2_buf_1 _23227_ (.A(_03204_),
    .X(_03205_));
 sg13g2_buf_1 _23228_ (.A(_03205_),
    .X(_03206_));
 sg13g2_nor2_1 _23229_ (.A(_02978_),
    .B(_03064_),
    .Y(_03207_));
 sg13g2_a21oi_2 _23230_ (.B1(_03207_),
    .Y(_03208_),
    .A2(net78),
    .A1(_03066_));
 sg13g2_nand2b_1 _23231_ (.Y(_03209_),
    .B(_02959_),
    .A_N(_02944_));
 sg13g2_xnor2_1 _23232_ (.Y(_03210_),
    .A(_02958_),
    .B(_03209_));
 sg13g2_buf_1 _23233_ (.A(_03210_),
    .X(_03211_));
 sg13g2_inv_1 _23234_ (.Y(_03212_),
    .A(net77));
 sg13g2_nand2_1 _23235_ (.Y(_03213_),
    .A(_03208_),
    .B(_03212_));
 sg13g2_nor2_1 _23236_ (.A(net74),
    .B(_03213_),
    .Y(_03214_));
 sg13g2_a21o_1 _23237_ (.A2(_02972_),
    .A1(_02813_),
    .B1(_03214_),
    .X(_03215_));
 sg13g2_nand3_1 _23238_ (.B(_02758_),
    .C(net243),
    .A(_02710_),
    .Y(_03216_));
 sg13g2_o21ai_1 _23239_ (.B1(_02454_),
    .Y(_03217_),
    .A1(net253),
    .A2(net245));
 sg13g2_nor2_1 _23240_ (.A(net225),
    .B(_02689_),
    .Y(_03218_));
 sg13g2_a22oi_1 _23241_ (.Y(_03219_),
    .B1(_03217_),
    .B2(_03218_),
    .A2(_03216_),
    .A1(net198));
 sg13g2_nand4_1 _23242_ (.B(_02758_),
    .C(net226),
    .A(net225),
    .Y(_03220_),
    .D(_03175_));
 sg13g2_a22oi_1 _23243_ (.Y(_03221_),
    .B1(_03145_),
    .B2(net226),
    .A2(_03175_),
    .A1(_02845_));
 sg13g2_a22oi_1 _23244_ (.Y(_03222_),
    .B1(_03076_),
    .B2(_02668_),
    .A2(_03000_),
    .A1(net253));
 sg13g2_nand3_1 _23245_ (.B(net226),
    .C(_02668_),
    .A(net227),
    .Y(_03223_));
 sg13g2_nand4_1 _23246_ (.B(_03221_),
    .C(_03222_),
    .A(_03220_),
    .Y(_03224_),
    .D(_03223_));
 sg13g2_and2_1 _23247_ (.A(net253),
    .B(_02765_),
    .X(_03225_));
 sg13g2_o21ai_1 _23248_ (.B1(_02703_),
    .Y(_03226_),
    .A1(_03048_),
    .A2(_03225_));
 sg13g2_a221oi_1 _23249_ (.B2(_03226_),
    .C1(net199),
    .B1(_03181_),
    .A1(_02755_),
    .Y(_03227_),
    .A2(_02756_));
 sg13g2_a221oi_1 _23250_ (.B2(net214),
    .C1(_03227_),
    .B1(_03224_),
    .A1(net274),
    .Y(_03228_),
    .A2(_03219_));
 sg13g2_buf_1 _23251_ (.A(_03228_),
    .X(_03229_));
 sg13g2_xor2_1 _23252_ (.B(net250),
    .A(_02673_),
    .X(_03230_));
 sg13g2_buf_1 _23253_ (.A(_03230_),
    .X(_03231_));
 sg13g2_nor2_1 _23254_ (.A(net201),
    .B(_03231_),
    .Y(_03232_));
 sg13g2_a221oi_1 _23255_ (.B2(_02765_),
    .C1(net271),
    .B1(_02763_),
    .A1(net249),
    .Y(_03233_),
    .A2(net275));
 sg13g2_mux2_1 _23256_ (.A0(_02547_),
    .A1(_03233_),
    .S(_03231_),
    .X(_03234_));
 sg13g2_mux2_1 _23257_ (.A0(_02720_),
    .A1(_02905_),
    .S(_02769_),
    .X(_03235_));
 sg13g2_mux2_1 _23258_ (.A0(_03234_),
    .A1(_03235_),
    .S(_02894_),
    .X(_03236_));
 sg13g2_nor2_1 _23259_ (.A(_02720_),
    .B(net245),
    .Y(_03237_));
 sg13g2_a21oi_1 _23260_ (.A1(_02699_),
    .A2(_02701_),
    .Y(_03238_),
    .B1(net248));
 sg13g2_xnor2_1 _23261_ (.Y(_03239_),
    .A(_02545_),
    .B(net285));
 sg13g2_nor3_1 _23262_ (.A(_03000_),
    .B(_03238_),
    .C(_03239_),
    .Y(_03240_));
 sg13g2_nor4_1 _23263_ (.A(_02454_),
    .B(_02720_),
    .C(net248),
    .D(_03151_),
    .Y(_03241_));
 sg13g2_a221oi_1 _23264_ (.B2(_03240_),
    .C1(_03241_),
    .B1(_03237_),
    .A1(_03156_),
    .Y(_03242_),
    .A2(net200));
 sg13g2_or3_1 _23265_ (.A(_03232_),
    .B(_03236_),
    .C(_03242_),
    .X(_03243_));
 sg13g2_buf_2 _23266_ (.A(_03243_),
    .X(_03244_));
 sg13g2_o21ai_1 _23267_ (.B1(_03242_),
    .Y(_03245_),
    .A1(_03232_),
    .A2(_03236_));
 sg13g2_buf_1 _23268_ (.A(_03245_),
    .X(_03246_));
 sg13g2_and3_1 _23269_ (.X(_03247_),
    .A(_03229_),
    .B(_03244_),
    .C(_03246_));
 sg13g2_buf_1 _23270_ (.A(_03247_),
    .X(_03248_));
 sg13g2_a21oi_1 _23271_ (.A1(_03244_),
    .A2(_03246_),
    .Y(_03249_),
    .B1(_03229_));
 sg13g2_nor2_1 _23272_ (.A(_03248_),
    .B(_03249_),
    .Y(_03250_));
 sg13g2_nand3_1 _23273_ (.B(net228),
    .C(_02668_),
    .A(_02547_),
    .Y(_03251_));
 sg13g2_buf_1 _23274_ (.A(_03251_),
    .X(_03252_));
 sg13g2_inv_1 _23275_ (.Y(_03253_),
    .A(_02593_));
 sg13g2_a221oi_1 _23276_ (.B2(_03253_),
    .C1(_02718_),
    .B1(net291),
    .A1(_02699_),
    .Y(_03254_),
    .A2(_02701_));
 sg13g2_nand2_1 _23277_ (.Y(_03255_),
    .A(net189),
    .B(_03254_));
 sg13g2_a221oi_1 _23278_ (.B2(_02769_),
    .C1(_03000_),
    .B1(_03254_),
    .A1(_02614_),
    .Y(_03256_),
    .A2(_02668_));
 sg13g2_nand3_1 _23279_ (.B(_03255_),
    .C(_03256_),
    .A(_03252_),
    .Y(_03257_));
 sg13g2_buf_1 _23280_ (.A(_03257_),
    .X(_03258_));
 sg13g2_nand2_1 _23281_ (.Y(_03259_),
    .A(net242),
    .B(net119));
 sg13g2_nor3_1 _23282_ (.A(net271),
    .B(_02892_),
    .C(net285),
    .Y(_03260_));
 sg13g2_buf_1 _23283_ (.A(_03260_),
    .X(_03261_));
 sg13g2_nor3_1 _23284_ (.A(_02421_),
    .B(_02452_),
    .C(net226),
    .Y(_03262_));
 sg13g2_a21oi_1 _23285_ (.A1(net228),
    .A2(_03261_),
    .Y(_03263_),
    .B1(_03262_));
 sg13g2_o21ai_1 _23286_ (.B1(net194),
    .Y(_03264_),
    .A1(_03261_),
    .A2(_03262_));
 sg13g2_nor2_1 _23287_ (.A(net226),
    .B(net252),
    .Y(_03265_));
 sg13g2_nand3_1 _23288_ (.B(_02871_),
    .C(_03265_),
    .A(_02759_),
    .Y(_03266_));
 sg13g2_o21ai_1 _23289_ (.B1(net220),
    .Y(_03267_),
    .A1(net229),
    .A2(_02685_));
 sg13g2_nand4_1 _23290_ (.B(_03264_),
    .C(_03266_),
    .A(net170),
    .Y(_03268_),
    .D(_03267_));
 sg13g2_o21ai_1 _23291_ (.B1(_03268_),
    .Y(_03269_),
    .A1(net170),
    .A2(_03263_));
 sg13g2_xnor2_1 _23292_ (.Y(_03270_),
    .A(_03259_),
    .B(_03269_));
 sg13g2_buf_2 _23293_ (.A(_03270_),
    .X(_03271_));
 sg13g2_a21oi_1 _23294_ (.A1(net273),
    .A2(net272),
    .Y(_03272_),
    .B1(_02767_));
 sg13g2_nor4_1 _23295_ (.A(_02892_),
    .B(_02561_),
    .C(_02673_),
    .D(net250),
    .Y(_03273_));
 sg13g2_mux2_1 _23296_ (.A0(_03089_),
    .A1(_03272_),
    .S(_03273_),
    .X(_03274_));
 sg13g2_nand3_1 _23297_ (.B(_02687_),
    .C(net189),
    .A(_02720_),
    .Y(_03275_));
 sg13g2_a221oi_1 _23298_ (.B2(_02614_),
    .C1(net226),
    .B1(net228),
    .A1(_02758_),
    .Y(_03276_),
    .A2(net269));
 sg13g2_o21ai_1 _23299_ (.B1(_02765_),
    .Y(_03277_),
    .A1(net287),
    .A2(net286));
 sg13g2_a221oi_1 _23300_ (.B2(net189),
    .C1(_03277_),
    .B1(net243),
    .A1(net249),
    .Y(_03278_),
    .A2(net275));
 sg13g2_a221oi_1 _23301_ (.B2(_03276_),
    .C1(_03278_),
    .B1(_03275_),
    .A1(net269),
    .Y(_03279_),
    .A2(_03274_));
 sg13g2_buf_1 _23302_ (.A(_03279_),
    .X(_03280_));
 sg13g2_nand3b_1 _23303_ (.B(net119),
    .C(_03171_),
    .Y(_03281_),
    .A_N(_03280_));
 sg13g2_nor2_1 _23304_ (.A(net199),
    .B(net274),
    .Y(_03282_));
 sg13g2_buf_2 _23305_ (.A(_03282_),
    .X(_03283_));
 sg13g2_xnor2_1 _23306_ (.Y(_03284_),
    .A(net196),
    .B(_02590_));
 sg13g2_nand3_1 _23307_ (.B(_03283_),
    .C(_03284_),
    .A(_02760_),
    .Y(_03285_));
 sg13g2_nand3_1 _23308_ (.B(_03281_),
    .C(_03285_),
    .A(net143),
    .Y(_03286_));
 sg13g2_buf_2 _23309_ (.A(_03286_),
    .X(_03287_));
 sg13g2_nor2_1 _23310_ (.A(_03271_),
    .B(_03287_),
    .Y(_03288_));
 sg13g2_nor2_1 _23311_ (.A(_02683_),
    .B(_02765_),
    .Y(_03289_));
 sg13g2_o21ai_1 _23312_ (.B1(_03000_),
    .Y(_03290_),
    .A1(_03261_),
    .A2(_03289_));
 sg13g2_nand3_1 _23313_ (.B(_02758_),
    .C(_03180_),
    .A(net225),
    .Y(_03291_));
 sg13g2_nor2_1 _23314_ (.A(net271),
    .B(net270),
    .Y(_03292_));
 sg13g2_nand3_1 _23315_ (.B(_02758_),
    .C(_03292_),
    .A(_02782_),
    .Y(_03293_));
 sg13g2_nor2_1 _23316_ (.A(net248),
    .B(_02763_),
    .Y(_03294_));
 sg13g2_nor3_1 _23317_ (.A(_02780_),
    .B(_02666_),
    .C(net248),
    .Y(_03295_));
 sg13g2_nor3_1 _23318_ (.A(net287),
    .B(net286),
    .C(_02687_),
    .Y(_03296_));
 sg13g2_nor3_1 _23319_ (.A(net248),
    .B(net246),
    .C(net285),
    .Y(_03297_));
 sg13g2_a221oi_1 _23320_ (.B2(_03296_),
    .C1(_03297_),
    .B1(_03295_),
    .A1(_02454_),
    .Y(_03298_),
    .A2(_03294_));
 sg13g2_and4_1 _23321_ (.A(_03290_),
    .B(_03291_),
    .C(_03293_),
    .D(_03298_),
    .X(_03299_));
 sg13g2_nor2_1 _23322_ (.A(net201),
    .B(net245),
    .Y(_03300_));
 sg13g2_nand4_1 _23323_ (.B(_02701_),
    .C(net273),
    .A(_02699_),
    .Y(_03301_),
    .D(net272));
 sg13g2_o21ai_1 _23324_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_02782_),
    .A2(_03277_));
 sg13g2_a21oi_1 _23325_ (.A1(_02699_),
    .A2(_02701_),
    .Y(_03303_),
    .B1(net245));
 sg13g2_a21oi_1 _23326_ (.A1(net249),
    .A2(net275),
    .Y(_03304_),
    .B1(net226));
 sg13g2_nor3_1 _23327_ (.A(net287),
    .B(net286),
    .C(net246),
    .Y(_03305_));
 sg13g2_nor4_1 _23328_ (.A(_03303_),
    .B(_03262_),
    .C(_03304_),
    .D(_03305_),
    .Y(_03306_));
 sg13g2_a22oi_1 _23329_ (.Y(_03307_),
    .B1(_03306_),
    .B2(net274),
    .A2(_03302_),
    .A1(_03300_));
 sg13g2_o21ai_1 _23330_ (.B1(_03307_),
    .Y(_03308_),
    .A1(net196),
    .A2(_03299_));
 sg13g2_buf_1 _23331_ (.A(_03308_),
    .X(_03309_));
 sg13g2_nor2_1 _23332_ (.A(_02548_),
    .B(_02745_),
    .Y(_03310_));
 sg13g2_xnor2_1 _23333_ (.Y(_03311_),
    .A(_03009_),
    .B(_03310_));
 sg13g2_nor3_1 _23334_ (.A(_02454_),
    .B(net245),
    .C(_03239_),
    .Y(_03312_));
 sg13g2_a21oi_1 _23335_ (.A1(_03045_),
    .A2(_03055_),
    .Y(_03313_),
    .B1(net196));
 sg13g2_o21ai_1 _23336_ (.B1(_02829_),
    .Y(_03314_),
    .A1(_03312_),
    .A2(_03313_));
 sg13g2_nor2_1 _23337_ (.A(net229),
    .B(net183),
    .Y(_03315_));
 sg13g2_nand2_1 _23338_ (.Y(_03316_),
    .A(net201),
    .B(_03315_));
 sg13g2_nand3_1 _23339_ (.B(_03314_),
    .C(_03316_),
    .A(_03311_),
    .Y(_03317_));
 sg13g2_a21oi_1 _23340_ (.A1(_03314_),
    .A2(_03316_),
    .Y(_03318_),
    .B1(_03311_));
 sg13g2_a21o_1 _23341_ (.A2(_03317_),
    .A1(_03309_),
    .B1(_03318_),
    .X(_03319_));
 sg13g2_buf_1 _23342_ (.A(_03319_),
    .X(_03320_));
 sg13g2_nor3_1 _23343_ (.A(_03248_),
    .B(_03249_),
    .C(_03320_),
    .Y(_03321_));
 sg13g2_a21oi_1 _23344_ (.A1(_03281_),
    .A2(_03285_),
    .Y(_03322_),
    .B1(net143));
 sg13g2_a21oi_1 _23345_ (.A1(_03271_),
    .A2(_03287_),
    .Y(_03323_),
    .B1(_03322_));
 sg13g2_nor3_1 _23346_ (.A(_03271_),
    .B(_03287_),
    .C(_03320_),
    .Y(_03324_));
 sg13g2_a221oi_1 _23347_ (.B2(_03323_),
    .C1(_03324_),
    .B1(_03321_),
    .A1(_03250_),
    .Y(_03325_),
    .A2(_03288_));
 sg13g2_buf_1 _23348_ (.A(_03325_),
    .X(_03326_));
 sg13g2_inv_1 _23349_ (.Y(_03327_),
    .A(_03326_));
 sg13g2_nor2_1 _23350_ (.A(_03049_),
    .B(net95),
    .Y(_03328_));
 sg13g2_nor2_1 _23351_ (.A(net244),
    .B(net120),
    .Y(_03329_));
 sg13g2_xnor2_1 _23352_ (.Y(_03330_),
    .A(_03328_),
    .B(_03329_));
 sg13g2_buf_2 _23353_ (.A(_03330_),
    .X(_03331_));
 sg13g2_nand3_1 _23354_ (.B(_03080_),
    .C(_03068_),
    .A(_02711_),
    .Y(_03332_));
 sg13g2_a22oi_1 _23355_ (.Y(_03333_),
    .B1(_03148_),
    .B2(_03332_),
    .A2(net165),
    .A1(_02774_));
 sg13g2_nand2_1 _23356_ (.Y(_03334_),
    .A(net144),
    .B(_02669_));
 sg13g2_a22oi_1 _23357_ (.Y(_03335_),
    .B1(_03143_),
    .B2(_03173_),
    .A2(_03252_),
    .A1(_03334_));
 sg13g2_nor4_1 _23358_ (.A(net193),
    .B(_03081_),
    .C(net214),
    .D(net244),
    .Y(_03336_));
 sg13g2_or4_1 _23359_ (.A(_03051_),
    .B(_03333_),
    .C(_03335_),
    .D(_03336_),
    .X(_03337_));
 sg13g2_buf_2 _23360_ (.A(_03337_),
    .X(_03338_));
 sg13g2_o21ai_1 _23361_ (.B1(_02758_),
    .Y(_03339_),
    .A1(_02614_),
    .A2(net228));
 sg13g2_mux2_1 _23362_ (.A0(_03295_),
    .A1(_03238_),
    .S(_03339_),
    .X(_03340_));
 sg13g2_a221oi_1 _23363_ (.B2(_02725_),
    .C1(net251),
    .B1(_02723_),
    .A1(_02545_),
    .Y(_03341_),
    .A2(net270));
 sg13g2_buf_1 _23364_ (.A(_03341_),
    .X(_03342_));
 sg13g2_or4_1 _23365_ (.A(_02758_),
    .B(net252),
    .C(net219),
    .D(_03342_),
    .X(_03343_));
 sg13g2_a21oi_1 _23366_ (.A1(net273),
    .A2(net272),
    .Y(_03344_),
    .B1(net252));
 sg13g2_nand3_1 _23367_ (.B(_03342_),
    .C(_03344_),
    .A(net201),
    .Y(_03345_));
 sg13g2_nor3_1 _23368_ (.A(net287),
    .B(net286),
    .C(net252),
    .Y(_03346_));
 sg13g2_and2_1 _23369_ (.A(_02581_),
    .B(_02586_),
    .X(_03347_));
 sg13g2_buf_1 _23370_ (.A(_03347_),
    .X(_03348_));
 sg13g2_a221oi_1 _23371_ (.B2(net275),
    .C1(_03348_),
    .B1(net249),
    .A1(_02403_),
    .Y(_03349_),
    .A2(net291));
 sg13g2_a221oi_1 _23372_ (.B2(_02826_),
    .C1(_02894_),
    .B1(_02825_),
    .A1(net249),
    .Y(_03350_),
    .A2(net275));
 sg13g2_a221oi_1 _23373_ (.B2(_03349_),
    .C1(_03350_),
    .B1(_03344_),
    .A1(_02720_),
    .Y(_03351_),
    .A2(_03346_));
 sg13g2_nand3_1 _23374_ (.B(_03345_),
    .C(_03351_),
    .A(_03343_),
    .Y(_03352_));
 sg13g2_xnor2_1 _23375_ (.Y(_03353_),
    .A(net167),
    .B(_03342_));
 sg13g2_and2_1 _23376_ (.A(net164),
    .B(_02915_),
    .X(_03354_));
 sg13g2_a22oi_1 _23377_ (.Y(_03355_),
    .B1(_03353_),
    .B2(_03354_),
    .A2(_03352_),
    .A1(_03340_));
 sg13g2_buf_2 _23378_ (.A(_03355_),
    .X(_03356_));
 sg13g2_xor2_1 _23379_ (.B(_03094_),
    .A(_03100_),
    .X(_03357_));
 sg13g2_buf_2 _23380_ (.A(_03357_),
    .X(_03358_));
 sg13g2_nand2_1 _23381_ (.Y(_03359_),
    .A(net220),
    .B(net219));
 sg13g2_nor2_1 _23382_ (.A(net202),
    .B(_03359_),
    .Y(_03360_));
 sg13g2_a21o_1 _23383_ (.A2(_02937_),
    .A1(_02759_),
    .B1(_02746_),
    .X(_03361_));
 sg13g2_a22oi_1 _23384_ (.Y(_03362_),
    .B1(_03361_),
    .B2(_02930_),
    .A2(_03360_),
    .A1(net187));
 sg13g2_buf_2 _23385_ (.A(_03362_),
    .X(_03363_));
 sg13g2_xor2_1 _23386_ (.B(_03363_),
    .A(_03358_),
    .X(_03364_));
 sg13g2_xnor2_1 _23387_ (.Y(_03365_),
    .A(_03356_),
    .B(_03364_));
 sg13g2_xnor2_1 _23388_ (.Y(_03366_),
    .A(_02455_),
    .B(net194));
 sg13g2_nor2_1 _23389_ (.A(net229),
    .B(_02894_),
    .Y(_03367_));
 sg13g2_a22oi_1 _23390_ (.Y(_03368_),
    .B1(_03367_),
    .B2(net190),
    .A2(_03366_),
    .A1(net223));
 sg13g2_nand2_1 _23391_ (.Y(_03369_),
    .A(net170),
    .B(_02839_));
 sg13g2_xnor2_1 _23392_ (.Y(_03370_),
    .A(_03368_),
    .B(_03369_));
 sg13g2_mux2_1 _23393_ (.A0(_03175_),
    .A1(_03145_),
    .S(net243),
    .X(_03371_));
 sg13g2_a22oi_1 _23394_ (.Y(_03372_),
    .B1(_03371_),
    .B2(net203),
    .A2(_03184_),
    .A1(_02710_));
 sg13g2_nor2_1 _23395_ (.A(_03148_),
    .B(_03272_),
    .Y(_03373_));
 sg13g2_a21o_1 _23396_ (.A2(net274),
    .A1(_02641_),
    .B1(net243),
    .X(_03374_));
 sg13g2_o21ai_1 _23397_ (.B1(_03374_),
    .Y(_03375_),
    .A1(net227),
    .A2(net188));
 sg13g2_a22oi_1 _23398_ (.Y(_03376_),
    .B1(_03375_),
    .B2(net217),
    .A2(_03373_),
    .A1(net168));
 sg13g2_o21ai_1 _23399_ (.B1(_03376_),
    .Y(_03377_),
    .A1(net168),
    .A2(_03372_));
 sg13g2_nand4_1 _23400_ (.B(net164),
    .C(net243),
    .A(_02710_),
    .Y(_03378_),
    .D(_03043_));
 sg13g2_nand2_1 _23401_ (.Y(_03379_),
    .A(_03292_),
    .B(_03225_));
 sg13g2_a21oi_1 _23402_ (.A1(_03378_),
    .A2(_03379_),
    .Y(_03380_),
    .B1(net168));
 sg13g2_nand4_1 _23403_ (.B(net164),
    .C(_03180_),
    .A(net168),
    .Y(_03381_),
    .D(_03145_));
 sg13g2_nor2b_1 _23404_ (.A(_03380_),
    .B_N(_03381_),
    .Y(_03382_));
 sg13g2_o21ai_1 _23405_ (.B1(_03382_),
    .Y(_03383_),
    .A1(_03370_),
    .A2(_03377_));
 sg13g2_buf_1 _23406_ (.A(_03383_),
    .X(_03384_));
 sg13g2_xor2_1 _23407_ (.B(_03170_),
    .A(_03161_),
    .X(_03385_));
 sg13g2_xor2_1 _23408_ (.B(_03385_),
    .A(_03384_),
    .X(_03386_));
 sg13g2_xnor2_1 _23409_ (.Y(_03387_),
    .A(_03365_),
    .B(_03386_));
 sg13g2_xnor2_1 _23410_ (.Y(_03388_),
    .A(_03338_),
    .B(_03387_));
 sg13g2_nand2_1 _23411_ (.Y(_03389_),
    .A(net220),
    .B(_03234_));
 sg13g2_a21oi_1 _23412_ (.A1(net247),
    .A2(_03235_),
    .Y(_03390_),
    .B1(_03232_));
 sg13g2_a21o_1 _23413_ (.A2(net200),
    .A1(_03156_),
    .B1(_03241_),
    .X(_03391_));
 sg13g2_a221oi_1 _23414_ (.B2(_03237_),
    .C1(_03391_),
    .B1(_03240_),
    .A1(_03389_),
    .Y(_03392_),
    .A2(_03390_));
 sg13g2_o21ai_1 _23415_ (.B1(_03244_),
    .Y(_03393_),
    .A1(_03229_),
    .A2(_03392_));
 sg13g2_buf_1 _23416_ (.A(_03393_),
    .X(_03394_));
 sg13g2_nand3_1 _23417_ (.B(_03231_),
    .C(_03233_),
    .A(net220),
    .Y(_03395_));
 sg13g2_nand2_1 _23418_ (.Y(_03396_),
    .A(net143),
    .B(_03395_));
 sg13g2_buf_1 _23419_ (.A(_03396_),
    .X(_03397_));
 sg13g2_nand3_1 _23420_ (.B(net191),
    .C(net246),
    .A(net198),
    .Y(_03398_));
 sg13g2_o21ai_1 _23421_ (.B1(net274),
    .Y(_03399_),
    .A1(net227),
    .A2(net246));
 sg13g2_a21oi_1 _23422_ (.A1(_03398_),
    .A2(_03399_),
    .Y(_03400_),
    .B1(net243));
 sg13g2_mux2_1 _23423_ (.A0(_02782_),
    .A1(_03303_),
    .S(net191),
    .X(_03401_));
 sg13g2_nor2b_1 _23424_ (.A(_03401_),
    .B_N(_03145_),
    .Y(_03402_));
 sg13g2_a21oi_1 _23425_ (.A1(_02845_),
    .A2(_03294_),
    .Y(_03403_),
    .B1(_03303_));
 sg13g2_a221oi_1 _23426_ (.B2(net272),
    .C1(net245),
    .B1(net273),
    .A1(_02707_),
    .Y(_03404_),
    .A2(_02708_));
 sg13g2_o21ai_1 _23427_ (.B1(net269),
    .Y(_03405_),
    .A1(_03295_),
    .A2(_03404_));
 sg13g2_o21ai_1 _23428_ (.B1(_03405_),
    .Y(_03406_),
    .A1(net227),
    .A2(_03403_));
 sg13g2_or3_1 _23429_ (.A(_03400_),
    .B(_03402_),
    .C(_03406_),
    .X(_03407_));
 sg13g2_xnor2_1 _23430_ (.Y(_03408_),
    .A(_03370_),
    .B(_03407_));
 sg13g2_buf_1 _23431_ (.A(_03408_),
    .X(_03409_));
 sg13g2_xor2_1 _23432_ (.B(_03352_),
    .A(_03340_),
    .X(_03410_));
 sg13g2_buf_2 _23433_ (.A(_03410_),
    .X(_03411_));
 sg13g2_a21oi_1 _23434_ (.A1(net202),
    .A2(net194),
    .Y(_03412_),
    .B1(_02720_));
 sg13g2_nor3_1 _23435_ (.A(net201),
    .B(_03039_),
    .C(_02871_),
    .Y(_03413_));
 sg13g2_o21ai_1 _23436_ (.B1(net247),
    .Y(_03414_),
    .A1(_03412_),
    .A2(_03413_));
 sg13g2_nand3_1 _23437_ (.B(net196),
    .C(net189),
    .A(net191),
    .Y(_03415_));
 sg13g2_a21oi_1 _23438_ (.A1(net229),
    .A2(_02615_),
    .Y(_03416_),
    .B1(_02684_));
 sg13g2_nand2_1 _23439_ (.Y(_03417_),
    .A(_03415_),
    .B(_03416_));
 sg13g2_nor2_1 _23440_ (.A(_02454_),
    .B(_03014_),
    .Y(_03418_));
 sg13g2_xnor2_1 _23441_ (.Y(_03419_),
    .A(_02720_),
    .B(net194));
 sg13g2_nand2_1 _23442_ (.Y(_03420_),
    .A(_03418_),
    .B(_03419_));
 sg13g2_and3_1 _23443_ (.X(_03421_),
    .A(_03252_),
    .B(_03255_),
    .C(_03256_));
 sg13g2_buf_8 _23444_ (.A(_03421_),
    .X(_03422_));
 sg13g2_a21oi_1 _23445_ (.A1(_03418_),
    .A2(_03419_),
    .Y(_03423_),
    .B1(net242));
 sg13g2_a221oi_1 _23446_ (.B2(_03422_),
    .C1(_03423_),
    .B1(_03420_),
    .A1(_03414_),
    .Y(_03424_),
    .A2(_03417_));
 sg13g2_buf_8 _23447_ (.A(_03424_),
    .X(_03425_));
 sg13g2_or2_1 _23448_ (.X(_03426_),
    .B(_03425_),
    .A(_03411_));
 sg13g2_buf_1 _23449_ (.A(_03426_),
    .X(_03427_));
 sg13g2_and4_1 _23450_ (.A(net88),
    .B(net105),
    .C(net94),
    .D(_03427_),
    .X(_03428_));
 sg13g2_nor3_1 _23451_ (.A(net88),
    .B(net105),
    .C(_03427_),
    .Y(_03429_));
 sg13g2_nor3_1 _23452_ (.A(net88),
    .B(net94),
    .C(_03427_),
    .Y(_03430_));
 sg13g2_and2_1 _23453_ (.A(_03411_),
    .B(_03425_),
    .X(_03431_));
 sg13g2_buf_1 _23454_ (.A(_03431_),
    .X(_03432_));
 sg13g2_nor4_1 _23455_ (.A(net88),
    .B(net105),
    .C(net94),
    .D(_03432_),
    .Y(_03433_));
 sg13g2_nor4_1 _23456_ (.A(_03428_),
    .B(_03429_),
    .C(_03430_),
    .D(_03433_),
    .Y(_03434_));
 sg13g2_and2_1 _23457_ (.A(_03394_),
    .B(net94),
    .X(_03435_));
 sg13g2_buf_1 _23458_ (.A(_03435_),
    .X(_03436_));
 sg13g2_nand2_1 _23459_ (.Y(_03437_),
    .A(_03436_),
    .B(_03432_));
 sg13g2_nand3_1 _23460_ (.B(_03409_),
    .C(_03432_),
    .A(net105),
    .Y(_03438_));
 sg13g2_or3_1 _23461_ (.A(net105),
    .B(_03409_),
    .C(_03427_),
    .X(_03439_));
 sg13g2_nand4_1 _23462_ (.B(_03437_),
    .C(_03438_),
    .A(_03434_),
    .Y(_03440_),
    .D(_03439_));
 sg13g2_buf_2 _23463_ (.A(_03440_),
    .X(_03441_));
 sg13g2_nor4_2 _23464_ (.A(_03327_),
    .B(_03331_),
    .C(_03388_),
    .Y(_03442_),
    .D(_03441_));
 sg13g2_xor2_1 _23465_ (.B(_03329_),
    .A(_03328_),
    .X(_03443_));
 sg13g2_and4_1 _23466_ (.A(_03326_),
    .B(_03443_),
    .C(_03388_),
    .D(_03441_),
    .X(_03444_));
 sg13g2_xnor2_1 _23467_ (.Y(_03445_),
    .A(_03411_),
    .B(_03425_));
 sg13g2_xnor2_1 _23468_ (.Y(_03446_),
    .A(net105),
    .B(_03445_));
 sg13g2_xor2_1 _23469_ (.B(net94),
    .A(net88),
    .X(_03447_));
 sg13g2_xnor2_1 _23470_ (.Y(_03448_),
    .A(_03446_),
    .B(_03447_));
 sg13g2_buf_1 _23471_ (.A(_03448_),
    .X(_03449_));
 sg13g2_nor4_1 _23472_ (.A(_03331_),
    .B(_03449_),
    .C(_03388_),
    .D(_03441_),
    .Y(_03450_));
 sg13g2_nor2_1 _23473_ (.A(_03331_),
    .B(_03449_),
    .Y(_03451_));
 sg13g2_and3_1 _23474_ (.X(_03452_),
    .A(_03451_),
    .B(_03388_),
    .C(_03441_));
 sg13g2_or4_1 _23475_ (.A(_03442_),
    .B(_03444_),
    .C(_03450_),
    .D(_03452_),
    .X(_03453_));
 sg13g2_buf_1 _23476_ (.A(_03453_),
    .X(_03454_));
 sg13g2_xnor2_1 _23477_ (.Y(_03455_),
    .A(_03388_),
    .B(_03441_));
 sg13g2_buf_8 _23478_ (.A(_03455_),
    .X(_03456_));
 sg13g2_xor2_1 _23479_ (.B(_03269_),
    .A(_03259_),
    .X(_03457_));
 sg13g2_buf_1 _23480_ (.A(_03280_),
    .X(_03458_));
 sg13g2_nor3_1 _23481_ (.A(_03049_),
    .B(net104),
    .C(_03422_),
    .Y(_03459_));
 sg13g2_xnor2_1 _23482_ (.Y(_03460_),
    .A(net201),
    .B(net228));
 sg13g2_nor4_1 _23483_ (.A(net203),
    .B(_02686_),
    .C(_03068_),
    .D(_03460_),
    .Y(_03461_));
 sg13g2_o21ai_1 _23484_ (.B1(net145),
    .Y(_03462_),
    .A1(_03459_),
    .A2(_03461_));
 sg13g2_or3_1 _23485_ (.A(_03457_),
    .B(_03462_),
    .C(_03321_),
    .X(_03463_));
 sg13g2_buf_1 _23486_ (.A(_03463_),
    .X(_03464_));
 sg13g2_o21ai_1 _23487_ (.B1(_03320_),
    .Y(_03465_),
    .A1(_03248_),
    .A2(_03249_));
 sg13g2_or2_1 _23488_ (.X(_03466_),
    .B(_03465_),
    .A(_03323_));
 sg13g2_buf_1 _23489_ (.A(_03466_),
    .X(_03467_));
 sg13g2_and2_1 _23490_ (.A(_03464_),
    .B(_03467_),
    .X(_03468_));
 sg13g2_o21ai_1 _23491_ (.B1(_03468_),
    .Y(_03469_),
    .A1(_03327_),
    .A2(_03449_));
 sg13g2_buf_1 _23492_ (.A(_03469_),
    .X(_03470_));
 sg13g2_and2_1 _23493_ (.A(_03456_),
    .B(_03470_),
    .X(_03471_));
 sg13g2_nor2_1 _23494_ (.A(_03454_),
    .B(_03471_),
    .Y(_03472_));
 sg13g2_nor2_1 _23495_ (.A(_03356_),
    .B(_03358_),
    .Y(_03473_));
 sg13g2_nand2_1 _23496_ (.Y(_03474_),
    .A(_03356_),
    .B(_03358_));
 sg13g2_inv_1 _23497_ (.Y(_03475_),
    .A(_03363_));
 sg13g2_nor2_1 _23498_ (.A(_03474_),
    .B(_03475_),
    .Y(_03476_));
 sg13g2_nand2_1 _23499_ (.Y(_03477_),
    .A(_03384_),
    .B(_03385_));
 sg13g2_mux2_1 _23500_ (.A0(_03473_),
    .A1(_03476_),
    .S(_03477_),
    .X(_03478_));
 sg13g2_or2_1 _23501_ (.X(_03479_),
    .B(_03363_),
    .A(_03356_));
 sg13g2_or2_1 _23502_ (.X(_03480_),
    .B(_03363_),
    .A(_03358_));
 sg13g2_a21oi_1 _23503_ (.A1(_03479_),
    .A2(_03480_),
    .Y(_03481_),
    .B1(_03477_));
 sg13g2_or2_1 _23504_ (.X(_03482_),
    .B(_03385_),
    .A(_03384_));
 sg13g2_buf_1 _23505_ (.A(_03482_),
    .X(_03483_));
 sg13g2_nor3_1 _23506_ (.A(_03356_),
    .B(_03358_),
    .C(_03363_),
    .Y(_03484_));
 sg13g2_nor3_1 _23507_ (.A(_03474_),
    .B(_03384_),
    .C(_03385_),
    .Y(_03485_));
 sg13g2_a21o_1 _23508_ (.A2(_03484_),
    .A1(_03483_),
    .B1(_03485_),
    .X(_03486_));
 sg13g2_nand2_1 _23509_ (.Y(_03487_),
    .A(_03356_),
    .B(_03363_));
 sg13g2_nand2_1 _23510_ (.Y(_03488_),
    .A(_03358_),
    .B(_03363_));
 sg13g2_a21oi_1 _23511_ (.A1(_03487_),
    .A2(_03488_),
    .Y(_03489_),
    .B1(_03483_));
 sg13g2_nor4_1 _23512_ (.A(_03478_),
    .B(_03481_),
    .C(_03486_),
    .D(_03489_),
    .Y(_03490_));
 sg13g2_a21oi_1 _23513_ (.A1(net202),
    .A2(_02917_),
    .Y(_03491_),
    .B1(net120));
 sg13g2_nor3_1 _23514_ (.A(net182),
    .B(_03283_),
    .C(_03491_),
    .Y(_03492_));
 sg13g2_nor2_1 _23515_ (.A(_03127_),
    .B(net120),
    .Y(_03493_));
 sg13g2_nand2_1 _23516_ (.Y(_03494_),
    .A(net193),
    .B(_03023_));
 sg13g2_a221oi_1 _23517_ (.B2(_03494_),
    .C1(net218),
    .B1(_03289_),
    .A1(_03261_),
    .Y(_03495_),
    .A2(_03493_));
 sg13g2_nand2_1 _23518_ (.Y(_03496_),
    .A(net181),
    .B(net120));
 sg13g2_o21ai_1 _23519_ (.B1(_03496_),
    .Y(_03497_),
    .A1(_03492_),
    .A2(_03495_));
 sg13g2_xor2_1 _23520_ (.B(_03191_),
    .A(_03179_),
    .X(_03498_));
 sg13g2_xnor2_1 _23521_ (.Y(_03499_),
    .A(_03192_),
    .B(_03498_));
 sg13g2_xnor2_1 _23522_ (.Y(_03500_),
    .A(_03497_),
    .B(_03499_));
 sg13g2_xnor2_1 _23523_ (.Y(_03501_),
    .A(_03490_),
    .B(_03500_));
 sg13g2_buf_1 _23524_ (.A(_03501_),
    .X(_03502_));
 sg13g2_or2_1 _23525_ (.X(_03503_),
    .B(net94),
    .A(net88));
 sg13g2_o21ai_1 _23526_ (.B1(_03397_),
    .Y(_03504_),
    .A1(_03411_),
    .A2(_03425_));
 sg13g2_and2_1 _23527_ (.A(net143),
    .B(_03395_),
    .X(_03505_));
 sg13g2_buf_1 _23528_ (.A(_03505_),
    .X(_03506_));
 sg13g2_nand2_1 _23529_ (.Y(_03507_),
    .A(_03506_),
    .B(_03445_));
 sg13g2_nand4_1 _23530_ (.B(_03338_),
    .C(_03504_),
    .A(_03503_),
    .Y(_03508_),
    .D(_03507_));
 sg13g2_nand2_1 _23531_ (.Y(_03509_),
    .A(_03411_),
    .B(_03425_));
 sg13g2_a21oi_1 _23532_ (.A1(_03509_),
    .A2(_03504_),
    .Y(_03510_),
    .B1(_03338_));
 sg13g2_nor4_2 _23533_ (.A(_03051_),
    .B(_03333_),
    .C(_03335_),
    .Y(_03511_),
    .D(_03336_));
 sg13g2_nor3_1 _23534_ (.A(_03397_),
    .B(_03411_),
    .C(_03511_),
    .Y(_03512_));
 sg13g2_o21ai_1 _23535_ (.B1(_03436_),
    .Y(_03513_),
    .A1(_03510_),
    .A2(_03512_));
 sg13g2_nand3_1 _23536_ (.B(_03508_),
    .C(_03513_),
    .A(_03387_),
    .Y(_03514_));
 sg13g2_buf_1 _23537_ (.A(_03514_),
    .X(_03515_));
 sg13g2_nor2_1 _23538_ (.A(net88),
    .B(net94),
    .Y(_03516_));
 sg13g2_nand2_1 _23539_ (.Y(_03517_),
    .A(net105),
    .B(_03425_));
 sg13g2_a21oi_1 _23540_ (.A1(_03338_),
    .A2(_03517_),
    .Y(_03518_),
    .B1(_03510_));
 sg13g2_and3_1 _23541_ (.X(_03519_),
    .A(_03411_),
    .B(_03425_),
    .C(_03338_));
 sg13g2_nor3_1 _23542_ (.A(_03411_),
    .B(_03425_),
    .C(_03338_),
    .Y(_03520_));
 sg13g2_o21ai_1 _23543_ (.B1(_03506_),
    .Y(_03521_),
    .A1(_03519_),
    .A2(_03520_));
 sg13g2_or3_1 _23544_ (.A(_03506_),
    .B(_03445_),
    .C(_03511_),
    .X(_03522_));
 sg13g2_a21oi_1 _23545_ (.A1(_03521_),
    .A2(_03522_),
    .Y(_03523_),
    .B1(_03436_));
 sg13g2_a21oi_2 _23546_ (.B1(_03523_),
    .Y(_03524_),
    .A2(_03518_),
    .A1(_03516_));
 sg13g2_nand2_2 _23547_ (.Y(_03525_),
    .A(_03515_),
    .B(_03524_));
 sg13g2_buf_1 _23548_ (.A(net217),
    .X(_03526_));
 sg13g2_nand2_1 _23549_ (.Y(_03527_),
    .A(net164),
    .B(_03156_));
 sg13g2_nand2_2 _23550_ (.Y(_03528_),
    .A(net221),
    .B(net195));
 sg13g2_o21ai_1 _23551_ (.B1(_03528_),
    .Y(_03529_),
    .A1(_03460_),
    .A2(_03527_));
 sg13g2_xnor2_1 _23552_ (.Y(_03530_),
    .A(net104),
    .B(net119));
 sg13g2_nand2_1 _23553_ (.Y(_03531_),
    .A(_03284_),
    .B(_03315_));
 sg13g2_nor2_1 _23554_ (.A(_03528_),
    .B(_03531_),
    .Y(_03532_));
 sg13g2_a21oi_1 _23555_ (.A1(_03529_),
    .A2(_03530_),
    .Y(_03533_),
    .B1(_03532_));
 sg13g2_nor3_1 _23556_ (.A(_03526_),
    .B(_03083_),
    .C(_03533_),
    .Y(_03534_));
 sg13g2_buf_2 _23557_ (.A(_03534_),
    .X(_03535_));
 sg13g2_nand3_1 _23558_ (.B(_03464_),
    .C(_03467_),
    .A(_03326_),
    .Y(_03536_));
 sg13g2_xnor2_1 _23559_ (.Y(_03537_),
    .A(_03443_),
    .B(_03449_));
 sg13g2_xnor2_1 _23560_ (.Y(_03538_),
    .A(_03536_),
    .B(_03537_));
 sg13g2_or2_1 _23561_ (.X(_03539_),
    .B(_03538_),
    .A(_03535_));
 sg13g2_buf_1 _23562_ (.A(_03539_),
    .X(_03540_));
 sg13g2_nand2_1 _23563_ (.Y(_03541_),
    .A(_03464_),
    .B(_03467_));
 sg13g2_a21o_1 _23564_ (.A2(_03331_),
    .A1(_03323_),
    .B1(_03465_),
    .X(_03542_));
 sg13g2_a21oi_1 _23565_ (.A1(_03462_),
    .A2(_03287_),
    .Y(_03543_),
    .B1(_03271_));
 sg13g2_nor3_1 _23566_ (.A(net145),
    .B(_03459_),
    .C(_03461_),
    .Y(_03544_));
 sg13g2_nor3_1 _23567_ (.A(_03457_),
    .B(_03322_),
    .C(_03544_),
    .Y(_03545_));
 sg13g2_or4_1 _23568_ (.A(_03543_),
    .B(_03545_),
    .C(_03321_),
    .D(_03331_),
    .X(_03546_));
 sg13g2_nand2b_1 _23569_ (.Y(_03547_),
    .B(_03443_),
    .A_N(_03323_));
 sg13g2_and4_1 _23570_ (.A(_03464_),
    .B(_03542_),
    .C(_03546_),
    .D(_03547_),
    .X(_03548_));
 sg13g2_nor2_1 _23571_ (.A(_03326_),
    .B(_03443_),
    .Y(_03549_));
 sg13g2_a221oi_1 _23572_ (.B2(_03449_),
    .C1(_03549_),
    .B1(_03548_),
    .A1(_03541_),
    .Y(_03550_),
    .A2(_03451_));
 sg13g2_xor2_1 _23573_ (.B(_03550_),
    .A(_03456_),
    .X(_03551_));
 sg13g2_buf_2 _23574_ (.A(_03551_),
    .X(_03552_));
 sg13g2_o21ai_1 _23575_ (.B1(_03457_),
    .Y(_03553_),
    .A1(_03322_),
    .A2(_03544_));
 sg13g2_nand3_1 _23576_ (.B(_03462_),
    .C(_03287_),
    .A(_03271_),
    .Y(_03554_));
 sg13g2_nand3_1 _23577_ (.B(_03244_),
    .C(_03246_),
    .A(_03229_),
    .Y(_03555_));
 sg13g2_a21o_1 _23578_ (.A2(_03246_),
    .A1(_03244_),
    .B1(_03229_),
    .X(_03556_));
 sg13g2_nand3_1 _23579_ (.B(_03556_),
    .C(_03320_),
    .A(_03555_),
    .Y(_03557_));
 sg13g2_a21o_1 _23580_ (.A2(_03556_),
    .A1(_03555_),
    .B1(_03320_),
    .X(_03558_));
 sg13g2_a22oi_1 _23581_ (.Y(_03559_),
    .B1(_03557_),
    .B2(_03558_),
    .A2(_03554_),
    .A1(_03553_));
 sg13g2_and4_1 _23582_ (.A(_03553_),
    .B(_03554_),
    .C(_03557_),
    .D(_03558_),
    .X(_03560_));
 sg13g2_buf_1 _23583_ (.A(_03560_),
    .X(_03561_));
 sg13g2_nor2_1 _23584_ (.A(_03460_),
    .B(_03527_),
    .Y(_03562_));
 sg13g2_o21ai_1 _23585_ (.B1(_03562_),
    .Y(_03563_),
    .A1(net104),
    .A2(_03422_));
 sg13g2_nor3_1 _23586_ (.A(_03562_),
    .B(net104),
    .C(_03422_),
    .Y(_03564_));
 sg13g2_a21o_1 _23587_ (.A2(_03563_),
    .A1(_03528_),
    .B1(_03564_),
    .X(_03565_));
 sg13g2_nand2_1 _23588_ (.Y(_03566_),
    .A(net106),
    .B(_03422_));
 sg13g2_nand3_1 _23589_ (.B(net119),
    .C(_03529_),
    .A(net120),
    .Y(_03567_));
 sg13g2_o21ai_1 _23590_ (.B1(_03567_),
    .Y(_03568_),
    .A1(_03532_),
    .A2(_03566_));
 sg13g2_a22oi_1 _23591_ (.Y(_03569_),
    .B1(_03568_),
    .B2(_03458_),
    .A2(_03565_),
    .A1(net106));
 sg13g2_o21ai_1 _23592_ (.B1(_03531_),
    .Y(_03570_),
    .A1(net104),
    .A2(net119));
 sg13g2_nor3_1 _23593_ (.A(_03531_),
    .B(net104),
    .C(net119),
    .Y(_03571_));
 sg13g2_a21o_1 _23594_ (.A2(_03570_),
    .A1(_02930_),
    .B1(_03571_),
    .X(_03572_));
 sg13g2_buf_1 _23595_ (.A(net214),
    .X(_03573_));
 sg13g2_nor3_1 _23596_ (.A(net179),
    .B(_03528_),
    .C(_03458_),
    .Y(_03574_));
 sg13g2_a21oi_1 _23597_ (.A1(net120),
    .A2(_03572_),
    .Y(_03575_),
    .B1(_03574_));
 sg13g2_o21ai_1 _23598_ (.B1(_03575_),
    .Y(_03576_),
    .A1(_03526_),
    .A2(_03569_));
 sg13g2_buf_1 _23599_ (.A(_03576_),
    .X(_03577_));
 sg13g2_nor3_1 _23600_ (.A(_03559_),
    .B(_03561_),
    .C(_03577_),
    .Y(_03578_));
 sg13g2_nor2b_1 _23601_ (.A(_03318_),
    .B_N(_03317_),
    .Y(_03579_));
 sg13g2_xnor2_1 _23602_ (.Y(_03580_),
    .A(_03309_),
    .B(_03579_));
 sg13g2_nand3_1 _23603_ (.B(_02746_),
    .C(_03292_),
    .A(net147),
    .Y(_03581_));
 sg13g2_nand3_1 _23604_ (.B(_02746_),
    .C(_03180_),
    .A(net203),
    .Y(_03582_));
 sg13g2_nand3_1 _23605_ (.B(_03089_),
    .C(_03261_),
    .A(_02829_),
    .Y(_03583_));
 sg13g2_nor3_1 _23606_ (.A(net287),
    .B(net286),
    .C(net186),
    .Y(_03584_));
 sg13g2_nor4_1 _23607_ (.A(_02716_),
    .B(_02718_),
    .C(net199),
    .D(net214),
    .Y(_03585_));
 sg13g2_nor4_1 _23608_ (.A(net199),
    .B(net214),
    .C(net274),
    .D(net186),
    .Y(_03586_));
 sg13g2_a221oi_1 _23609_ (.B2(_02829_),
    .C1(_03586_),
    .B1(_03585_),
    .A1(_03584_),
    .Y(_03587_),
    .A2(_03184_));
 sg13g2_nand4_1 _23610_ (.B(_03582_),
    .C(_03583_),
    .A(_03581_),
    .Y(_03588_),
    .D(_03587_));
 sg13g2_a21oi_1 _23611_ (.A1(net273),
    .A2(net272),
    .Y(_03589_),
    .B1(net242));
 sg13g2_nand3_1 _23612_ (.B(net163),
    .C(_03589_),
    .A(net170),
    .Y(_03590_));
 sg13g2_nand4_1 _23613_ (.B(net167),
    .C(net214),
    .A(net164),
    .Y(_03591_),
    .D(net163));
 sg13g2_nand3_1 _23614_ (.B(net167),
    .C(_03051_),
    .A(net164),
    .Y(_03592_));
 sg13g2_nand3_1 _23615_ (.B(net244),
    .C(_03292_),
    .A(net164),
    .Y(_03593_));
 sg13g2_nand4_1 _23616_ (.B(_03591_),
    .C(_03592_),
    .A(_03590_),
    .Y(_03594_),
    .D(_03593_));
 sg13g2_o21ai_1 _23617_ (.B1(_03043_),
    .Y(_03595_),
    .A1(_02686_),
    .A2(net163));
 sg13g2_nand4_1 _23618_ (.B(net214),
    .C(_03129_),
    .A(net203),
    .Y(_03596_),
    .D(net163));
 sg13g2_a21oi_1 _23619_ (.A1(_03595_),
    .A2(_03596_),
    .Y(_03597_),
    .B1(_02722_));
 sg13g2_nor3_2 _23620_ (.A(_03588_),
    .B(_03594_),
    .C(_03597_),
    .Y(_03598_));
 sg13g2_nor2_1 _23621_ (.A(_02871_),
    .B(_03151_),
    .Y(_03599_));
 sg13g2_o21ai_1 _23622_ (.B1(net186),
    .Y(_03600_),
    .A1(_03079_),
    .A2(net219));
 sg13g2_nor3_1 _23623_ (.A(_03079_),
    .B(net186),
    .C(net184),
    .Y(_03601_));
 sg13g2_a21o_1 _23624_ (.A2(_03600_),
    .A1(net170),
    .B1(_03601_),
    .X(_03602_));
 sg13g2_nor4_1 _23625_ (.A(net167),
    .B(net169),
    .C(net217),
    .D(_03131_),
    .Y(_03603_));
 sg13g2_a221oi_1 _23626_ (.B2(_03156_),
    .C1(_03603_),
    .B1(_03602_),
    .A1(net215),
    .Y(_03604_),
    .A2(_03599_));
 sg13g2_buf_1 _23627_ (.A(_03604_),
    .X(_03605_));
 sg13g2_nand2_1 _23628_ (.Y(_03606_),
    .A(_03598_),
    .B(_03605_));
 sg13g2_a221oi_1 _23629_ (.B2(_02770_),
    .C1(net247),
    .B1(net221),
    .A1(net215),
    .Y(_03607_),
    .A2(net163));
 sg13g2_a221oi_1 _23630_ (.B2(_03080_),
    .C1(_02913_),
    .B1(_02730_),
    .A1(net190),
    .Y(_03608_),
    .A2(net184));
 sg13g2_nand2_1 _23631_ (.Y(_03609_),
    .A(net215),
    .B(_03106_));
 sg13g2_o21ai_1 _23632_ (.B1(_03609_),
    .Y(_03610_),
    .A1(_03607_),
    .A2(_03608_));
 sg13g2_inv_1 _23633_ (.Y(_03611_),
    .A(_03610_));
 sg13g2_o21ai_1 _23634_ (.B1(_03611_),
    .Y(_03612_),
    .A1(_03598_),
    .A2(_03605_));
 sg13g2_nand2_1 _23635_ (.Y(_03613_),
    .A(net214),
    .B(net119));
 sg13g2_a21oi_1 _23636_ (.A1(_03284_),
    .A2(_03315_),
    .Y(_03614_),
    .B1(_03528_));
 sg13g2_nor3_1 _23637_ (.A(_02930_),
    .B(_03460_),
    .C(_03527_),
    .Y(_03615_));
 sg13g2_or3_1 _23638_ (.A(_03614_),
    .B(_03615_),
    .C(net104),
    .X(_03616_));
 sg13g2_o21ai_1 _23639_ (.B1(net104),
    .Y(_03617_),
    .A1(_03614_),
    .A2(_03615_));
 sg13g2_nand3_1 _23640_ (.B(_03616_),
    .C(_03617_),
    .A(_03613_),
    .Y(_03618_));
 sg13g2_buf_1 _23641_ (.A(_03618_),
    .X(_03619_));
 sg13g2_a21o_1 _23642_ (.A2(_03617_),
    .A1(_03616_),
    .B1(_03613_),
    .X(_03620_));
 sg13g2_buf_1 _23643_ (.A(_03620_),
    .X(_03621_));
 sg13g2_nand4_1 _23644_ (.B(_03612_),
    .C(_03619_),
    .A(_03606_),
    .Y(_03622_),
    .D(_03621_));
 sg13g2_a22oi_1 _23645_ (.Y(_03623_),
    .B1(_03619_),
    .B2(_03621_),
    .A2(_03612_),
    .A1(_03606_));
 sg13g2_a21o_1 _23646_ (.A2(_03622_),
    .A1(_03580_),
    .B1(_03623_),
    .X(_03624_));
 sg13g2_buf_2 _23647_ (.A(_03624_),
    .X(_03625_));
 sg13g2_o21ai_1 _23648_ (.B1(_03577_),
    .Y(_03626_),
    .A1(_03559_),
    .A2(_03561_));
 sg13g2_o21ai_1 _23649_ (.B1(_03626_),
    .Y(_03627_),
    .A1(_03578_),
    .A2(_03625_));
 sg13g2_buf_1 _23650_ (.A(_03627_),
    .X(_03628_));
 sg13g2_a21o_1 _23651_ (.A2(_03538_),
    .A1(_03535_),
    .B1(_03628_),
    .X(_03629_));
 sg13g2_buf_1 _23652_ (.A(_03629_),
    .X(_03630_));
 sg13g2_nand3_1 _23653_ (.B(_03552_),
    .C(_03630_),
    .A(_03540_),
    .Y(_03631_));
 sg13g2_nand4_1 _23654_ (.B(net79),
    .C(_03525_),
    .A(_03472_),
    .Y(_03632_),
    .D(_03631_));
 sg13g2_and2_1 _23655_ (.A(_03509_),
    .B(_03504_),
    .X(_03633_));
 sg13g2_or2_1 _23656_ (.X(_03634_),
    .B(_03633_),
    .A(_03511_));
 sg13g2_buf_1 _23657_ (.A(_03634_),
    .X(_03635_));
 sg13g2_xnor2_1 _23658_ (.Y(_03636_),
    .A(_03198_),
    .B(_03199_));
 sg13g2_xor2_1 _23659_ (.B(_03636_),
    .A(_03195_),
    .X(_03637_));
 sg13g2_buf_2 _23660_ (.A(_03637_),
    .X(_03638_));
 sg13g2_a21oi_1 _23661_ (.A1(_03474_),
    .A2(_03475_),
    .Y(_03639_),
    .B1(_03473_));
 sg13g2_xor2_1 _23662_ (.B(_03497_),
    .A(_03639_),
    .X(_03640_));
 sg13g2_and2_1 _23663_ (.A(_03384_),
    .B(_03385_),
    .X(_03641_));
 sg13g2_o21ai_1 _23664_ (.B1(_03483_),
    .Y(_03642_),
    .A1(_03365_),
    .A2(_03641_));
 sg13g2_nor2_1 _23665_ (.A(_03640_),
    .B(_03642_),
    .Y(_03643_));
 sg13g2_a21oi_1 _23666_ (.A1(_03640_),
    .A2(_03642_),
    .Y(_03644_),
    .B1(_03499_));
 sg13g2_buf_1 _23667_ (.A(net242),
    .X(_03645_));
 sg13g2_nor2_1 _23668_ (.A(_03645_),
    .B(_03023_),
    .Y(_03646_));
 sg13g2_a22oi_1 _23669_ (.Y(_03647_),
    .B1(_03265_),
    .B2(_03646_),
    .A2(_03023_),
    .A1(net141));
 sg13g2_inv_1 _23670_ (.Y(_03648_),
    .A(_03647_));
 sg13g2_nand2_1 _23671_ (.Y(_03649_),
    .A(_03261_),
    .B(_03493_));
 sg13g2_nand2_1 _23672_ (.Y(_03650_),
    .A(_03010_),
    .B(_03023_));
 sg13g2_o21ai_1 _23673_ (.B1(_03650_),
    .Y(_03651_),
    .A1(net141),
    .A2(_03023_));
 sg13g2_a21oi_1 _23674_ (.A1(_02801_),
    .A2(_03175_),
    .Y(_03652_),
    .B1(net141));
 sg13g2_nand2b_1 _23675_ (.Y(_03653_),
    .B(_03074_),
    .A_N(_03652_));
 sg13g2_o21ai_1 _23676_ (.B1(_03653_),
    .Y(_03654_),
    .A1(net224),
    .A2(_03651_));
 sg13g2_a221oi_1 _23677_ (.B2(_03649_),
    .C1(_03654_),
    .B1(_03639_),
    .A1(net197),
    .Y(_03655_),
    .A2(_03648_));
 sg13g2_buf_1 _23678_ (.A(_03655_),
    .X(_03656_));
 sg13g2_inv_1 _23679_ (.Y(_03657_),
    .A(_03656_));
 sg13g2_o21ai_1 _23680_ (.B1(_03657_),
    .Y(_03658_),
    .A1(_03643_),
    .A2(_03644_));
 sg13g2_buf_1 _23681_ (.A(_03658_),
    .X(_03659_));
 sg13g2_or3_1 _23682_ (.A(_03657_),
    .B(_03643_),
    .C(_03644_),
    .X(_03660_));
 sg13g2_buf_2 _23683_ (.A(_03660_),
    .X(_03661_));
 sg13g2_and3_1 _23684_ (.X(_03662_),
    .A(_03638_),
    .B(_03659_),
    .C(_03661_));
 sg13g2_buf_2 _23685_ (.A(_03662_),
    .X(_03663_));
 sg13g2_a21oi_2 _23686_ (.B1(_03638_),
    .Y(_03664_),
    .A2(_03661_),
    .A1(_03659_));
 sg13g2_nor3_1 _23687_ (.A(_03635_),
    .B(_03663_),
    .C(_03664_),
    .Y(_03665_));
 sg13g2_inv_1 _23688_ (.Y(_03666_),
    .A(net79));
 sg13g2_nand3_1 _23689_ (.B(_03659_),
    .C(_03661_),
    .A(_03638_),
    .Y(_03667_));
 sg13g2_a21o_1 _23690_ (.A2(_03661_),
    .A1(_03659_),
    .B1(_03638_),
    .X(_03668_));
 sg13g2_nand4_1 _23691_ (.B(_03666_),
    .C(_03667_),
    .A(_03635_),
    .Y(_03669_),
    .D(_03668_));
 sg13g2_or4_1 _23692_ (.A(_03666_),
    .B(_03525_),
    .C(_03663_),
    .D(_03664_),
    .X(_03670_));
 sg13g2_a22oi_1 _23693_ (.Y(_03671_),
    .B1(_03669_),
    .B2(_03670_),
    .A2(_03631_),
    .A1(_03472_));
 sg13g2_a21oi_2 _23694_ (.B1(_03671_),
    .Y(_03672_),
    .A2(_03665_),
    .A1(_03632_));
 sg13g2_nor4_2 _23695_ (.A(_03442_),
    .B(_03444_),
    .C(_03450_),
    .Y(_03673_),
    .D(_03452_));
 sg13g2_nand2_1 _23696_ (.Y(_03674_),
    .A(_03456_),
    .B(_03470_));
 sg13g2_nand2_1 _23697_ (.Y(_03675_),
    .A(_03673_),
    .B(_03674_));
 sg13g2_buf_2 _23698_ (.A(_03675_),
    .X(_03676_));
 sg13g2_nor2_1 _23699_ (.A(_03663_),
    .B(_03664_),
    .Y(_03677_));
 sg13g2_buf_2 _23700_ (.A(_03677_),
    .X(_03678_));
 sg13g2_and3_1 _23701_ (.X(_03679_),
    .A(_03540_),
    .B(_03552_),
    .C(_03630_));
 sg13g2_buf_8 _23702_ (.A(_03679_),
    .X(_03680_));
 sg13g2_nand2_1 _23703_ (.Y(_03681_),
    .A(_03635_),
    .B(net79));
 sg13g2_nor4_2 _23704_ (.A(_03676_),
    .B(_03678_),
    .C(_03680_),
    .Y(_03682_),
    .D(_03681_));
 sg13g2_nand2_1 _23705_ (.Y(_03683_),
    .A(net79),
    .B(_03525_));
 sg13g2_nor4_2 _23706_ (.A(_03676_),
    .B(_03683_),
    .C(_03678_),
    .Y(_03684_),
    .D(_03680_));
 sg13g2_nor2_1 _23707_ (.A(_03511_),
    .B(_03633_),
    .Y(_03685_));
 sg13g2_a21oi_1 _23708_ (.A1(_03515_),
    .A2(_03524_),
    .Y(_03686_),
    .B1(_03685_));
 sg13g2_o21ai_1 _23709_ (.B1(_03686_),
    .Y(_03687_),
    .A1(_03663_),
    .A2(_03664_));
 sg13g2_nor3_1 _23710_ (.A(_03676_),
    .B(_03680_),
    .C(_03687_),
    .Y(_03688_));
 sg13g2_nor2_1 _23711_ (.A(_03685_),
    .B(_03683_),
    .Y(_03689_));
 sg13g2_nor3_1 _23712_ (.A(_03685_),
    .B(net79),
    .C(_03525_),
    .Y(_03690_));
 sg13g2_mux2_1 _23713_ (.A0(_03689_),
    .A1(_03690_),
    .S(_03678_),
    .X(_03691_));
 sg13g2_nor4_2 _23714_ (.A(_03682_),
    .B(_03684_),
    .C(_03688_),
    .Y(_03692_),
    .D(_03691_));
 sg13g2_xnor2_1 _23715_ (.Y(_03693_),
    .A(_03139_),
    .B(_03141_));
 sg13g2_xnor2_1 _23716_ (.Y(_03694_),
    .A(_03202_),
    .B(_03693_));
 sg13g2_or2_1 _23717_ (.X(_03695_),
    .B(_03644_),
    .A(_03643_));
 sg13g2_buf_1 _23718_ (.A(_03695_),
    .X(_03696_));
 sg13g2_nor2_1 _23719_ (.A(_03638_),
    .B(_03696_),
    .Y(_03697_));
 sg13g2_a21oi_1 _23720_ (.A1(_03638_),
    .A2(_03696_),
    .Y(_03698_),
    .B1(_03656_));
 sg13g2_nor2_2 _23721_ (.A(_03697_),
    .B(_03698_),
    .Y(_03699_));
 sg13g2_xnor2_1 _23722_ (.Y(_03700_),
    .A(_03694_),
    .B(_03699_));
 sg13g2_buf_1 _23723_ (.A(_03700_),
    .X(_03701_));
 sg13g2_nor2_1 _23724_ (.A(net242),
    .B(net142),
    .Y(_03702_));
 sg13g2_xnor2_1 _23725_ (.Y(_03703_),
    .A(_03134_),
    .B(_03702_));
 sg13g2_or2_1 _23726_ (.X(_03704_),
    .B(net163),
    .A(net244));
 sg13g2_o21ai_1 _23727_ (.B1(net242),
    .Y(_03705_),
    .A1(net163),
    .A2(net184));
 sg13g2_and3_1 _23728_ (.X(_03706_),
    .A(net215),
    .B(net242),
    .C(net142));
 sg13g2_a221oi_1 _23729_ (.B2(net169),
    .C1(_03706_),
    .B1(_03705_),
    .A1(net184),
    .Y(_03707_),
    .A2(_03704_));
 sg13g2_mux2_1 _23730_ (.A0(_03300_),
    .A1(_03237_),
    .S(_03707_),
    .X(_03708_));
 sg13g2_a21o_1 _23731_ (.A2(_03703_),
    .A1(net180),
    .B1(_03708_),
    .X(_03709_));
 sg13g2_nand2_1 _23732_ (.Y(_03710_),
    .A(net244),
    .B(net162));
 sg13g2_a22oi_1 _23733_ (.Y(_03711_),
    .B1(_03710_),
    .B2(net121),
    .A2(_03283_),
    .A1(net185));
 sg13g2_nand2_1 _23734_ (.Y(_03712_),
    .A(net121),
    .B(_03283_));
 sg13g2_o21ai_1 _23735_ (.B1(_03712_),
    .Y(_03713_),
    .A1(net180),
    .A2(_03711_));
 sg13g2_nor3_1 _23736_ (.A(net180),
    .B(net213),
    .C(net182),
    .Y(_03714_));
 sg13g2_o21ai_1 _23737_ (.B1(_02829_),
    .Y(_03715_),
    .A1(net141),
    .A2(_03714_));
 sg13g2_nand2_1 _23738_ (.Y(_03716_),
    .A(_03712_),
    .B(_03715_));
 sg13g2_a21oi_1 _23739_ (.A1(net217),
    .A2(_02829_),
    .Y(_03717_),
    .B1(net216));
 sg13g2_nor2_1 _23740_ (.A(net141),
    .B(_03124_),
    .Y(_03718_));
 sg13g2_nor2_1 _23741_ (.A(_03717_),
    .B(_03718_),
    .Y(_03719_));
 sg13g2_a221oi_1 _23742_ (.B2(net162),
    .C1(_03719_),
    .B1(_03716_),
    .A1(net218),
    .Y(_03720_),
    .A2(_03713_));
 sg13g2_xnor2_1 _23743_ (.Y(_03721_),
    .A(_03709_),
    .B(_03720_));
 sg13g2_nand2_1 _23744_ (.Y(_03722_),
    .A(net179),
    .B(net218));
 sg13g2_a22oi_1 _23745_ (.Y(_03723_),
    .B1(_02905_),
    .B2(net181),
    .A2(net194),
    .A1(_03645_));
 sg13g2_and4_1 _23746_ (.A(net213),
    .B(net182),
    .C(net142),
    .D(net162),
    .X(_03724_));
 sg13g2_a22oi_1 _23747_ (.Y(_03725_),
    .B1(_03724_),
    .B2(net179),
    .A2(_03283_),
    .A1(_02915_));
 sg13g2_o21ai_1 _23748_ (.B1(_03725_),
    .Y(_03726_),
    .A1(_03722_),
    .A2(_03723_));
 sg13g2_nor3_1 _23749_ (.A(net180),
    .B(net122),
    .C(_02692_),
    .Y(_03727_));
 sg13g2_xnor2_1 _23750_ (.Y(_03728_),
    .A(_03726_),
    .B(_03727_));
 sg13g2_nand2b_1 _23751_ (.Y(_03729_),
    .B(net121),
    .A_N(net162));
 sg13g2_a21oi_1 _23752_ (.A1(net179),
    .A2(_03729_),
    .Y(_03730_),
    .B1(net213));
 sg13g2_a21oi_1 _23753_ (.A1(net179),
    .A2(_03704_),
    .Y(_03731_),
    .B1(net185));
 sg13g2_or2_1 _23754_ (.X(_03732_),
    .B(_03731_),
    .A(_03730_));
 sg13g2_a221oi_1 _23755_ (.B2(net142),
    .C1(_03348_),
    .B1(net141),
    .A1(_02403_),
    .Y(_03733_),
    .A2(net291));
 sg13g2_o21ai_1 _23756_ (.B1(_03729_),
    .Y(_03734_),
    .A1(net182),
    .A2(_03733_));
 sg13g2_and2_1 _23757_ (.A(_02403_),
    .B(net291),
    .X(_03735_));
 sg13g2_or4_1 _23758_ (.A(net244),
    .B(net142),
    .C(_03735_),
    .D(_03348_),
    .X(_03736_));
 sg13g2_or3_1 _23759_ (.A(net141),
    .B(net213),
    .C(net162),
    .X(_03737_));
 sg13g2_a21oi_1 _23760_ (.A1(_03736_),
    .A2(_03737_),
    .Y(_03738_),
    .B1(net218));
 sg13g2_a21o_1 _23761_ (.A2(_03734_),
    .A1(net213),
    .B1(_03738_),
    .X(_03739_));
 sg13g2_a22oi_1 _23762_ (.Y(_03740_),
    .B1(_03739_),
    .B2(net179),
    .A2(_03732_),
    .A1(_03265_));
 sg13g2_buf_1 _23763_ (.A(_03740_),
    .X(_03741_));
 sg13g2_xnor2_1 _23764_ (.Y(_03742_),
    .A(_03728_),
    .B(_03741_));
 sg13g2_xnor2_1 _23765_ (.Y(_03743_),
    .A(_03721_),
    .B(_03742_));
 sg13g2_buf_1 _23766_ (.A(net213),
    .X(_03744_));
 sg13g2_nor3_1 _23767_ (.A(net180),
    .B(net178),
    .C(_03359_),
    .Y(_03745_));
 sg13g2_nand3_1 _23768_ (.B(_03743_),
    .C(_03745_),
    .A(net181),
    .Y(_03746_));
 sg13g2_nor4_1 _23769_ (.A(net179),
    .B(net216),
    .C(net182),
    .D(net162),
    .Y(_03747_));
 sg13g2_nand3_1 _23770_ (.B(_03743_),
    .C(_03747_),
    .A(net181),
    .Y(_03748_));
 sg13g2_and2_1 _23771_ (.A(_03746_),
    .B(_03748_),
    .X(_03749_));
 sg13g2_nor2_1 _23772_ (.A(net217),
    .B(net185),
    .Y(_03750_));
 sg13g2_nand3_1 _23773_ (.B(net218),
    .C(_03750_),
    .A(net178),
    .Y(_03751_));
 sg13g2_o21ai_1 _23774_ (.B1(_03609_),
    .Y(_03752_),
    .A1(_03231_),
    .A2(_03722_));
 sg13g2_a22oi_1 _23775_ (.Y(_03753_),
    .B1(_03752_),
    .B2(net178),
    .A2(_03134_),
    .A1(net218));
 sg13g2_buf_1 _23776_ (.A(_03753_),
    .X(_03754_));
 sg13g2_nand2_1 _23777_ (.Y(_03755_),
    .A(_02774_),
    .B(_02713_));
 sg13g2_buf_2 _23778_ (.A(_03755_),
    .X(_03756_));
 sg13g2_o21ai_1 _23779_ (.B1(_03296_),
    .Y(_03757_),
    .A1(_02722_),
    .A2(_02772_));
 sg13g2_nand2_1 _23780_ (.Y(_03758_),
    .A(net144),
    .B(_03589_));
 sg13g2_nand2_1 _23781_ (.Y(_03759_),
    .A(_03757_),
    .B(_03758_));
 sg13g2_a221oi_1 _23782_ (.B2(net145),
    .C1(_03759_),
    .B1(_03589_),
    .A1(_03756_),
    .Y(_03760_),
    .A2(_02618_));
 sg13g2_nand3_1 _23783_ (.B(net213),
    .C(_02694_),
    .A(net180),
    .Y(_03761_));
 sg13g2_o21ai_1 _23784_ (.B1(_03761_),
    .Y(_03762_),
    .A1(net180),
    .A2(_03760_));
 sg13g2_buf_1 _23785_ (.A(_03762_),
    .X(_03763_));
 sg13g2_xnor2_1 _23786_ (.Y(_03764_),
    .A(_03754_),
    .B(_03763_));
 sg13g2_xor2_1 _23787_ (.B(_03610_),
    .A(_03605_),
    .X(_03765_));
 sg13g2_xnor2_1 _23788_ (.Y(_03766_),
    .A(_03598_),
    .B(_03765_));
 sg13g2_buf_1 _23789_ (.A(_03766_),
    .X(_03767_));
 sg13g2_o21ai_1 _23790_ (.B1(_03289_),
    .Y(_03768_),
    .A1(net217),
    .A2(net162));
 sg13g2_o21ai_1 _23791_ (.B1(_03768_),
    .Y(_03769_),
    .A1(net181),
    .A2(_03750_));
 sg13g2_nand2_1 _23792_ (.Y(_03770_),
    .A(net162),
    .B(_03283_));
 sg13g2_o21ai_1 _23793_ (.B1(_03770_),
    .Y(_03771_),
    .A1(net182),
    .A2(_03769_));
 sg13g2_mux2_1 _23794_ (.A0(net194),
    .A1(_03231_),
    .S(net169),
    .X(_03772_));
 sg13g2_a22oi_1 _23795_ (.Y(_03773_),
    .B1(_03772_),
    .B2(net213),
    .A2(_03289_),
    .A1(_03091_));
 sg13g2_or2_1 _23796_ (.X(_03774_),
    .B(_03773_),
    .A(_03722_));
 sg13g2_nand3_1 _23797_ (.B(net182),
    .C(_03091_),
    .A(net141),
    .Y(_03775_));
 sg13g2_nand2b_1 _23798_ (.Y(_03776_),
    .B(_03775_),
    .A_N(_03719_));
 sg13g2_a221oi_1 _23799_ (.B2(_03709_),
    .C1(_03776_),
    .B1(_03774_),
    .A1(net121),
    .Y(_03777_),
    .A2(_03771_));
 sg13g2_buf_1 _23800_ (.A(_03777_),
    .X(_03778_));
 sg13g2_xnor2_1 _23801_ (.Y(_03779_),
    .A(_03767_),
    .B(_03778_));
 sg13g2_xnor2_1 _23802_ (.Y(_03780_),
    .A(_03764_),
    .B(_03779_));
 sg13g2_buf_1 _23803_ (.A(_03780_),
    .X(_03781_));
 sg13g2_nor2_1 _23804_ (.A(_03728_),
    .B(_03741_),
    .Y(_03782_));
 sg13g2_nand2_1 _23805_ (.Y(_03783_),
    .A(_03728_),
    .B(_03741_));
 sg13g2_o21ai_1 _23806_ (.B1(_03783_),
    .Y(_03784_),
    .A1(_03721_),
    .A2(_03782_));
 sg13g2_buf_1 _23807_ (.A(_03784_),
    .X(_03785_));
 sg13g2_xnor2_1 _23808_ (.Y(_03786_),
    .A(_03781_),
    .B(_03785_));
 sg13g2_nand2_1 _23809_ (.Y(_03787_),
    .A(_03726_),
    .B(_03727_));
 sg13g2_a21oi_1 _23810_ (.A1(_03781_),
    .A2(_03785_),
    .Y(_03788_),
    .B1(_03787_));
 sg13g2_a221oi_1 _23811_ (.B2(_03787_),
    .C1(_03788_),
    .B1(_03786_),
    .A1(_03749_),
    .Y(_03789_),
    .A2(_03751_));
 sg13g2_nand3b_1 _23812_ (.B(_03622_),
    .C(_03580_),
    .Y(_03790_),
    .A_N(_03623_));
 sg13g2_buf_1 _23813_ (.A(_03790_),
    .X(_03791_));
 sg13g2_and4_1 _23814_ (.A(_03606_),
    .B(_03612_),
    .C(_03619_),
    .D(_03621_),
    .X(_03792_));
 sg13g2_xor2_1 _23815_ (.B(_03579_),
    .A(_03309_),
    .X(_03793_));
 sg13g2_o21ai_1 _23816_ (.B1(_03793_),
    .Y(_03794_),
    .A1(_03623_),
    .A2(_03792_));
 sg13g2_buf_1 _23817_ (.A(_03794_),
    .X(_03795_));
 sg13g2_nand2b_1 _23818_ (.Y(_03796_),
    .B(_03778_),
    .A_N(_03754_));
 sg13g2_buf_1 _23819_ (.A(_03796_),
    .X(_03797_));
 sg13g2_nand2b_1 _23820_ (.Y(_03798_),
    .B(_03763_),
    .A_N(_03767_));
 sg13g2_buf_1 _23821_ (.A(_03798_),
    .X(_03799_));
 sg13g2_or2_1 _23822_ (.X(_03800_),
    .B(_03799_),
    .A(_03797_));
 sg13g2_and3_1 _23823_ (.X(_03801_),
    .A(_03791_),
    .B(_03795_),
    .C(_03800_));
 sg13g2_nand2_1 _23824_ (.Y(_03802_),
    .A(_03791_),
    .B(_03795_));
 sg13g2_nor2b_1 _23825_ (.A(_03778_),
    .B_N(_03754_),
    .Y(_03803_));
 sg13g2_a21oi_1 _23826_ (.A1(_03767_),
    .A2(_03797_),
    .Y(_03804_),
    .B1(_03803_));
 sg13g2_nand2_1 _23827_ (.Y(_03805_),
    .A(_03767_),
    .B(_03803_));
 sg13g2_o21ai_1 _23828_ (.B1(_03805_),
    .Y(_03806_),
    .A1(_03763_),
    .A2(_03804_));
 sg13g2_mux2_1 _23829_ (.A0(_03801_),
    .A1(_03802_),
    .S(_03806_),
    .X(_03807_));
 sg13g2_nand2b_1 _23830_ (.Y(_03808_),
    .B(_03754_),
    .A_N(_03778_));
 sg13g2_or2_1 _23831_ (.X(_03809_),
    .B(_03785_),
    .A(_03787_));
 sg13g2_and2_1 _23832_ (.A(_03787_),
    .B(_03785_),
    .X(_03810_));
 sg13g2_a21oi_1 _23833_ (.A1(_03781_),
    .A2(_03809_),
    .Y(_03811_),
    .B1(_03810_));
 sg13g2_a21oi_1 _23834_ (.A1(_03802_),
    .A2(_03808_),
    .Y(_03812_),
    .B1(_03811_));
 sg13g2_nor2_1 _23835_ (.A(_03802_),
    .B(_03808_),
    .Y(_03813_));
 sg13g2_o21ai_1 _23836_ (.B1(_03799_),
    .Y(_03814_),
    .A1(_03812_),
    .A2(_03813_));
 sg13g2_nand2b_1 _23837_ (.Y(_03815_),
    .B(_03767_),
    .A_N(_03763_));
 sg13g2_a21oi_1 _23838_ (.A1(_03811_),
    .A2(_03815_),
    .Y(_03816_),
    .B1(_03802_));
 sg13g2_nor2_1 _23839_ (.A(_03811_),
    .B(_03815_),
    .Y(_03817_));
 sg13g2_o21ai_1 _23840_ (.B1(_03797_),
    .Y(_03818_),
    .A1(_03816_),
    .A2(_03817_));
 sg13g2_a22oi_1 _23841_ (.Y(_03819_),
    .B1(_03814_),
    .B2(_03818_),
    .A2(_03807_),
    .A1(_03789_));
 sg13g2_xnor2_1 _23842_ (.Y(_03820_),
    .A(net105),
    .B(net94));
 sg13g2_xnor2_1 _23843_ (.Y(_03821_),
    .A(net88),
    .B(_03820_));
 sg13g2_xnor2_1 _23844_ (.Y(_03822_),
    .A(_03331_),
    .B(_03445_));
 sg13g2_xnor2_1 _23845_ (.Y(_03823_),
    .A(_03822_),
    .B(_03535_));
 sg13g2_xnor2_1 _23846_ (.Y(_03824_),
    .A(_03821_),
    .B(_03823_));
 sg13g2_xnor2_1 _23847_ (.Y(_03825_),
    .A(_03536_),
    .B(_03824_));
 sg13g2_xnor2_1 _23848_ (.Y(_03826_),
    .A(_03628_),
    .B(_03825_));
 sg13g2_or2_1 _23849_ (.X(_03827_),
    .B(_03561_),
    .A(_03559_));
 sg13g2_xor2_1 _23850_ (.B(_03625_),
    .A(_03577_),
    .X(_03828_));
 sg13g2_xnor2_1 _23851_ (.Y(_03829_),
    .A(_03827_),
    .B(_03828_));
 sg13g2_nand3b_1 _23852_ (.B(_03826_),
    .C(_03829_),
    .Y(_03830_),
    .A_N(_03819_));
 sg13g2_xnor2_1 _23853_ (.Y(_03831_),
    .A(_03635_),
    .B(_03525_));
 sg13g2_xnor2_1 _23854_ (.Y(_03832_),
    .A(net79),
    .B(_03831_));
 sg13g2_xnor2_1 _23855_ (.Y(_03833_),
    .A(_03472_),
    .B(_03832_));
 sg13g2_buf_2 _23856_ (.A(_03833_),
    .X(_03834_));
 sg13g2_a21oi_1 _23857_ (.A1(_03540_),
    .A2(_03630_),
    .Y(_03835_),
    .B1(_03552_));
 sg13g2_or4_1 _23858_ (.A(_03701_),
    .B(_03830_),
    .C(_03834_),
    .D(_03835_),
    .X(_03836_));
 sg13g2_a21o_1 _23859_ (.A2(_03692_),
    .A1(_03672_),
    .B1(_03836_),
    .X(_03837_));
 sg13g2_buf_8 _23860_ (.A(_03837_),
    .X(_03838_));
 sg13g2_nor2_1 _23861_ (.A(_03676_),
    .B(_03680_),
    .Y(_03839_));
 sg13g2_nand3_1 _23862_ (.B(_03515_),
    .C(_03524_),
    .A(_03685_),
    .Y(_03840_));
 sg13g2_a21o_1 _23863_ (.A2(_03840_),
    .A1(net79),
    .B1(_03686_),
    .X(_03841_));
 sg13g2_buf_1 _23864_ (.A(_03841_),
    .X(_03842_));
 sg13g2_xnor2_1 _23865_ (.Y(_03843_),
    .A(_03678_),
    .B(_03842_));
 sg13g2_nor4_1 _23866_ (.A(_03701_),
    .B(_03832_),
    .C(_03839_),
    .D(_03843_),
    .Y(_03844_));
 sg13g2_buf_1 _23867_ (.A(_03844_),
    .X(_03845_));
 sg13g2_xnor2_1 _23868_ (.Y(_03846_),
    .A(_03017_),
    .B(_03063_));
 sg13g2_and2_1 _23869_ (.A(_03018_),
    .B(_03063_),
    .X(_03847_));
 sg13g2_mux2_1 _23870_ (.A0(_03846_),
    .A1(_03847_),
    .S(_02978_),
    .X(_03848_));
 sg13g2_buf_1 _23871_ (.A(_03848_),
    .X(_03849_));
 sg13g2_xor2_1 _23872_ (.B(_03849_),
    .A(_03205_),
    .X(_03850_));
 sg13g2_nor2_1 _23873_ (.A(_03656_),
    .B(_03696_),
    .Y(_03851_));
 sg13g2_o21ai_1 _23874_ (.B1(_03842_),
    .Y(_03852_),
    .A1(_03697_),
    .A2(_03851_));
 sg13g2_nand2_1 _23875_ (.Y(_03853_),
    .A(_03657_),
    .B(_03697_));
 sg13g2_nand3b_1 _23876_ (.B(_03657_),
    .C(_03842_),
    .Y(_03854_),
    .A_N(_03638_));
 sg13g2_nand4_1 _23877_ (.B(_03852_),
    .C(_03853_),
    .A(_03694_),
    .Y(_03855_),
    .D(_03854_));
 sg13g2_buf_1 _23878_ (.A(_03855_),
    .X(_03856_));
 sg13g2_nor2_1 _23879_ (.A(_03850_),
    .B(_03856_),
    .Y(_03857_));
 sg13g2_nor2_1 _23880_ (.A(_03845_),
    .B(_03857_),
    .Y(_03858_));
 sg13g2_a22oi_1 _23881_ (.Y(_03859_),
    .B1(_02812_),
    .B2(_02970_),
    .A2(_02694_),
    .A1(_02679_));
 sg13g2_nand2_1 _23882_ (.Y(_03860_),
    .A(_02962_),
    .B(_03859_));
 sg13g2_nor2_1 _23883_ (.A(_03066_),
    .B(net77),
    .Y(_03861_));
 sg13g2_nor2_1 _23884_ (.A(_02961_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_or3_1 _23885_ (.A(_02887_),
    .B(_03859_),
    .C(_03862_),
    .X(_03863_));
 sg13g2_xnor2_1 _23886_ (.Y(_03864_),
    .A(_03208_),
    .B(_03212_));
 sg13g2_buf_2 _23887_ (.A(_03864_),
    .X(_03865_));
 sg13g2_nor2_1 _23888_ (.A(net74),
    .B(_03865_),
    .Y(_03866_));
 sg13g2_nand2_1 _23889_ (.Y(_03867_),
    .A(_03850_),
    .B(_03856_));
 sg13g2_nand4_1 _23890_ (.B(_03863_),
    .C(_03866_),
    .A(_03860_),
    .Y(_03868_),
    .D(_03867_));
 sg13g2_a21oi_1 _23891_ (.A1(_03838_),
    .A2(_03858_),
    .Y(_03869_),
    .B1(_03868_));
 sg13g2_and2_1 _23892_ (.A(_02737_),
    .B(_02809_),
    .X(_03870_));
 sg13g2_o21ai_1 _23893_ (.B1(net192),
    .Y(_03871_),
    .A1(_02737_),
    .A2(_02809_));
 sg13g2_nor3_1 _23894_ (.A(_02798_),
    .B(_03870_),
    .C(_03871_),
    .Y(_03872_));
 sg13g2_inv_1 _23895_ (.Y(_03873_),
    .A(_03872_));
 sg13g2_a22oi_1 _23896_ (.Y(_03874_),
    .B1(_03000_),
    .B2(_02784_),
    .A2(_02785_),
    .A1(net165));
 sg13g2_inv_1 _23897_ (.Y(_03875_),
    .A(_03874_));
 sg13g2_a21oi_1 _23898_ (.A1(net197),
    .A2(_03023_),
    .Y(_03876_),
    .B1(_02834_));
 sg13g2_o21ai_1 _23899_ (.B1(_03876_),
    .Y(_03877_),
    .A1(_02743_),
    .A2(_03875_));
 sg13g2_a21oi_1 _23900_ (.A1(_03873_),
    .A2(_03877_),
    .Y(_03878_),
    .B1(_02679_));
 sg13g2_nor3_1 _23901_ (.A(_03215_),
    .B(_03869_),
    .C(_03878_),
    .Y(_03879_));
 sg13g2_buf_1 _23902_ (.A(_03879_),
    .X(_03880_));
 sg13g2_inv_2 _23903_ (.Y(_03881_),
    .A(_03850_));
 sg13g2_inv_1 _23904_ (.Y(_03882_),
    .A(_03694_));
 sg13g2_o21ai_1 _23905_ (.B1(net79),
    .Y(_03883_),
    .A1(_03454_),
    .A2(_03471_));
 sg13g2_nand3_1 _23906_ (.B(_03674_),
    .C(_03666_),
    .A(_03673_),
    .Y(_03884_));
 sg13g2_nand3b_1 _23907_ (.B(_03668_),
    .C(_03667_),
    .Y(_03885_),
    .A_N(_03840_));
 sg13g2_a22oi_1 _23908_ (.Y(_03886_),
    .B1(_03885_),
    .B2(_03687_),
    .A2(_03884_),
    .A1(_03883_));
 sg13g2_a221oi_1 _23909_ (.B2(_03681_),
    .C1(_03454_),
    .B1(_03683_),
    .A1(_03456_),
    .Y(_03887_),
    .A2(_03470_));
 sg13g2_and3_1 _23910_ (.X(_03888_),
    .A(_03673_),
    .B(_03674_),
    .C(_03686_));
 sg13g2_nor4_1 _23911_ (.A(_03678_),
    .B(_03689_),
    .C(_03887_),
    .D(_03888_),
    .Y(_03889_));
 sg13g2_nor4_1 _23912_ (.A(_03502_),
    .B(_03831_),
    .C(_03663_),
    .D(_03664_),
    .Y(_03890_));
 sg13g2_and2_1 _23913_ (.A(_03676_),
    .B(_03890_),
    .X(_03891_));
 sg13g2_nor4_1 _23914_ (.A(_03676_),
    .B(_03666_),
    .C(_03831_),
    .D(_03678_),
    .Y(_03892_));
 sg13g2_or4_1 _23915_ (.A(_03886_),
    .B(_03889_),
    .C(_03891_),
    .D(_03892_),
    .X(_03893_));
 sg13g2_buf_1 _23916_ (.A(_03893_),
    .X(_03894_));
 sg13g2_nor2b_1 _23917_ (.A(_03754_),
    .B_N(_03778_),
    .Y(_03895_));
 sg13g2_a21oi_1 _23918_ (.A1(_03808_),
    .A2(_03815_),
    .Y(_03896_),
    .B1(_03895_));
 sg13g2_a21o_1 _23919_ (.A2(_03795_),
    .A1(_03791_),
    .B1(_03896_),
    .X(_03897_));
 sg13g2_nor3_1 _23920_ (.A(_03626_),
    .B(_03625_),
    .C(_03897_),
    .Y(_03898_));
 sg13g2_and3_1 _23921_ (.X(_03899_),
    .A(_03791_),
    .B(_03795_),
    .C(_03797_));
 sg13g2_nor4_1 _23922_ (.A(_03899_),
    .B(_03799_),
    .C(_03626_),
    .D(_03625_),
    .Y(_03900_));
 sg13g2_nor4_2 _23923_ (.A(_03535_),
    .B(_03538_),
    .C(_03898_),
    .Y(_03901_),
    .D(_03900_));
 sg13g2_o21ai_1 _23924_ (.B1(_03897_),
    .Y(_03902_),
    .A1(_03899_),
    .A2(_03799_));
 sg13g2_a221oi_1 _23925_ (.B2(_03902_),
    .C1(_03628_),
    .B1(_03829_),
    .A1(_03535_),
    .Y(_03903_),
    .A2(_03538_));
 sg13g2_nor2_2 _23926_ (.A(_03901_),
    .B(_03903_),
    .Y(_03904_));
 sg13g2_and2_1 _23927_ (.A(_03807_),
    .B(_03829_),
    .X(_03905_));
 sg13g2_nand2_1 _23928_ (.Y(_03906_),
    .A(_03781_),
    .B(_03785_));
 sg13g2_o21ai_1 _23929_ (.B1(_03787_),
    .Y(_03907_),
    .A1(_03781_),
    .A2(_03785_));
 sg13g2_nand3_1 _23930_ (.B(_03748_),
    .C(_03751_),
    .A(_03746_),
    .Y(_03908_));
 sg13g2_a21oi_1 _23931_ (.A1(_03906_),
    .A2(_03907_),
    .Y(_03909_),
    .B1(_03908_));
 sg13g2_a21oi_1 _23932_ (.A1(_03781_),
    .A2(_03810_),
    .Y(_03910_),
    .B1(_03909_));
 sg13g2_and3_1 _23933_ (.X(_03911_),
    .A(_03826_),
    .B(_03905_),
    .C(_03910_));
 sg13g2_o21ai_1 _23934_ (.B1(_03552_),
    .Y(_03912_),
    .A1(_03904_),
    .A2(_03911_));
 sg13g2_nand2b_1 _23935_ (.Y(_03913_),
    .B(_03912_),
    .A_N(_03889_));
 sg13g2_buf_2 _23936_ (.A(_03913_),
    .X(_03914_));
 sg13g2_a21oi_1 _23937_ (.A1(_03894_),
    .A2(_03914_),
    .Y(_03915_),
    .B1(_03699_));
 sg13g2_nand3_1 _23938_ (.B(_03894_),
    .C(_03914_),
    .A(_03699_),
    .Y(_03916_));
 sg13g2_o21ai_1 _23939_ (.B1(_03916_),
    .Y(_03917_),
    .A1(_03882_),
    .A2(_03915_));
 sg13g2_buf_1 _23940_ (.A(_03917_),
    .X(_03918_));
 sg13g2_a21oi_2 _23941_ (.B1(_03865_),
    .Y(_03919_),
    .A2(_03918_),
    .A1(_03881_));
 sg13g2_and3_1 _23942_ (.X(_03920_),
    .A(_03881_),
    .B(_03865_),
    .C(_03918_));
 sg13g2_buf_1 _23943_ (.A(_03920_),
    .X(_03921_));
 sg13g2_nand2b_1 _23944_ (.Y(_03922_),
    .B(_03063_),
    .A_N(_02978_));
 sg13g2_inv_1 _23945_ (.Y(_03923_),
    .A(_03922_));
 sg13g2_a21oi_1 _23946_ (.A1(_03923_),
    .A2(_03206_),
    .Y(_03924_),
    .B1(net77));
 sg13g2_nor2b_1 _23947_ (.A(net77),
    .B_N(net74),
    .Y(_03925_));
 sg13g2_nor2_1 _23948_ (.A(_03018_),
    .B(net78),
    .Y(_03926_));
 sg13g2_o21ai_1 _23949_ (.B1(_03922_),
    .Y(_03927_),
    .A1(_03925_),
    .A2(_03926_));
 sg13g2_o21ai_1 _23950_ (.B1(_03927_),
    .Y(_03928_),
    .A1(net74),
    .A2(_03924_));
 sg13g2_nand2b_1 _23951_ (.Y(_03929_),
    .B(_02978_),
    .A_N(_03063_));
 sg13g2_a21oi_1 _23952_ (.A1(_03018_),
    .A2(net78),
    .Y(_03930_),
    .B1(_03929_));
 sg13g2_nor2_1 _23953_ (.A(_03207_),
    .B(_03925_),
    .Y(_03931_));
 sg13g2_nand2_1 _23954_ (.Y(_03932_),
    .A(net78),
    .B(_03849_));
 sg13g2_o21ai_1 _23955_ (.B1(_03932_),
    .Y(_03933_),
    .A1(net78),
    .A2(_03931_));
 sg13g2_nor3_1 _23956_ (.A(_03928_),
    .B(_03930_),
    .C(_03933_),
    .Y(_03934_));
 sg13g2_nor2b_1 _23957_ (.A(_03208_),
    .B_N(net74),
    .Y(_03935_));
 sg13g2_a221oi_1 _23958_ (.B2(net77),
    .C1(_03214_),
    .B1(_03935_),
    .A1(_03856_),
    .Y(_03936_),
    .A2(_03934_));
 sg13g2_inv_1 _23959_ (.Y(_03937_),
    .A(_03856_));
 sg13g2_xnor2_1 _23960_ (.Y(_03938_),
    .A(_02978_),
    .B(net78));
 sg13g2_nor2_1 _23961_ (.A(_03064_),
    .B(net77),
    .Y(_03939_));
 sg13g2_nand2b_1 _23962_ (.Y(_03940_),
    .B(net78),
    .A_N(_02978_));
 sg13g2_nand3b_1 _23963_ (.B(net77),
    .C(_02978_),
    .Y(_03941_),
    .A_N(net78));
 sg13g2_o21ai_1 _23964_ (.B1(_03941_),
    .Y(_03942_),
    .A1(net77),
    .A2(_03940_));
 sg13g2_a22oi_1 _23965_ (.Y(_03943_),
    .B1(_03942_),
    .B2(_03846_),
    .A2(_03939_),
    .A1(_03938_));
 sg13g2_nor2_1 _23966_ (.A(net74),
    .B(_03943_),
    .Y(_03944_));
 sg13g2_o21ai_1 _23967_ (.B1(_03944_),
    .Y(_03945_),
    .A1(_03845_),
    .A2(_03937_));
 sg13g2_nand2_1 _23968_ (.Y(_03946_),
    .A(_03866_),
    .B(_03867_));
 sg13g2_xor2_1 _23969_ (.B(_03213_),
    .A(net74),
    .X(_03947_));
 sg13g2_or3_1 _23970_ (.A(_03845_),
    .B(_03857_),
    .C(_03947_),
    .X(_03948_));
 sg13g2_mux2_1 _23971_ (.A0(_03946_),
    .A1(_03948_),
    .S(_03838_),
    .X(_03949_));
 sg13g2_and3_1 _23972_ (.X(_03950_),
    .A(_03936_),
    .B(_03945_),
    .C(_03949_));
 sg13g2_buf_2 _23973_ (.A(_03950_),
    .X(_03951_));
 sg13g2_or4_1 _23974_ (.A(_03701_),
    .B(_03832_),
    .C(_03839_),
    .D(_03843_),
    .X(_03952_));
 sg13g2_xnor2_1 _23975_ (.Y(_03953_),
    .A(_03881_),
    .B(_03856_));
 sg13g2_inv_1 _23976_ (.Y(_03954_),
    .A(_03953_));
 sg13g2_a21oi_2 _23977_ (.B1(_03954_),
    .Y(_03955_),
    .A2(_03952_),
    .A1(_03838_));
 sg13g2_a21oi_1 _23978_ (.A1(_03672_),
    .A2(_03692_),
    .Y(_03956_),
    .B1(_03836_));
 sg13g2_nor3_2 _23979_ (.A(_03956_),
    .B(_03845_),
    .C(_03953_),
    .Y(_03957_));
 sg13g2_a21o_1 _23980_ (.A2(_03665_),
    .A1(_03632_),
    .B1(_03671_),
    .X(_03958_));
 sg13g2_or4_1 _23981_ (.A(_03682_),
    .B(_03684_),
    .C(_03688_),
    .D(_03691_),
    .X(_03959_));
 sg13g2_xnor2_1 _23982_ (.Y(_03960_),
    .A(_03456_),
    .B(_03550_));
 sg13g2_xnor2_1 _23983_ (.Y(_03961_),
    .A(_03960_),
    .B(_03904_));
 sg13g2_nand3_1 _23984_ (.B(_03905_),
    .C(_03910_),
    .A(_03826_),
    .Y(_03962_));
 sg13g2_buf_1 _23985_ (.A(_03962_),
    .X(_03963_));
 sg13g2_nand2b_1 _23986_ (.Y(_03964_),
    .B(_03825_),
    .A_N(_03628_));
 sg13g2_o21ai_1 _23987_ (.B1(_03628_),
    .Y(_03965_),
    .A1(_03535_),
    .A2(_03538_));
 sg13g2_and2_1 _23988_ (.A(_03829_),
    .B(_03902_),
    .X(_03966_));
 sg13g2_nand4_1 _23989_ (.B(_03552_),
    .C(_03965_),
    .A(_03964_),
    .Y(_03967_),
    .D(_03966_));
 sg13g2_buf_1 _23990_ (.A(_03967_),
    .X(_03968_));
 sg13g2_o21ai_1 _23991_ (.B1(_03968_),
    .Y(_03969_),
    .A1(_03552_),
    .A2(_03963_));
 sg13g2_xnor2_1 _23992_ (.Y(_03970_),
    .A(_03676_),
    .B(_03832_));
 sg13g2_o21ai_1 _23993_ (.B1(_03970_),
    .Y(_03971_),
    .A1(_03961_),
    .A2(_03969_));
 sg13g2_buf_2 _23994_ (.A(_03971_),
    .X(_03972_));
 sg13g2_nor3_2 _23995_ (.A(_03958_),
    .B(_03959_),
    .C(_03972_),
    .Y(_03973_));
 sg13g2_nor3_2 _23996_ (.A(_03830_),
    .B(_03834_),
    .C(_03835_),
    .Y(_03974_));
 sg13g2_a21oi_2 _23997_ (.B1(_03974_),
    .Y(_03975_),
    .A2(_03692_),
    .A1(_03672_));
 sg13g2_a21oi_1 _23998_ (.A1(_03894_),
    .A2(_03914_),
    .Y(_03976_),
    .B1(_03701_));
 sg13g2_and3_1 _23999_ (.X(_03977_),
    .A(_03701_),
    .B(_03894_),
    .C(_03914_));
 sg13g2_buf_1 _24000_ (.A(_03977_),
    .X(_03978_));
 sg13g2_nor4_1 _24001_ (.A(_03973_),
    .B(_03975_),
    .C(_03976_),
    .D(_03978_),
    .Y(_03979_));
 sg13g2_buf_2 _24002_ (.A(_03979_),
    .X(_03980_));
 sg13g2_o21ai_1 _24003_ (.B1(_03980_),
    .Y(_03981_),
    .A1(_03955_),
    .A2(_03957_));
 sg13g2_buf_1 _24004_ (.A(_03981_),
    .X(_03982_));
 sg13g2_nor4_1 _24005_ (.A(_03919_),
    .B(_03921_),
    .C(_03951_),
    .D(_03982_),
    .Y(_03983_));
 sg13g2_buf_2 _24006_ (.A(_03983_),
    .X(_03984_));
 sg13g2_nor2_1 _24007_ (.A(net48),
    .B(_03984_),
    .Y(_03985_));
 sg13g2_buf_2 _24008_ (.A(_03985_),
    .X(_03986_));
 sg13g2_buf_1 _24009_ (.A(_03986_),
    .X(_03987_));
 sg13g2_nor3_2 _24010_ (.A(_03875_),
    .B(_02834_),
    .C(net96),
    .Y(_03988_));
 sg13g2_o21ai_1 _24011_ (.B1(_03875_),
    .Y(_03989_),
    .A1(_02738_),
    .A2(net96));
 sg13g2_a21oi_1 _24012_ (.A1(_02815_),
    .A2(_03989_),
    .Y(_03990_),
    .B1(_02817_));
 sg13g2_and2_1 _24013_ (.A(_03872_),
    .B(_03877_),
    .X(_03991_));
 sg13g2_nor4_2 _24014_ (.A(_03215_),
    .B(_03869_),
    .C(_03990_),
    .Y(_03992_),
    .D(_03991_));
 sg13g2_nor2_1 _24015_ (.A(_03984_),
    .B(_03992_),
    .Y(_03993_));
 sg13g2_nor2_1 _24016_ (.A(_03988_),
    .B(_03993_),
    .Y(_03994_));
 sg13g2_buf_2 _24017_ (.A(_03994_),
    .X(_03995_));
 sg13g2_buf_1 _24018_ (.A(_02695_),
    .X(_03996_));
 sg13g2_nand4_1 _24019_ (.B(_02815_),
    .C(_03874_),
    .A(_02807_),
    .Y(_03997_),
    .D(net95));
 sg13g2_buf_1 _24020_ (.A(_03997_),
    .X(_03998_));
 sg13g2_nand2_1 _24021_ (.Y(_03999_),
    .A(net192),
    .B(_03998_));
 sg13g2_a221oi_1 _24022_ (.B2(net80),
    .C1(_03999_),
    .B1(_03995_),
    .A1(net107),
    .Y(_04000_),
    .A2(net32));
 sg13g2_buf_1 _24023_ (.A(net120),
    .X(_04001_));
 sg13g2_or4_1 _24024_ (.A(_03919_),
    .B(_03921_),
    .C(_03951_),
    .D(_03982_),
    .X(_04002_));
 sg13g2_buf_1 _24025_ (.A(_04002_),
    .X(_04003_));
 sg13g2_buf_1 _24026_ (.A(net38),
    .X(_04004_));
 sg13g2_nand2_1 _24027_ (.Y(_04005_),
    .A(_03694_),
    .B(_03699_));
 sg13g2_nand2_1 _24028_ (.Y(_04006_),
    .A(_03206_),
    .B(_04005_));
 sg13g2_or2_1 _24029_ (.X(_04007_),
    .B(_03211_),
    .A(_02974_));
 sg13g2_nor2b_1 _24030_ (.A(_04007_),
    .B_N(_03849_),
    .Y(_04008_));
 sg13g2_nor4_1 _24031_ (.A(net74),
    .B(_03701_),
    .C(_03850_),
    .D(_03865_),
    .Y(_04009_));
 sg13g2_and2_1 _24032_ (.A(_03894_),
    .B(_03914_),
    .X(_04010_));
 sg13g2_nand2_1 _24033_ (.Y(_04011_),
    .A(_03860_),
    .B(_03863_));
 sg13g2_a221oi_1 _24034_ (.B2(_04010_),
    .C1(_04011_),
    .B1(_04009_),
    .A1(_04006_),
    .Y(_04012_),
    .A2(_04008_));
 sg13g2_buf_1 _24035_ (.A(_04012_),
    .X(_04013_));
 sg13g2_inv_1 _24036_ (.Y(_04014_),
    .A(_04013_));
 sg13g2_nand2_1 _24037_ (.Y(_04015_),
    .A(net37),
    .B(_04014_));
 sg13g2_nor2_1 _24038_ (.A(net103),
    .B(_04015_),
    .Y(_04016_));
 sg13g2_buf_1 _24039_ (.A(net119),
    .X(_04017_));
 sg13g2_buf_1 _24040_ (.A(_03951_),
    .X(_04018_));
 sg13g2_a21o_1 _24041_ (.A2(_03918_),
    .A1(_03881_),
    .B1(_03865_),
    .X(_04019_));
 sg13g2_buf_2 _24042_ (.A(_04019_),
    .X(_04020_));
 sg13g2_nand3_1 _24043_ (.B(_03865_),
    .C(_03918_),
    .A(_03881_),
    .Y(_04021_));
 sg13g2_buf_2 _24044_ (.A(_04021_),
    .X(_04022_));
 sg13g2_nand2_1 _24045_ (.Y(_04023_),
    .A(_03672_),
    .B(_03692_));
 sg13g2_buf_2 _24046_ (.A(_04023_),
    .X(_04024_));
 sg13g2_nand2_1 _24047_ (.Y(_04025_),
    .A(_03974_),
    .B(_04024_));
 sg13g2_nor2_1 _24048_ (.A(_03958_),
    .B(_03959_),
    .Y(_04026_));
 sg13g2_nand2_1 _24049_ (.Y(_04027_),
    .A(_04026_),
    .B(_03972_));
 sg13g2_o21ai_1 _24050_ (.B1(_03953_),
    .Y(_04028_),
    .A1(_03956_),
    .A2(_03845_));
 sg13g2_buf_2 _24051_ (.A(_04028_),
    .X(_04029_));
 sg13g2_nand3_1 _24052_ (.B(_03952_),
    .C(_03954_),
    .A(_03838_),
    .Y(_04030_));
 sg13g2_buf_1 _24053_ (.A(_04030_),
    .X(_04031_));
 sg13g2_or2_1 _24054_ (.X(_04032_),
    .B(_03978_),
    .A(_03976_));
 sg13g2_buf_1 _24055_ (.A(_04032_),
    .X(_04033_));
 sg13g2_a221oi_1 _24056_ (.B2(_04031_),
    .C1(net52),
    .B1(_04029_),
    .A1(_04025_),
    .Y(_04034_),
    .A2(_04027_));
 sg13g2_buf_1 _24057_ (.A(_04034_),
    .X(_04035_));
 sg13g2_buf_8 _24058_ (.A(_04035_),
    .X(_04036_));
 sg13g2_nand3_1 _24059_ (.B(_04022_),
    .C(net42),
    .A(_04020_),
    .Y(_04037_));
 sg13g2_buf_1 _24060_ (.A(_04037_),
    .X(_04038_));
 sg13g2_buf_8 _24061_ (.A(_04038_),
    .X(_04039_));
 sg13g2_nand2_1 _24062_ (.Y(_04040_),
    .A(net46),
    .B(net33));
 sg13g2_buf_1 _24063_ (.A(_04040_),
    .X(_04041_));
 sg13g2_o21ai_1 _24064_ (.B1(net32),
    .Y(_04042_),
    .A1(net102),
    .A2(_04041_));
 sg13g2_buf_1 _24065_ (.A(net106),
    .X(_04043_));
 sg13g2_o21ai_1 _24066_ (.B1(_03986_),
    .Y(_04044_),
    .A1(net93),
    .A2(net102));
 sg13g2_buf_1 _24067_ (.A(_03422_),
    .X(_04045_));
 sg13g2_nor2_2 _24068_ (.A(net103),
    .B(net101),
    .Y(_04046_));
 sg13g2_buf_8 _24069_ (.A(_03984_),
    .X(_04047_));
 sg13g2_buf_1 _24070_ (.A(_04013_),
    .X(_04048_));
 sg13g2_nor2_1 _24071_ (.A(net36),
    .B(net51),
    .Y(_04049_));
 sg13g2_and2_1 _24072_ (.A(_04046_),
    .B(_04049_),
    .X(_04050_));
 sg13g2_a21o_1 _24073_ (.A2(_04044_),
    .A1(net96),
    .B1(_04050_),
    .X(_04051_));
 sg13g2_a21oi_1 _24074_ (.A1(_03951_),
    .A2(_04038_),
    .Y(_04052_),
    .B1(_03984_));
 sg13g2_buf_2 _24075_ (.A(_04052_),
    .X(_04053_));
 sg13g2_buf_1 _24076_ (.A(net46),
    .X(_04054_));
 sg13g2_o21ai_1 _24077_ (.B1(net41),
    .Y(_04055_),
    .A1(net93),
    .A2(net33));
 sg13g2_nand2_1 _24078_ (.Y(_04056_),
    .A(net93),
    .B(net33));
 sg13g2_and2_1 _24079_ (.A(_04055_),
    .B(_04056_),
    .X(_04057_));
 sg13g2_nor4_1 _24080_ (.A(net101),
    .B(net48),
    .C(_04057_),
    .D(_04016_),
    .Y(_04058_));
 sg13g2_a221oi_1 _24081_ (.B2(_04053_),
    .C1(_04058_),
    .B1(_04051_),
    .A1(_04016_),
    .Y(_04059_),
    .A2(_04042_));
 sg13g2_inv_2 _24082_ (.Y(_04060_),
    .A(net48));
 sg13g2_nand3_1 _24083_ (.B(net33),
    .C(net51),
    .A(net41),
    .Y(_04061_));
 sg13g2_a21oi_1 _24084_ (.A1(net41),
    .A2(net33),
    .Y(_04062_),
    .B1(net51));
 sg13g2_a21o_1 _24085_ (.A2(_04061_),
    .A1(_04060_),
    .B1(_04062_),
    .X(_04063_));
 sg13g2_and2_1 _24086_ (.A(_03881_),
    .B(_03918_),
    .X(_04064_));
 sg13g2_buf_1 _24087_ (.A(_04064_),
    .X(_04065_));
 sg13g2_xnor2_1 _24088_ (.Y(_04066_),
    .A(_03865_),
    .B(_04035_));
 sg13g2_xor2_1 _24089_ (.B(_04066_),
    .A(_04065_),
    .X(_04067_));
 sg13g2_buf_2 _24090_ (.A(_04067_),
    .X(_04068_));
 sg13g2_nor3_1 _24091_ (.A(_03128_),
    .B(_04068_),
    .C(_04048_),
    .Y(_04069_));
 sg13g2_a21oi_1 _24092_ (.A1(net93),
    .A2(_04063_),
    .Y(_04070_),
    .B1(_04069_));
 sg13g2_nor3_1 _24093_ (.A(net101),
    .B(net36),
    .C(_04070_),
    .Y(_04071_));
 sg13g2_nor2_1 _24094_ (.A(_04059_),
    .B(_04071_),
    .Y(_04072_));
 sg13g2_xnor2_1 _24095_ (.Y(_04073_),
    .A(_04000_),
    .B(_04072_));
 sg13g2_and3_1 _24096_ (.X(_04074_),
    .A(_03980_),
    .B(_04029_),
    .C(_04031_));
 sg13g2_buf_1 _24097_ (.A(_04074_),
    .X(_04075_));
 sg13g2_a21oi_1 _24098_ (.A1(_04029_),
    .A2(_04031_),
    .Y(_04076_),
    .B1(_03980_));
 sg13g2_nor2_2 _24099_ (.A(_04075_),
    .B(_04076_),
    .Y(_04077_));
 sg13g2_nor2_1 _24100_ (.A(net101),
    .B(_04077_),
    .Y(_04078_));
 sg13g2_nor2_2 _24101_ (.A(net103),
    .B(_04077_),
    .Y(_04079_));
 sg13g2_xnor2_1 _24102_ (.Y(_04080_),
    .A(_04065_),
    .B(_04066_));
 sg13g2_buf_1 _24103_ (.A(_04080_),
    .X(_04081_));
 sg13g2_a22oi_1 _24104_ (.Y(_04082_),
    .B1(_04079_),
    .B2(net35),
    .A2(_04078_),
    .A1(_04053_));
 sg13g2_nand3b_1 _24105_ (.B(net35),
    .C(_04046_),
    .Y(_04083_),
    .A_N(net41));
 sg13g2_o21ai_1 _24106_ (.B1(_04083_),
    .Y(_04084_),
    .A1(_03128_),
    .A2(_04082_));
 sg13g2_and3_1 _24107_ (.X(_04085_),
    .A(_03986_),
    .B(_04046_),
    .C(_04061_));
 sg13g2_nor3_2 _24108_ (.A(_03919_),
    .B(_03921_),
    .C(_03982_),
    .Y(_04086_));
 sg13g2_xnor2_1 _24109_ (.Y(_04087_),
    .A(_04018_),
    .B(_04086_));
 sg13g2_a22oi_1 _24110_ (.Y(_04088_),
    .B1(_04087_),
    .B2(net93),
    .A2(net35),
    .A1(net96));
 sg13g2_nor2_1 _24111_ (.A(net101),
    .B(_04015_),
    .Y(_04089_));
 sg13g2_o21ai_1 _24112_ (.B1(_04089_),
    .Y(_04090_),
    .A1(_04085_),
    .A2(_04088_));
 sg13g2_or3_1 _24113_ (.A(_04085_),
    .B(_04088_),
    .C(_04089_),
    .X(_04091_));
 sg13g2_buf_1 _24114_ (.A(_02986_),
    .X(_04092_));
 sg13g2_buf_1 _24115_ (.A(net92),
    .X(_04093_));
 sg13g2_xnor2_1 _24116_ (.Y(_04094_),
    .A(net147),
    .B(_02692_));
 sg13g2_a22oi_1 _24117_ (.Y(_04095_),
    .B1(_04094_),
    .B2(_03987_),
    .A2(_03995_),
    .A1(net87));
 sg13g2_a21oi_1 _24118_ (.A1(_04090_),
    .A2(_04091_),
    .Y(_04096_),
    .B1(_04095_));
 sg13g2_or2_1 _24119_ (.X(_04097_),
    .B(_04096_),
    .A(_04084_));
 sg13g2_buf_1 _24120_ (.A(_04097_),
    .X(_04098_));
 sg13g2_nand2_1 _24121_ (.Y(_04099_),
    .A(_04073_),
    .B(_04098_));
 sg13g2_buf_1 _24122_ (.A(_02815_),
    .X(_04100_));
 sg13g2_nand2_1 _24123_ (.Y(_04101_),
    .A(net37),
    .B(_04041_));
 sg13g2_a21oi_1 _24124_ (.A1(net32),
    .A2(_04046_),
    .Y(_04102_),
    .B1(_04101_));
 sg13g2_nor2_1 _24125_ (.A(_02738_),
    .B(_02815_),
    .Y(_04103_));
 sg13g2_buf_1 _24126_ (.A(_04103_),
    .X(_04104_));
 sg13g2_a221oi_1 _24127_ (.B2(net96),
    .C1(_04104_),
    .B1(_04102_),
    .A1(net107),
    .Y(_04105_),
    .A2(_03995_));
 sg13g2_nor2_1 _24128_ (.A(_04000_),
    .B(_04059_),
    .Y(_04106_));
 sg13g2_nor2_1 _24129_ (.A(_04071_),
    .B(_04106_),
    .Y(_04107_));
 sg13g2_xnor2_1 _24130_ (.Y(_04108_),
    .A(_04105_),
    .B(_04107_));
 sg13g2_a21oi_1 _24131_ (.A1(net241),
    .A2(_04108_),
    .Y(_04109_),
    .B1(_04104_));
 sg13g2_nor2b_1 _24132_ (.A(_04099_),
    .B_N(_04109_),
    .Y(_04110_));
 sg13g2_nand2b_1 _24133_ (.Y(_04111_),
    .B(_04106_),
    .A_N(_04071_));
 sg13g2_and2_1 _24134_ (.A(net32),
    .B(_04061_),
    .X(_04112_));
 sg13g2_nand2_1 _24135_ (.Y(_04113_),
    .A(_04060_),
    .B(net37));
 sg13g2_o21ai_1 _24136_ (.B1(net103),
    .Y(_04114_),
    .A1(net102),
    .A2(_04113_));
 sg13g2_o21ai_1 _24137_ (.B1(_04114_),
    .Y(_04115_),
    .A1(net32),
    .A2(_03995_));
 sg13g2_a22oi_1 _24138_ (.Y(_04116_),
    .B1(_04115_),
    .B2(_03998_),
    .A2(_04112_),
    .A1(_04046_));
 sg13g2_nand2_1 _24139_ (.Y(_04117_),
    .A(_04111_),
    .B(_04116_));
 sg13g2_o21ai_1 _24140_ (.B1(_04100_),
    .Y(_04118_),
    .A1(_04110_),
    .A2(_04117_));
 sg13g2_buf_1 _24141_ (.A(_04118_),
    .X(_04119_));
 sg13g2_nand2_1 _24142_ (.Y(_04120_),
    .A(_02761_),
    .B(net83));
 sg13g2_nand2b_1 _24143_ (.Y(_04121_),
    .B(net32),
    .A_N(_04120_));
 sg13g2_buf_1 _24144_ (.A(_04121_),
    .X(_04122_));
 sg13g2_buf_1 _24145_ (.A(_03982_),
    .X(_04123_));
 sg13g2_nor2_2 _24146_ (.A(_03973_),
    .B(_03975_),
    .Y(_04124_));
 sg13g2_nor2_1 _24147_ (.A(_03976_),
    .B(_03978_),
    .Y(_04125_));
 sg13g2_buf_2 _24148_ (.A(_04125_),
    .X(_04126_));
 sg13g2_xnor2_1 _24149_ (.Y(_04127_),
    .A(_04124_),
    .B(_04126_));
 sg13g2_buf_1 _24150_ (.A(_04127_),
    .X(_04128_));
 sg13g2_nor2_1 _24151_ (.A(net95),
    .B(net45),
    .Y(_04129_));
 sg13g2_a21oi_1 _24152_ (.A1(_04123_),
    .A2(_04129_),
    .Y(_04130_),
    .B1(_04079_));
 sg13g2_nor2_1 _24153_ (.A(_03919_),
    .B(_03921_),
    .Y(_04131_));
 sg13g2_buf_2 _24154_ (.A(_04131_),
    .X(_04132_));
 sg13g2_nand2_1 _24155_ (.Y(_04133_),
    .A(net102),
    .B(_04132_));
 sg13g2_nand2_1 _24156_ (.Y(_04134_),
    .A(_04129_),
    .B(_04079_));
 sg13g2_o21ai_1 _24157_ (.B1(_04134_),
    .Y(_04135_),
    .A1(_04130_),
    .A2(_04133_));
 sg13g2_buf_1 _24158_ (.A(_04135_),
    .X(_04136_));
 sg13g2_inv_1 _24159_ (.Y(_04137_),
    .A(_04136_));
 sg13g2_buf_1 _24160_ (.A(_03756_),
    .X(_04138_));
 sg13g2_buf_1 _24161_ (.A(_02800_),
    .X(_04139_));
 sg13g2_nor2_1 _24162_ (.A(net85),
    .B(net51),
    .Y(_04140_));
 sg13g2_nand2_1 _24163_ (.Y(_04141_),
    .A(net86),
    .B(_04140_));
 sg13g2_nand3b_1 _24164_ (.B(net80),
    .C(net85),
    .Y(_04142_),
    .A_N(net48));
 sg13g2_a21oi_1 _24165_ (.A1(_04141_),
    .A2(_04142_),
    .Y(_04143_),
    .B1(net87));
 sg13g2_o21ai_1 _24166_ (.B1(net86),
    .Y(_04144_),
    .A1(net85),
    .A2(net51));
 sg13g2_buf_1 _24167_ (.A(_02832_),
    .X(_04145_));
 sg13g2_a21oi_1 _24168_ (.A1(_04120_),
    .A2(_04144_),
    .Y(_04146_),
    .B1(net91));
 sg13g2_mux2_1 _24169_ (.A0(_04140_),
    .A1(_04146_),
    .S(_04060_),
    .X(_04147_));
 sg13g2_o21ai_1 _24170_ (.B1(net37),
    .Y(_04148_),
    .A1(_04143_),
    .A2(_04147_));
 sg13g2_buf_1 _24171_ (.A(_04148_),
    .X(_04149_));
 sg13g2_inv_1 _24172_ (.Y(_04150_),
    .A(_04149_));
 sg13g2_or2_1 _24173_ (.X(_04151_),
    .B(_04076_),
    .A(_04075_));
 sg13g2_buf_1 _24174_ (.A(_04151_),
    .X(_04152_));
 sg13g2_buf_1 _24175_ (.A(_04152_),
    .X(_04153_));
 sg13g2_nor3_2 _24176_ (.A(_03980_),
    .B(_03955_),
    .C(_03957_),
    .Y(_04154_));
 sg13g2_a21oi_1 _24177_ (.A1(_04020_),
    .A2(_04022_),
    .Y(_04155_),
    .B1(_04154_));
 sg13g2_mux2_1 _24178_ (.A0(net34),
    .A1(_04155_),
    .S(_04043_),
    .X(_04156_));
 sg13g2_nand3b_1 _24179_ (.B(_04029_),
    .C(_04031_),
    .Y(_04157_),
    .A_N(_03980_));
 sg13g2_buf_1 _24180_ (.A(_04157_),
    .X(_04158_));
 sg13g2_o21ai_1 _24181_ (.B1(_04158_),
    .Y(_04159_),
    .A1(_03070_),
    .A2(net42));
 sg13g2_mux2_1 _24182_ (.A0(net42),
    .A1(_04159_),
    .S(_04132_),
    .X(_04160_));
 sg13g2_a22oi_1 _24183_ (.Y(_04161_),
    .B1(_04160_),
    .B2(_04043_),
    .A2(_04156_),
    .A1(_03070_));
 sg13g2_nand2_1 _24184_ (.Y(_04162_),
    .A(net102),
    .B(_04053_));
 sg13g2_xor2_1 _24185_ (.B(_04162_),
    .A(_04161_),
    .X(_04163_));
 sg13g2_o21ai_1 _24186_ (.B1(_04163_),
    .Y(_04164_),
    .A1(_04136_),
    .A2(_04150_));
 sg13g2_o21ai_1 _24187_ (.B1(_04164_),
    .Y(_04165_),
    .A1(_04137_),
    .A2(_04149_));
 sg13g2_a21oi_1 _24188_ (.A1(_04090_),
    .A2(_04091_),
    .Y(_04166_),
    .B1(_04084_));
 sg13g2_xnor2_1 _24189_ (.Y(_04167_),
    .A(_04095_),
    .B(_04166_));
 sg13g2_nand2_1 _24190_ (.Y(_04168_),
    .A(_04165_),
    .B(_04167_));
 sg13g2_nand2_1 _24191_ (.Y(_04169_),
    .A(_02807_),
    .B(net254));
 sg13g2_buf_1 _24192_ (.A(_04169_),
    .X(_04170_));
 sg13g2_xor2_1 _24193_ (.B(_04098_),
    .A(_04073_),
    .X(_04171_));
 sg13g2_nor2_1 _24194_ (.A(_04122_),
    .B(_04168_),
    .Y(_04172_));
 sg13g2_a21oi_1 _24195_ (.A1(_04170_),
    .A2(_04171_),
    .Y(_04173_),
    .B1(_04172_));
 sg13g2_a21oi_1 _24196_ (.A1(_04122_),
    .A2(_04168_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_nor2_1 _24197_ (.A(_04104_),
    .B(_04174_),
    .Y(_04175_));
 sg13g2_nor2b_1 _24198_ (.A(_04119_),
    .B_N(_04174_),
    .Y(_04176_));
 sg13g2_a21oi_1 _24199_ (.A1(_04119_),
    .A2(_04175_),
    .Y(_04177_),
    .B1(_04176_));
 sg13g2_xnor2_1 _24200_ (.Y(_04178_),
    .A(_04122_),
    .B(_04168_));
 sg13g2_xnor2_1 _24201_ (.Y(_04179_),
    .A(_04171_),
    .B(_04178_));
 sg13g2_and2_1 _24202_ (.A(_04170_),
    .B(_04179_),
    .X(_04180_));
 sg13g2_buf_1 _24203_ (.A(_04180_),
    .X(_04181_));
 sg13g2_xnor2_1 _24204_ (.Y(_04182_),
    .A(_04136_),
    .B(_04149_));
 sg13g2_xnor2_1 _24205_ (.Y(_04183_),
    .A(_04163_),
    .B(_04182_));
 sg13g2_o21ai_1 _24206_ (.B1(_03996_),
    .Y(_04184_),
    .A1(_04060_),
    .A2(_04062_));
 sg13g2_nand2_1 _24207_ (.Y(_04185_),
    .A(net87),
    .B(_04060_));
 sg13g2_a21oi_1 _24208_ (.A1(_04184_),
    .A2(_04185_),
    .Y(_04186_),
    .B1(net36));
 sg13g2_nand2_1 _24209_ (.Y(_04187_),
    .A(net107),
    .B(_04053_));
 sg13g2_o21ai_1 _24210_ (.B1(net80),
    .Y(_04188_),
    .A1(net87),
    .A2(net51));
 sg13g2_a221oi_1 _24211_ (.B2(net107),
    .C1(net36),
    .B1(_04188_),
    .A1(net41),
    .Y(_04189_),
    .A2(net33));
 sg13g2_a21oi_1 _24212_ (.A1(net87),
    .A2(net80),
    .Y(_04190_),
    .B1(_04041_));
 sg13g2_nor3_1 _24213_ (.A(net91),
    .B(net86),
    .C(_04140_),
    .Y(_04191_));
 sg13g2_nor2_1 _24214_ (.A(net87),
    .B(net80),
    .Y(_04192_));
 sg13g2_nor3_1 _24215_ (.A(net48),
    .B(_04191_),
    .C(_04192_),
    .Y(_04193_));
 sg13g2_o21ai_1 _24216_ (.B1(_04193_),
    .Y(_04194_),
    .A1(_04189_),
    .A2(_04190_));
 sg13g2_o21ai_1 _24217_ (.B1(_04194_),
    .Y(_04195_),
    .A1(_04186_),
    .A2(_04187_));
 sg13g2_a21oi_1 _24218_ (.A1(_03972_),
    .A2(_03975_),
    .Y(_04196_),
    .B1(_03973_));
 sg13g2_buf_1 _24219_ (.A(_04196_),
    .X(_04197_));
 sg13g2_nand2b_1 _24220_ (.Y(_04198_),
    .B(_04126_),
    .A_N(net50));
 sg13g2_nand4_1 _24221_ (.B(_04024_),
    .C(_03972_),
    .A(_03974_),
    .Y(_04199_),
    .D(net52));
 sg13g2_a21oi_1 _24222_ (.A1(_04198_),
    .A2(_04199_),
    .Y(_04200_),
    .B1(_03071_));
 sg13g2_nand2_1 _24223_ (.Y(_04201_),
    .A(_03258_),
    .B(_04152_));
 sg13g2_xnor2_1 _24224_ (.Y(_04202_),
    .A(_04124_),
    .B(net52));
 sg13g2_buf_1 _24225_ (.A(_04202_),
    .X(_04203_));
 sg13g2_nor2_1 _24226_ (.A(net95),
    .B(net50),
    .Y(_04204_));
 sg13g2_a21oi_1 _24227_ (.A1(_02926_),
    .A2(_04203_),
    .Y(_04205_),
    .B1(_04204_));
 sg13g2_nor2_1 _24228_ (.A(_04201_),
    .B(_04205_),
    .Y(_04206_));
 sg13g2_nor2_1 _24229_ (.A(_04200_),
    .B(_04206_),
    .Y(_04207_));
 sg13g2_nand2_1 _24230_ (.Y(_04208_),
    .A(_04020_),
    .B(_04022_));
 sg13g2_buf_1 _24231_ (.A(_04208_),
    .X(_04209_));
 sg13g2_a21oi_1 _24232_ (.A1(net103),
    .A2(net40),
    .Y(_04210_),
    .B1(_04154_));
 sg13g2_xnor2_1 _24233_ (.Y(_04211_),
    .A(net39),
    .B(_04210_));
 sg13g2_mux2_1 _24234_ (.A0(_04079_),
    .A1(_04211_),
    .S(net102),
    .X(_04212_));
 sg13g2_xnor2_1 _24235_ (.Y(_04213_),
    .A(_04129_),
    .B(_04212_));
 sg13g2_nand2_1 _24236_ (.Y(_04214_),
    .A(_04207_),
    .B(_04213_));
 sg13g2_nor2_1 _24237_ (.A(_04207_),
    .B(_04213_),
    .Y(_04215_));
 sg13g2_a21oi_1 _24238_ (.A1(_04195_),
    .A2(_04214_),
    .Y(_04216_),
    .B1(_04215_));
 sg13g2_nor2_1 _24239_ (.A(_04183_),
    .B(_04216_),
    .Y(_04217_));
 sg13g2_nor2_2 _24240_ (.A(net254),
    .B(_03988_),
    .Y(_04218_));
 sg13g2_a21oi_1 _24241_ (.A1(_02457_),
    .A2(net91),
    .Y(_04219_),
    .B1(net86));
 sg13g2_nor3_1 _24242_ (.A(net91),
    .B(net85),
    .C(_04015_),
    .Y(_04220_));
 sg13g2_o21ai_1 _24243_ (.B1(net32),
    .Y(_04221_),
    .A1(_04219_),
    .A2(_04220_));
 sg13g2_a21oi_2 _24244_ (.B1(_02817_),
    .Y(_04222_),
    .A2(_04221_),
    .A1(_04218_));
 sg13g2_buf_1 _24245_ (.A(_02839_),
    .X(_04223_));
 sg13g2_a21oi_1 _24246_ (.A1(net140),
    .A2(_03986_),
    .Y(_04224_),
    .B1(_04104_));
 sg13g2_a21oi_1 _24247_ (.A1(net46),
    .A2(net33),
    .Y(_04225_),
    .B1(net86));
 sg13g2_a21oi_1 _24248_ (.A1(net107),
    .A2(net35),
    .Y(_04226_),
    .B1(_04225_));
 sg13g2_nor2_1 _24249_ (.A(net91),
    .B(_04013_),
    .Y(_04227_));
 sg13g2_nand2_1 _24250_ (.Y(_04228_),
    .A(net37),
    .B(_04227_));
 sg13g2_or3_1 _24251_ (.A(_04224_),
    .B(_04226_),
    .C(_04228_),
    .X(_04229_));
 sg13g2_buf_1 _24252_ (.A(_04229_),
    .X(_04230_));
 sg13g2_buf_1 _24253_ (.A(_02991_),
    .X(_04231_));
 sg13g2_nor2_1 _24254_ (.A(_02817_),
    .B(net139),
    .Y(_04232_));
 sg13g2_a21o_1 _24255_ (.A2(_04041_),
    .A1(net107),
    .B1(net80),
    .X(_04233_));
 sg13g2_nor2_1 _24256_ (.A(net91),
    .B(_04113_),
    .Y(_04234_));
 sg13g2_and4_1 _24257_ (.A(net147),
    .B(net80),
    .C(_04014_),
    .D(_04053_),
    .X(_04235_));
 sg13g2_a221oi_1 _24258_ (.B2(_04234_),
    .C1(_04235_),
    .B1(_04233_),
    .A1(_04232_),
    .Y(_04236_),
    .A2(_03995_));
 sg13g2_or2_1 _24259_ (.X(_04237_),
    .B(_04236_),
    .A(_04230_));
 sg13g2_inv_1 _24260_ (.Y(_04238_),
    .A(_04237_));
 sg13g2_a21o_1 _24261_ (.A2(_04222_),
    .A1(_04217_),
    .B1(_04238_),
    .X(_04239_));
 sg13g2_o21ai_1 _24262_ (.B1(_04239_),
    .Y(_04240_),
    .A1(_04217_),
    .A2(_04222_));
 sg13g2_buf_1 _24263_ (.A(_04240_),
    .X(_04241_));
 sg13g2_inv_1 _24264_ (.Y(_04242_),
    .A(_04241_));
 sg13g2_nand2_1 _24265_ (.Y(_04243_),
    .A(_04181_),
    .B(_04242_));
 sg13g2_nand2_1 _24266_ (.Y(_04244_),
    .A(_04170_),
    .B(_04167_));
 sg13g2_xor2_1 _24267_ (.B(_04244_),
    .A(_04165_),
    .X(_04245_));
 sg13g2_xnor2_1 _24268_ (.Y(_04246_),
    .A(_04237_),
    .B(_04222_));
 sg13g2_xnor2_1 _24269_ (.Y(_04247_),
    .A(_04217_),
    .B(_04246_));
 sg13g2_o21ai_1 _24270_ (.B1(net192),
    .Y(_04248_),
    .A1(_04245_),
    .A2(_04247_));
 sg13g2_buf_1 _24271_ (.A(_04248_),
    .X(_04249_));
 sg13g2_nand2_2 _24272_ (.Y(_04250_),
    .A(_04170_),
    .B(_04179_));
 sg13g2_nand2_1 _24273_ (.Y(_04251_),
    .A(_04250_),
    .B(_04241_));
 sg13g2_nand2_1 _24274_ (.Y(_04252_),
    .A(_04249_),
    .B(_04251_));
 sg13g2_nand2_1 _24275_ (.Y(_04253_),
    .A(_04122_),
    .B(_04168_));
 sg13g2_o21ai_1 _24276_ (.B1(_04253_),
    .Y(_04254_),
    .A1(_04171_),
    .A2(_04172_));
 sg13g2_and2_1 _24277_ (.A(_04170_),
    .B(_04254_),
    .X(_04255_));
 sg13g2_nor2_1 _24278_ (.A(net254),
    .B(_04099_),
    .Y(_04256_));
 sg13g2_xor2_1 _24279_ (.B(_04256_),
    .A(_04109_),
    .X(_04257_));
 sg13g2_nand2_1 _24280_ (.Y(_04258_),
    .A(_04255_),
    .B(_04257_));
 sg13g2_buf_1 _24281_ (.A(_04258_),
    .X(_04259_));
 sg13g2_a21oi_1 _24282_ (.A1(_04243_),
    .A2(_04252_),
    .Y(_04260_),
    .B1(net28));
 sg13g2_xnor2_1 _24283_ (.Y(_04261_),
    .A(_04177_),
    .B(_04260_));
 sg13g2_inv_1 _24284_ (.Y(_04262_),
    .A(_04261_));
 sg13g2_xnor2_1 _24285_ (.Y(_04263_),
    .A(_04230_),
    .B(_04236_));
 sg13g2_nand2b_1 _24286_ (.Y(_04264_),
    .B(_04263_),
    .A_N(_03999_));
 sg13g2_and2_1 _24287_ (.A(net95),
    .B(net50),
    .X(_04265_));
 sg13g2_buf_1 _24288_ (.A(_04265_),
    .X(_04266_));
 sg13g2_nor2_1 _24289_ (.A(_03422_),
    .B(net45),
    .Y(_04267_));
 sg13g2_o21ai_1 _24290_ (.B1(_03083_),
    .Y(_04268_),
    .A1(_03834_),
    .A2(_03968_));
 sg13g2_nor2_1 _24291_ (.A(_03552_),
    .B(_03904_),
    .Y(_04269_));
 sg13g2_mux2_1 _24292_ (.A0(_03680_),
    .A1(_04269_),
    .S(_03834_),
    .X(_04270_));
 sg13g2_nand2_1 _24293_ (.Y(_04271_),
    .A(_03963_),
    .B(_04270_));
 sg13g2_nand3_1 _24294_ (.B(_04268_),
    .C(_04271_),
    .A(_04024_),
    .Y(_04272_));
 sg13g2_nand3b_1 _24295_ (.B(_03963_),
    .C(_03960_),
    .Y(_04273_),
    .A_N(_03904_));
 sg13g2_buf_1 _24296_ (.A(_04273_),
    .X(_04274_));
 sg13g2_xnor2_1 _24297_ (.Y(_04275_),
    .A(_03834_),
    .B(_04274_));
 sg13g2_o21ai_1 _24298_ (.B1(net96),
    .Y(_04276_),
    .A1(_02926_),
    .A2(_04275_));
 sg13g2_nor2_1 _24299_ (.A(_04024_),
    .B(_04271_),
    .Y(_04277_));
 sg13g2_nor2_1 _24300_ (.A(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sg13g2_nand2_1 _24301_ (.Y(_04279_),
    .A(_04272_),
    .B(_04278_));
 sg13g2_buf_1 _24302_ (.A(net50),
    .X(_04280_));
 sg13g2_buf_1 _24303_ (.A(_04275_),
    .X(_04281_));
 sg13g2_nor2_1 _24304_ (.A(net47),
    .B(net54),
    .Y(_04282_));
 sg13g2_a22oi_1 _24305_ (.Y(_04283_),
    .B1(_04282_),
    .B2(_03493_),
    .A2(_04279_),
    .A1(_04267_));
 sg13g2_nor2_1 _24306_ (.A(_04266_),
    .B(_04283_),
    .Y(_04284_));
 sg13g2_nor2_1 _24307_ (.A(_04200_),
    .B(_04205_),
    .Y(_04285_));
 sg13g2_xnor2_1 _24308_ (.Y(_04286_),
    .A(_04201_),
    .B(_04285_));
 sg13g2_nor2_1 _24309_ (.A(_04284_),
    .B(_04286_),
    .Y(_04287_));
 sg13g2_a21o_1 _24310_ (.A2(net35),
    .A1(net107),
    .B1(_04225_),
    .X(_04288_));
 sg13g2_o21ai_1 _24311_ (.B1(net37),
    .Y(_04289_),
    .A1(_04225_),
    .A2(_04227_));
 sg13g2_nand2_1 _24312_ (.Y(_04290_),
    .A(net107),
    .B(net35));
 sg13g2_a22oi_1 _24313_ (.Y(_04291_),
    .B1(_04289_),
    .B2(_04290_),
    .A2(_04227_),
    .A1(_04288_));
 sg13g2_a21o_1 _24314_ (.A2(_04286_),
    .A1(_04284_),
    .B1(_04291_),
    .X(_04292_));
 sg13g2_nor2b_1 _24315_ (.A(_04287_),
    .B_N(_04292_),
    .Y(_04293_));
 sg13g2_xnor2_1 _24316_ (.Y(_04294_),
    .A(_04207_),
    .B(_04213_));
 sg13g2_xnor2_1 _24317_ (.Y(_04295_),
    .A(_04195_),
    .B(_04294_));
 sg13g2_and3_1 _24318_ (.X(_04296_),
    .A(_04264_),
    .B(_04293_),
    .C(_04295_));
 sg13g2_a21oi_1 _24319_ (.A1(_04293_),
    .A2(_04295_),
    .Y(_04297_),
    .B1(_04264_));
 sg13g2_nand3_1 _24320_ (.B(_04132_),
    .C(net40),
    .A(net83),
    .Y(_04298_));
 sg13g2_nand2_1 _24321_ (.Y(_04299_),
    .A(_04029_),
    .B(_04031_));
 sg13g2_buf_2 _24322_ (.A(_04299_),
    .X(_04300_));
 sg13g2_nand2_1 _24323_ (.Y(_04301_),
    .A(net92),
    .B(_04300_));
 sg13g2_or4_1 _24324_ (.A(_02800_),
    .B(_03951_),
    .C(_03980_),
    .D(_04301_),
    .X(_04302_));
 sg13g2_a221oi_1 _24325_ (.B2(_04031_),
    .C1(_03756_),
    .B1(_04029_),
    .A1(_04020_),
    .Y(_04303_),
    .A2(_04022_));
 sg13g2_nor4_1 _24326_ (.A(_02832_),
    .B(_02800_),
    .C(_03951_),
    .D(_04300_),
    .Y(_04304_));
 sg13g2_o21ai_1 _24327_ (.B1(_03980_),
    .Y(_04305_),
    .A1(_04303_),
    .A2(_04304_));
 sg13g2_and3_1 _24328_ (.X(_04306_),
    .A(_04298_),
    .B(_04302_),
    .C(_04305_));
 sg13g2_buf_1 _24329_ (.A(_04306_),
    .X(_04307_));
 sg13g2_nor2_1 _24330_ (.A(net85),
    .B(_04077_),
    .Y(_04308_));
 sg13g2_a21oi_1 _24331_ (.A1(net92),
    .A2(_04087_),
    .Y(_04309_),
    .B1(_04308_));
 sg13g2_a21oi_1 _24332_ (.A1(net140),
    .A2(_03986_),
    .Y(_04310_),
    .B1(_03999_));
 sg13g2_nor3_1 _24333_ (.A(_04307_),
    .B(_04309_),
    .C(_04310_),
    .Y(_04311_));
 sg13g2_o21ai_1 _24334_ (.B1(_04224_),
    .Y(_04312_),
    .A1(_04226_),
    .A2(_04228_));
 sg13g2_nand3_1 _24335_ (.B(_04311_),
    .C(_04312_),
    .A(_04230_),
    .Y(_04313_));
 sg13g2_o21ai_1 _24336_ (.B1(_04313_),
    .Y(_04314_),
    .A1(_04296_),
    .A2(_04297_));
 sg13g2_xor2_1 _24337_ (.B(_04216_),
    .A(_04183_),
    .X(_04315_));
 sg13g2_xnor2_1 _24338_ (.Y(_04316_),
    .A(_04314_),
    .B(_04315_));
 sg13g2_nor2_1 _24339_ (.A(_02817_),
    .B(_04316_),
    .Y(_04317_));
 sg13g2_and3_1 _24340_ (.X(_04318_),
    .A(_04230_),
    .B(_04311_),
    .C(_04312_));
 sg13g2_a21oi_1 _24341_ (.A1(_04230_),
    .A2(_04312_),
    .Y(_04319_),
    .B1(_04311_));
 sg13g2_nor2_1 _24342_ (.A(_02896_),
    .B(_02900_),
    .Y(_04320_));
 sg13g2_buf_1 _24343_ (.A(_04320_),
    .X(_04321_));
 sg13g2_nand2_1 _24344_ (.Y(_04322_),
    .A(net138),
    .B(_03995_));
 sg13g2_o21ai_1 _24345_ (.B1(_04322_),
    .Y(_04323_),
    .A1(_04318_),
    .A2(_04319_));
 sg13g2_xor2_1 _24346_ (.B(_04286_),
    .A(_04284_),
    .X(_04324_));
 sg13g2_xnor2_1 _24347_ (.Y(_04325_),
    .A(_04291_),
    .B(_04324_));
 sg13g2_nor3_1 _24348_ (.A(_03919_),
    .B(_03921_),
    .C(_04154_),
    .Y(_04326_));
 sg13g2_a221oi_1 _24349_ (.B2(_02619_),
    .C1(net42),
    .B1(_04158_),
    .A1(_04020_),
    .Y(_04327_),
    .A2(_04022_));
 sg13g2_nand4_1 _24350_ (.B(_04020_),
    .C(_04022_),
    .A(_04139_),
    .Y(_04328_),
    .D(net40));
 sg13g2_o21ai_1 _24351_ (.B1(_04328_),
    .Y(_04329_),
    .A1(_04326_),
    .A2(_04327_));
 sg13g2_mux2_1 _24352_ (.A0(_04308_),
    .A1(_04329_),
    .S(net80),
    .X(_04330_));
 sg13g2_nand2_1 _24353_ (.Y(_04331_),
    .A(net92),
    .B(_04053_));
 sg13g2_xor2_1 _24354_ (.B(_04331_),
    .A(_04330_),
    .X(_04332_));
 sg13g2_nor2b_1 _24355_ (.A(_04266_),
    .B_N(_04279_),
    .Y(_04333_));
 sg13g2_xnor2_1 _24356_ (.Y(_04334_),
    .A(_04267_),
    .B(_04333_));
 sg13g2_nor2_1 _24357_ (.A(_03904_),
    .B(_03911_),
    .Y(_04335_));
 sg13g2_xnor2_1 _24358_ (.Y(_04336_),
    .A(_03960_),
    .B(_04335_));
 sg13g2_buf_1 _24359_ (.A(_04336_),
    .X(_04337_));
 sg13g2_nor2_2 _24360_ (.A(net95),
    .B(net62),
    .Y(_04338_));
 sg13g2_nor2_1 _24361_ (.A(_03422_),
    .B(net50),
    .Y(_04339_));
 sg13g2_xnor2_1 _24362_ (.Y(_04340_),
    .A(_03970_),
    .B(_04274_));
 sg13g2_buf_2 _24363_ (.A(_04340_),
    .X(_04341_));
 sg13g2_nor3_1 _24364_ (.A(_03960_),
    .B(_03901_),
    .C(_03903_),
    .Y(_04342_));
 sg13g2_xnor2_1 _24365_ (.Y(_04343_),
    .A(_03834_),
    .B(_04342_));
 sg13g2_a22oi_1 _24366_ (.Y(_04344_),
    .B1(_04343_),
    .B2(_04338_),
    .A2(_04339_),
    .A1(_04341_));
 sg13g2_inv_1 _24367_ (.Y(_04345_),
    .A(_04344_));
 sg13g2_a22oi_1 _24368_ (.Y(_04346_),
    .B1(_04345_),
    .B2(net93),
    .A2(_04339_),
    .A1(_04338_));
 sg13g2_and2_1 _24369_ (.A(_04334_),
    .B(_04346_),
    .X(_04347_));
 sg13g2_or2_1 _24370_ (.X(_04348_),
    .B(_04346_),
    .A(_04334_));
 sg13g2_o21ai_1 _24371_ (.B1(_04348_),
    .Y(_04349_),
    .A1(_04332_),
    .A2(_04347_));
 sg13g2_nand2b_1 _24372_ (.Y(_04350_),
    .B(_04349_),
    .A_N(_04325_));
 sg13g2_buf_1 _24373_ (.A(_04350_),
    .X(_04351_));
 sg13g2_a21o_1 _24374_ (.A2(_04323_),
    .A1(net192),
    .B1(_04351_),
    .X(_04352_));
 sg13g2_nand3_1 _24375_ (.B(_04351_),
    .C(_04323_),
    .A(net192),
    .Y(_04353_));
 sg13g2_nor2_1 _24376_ (.A(_03156_),
    .B(_03043_),
    .Y(_04354_));
 sg13g2_buf_1 _24377_ (.A(_04354_),
    .X(_04355_));
 sg13g2_nor2_1 _24378_ (.A(_03879_),
    .B(net137),
    .Y(_04356_));
 sg13g2_and2_1 _24379_ (.A(net38),
    .B(_04356_),
    .X(_04357_));
 sg13g2_buf_1 _24380_ (.A(_04357_),
    .X(_04358_));
 sg13g2_a21oi_2 _24381_ (.B1(_04231_),
    .Y(_04359_),
    .A2(_04038_),
    .A1(_03951_));
 sg13g2_and2_1 _24382_ (.A(_03573_),
    .B(_03992_),
    .X(_04360_));
 sg13g2_xor2_1 _24383_ (.B(_04360_),
    .A(_04359_),
    .X(_04361_));
 sg13g2_buf_1 _24384_ (.A(_03573_),
    .X(_04362_));
 sg13g2_and4_1 _24385_ (.A(net161),
    .B(_04223_),
    .C(_03992_),
    .D(_04053_),
    .X(_04363_));
 sg13g2_a21o_1 _24386_ (.A2(_04361_),
    .A1(_04358_),
    .B1(_04363_),
    .X(_04364_));
 sg13g2_nand2_1 _24387_ (.Y(_04365_),
    .A(net183),
    .B(_03151_));
 sg13g2_buf_2 _24388_ (.A(_04365_),
    .X(_04366_));
 sg13g2_nand3_1 _24389_ (.B(_03998_),
    .C(_04366_),
    .A(net192),
    .Y(_04367_));
 sg13g2_nand3_1 _24390_ (.B(_04014_),
    .C(_04232_),
    .A(net38),
    .Y(_04368_));
 sg13g2_o21ai_1 _24391_ (.B1(_04368_),
    .Y(_04369_),
    .A1(_03993_),
    .A2(_04367_));
 sg13g2_nand2_1 _24392_ (.Y(_04370_),
    .A(net83),
    .B(_04158_));
 sg13g2_nand2_1 _24393_ (.Y(_04371_),
    .A(_02619_),
    .B(net44));
 sg13g2_nor2_1 _24394_ (.A(_04370_),
    .B(_04371_),
    .Y(_04372_));
 sg13g2_nand3_1 _24395_ (.B(_04020_),
    .C(_04022_),
    .A(_04092_),
    .Y(_04373_));
 sg13g2_a21oi_1 _24396_ (.A1(_04370_),
    .A2(_04371_),
    .Y(_04374_),
    .B1(_04373_));
 sg13g2_o21ai_1 _24397_ (.B1(_03982_),
    .Y(_04375_),
    .A1(_04372_),
    .A2(_04374_));
 sg13g2_buf_1 _24398_ (.A(_04375_),
    .X(_04376_));
 sg13g2_nand2b_1 _24399_ (.Y(_04377_),
    .B(_04376_),
    .A_N(_04369_));
 sg13g2_nor2b_1 _24400_ (.A(_04376_),
    .B_N(_04369_),
    .Y(_04378_));
 sg13g2_a21o_1 _24401_ (.A2(_04377_),
    .A1(_04364_),
    .B1(_04378_),
    .X(_04379_));
 sg13g2_buf_1 _24402_ (.A(_03052_),
    .X(_04380_));
 sg13g2_a22oi_1 _24403_ (.Y(_04381_),
    .B1(_03995_),
    .B2(net100),
    .A2(_03986_),
    .A1(net138));
 sg13g2_buf_1 _24404_ (.A(_04381_),
    .X(_04382_));
 sg13g2_a21oi_1 _24405_ (.A1(net140),
    .A2(_03986_),
    .Y(_04383_),
    .B1(_03988_));
 sg13g2_o21ai_1 _24406_ (.B1(_04383_),
    .Y(_04384_),
    .A1(_04307_),
    .A2(_04309_));
 sg13g2_or3_1 _24407_ (.A(_04307_),
    .B(_04309_),
    .C(_04383_),
    .X(_04385_));
 sg13g2_a21oi_1 _24408_ (.A1(_04384_),
    .A2(_04385_),
    .Y(_04386_),
    .B1(_02817_));
 sg13g2_nand2_1 _24409_ (.Y(_04387_),
    .A(_04382_),
    .B(_04386_));
 sg13g2_nor2_1 _24410_ (.A(_04382_),
    .B(_04386_),
    .Y(_04388_));
 sg13g2_a21oi_1 _24411_ (.A1(_04379_),
    .A2(_04387_),
    .Y(_04389_),
    .B1(_04388_));
 sg13g2_a21o_1 _24412_ (.A2(_04353_),
    .A1(_04352_),
    .B1(_04389_),
    .X(_04390_));
 sg13g2_buf_1 _24413_ (.A(_04390_),
    .X(_04391_));
 sg13g2_nand3_1 _24414_ (.B(_04352_),
    .C(_04353_),
    .A(_04389_),
    .Y(_04392_));
 sg13g2_buf_1 _24415_ (.A(_04392_),
    .X(_04393_));
 sg13g2_nand2_1 _24416_ (.Y(_04394_),
    .A(_04391_),
    .B(_04393_));
 sg13g2_xnor2_1 _24417_ (.Y(_04395_),
    .A(_04293_),
    .B(_04295_));
 sg13g2_o21ai_1 _24418_ (.B1(_04170_),
    .Y(_04396_),
    .A1(_04394_),
    .A2(_04395_));
 sg13g2_buf_1 _24419_ (.A(_04396_),
    .X(_04397_));
 sg13g2_nand2_1 _24420_ (.Y(_04398_),
    .A(_02740_),
    .B(_04323_));
 sg13g2_o21ai_1 _24421_ (.B1(_04389_),
    .Y(_04399_),
    .A1(_04351_),
    .A2(_04398_));
 sg13g2_inv_1 _24422_ (.Y(_04400_),
    .A(_04399_));
 sg13g2_a21oi_1 _24423_ (.A1(_04351_),
    .A2(_04398_),
    .Y(_04401_),
    .B1(_04400_));
 sg13g2_xor2_1 _24424_ (.B(_04401_),
    .A(_04397_),
    .X(_04402_));
 sg13g2_xnor2_1 _24425_ (.Y(_04403_),
    .A(_04317_),
    .B(_04402_));
 sg13g2_nor2_2 _24426_ (.A(_02817_),
    .B(_04296_),
    .Y(_04404_));
 sg13g2_xnor2_1 _24427_ (.Y(_04405_),
    .A(_04245_),
    .B(_04247_));
 sg13g2_nand3_1 _24428_ (.B(_04314_),
    .C(_04315_),
    .A(_02740_),
    .Y(_04406_));
 sg13g2_buf_1 _24429_ (.A(_04406_),
    .X(_04407_));
 sg13g2_xnor2_1 _24430_ (.Y(_04408_),
    .A(_04405_),
    .B(_04407_));
 sg13g2_xnor2_1 _24431_ (.Y(_04409_),
    .A(_04404_),
    .B(_04408_));
 sg13g2_buf_1 _24432_ (.A(_04409_),
    .X(_04410_));
 sg13g2_or2_1 _24433_ (.X(_04411_),
    .B(_04401_),
    .A(_04317_));
 sg13g2_buf_1 _24434_ (.A(_04411_),
    .X(_04412_));
 sg13g2_and2_1 _24435_ (.A(_04317_),
    .B(_04401_),
    .X(_04413_));
 sg13g2_buf_1 _24436_ (.A(_04413_),
    .X(_04414_));
 sg13g2_a21oi_1 _24437_ (.A1(_04397_),
    .A2(_04412_),
    .Y(_04415_),
    .B1(_04414_));
 sg13g2_xnor2_1 _24438_ (.Y(_04416_),
    .A(_04410_),
    .B(_04415_));
 sg13g2_nor2_1 _24439_ (.A(_04403_),
    .B(_04416_),
    .Y(_04417_));
 sg13g2_nand2_1 _24440_ (.Y(_04418_),
    .A(net140),
    .B(_04081_));
 sg13g2_buf_1 _24441_ (.A(net180),
    .X(_04419_));
 sg13g2_nor2_1 _24442_ (.A(net160),
    .B(net48),
    .Y(_04420_));
 sg13g2_buf_2 _24443_ (.A(_04420_),
    .X(_04421_));
 sg13g2_nand2_1 _24444_ (.Y(_04422_),
    .A(_04004_),
    .B(_04421_));
 sg13g2_nand2_1 _24445_ (.Y(_04423_),
    .A(_03951_),
    .B(_04366_));
 sg13g2_a21oi_1 _24446_ (.A1(_04086_),
    .A2(_04423_),
    .Y(_04424_),
    .B1(_03880_));
 sg13g2_nand2_1 _24447_ (.Y(_04425_),
    .A(net179),
    .B(_02839_));
 sg13g2_a21oi_1 _24448_ (.A1(_04020_),
    .A2(_04022_),
    .Y(_04426_),
    .B1(net42));
 sg13g2_o21ai_1 _24449_ (.B1(net137),
    .Y(_04427_),
    .A1(_04425_),
    .A2(_04426_));
 sg13g2_nand2_1 _24450_ (.Y(_04428_),
    .A(_04424_),
    .B(_04427_));
 sg13g2_a221oi_1 _24451_ (.B2(_04422_),
    .C1(_04428_),
    .B1(_04418_),
    .A1(_04358_),
    .Y(_04429_),
    .A2(_04361_));
 sg13g2_nand2_1 _24452_ (.Y(_04430_),
    .A(net38),
    .B(_04356_));
 sg13g2_a221oi_1 _24453_ (.B2(_04004_),
    .C1(_04430_),
    .B1(_04421_),
    .A1(net140),
    .Y(_04431_),
    .A2(_04081_));
 sg13g2_nor2_1 _24454_ (.A(_03955_),
    .B(_03957_),
    .Y(_04432_));
 sg13g2_buf_1 _24455_ (.A(_04432_),
    .X(_04433_));
 sg13g2_nor2_1 _24456_ (.A(_02832_),
    .B(_04433_),
    .Y(_04434_));
 sg13g2_nand2b_1 _24457_ (.Y(_04435_),
    .B(_02618_),
    .A_N(net50));
 sg13g2_buf_1 _24458_ (.A(_04435_),
    .X(_04436_));
 sg13g2_o21ai_1 _24459_ (.B1(_04436_),
    .Y(_04437_),
    .A1(_03756_),
    .A2(_04127_));
 sg13g2_nor2_1 _24460_ (.A(_04120_),
    .B(_04198_),
    .Y(_04438_));
 sg13g2_a21oi_1 _24461_ (.A1(_04434_),
    .A2(_04437_),
    .Y(_04439_),
    .B1(_04438_));
 sg13g2_a21oi_1 _24462_ (.A1(_04361_),
    .A2(_04431_),
    .Y(_04440_),
    .B1(_04439_));
 sg13g2_and2_1 _24463_ (.A(_04003_),
    .B(_04360_),
    .X(_04441_));
 sg13g2_mux2_1 _24464_ (.A0(net160),
    .A1(_04441_),
    .S(_04359_),
    .X(_04442_));
 sg13g2_or2_1 _24465_ (.X(_04443_),
    .B(_03992_),
    .A(net36));
 sg13g2_nand2_1 _24466_ (.Y(_04444_),
    .A(net160),
    .B(_04047_));
 sg13g2_o21ai_1 _24467_ (.B1(_04444_),
    .Y(_04445_),
    .A1(_04443_),
    .A2(_04359_));
 sg13g2_a221oi_1 _24468_ (.B2(_04434_),
    .C1(_04438_),
    .B1(_04437_),
    .A1(net38),
    .Y(_04446_),
    .A2(_04356_));
 sg13g2_nand3b_1 _24469_ (.B(_04424_),
    .C(_04427_),
    .Y(_04447_),
    .A_N(_04446_));
 sg13g2_o21ai_1 _24470_ (.B1(_04447_),
    .Y(_04448_),
    .A1(_04442_),
    .A2(_04445_));
 sg13g2_o21ai_1 _24471_ (.B1(_04448_),
    .Y(_04449_),
    .A1(_04429_),
    .A2(_04440_));
 sg13g2_buf_1 _24472_ (.A(_04449_),
    .X(_04450_));
 sg13g2_or2_1 _24473_ (.X(_04451_),
    .B(_03051_),
    .A(net190));
 sg13g2_buf_1 _24474_ (.A(_04451_),
    .X(_04452_));
 sg13g2_xnor2_1 _24475_ (.Y(_04453_),
    .A(_04320_),
    .B(_04452_));
 sg13g2_nand2_2 _24476_ (.Y(_04454_),
    .A(_03986_),
    .B(_04453_));
 sg13g2_xnor2_1 _24477_ (.Y(_04455_),
    .A(_04369_),
    .B(_04376_));
 sg13g2_xnor2_1 _24478_ (.Y(_04456_),
    .A(_04364_),
    .B(_04455_));
 sg13g2_xnor2_1 _24479_ (.Y(_04457_),
    .A(_04454_),
    .B(_04456_));
 sg13g2_xnor2_1 _24480_ (.Y(_04458_),
    .A(_04450_),
    .B(_04457_));
 sg13g2_buf_1 _24481_ (.A(_04458_),
    .X(_04459_));
 sg13g2_o21ai_1 _24482_ (.B1(_04223_),
    .Y(_04460_),
    .A1(_04075_),
    .A2(_04076_));
 sg13g2_buf_1 _24483_ (.A(_04460_),
    .X(_04461_));
 sg13g2_nor2_1 _24484_ (.A(_04013_),
    .B(net137),
    .Y(_04462_));
 sg13g2_nand2_1 _24485_ (.Y(_04463_),
    .A(net38),
    .B(_04462_));
 sg13g2_nor2_1 _24486_ (.A(_04461_),
    .B(_04463_),
    .Y(_04464_));
 sg13g2_nand2_1 _24487_ (.Y(_04465_),
    .A(_04461_),
    .B(_04463_));
 sg13g2_o21ai_1 _24488_ (.B1(_04465_),
    .Y(_04466_),
    .A1(_04421_),
    .A2(_04464_));
 sg13g2_inv_1 _24489_ (.Y(_04467_),
    .A(_04466_));
 sg13g2_nor2_1 _24490_ (.A(net86),
    .B(net50),
    .Y(_04468_));
 sg13g2_nor2_1 _24491_ (.A(net91),
    .B(_04128_),
    .Y(_04469_));
 sg13g2_mux2_1 _24492_ (.A0(_04341_),
    .A1(_04469_),
    .S(net85),
    .X(_04470_));
 sg13g2_nand2_1 _24493_ (.Y(_04471_),
    .A(_04468_),
    .B(_04470_));
 sg13g2_o21ai_1 _24494_ (.B1(_03756_),
    .Y(_04472_),
    .A1(_03834_),
    .A2(_03968_));
 sg13g2_nand3_1 _24495_ (.B(_04271_),
    .C(_04472_),
    .A(_04024_),
    .Y(_04473_));
 sg13g2_a21oi_1 _24496_ (.A1(_03756_),
    .A2(_04341_),
    .Y(_04474_),
    .B1(_04277_));
 sg13g2_a21oi_1 _24497_ (.A1(_04473_),
    .A2(_04474_),
    .Y(_04475_),
    .B1(net85));
 sg13g2_nand2_1 _24498_ (.Y(_04476_),
    .A(_04469_),
    .B(_04475_));
 sg13g2_nand2_1 _24499_ (.Y(_04477_),
    .A(_04471_),
    .B(_04476_));
 sg13g2_nor2_1 _24500_ (.A(net178),
    .B(net48),
    .Y(_04478_));
 sg13g2_nor2_1 _24501_ (.A(net139),
    .B(_04426_),
    .Y(_04479_));
 sg13g2_or2_1 _24502_ (.X(_04480_),
    .B(_04479_),
    .A(_04478_));
 sg13g2_a21o_1 _24503_ (.A2(_04478_),
    .A1(_04018_),
    .B1(_04039_),
    .X(_04481_));
 sg13g2_nand3_1 _24504_ (.B(_04080_),
    .C(_04478_),
    .A(net140),
    .Y(_04482_));
 sg13g2_nand3_1 _24505_ (.B(_04481_),
    .C(_04482_),
    .A(_04480_),
    .Y(_04483_));
 sg13g2_buf_1 _24506_ (.A(_04483_),
    .X(_04484_));
 sg13g2_nand2b_1 _24507_ (.Y(_04485_),
    .B(_04484_),
    .A_N(_04477_));
 sg13g2_nor2b_1 _24508_ (.A(_04484_),
    .B_N(_04477_),
    .Y(_04486_));
 sg13g2_a21oi_2 _24509_ (.B1(_04486_),
    .Y(_04487_),
    .A2(_04485_),
    .A1(_04467_));
 sg13g2_nor2_1 _24510_ (.A(_04442_),
    .B(_04445_),
    .Y(_04488_));
 sg13g2_inv_1 _24511_ (.Y(_04489_),
    .A(_04428_));
 sg13g2_o21ai_1 _24512_ (.B1(net160),
    .Y(_04490_),
    .A1(_04231_),
    .A2(_04068_));
 sg13g2_inv_1 _24513_ (.Y(_04491_),
    .A(_04439_));
 sg13g2_a21oi_1 _24514_ (.A1(_04358_),
    .A2(_04490_),
    .Y(_04492_),
    .B1(_04491_));
 sg13g2_nor2_1 _24515_ (.A(_03880_),
    .B(_04425_),
    .Y(_04493_));
 sg13g2_nand3_1 _24516_ (.B(net137),
    .C(_04493_),
    .A(_04080_),
    .Y(_04494_));
 sg13g2_and2_1 _24517_ (.A(_04491_),
    .B(_04494_),
    .X(_04495_));
 sg13g2_or2_1 _24518_ (.X(_04496_),
    .B(_04490_),
    .A(_04430_));
 sg13g2_a22oi_1 _24519_ (.Y(_04497_),
    .B1(_04495_),
    .B2(_04496_),
    .A2(_04492_),
    .A1(_04489_));
 sg13g2_xor2_1 _24520_ (.B(_04497_),
    .A(_04488_),
    .X(_04498_));
 sg13g2_nand2_1 _24521_ (.Y(_04499_),
    .A(_04487_),
    .B(_04498_));
 sg13g2_buf_1 _24522_ (.A(_02988_),
    .X(_04500_));
 sg13g2_nor2_1 _24523_ (.A(net118),
    .B(net51),
    .Y(_04501_));
 sg13g2_nand2_1 _24524_ (.Y(_04502_),
    .A(net100),
    .B(_04060_));
 sg13g2_mux2_1 _24525_ (.A0(net118),
    .A1(_04501_),
    .S(_04502_),
    .X(_04503_));
 sg13g2_nand2_1 _24526_ (.Y(_04504_),
    .A(net37),
    .B(_04503_));
 sg13g2_o21ai_1 _24527_ (.B1(_04504_),
    .Y(_04505_),
    .A1(_04487_),
    .A2(_04498_));
 sg13g2_nor2_1 _24528_ (.A(_04092_),
    .B(_04138_),
    .Y(_04506_));
 sg13g2_o21ai_1 _24529_ (.B1(_04158_),
    .Y(_04507_),
    .A1(net83),
    .A2(net42));
 sg13g2_a21oi_1 _24530_ (.A1(net40),
    .A2(_04370_),
    .Y(_04508_),
    .B1(_04132_));
 sg13g2_a21o_1 _24531_ (.A2(_04507_),
    .A1(_04132_),
    .B1(_04508_),
    .X(_04509_));
 sg13g2_a22oi_1 _24532_ (.Y(_04510_),
    .B1(_04509_),
    .B2(net87),
    .A2(_04506_),
    .A1(net34));
 sg13g2_nor2_1 _24533_ (.A(_04138_),
    .B(_04154_),
    .Y(_04511_));
 sg13g2_mux2_1 _24534_ (.A0(_04511_),
    .A1(_04507_),
    .S(_04132_),
    .X(_04512_));
 sg13g2_a22oi_1 _24535_ (.Y(_04513_),
    .B1(_04512_),
    .B2(_04093_),
    .A2(_04506_),
    .A1(_04152_));
 sg13g2_nor2_1 _24536_ (.A(_04371_),
    .B(_04513_),
    .Y(_04514_));
 sg13g2_a21oi_1 _24537_ (.A1(_04371_),
    .A2(_04510_),
    .Y(_04515_),
    .B1(_04514_));
 sg13g2_or2_1 _24538_ (.X(_04516_),
    .B(_04204_),
    .A(_04266_));
 sg13g2_nor2_1 _24539_ (.A(net101),
    .B(net62),
    .Y(_04517_));
 sg13g2_inv_2 _24540_ (.Y(_04518_),
    .A(net62));
 sg13g2_inv_1 _24541_ (.Y(_04519_),
    .A(_04266_));
 sg13g2_o21ai_1 _24542_ (.B1(_04519_),
    .Y(_04520_),
    .A1(_04518_),
    .A2(_04339_));
 sg13g2_nand2_1 _24543_ (.Y(_04521_),
    .A(net93),
    .B(_04341_));
 sg13g2_nor3_1 _24544_ (.A(net101),
    .B(net47),
    .C(_04518_),
    .Y(_04522_));
 sg13g2_a21oi_1 _24545_ (.A1(net101),
    .A2(_04338_),
    .Y(_04523_),
    .B1(_04522_));
 sg13g2_nor2_1 _24546_ (.A(_04521_),
    .B(_04523_),
    .Y(_04524_));
 sg13g2_a221oi_1 _24547_ (.B2(_04521_),
    .C1(_04524_),
    .B1(_04520_),
    .A1(_04516_),
    .Y(_04525_),
    .A2(_04517_));
 sg13g2_xnor2_1 _24548_ (.Y(_04526_),
    .A(_04515_),
    .B(_04525_));
 sg13g2_buf_1 _24549_ (.A(_04124_),
    .X(_04527_));
 sg13g2_nor2_2 _24550_ (.A(_02800_),
    .B(net50),
    .Y(_04528_));
 sg13g2_nand4_1 _24551_ (.B(net86),
    .C(_04433_),
    .A(net92),
    .Y(_04529_),
    .D(_04528_));
 sg13g2_o21ai_1 _24552_ (.B1(_04529_),
    .Y(_04530_),
    .A1(_04433_),
    .A2(_04528_));
 sg13g2_nor3_1 _24553_ (.A(net49),
    .B(_04300_),
    .C(_04436_),
    .Y(_04531_));
 sg13g2_a21oi_1 _24554_ (.A1(_04434_),
    .A2(_04436_),
    .Y(_04532_),
    .B1(_04531_));
 sg13g2_o21ai_1 _24555_ (.B1(_04145_),
    .Y(_04533_),
    .A1(net49),
    .A2(_04528_));
 sg13g2_nand2_1 _24556_ (.Y(_04534_),
    .A(_04532_),
    .B(_04533_));
 sg13g2_a22oi_1 _24557_ (.Y(_04535_),
    .B1(_04534_),
    .B2(_03996_),
    .A2(_04530_),
    .A1(net49));
 sg13g2_o21ai_1 _24558_ (.B1(_04126_),
    .Y(_04536_),
    .A1(net83),
    .A2(net49));
 sg13g2_a22oi_1 _24559_ (.Y(_04537_),
    .B1(_04528_),
    .B2(_04536_),
    .A2(net49),
    .A1(net83));
 sg13g2_nand3_1 _24560_ (.B(_04527_),
    .C(_04126_),
    .A(net92),
    .Y(_04538_));
 sg13g2_nand2b_1 _24561_ (.Y(_04539_),
    .B(net52),
    .A_N(net49));
 sg13g2_a22oi_1 _24562_ (.Y(_04540_),
    .B1(_04539_),
    .B2(net83),
    .A2(_04300_),
    .A1(net92));
 sg13g2_nand3_1 _24563_ (.B(_04538_),
    .C(_04540_),
    .A(_04436_),
    .Y(_04541_));
 sg13g2_o21ai_1 _24564_ (.B1(_04541_),
    .Y(_04542_),
    .A1(_04301_),
    .A2(_04537_));
 sg13g2_inv_1 _24565_ (.Y(_04543_),
    .A(_04542_));
 sg13g2_o21ai_1 _24566_ (.B1(_04543_),
    .Y(_04544_),
    .A1(net52),
    .A2(_04535_));
 sg13g2_buf_1 _24567_ (.A(_04544_),
    .X(_04545_));
 sg13g2_nor2_1 _24568_ (.A(net103),
    .B(net62),
    .Y(_04546_));
 sg13g2_buf_1 _24569_ (.A(_04341_),
    .X(_04547_));
 sg13g2_nand2_1 _24570_ (.Y(_04548_),
    .A(net102),
    .B(net53));
 sg13g2_xnor2_1 _24571_ (.Y(_04549_),
    .A(_04546_),
    .B(_04548_));
 sg13g2_nand2b_1 _24572_ (.Y(_04550_),
    .B(_04549_),
    .A_N(_04545_));
 sg13g2_nor2_1 _24573_ (.A(_04526_),
    .B(_04550_),
    .Y(_04551_));
 sg13g2_a21oi_1 _24574_ (.A1(_04499_),
    .A2(_04505_),
    .Y(_04552_),
    .B1(_04551_));
 sg13g2_buf_1 _24575_ (.A(_04552_),
    .X(_04553_));
 sg13g2_nor2_1 _24576_ (.A(net30),
    .B(net29),
    .Y(_04554_));
 sg13g2_inv_1 _24577_ (.Y(_04555_),
    .A(_04338_));
 sg13g2_a22oi_1 _24578_ (.Y(_04556_),
    .B1(_04555_),
    .B2(net47),
    .A2(_04337_),
    .A1(_04045_));
 sg13g2_inv_1 _24579_ (.Y(_04557_),
    .A(_04556_));
 sg13g2_a221oi_1 _24580_ (.B2(_04557_),
    .C1(_04524_),
    .B1(_04521_),
    .A1(_04338_),
    .Y(_04558_),
    .A2(_04339_));
 sg13g2_nor4_1 _24581_ (.A(net103),
    .B(_04045_),
    .C(net54),
    .D(net62),
    .Y(_04559_));
 sg13g2_a22oi_1 _24582_ (.Y(_04560_),
    .B1(_04516_),
    .B2(_04559_),
    .A2(_04558_),
    .A1(_04515_));
 sg13g2_xnor2_1 _24583_ (.Y(_04561_),
    .A(_04334_),
    .B(_04346_));
 sg13g2_xnor2_1 _24584_ (.Y(_04562_),
    .A(_04332_),
    .B(_04561_));
 sg13g2_xor2_1 _24585_ (.B(_04562_),
    .A(_04560_),
    .X(_04563_));
 sg13g2_inv_1 _24586_ (.Y(_04564_),
    .A(_04563_));
 sg13g2_a21oi_1 _24587_ (.A1(net30),
    .A2(_04553_),
    .Y(_04565_),
    .B1(_04564_));
 sg13g2_nand2_1 _24588_ (.Y(_04566_),
    .A(_02807_),
    .B(_02743_));
 sg13g2_xor2_1 _24589_ (.B(_04325_),
    .A(_04349_),
    .X(_04567_));
 sg13g2_a21oi_2 _24590_ (.B1(_04104_),
    .Y(_04568_),
    .A2(_04567_),
    .A1(_04566_));
 sg13g2_o21ai_1 _24591_ (.B1(_04456_),
    .Y(_04569_),
    .A1(_04450_),
    .A2(_04454_));
 sg13g2_nand2_1 _24592_ (.Y(_04570_),
    .A(_04450_),
    .B(_04454_));
 sg13g2_nand2_1 _24593_ (.Y(_04571_),
    .A(_04569_),
    .B(_04570_));
 sg13g2_xor2_1 _24594_ (.B(_04571_),
    .A(_04568_),
    .X(_04572_));
 sg13g2_xnor2_1 _24595_ (.Y(_04573_),
    .A(_04379_),
    .B(_04386_));
 sg13g2_xor2_1 _24596_ (.B(_04573_),
    .A(_04382_),
    .X(_04574_));
 sg13g2_nor2_2 _24597_ (.A(_04560_),
    .B(_04562_),
    .Y(_04575_));
 sg13g2_xnor2_1 _24598_ (.Y(_04576_),
    .A(_04574_),
    .B(_04575_));
 sg13g2_xnor2_1 _24599_ (.Y(_04577_),
    .A(_04572_),
    .B(_04576_));
 sg13g2_buf_2 _24600_ (.A(_04577_),
    .X(_04578_));
 sg13g2_o21ai_1 _24601_ (.B1(_04578_),
    .Y(_04579_),
    .A1(_04554_),
    .A2(_04565_));
 sg13g2_nor2_1 _24602_ (.A(_04487_),
    .B(_04498_),
    .Y(_04580_));
 sg13g2_a21oi_1 _24603_ (.A1(_04487_),
    .A2(_04498_),
    .Y(_04581_),
    .B1(_04504_));
 sg13g2_o21ai_1 _24604_ (.B1(_04551_),
    .Y(_04582_),
    .A1(_04580_),
    .A2(_04581_));
 sg13g2_buf_1 _24605_ (.A(_04582_),
    .X(_04583_));
 sg13g2_nor2_1 _24606_ (.A(net29),
    .B(_04583_),
    .Y(_04584_));
 sg13g2_nand2b_1 _24607_ (.Y(_04585_),
    .B(_04563_),
    .A_N(net30));
 sg13g2_nor2_1 _24608_ (.A(_04583_),
    .B(_04585_),
    .Y(_04586_));
 sg13g2_a21oi_1 _24609_ (.A1(_04578_),
    .A2(_04584_),
    .Y(_04587_),
    .B1(_04586_));
 sg13g2_nor2_2 _24610_ (.A(_02988_),
    .B(_04452_),
    .Y(_04588_));
 sg13g2_and2_1 _24611_ (.A(_03987_),
    .B(_04588_),
    .X(_04589_));
 sg13g2_buf_1 _24612_ (.A(_04589_),
    .X(_04590_));
 sg13g2_a21oi_1 _24613_ (.A1(_04579_),
    .A2(_04587_),
    .Y(_04591_),
    .B1(net31));
 sg13g2_nand2_1 _24614_ (.Y(_04592_),
    .A(net30),
    .B(_04583_));
 sg13g2_nand2b_1 _24615_ (.Y(_04593_),
    .B(_04592_),
    .A_N(net29));
 sg13g2_a21oi_1 _24616_ (.A1(net31),
    .A2(_04593_),
    .Y(_04594_),
    .B1(_04586_));
 sg13g2_nor2b_1 _24617_ (.A(_04594_),
    .B_N(_04578_),
    .Y(_04595_));
 sg13g2_mux2_1 _24618_ (.A0(_04592_),
    .A1(net30),
    .S(net29),
    .X(_04596_));
 sg13g2_nand2_1 _24619_ (.Y(_04597_),
    .A(net31),
    .B(_04563_));
 sg13g2_inv_1 _24620_ (.Y(_04598_),
    .A(_04583_));
 sg13g2_o21ai_1 _24621_ (.B1(net31),
    .Y(_04599_),
    .A1(_04598_),
    .A2(_04554_));
 sg13g2_buf_1 _24622_ (.A(_04599_),
    .X(_04600_));
 sg13g2_o21ai_1 _24623_ (.B1(_04600_),
    .Y(_04601_),
    .A1(_04596_),
    .A2(_04597_));
 sg13g2_or2_1 _24624_ (.X(_04602_),
    .B(_04601_),
    .A(_04595_));
 sg13g2_and2_1 _24625_ (.A(net30),
    .B(_04583_),
    .X(_04603_));
 sg13g2_o21ai_1 _24626_ (.B1(_04578_),
    .Y(_04604_),
    .A1(net29),
    .A2(_04603_));
 sg13g2_nand2_1 _24627_ (.Y(_04605_),
    .A(_04586_),
    .B(_04578_));
 sg13g2_inv_1 _24628_ (.Y(_04606_),
    .A(_04585_));
 sg13g2_nor2_1 _24629_ (.A(_04564_),
    .B(net29),
    .Y(_04607_));
 sg13g2_a22oi_1 _24630_ (.Y(_04608_),
    .B1(_04603_),
    .B2(_04607_),
    .A2(_04606_),
    .A1(net29));
 sg13g2_and3_1 _24631_ (.X(_04609_),
    .A(_04604_),
    .B(_04605_),
    .C(_04608_));
 sg13g2_buf_1 _24632_ (.A(_04609_),
    .X(_04610_));
 sg13g2_nor2_1 _24633_ (.A(_04104_),
    .B(_04395_),
    .Y(_04611_));
 sg13g2_nand3_1 _24634_ (.B(_04393_),
    .C(_04611_),
    .A(_04391_),
    .Y(_04612_));
 sg13g2_a21o_1 _24635_ (.A2(_04393_),
    .A1(_04391_),
    .B1(_04611_),
    .X(_04613_));
 sg13g2_buf_1 _24636_ (.A(_04613_),
    .X(_04614_));
 sg13g2_and2_1 _24637_ (.A(_04612_),
    .B(_04614_),
    .X(_04615_));
 sg13g2_inv_1 _24638_ (.Y(_04616_),
    .A(_04575_));
 sg13g2_o21ai_1 _24639_ (.B1(_04450_),
    .Y(_04617_),
    .A1(_04454_),
    .A2(_04456_));
 sg13g2_nand2_1 _24640_ (.Y(_04618_),
    .A(_04454_),
    .B(_04456_));
 sg13g2_nand2_1 _24641_ (.Y(_04619_),
    .A(_04617_),
    .B(_04618_));
 sg13g2_nor2_1 _24642_ (.A(_04574_),
    .B(_04619_),
    .Y(_04620_));
 sg13g2_nand2_1 _24643_ (.Y(_04621_),
    .A(_04574_),
    .B(_04619_));
 sg13g2_o21ai_1 _24644_ (.B1(_04621_),
    .Y(_04622_),
    .A1(_04620_),
    .A2(_04568_));
 sg13g2_inv_1 _24645_ (.Y(_04623_),
    .A(_04568_));
 sg13g2_a21oi_1 _24646_ (.A1(_04620_),
    .A2(_04575_),
    .Y(_04624_),
    .B1(_04623_));
 sg13g2_a21oi_1 _24647_ (.A1(_04623_),
    .A2(_04621_),
    .Y(_04625_),
    .B1(_04624_));
 sg13g2_a21oi_1 _24648_ (.A1(_04616_),
    .A2(_04622_),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_xnor2_1 _24649_ (.Y(_04627_),
    .A(_04615_),
    .B(_04626_));
 sg13g2_buf_2 _24650_ (.A(_04627_),
    .X(_04628_));
 sg13g2_o21ai_1 _24651_ (.B1(_04628_),
    .Y(_04629_),
    .A1(_04600_),
    .A2(_04610_));
 sg13g2_o21ai_1 _24652_ (.B1(_04629_),
    .Y(_04630_),
    .A1(_04591_),
    .A2(_04602_));
 sg13g2_buf_1 _24653_ (.A(_04630_),
    .X(_04631_));
 sg13g2_nor2_1 _24654_ (.A(_04631_),
    .B(_04416_),
    .Y(_04632_));
 sg13g2_nand3_1 _24655_ (.B(net34),
    .C(_04588_),
    .A(net44),
    .Y(_04633_));
 sg13g2_buf_1 _24656_ (.A(_04633_),
    .X(_04634_));
 sg13g2_nand2_1 _24657_ (.Y(_04635_),
    .A(_04527_),
    .B(_04126_));
 sg13g2_nand2_1 _24658_ (.Y(_04636_),
    .A(_04433_),
    .B(_04366_));
 sg13g2_nor2_2 _24659_ (.A(net139),
    .B(_04275_),
    .Y(_04637_));
 sg13g2_nand2_1 _24660_ (.Y(_04638_),
    .A(_04300_),
    .B(_04637_));
 sg13g2_mux2_1 _24661_ (.A0(_04636_),
    .A1(_04638_),
    .S(net39),
    .X(_04639_));
 sg13g2_nor2_1 _24662_ (.A(_04635_),
    .B(_04639_),
    .Y(_04640_));
 sg13g2_nor2_1 _24663_ (.A(_04366_),
    .B(_04637_),
    .Y(_04641_));
 sg13g2_o21ai_1 _24664_ (.B1(net40),
    .Y(_04642_),
    .A1(_04300_),
    .A2(_04637_));
 sg13g2_nor3_1 _24665_ (.A(net39),
    .B(_04641_),
    .C(_04642_),
    .Y(_04643_));
 sg13g2_o21ai_1 _24666_ (.B1(_04362_),
    .Y(_04644_),
    .A1(_04640_),
    .A2(_04643_));
 sg13g2_nand3_1 _24667_ (.B(_04366_),
    .C(_04637_),
    .A(net34),
    .Y(_04645_));
 sg13g2_and2_1 _24668_ (.A(_04644_),
    .B(_04645_),
    .X(_04646_));
 sg13g2_nor2_2 _24669_ (.A(net139),
    .B(_04197_),
    .Y(_04647_));
 sg13g2_or2_1 _24670_ (.X(_04648_),
    .B(_04197_),
    .A(_02991_));
 sg13g2_buf_2 _24671_ (.A(_04648_),
    .X(_04649_));
 sg13g2_nand3_1 _24672_ (.B(net35),
    .C(_04649_),
    .A(net216),
    .Y(_04650_));
 sg13g2_o21ai_1 _24673_ (.B1(_04650_),
    .Y(_04651_),
    .A1(net216),
    .A2(_04649_));
 sg13g2_nand2_1 _24674_ (.Y(_04652_),
    .A(net46),
    .B(net42));
 sg13g2_o21ai_1 _24675_ (.B1(_04652_),
    .Y(_04653_),
    .A1(net39),
    .A2(_04036_));
 sg13g2_nand3_1 _24676_ (.B(_04649_),
    .C(_04653_),
    .A(net178),
    .Y(_04654_));
 sg13g2_a21oi_1 _24677_ (.A1(net216),
    .A2(_04647_),
    .Y(_04655_),
    .B1(_04087_));
 sg13g2_a21oi_1 _24678_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04656_),
    .B1(_04419_));
 sg13g2_a221oi_1 _24679_ (.B2(net160),
    .C1(_04656_),
    .B1(_04651_),
    .A1(_04068_),
    .Y(_04657_),
    .A2(_04647_));
 sg13g2_o21ai_1 _24680_ (.B1(net40),
    .Y(_04658_),
    .A1(net39),
    .A2(net137));
 sg13g2_a21oi_1 _24681_ (.A1(_04209_),
    .A2(net137),
    .Y(_04659_),
    .B1(_04649_));
 sg13g2_nand2_1 _24682_ (.Y(_04660_),
    .A(_04658_),
    .B(_04659_));
 sg13g2_o21ai_1 _24683_ (.B1(_04649_),
    .Y(_04661_),
    .A1(_04068_),
    .A2(net137));
 sg13g2_nand3b_1 _24684_ (.B(_04660_),
    .C(_04661_),
    .Y(_04662_),
    .A_N(net41));
 sg13g2_nand3_1 _24685_ (.B(_04086_),
    .C(_04647_),
    .A(net41),
    .Y(_04663_));
 sg13g2_a21oi_1 _24686_ (.A1(_04662_),
    .A2(_04663_),
    .Y(_04664_),
    .B1(_04419_));
 sg13g2_nor3_1 _24687_ (.A(_04646_),
    .B(_04657_),
    .C(_04664_),
    .Y(_04665_));
 sg13g2_buf_1 _24688_ (.A(_04665_),
    .X(_04666_));
 sg13g2_o21ai_1 _24689_ (.B1(_04646_),
    .Y(_04667_),
    .A1(_04657_),
    .A2(_04664_));
 sg13g2_nand2b_1 _24690_ (.Y(_04668_),
    .B(_04667_),
    .A_N(_04666_));
 sg13g2_nand2_1 _24691_ (.Y(_04669_),
    .A(net178),
    .B(_03980_));
 sg13g2_o21ai_1 _24692_ (.B1(net178),
    .Y(_04670_),
    .A1(_03955_),
    .A2(_03957_));
 sg13g2_nand3_1 _24693_ (.B(_04669_),
    .C(_04670_),
    .A(net40),
    .Y(_04671_));
 sg13g2_xnor2_1 _24694_ (.Y(_04672_),
    .A(net39),
    .B(_04671_));
 sg13g2_a22oi_1 _24695_ (.Y(_04673_),
    .B1(_04672_),
    .B2(net161),
    .A2(net34),
    .A1(_03043_));
 sg13g2_xor2_1 _24696_ (.B(_04673_),
    .A(_04637_),
    .X(_04674_));
 sg13g2_nand2_2 _24697_ (.Y(_04675_),
    .A(net140),
    .B(_04518_));
 sg13g2_a22oi_1 _24698_ (.Y(_04676_),
    .B1(_04366_),
    .B2(net44),
    .A2(net34),
    .A1(net161));
 sg13g2_nor2_1 _24699_ (.A(net183),
    .B(net45),
    .Y(_04677_));
 sg13g2_nand2_1 _24700_ (.Y(_04678_),
    .A(net34),
    .B(_04677_));
 sg13g2_o21ai_1 _24701_ (.B1(_04678_),
    .Y(_04679_),
    .A1(_04675_),
    .A2(_04676_));
 sg13g2_nand2b_1 _24702_ (.Y(_04680_),
    .B(_04679_),
    .A_N(_04674_));
 sg13g2_a22oi_1 _24703_ (.Y(_04681_),
    .B1(_04158_),
    .B2(net100),
    .A2(net44),
    .A1(net138));
 sg13g2_nand2_1 _24704_ (.Y(_04682_),
    .A(_02988_),
    .B(_04635_));
 sg13g2_nand4_1 _24705_ (.B(_04300_),
    .C(_04539_),
    .A(net100),
    .Y(_04683_),
    .D(_04682_));
 sg13g2_nand2b_1 _24706_ (.Y(_04684_),
    .B(_04683_),
    .A_N(_04681_));
 sg13g2_or2_1 _24707_ (.X(_04685_),
    .B(_04684_),
    .A(_04680_));
 sg13g2_buf_1 _24708_ (.A(_04685_),
    .X(_04686_));
 sg13g2_and2_1 _24709_ (.A(_04680_),
    .B(_04684_),
    .X(_04687_));
 sg13g2_buf_1 _24710_ (.A(_04687_),
    .X(_04688_));
 sg13g2_a21oi_1 _24711_ (.A1(_04668_),
    .A2(_04686_),
    .Y(_04689_),
    .B1(_04688_));
 sg13g2_nor2_1 _24712_ (.A(_04145_),
    .B(_04280_),
    .Y(_04690_));
 sg13g2_nand2_1 _24713_ (.Y(_04691_),
    .A(_02695_),
    .B(_04341_));
 sg13g2_nor2_1 _24714_ (.A(_04139_),
    .B(net62),
    .Y(_04692_));
 sg13g2_xor2_1 _24715_ (.B(_04692_),
    .A(_04691_),
    .X(_04693_));
 sg13g2_xnor2_1 _24716_ (.Y(_04694_),
    .A(_04690_),
    .B(_04693_));
 sg13g2_buf_1 _24717_ (.A(_04452_),
    .X(_04695_));
 sg13g2_a21oi_1 _24718_ (.A1(_02988_),
    .A2(_04123_),
    .Y(_04696_),
    .B1(_04154_));
 sg13g2_nor2_1 _24719_ (.A(net39),
    .B(_04696_),
    .Y(_04697_));
 sg13g2_a21oi_1 _24720_ (.A1(net39),
    .A2(_04036_),
    .Y(_04698_),
    .B1(_04697_));
 sg13g2_nand2_1 _24721_ (.Y(_04699_),
    .A(_04380_),
    .B(_04132_));
 sg13g2_nand3_1 _24722_ (.B(net34),
    .C(_04699_),
    .A(net138),
    .Y(_04700_));
 sg13g2_o21ai_1 _24723_ (.B1(_04700_),
    .Y(_04701_),
    .A1(net90),
    .A2(_04698_));
 sg13g2_buf_1 _24724_ (.A(_04701_),
    .X(_04702_));
 sg13g2_o21ai_1 _24725_ (.B1(net46),
    .Y(_04703_),
    .A1(_04208_),
    .A2(_04649_));
 sg13g2_nor2_1 _24726_ (.A(net42),
    .B(_04647_),
    .Y(_04704_));
 sg13g2_a21oi_1 _24727_ (.A1(_04209_),
    .A2(_04704_),
    .Y(_04705_),
    .B1(_04047_));
 sg13g2_nor2_1 _24728_ (.A(net46),
    .B(_04647_),
    .Y(_04706_));
 sg13g2_a22oi_1 _24729_ (.Y(_04707_),
    .B1(net137),
    .B2(_04706_),
    .A2(net40),
    .A1(net46));
 sg13g2_and4_1 _24730_ (.A(net161),
    .B(_04703_),
    .C(_04705_),
    .D(_04707_),
    .X(_04708_));
 sg13g2_buf_1 _24731_ (.A(_04708_),
    .X(_04709_));
 sg13g2_nor3_1 _24732_ (.A(_04068_),
    .B(_04355_),
    .C(_04649_),
    .Y(_04710_));
 sg13g2_nor2_1 _24733_ (.A(_04709_),
    .B(_04710_),
    .Y(_04711_));
 sg13g2_and2_1 _24734_ (.A(net38),
    .B(_04421_),
    .X(_04712_));
 sg13g2_nand3_1 _24735_ (.B(net38),
    .C(_04014_),
    .A(net161),
    .Y(_04713_));
 sg13g2_nor2_1 _24736_ (.A(net139),
    .B(net45),
    .Y(_04714_));
 sg13g2_mux2_1 _24737_ (.A0(_04712_),
    .A1(_04713_),
    .S(_04714_),
    .X(_04715_));
 sg13g2_nand2_1 _24738_ (.Y(_04716_),
    .A(net92),
    .B(_04518_));
 sg13g2_nor2_1 _24739_ (.A(_04691_),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_a221oi_1 _24740_ (.B2(net33),
    .C1(net36),
    .B1(net46),
    .A1(net183),
    .Y(_04718_),
    .A2(_03151_));
 sg13g2_xor2_1 _24741_ (.B(_04718_),
    .A(_04717_),
    .X(_04719_));
 sg13g2_xnor2_1 _24742_ (.Y(_04720_),
    .A(_04715_),
    .B(_04719_));
 sg13g2_xnor2_1 _24743_ (.Y(_04721_),
    .A(_04711_),
    .B(_04720_));
 sg13g2_xnor2_1 _24744_ (.Y(_04722_),
    .A(_04702_),
    .B(_04721_));
 sg13g2_xnor2_1 _24745_ (.Y(_04723_),
    .A(_04666_),
    .B(_04722_));
 sg13g2_xnor2_1 _24746_ (.Y(_04724_),
    .A(_04694_),
    .B(_04723_));
 sg13g2_xnor2_1 _24747_ (.Y(_04725_),
    .A(_04689_),
    .B(_04724_));
 sg13g2_buf_1 _24748_ (.A(net47),
    .X(_04726_));
 sg13g2_nor2_2 _24749_ (.A(net139),
    .B(net62),
    .Y(_04727_));
 sg13g2_xnor2_1 _24750_ (.Y(_04728_),
    .A(_04433_),
    .B(_04727_));
 sg13g2_nor4_2 _24751_ (.A(net183),
    .B(_04726_),
    .C(_04128_),
    .Y(_04729_),
    .D(_04728_));
 sg13g2_nor2_1 _24752_ (.A(_04500_),
    .B(_04280_),
    .Y(_04730_));
 sg13g2_a21oi_1 _24753_ (.A1(net100),
    .A2(_04539_),
    .Y(_04731_),
    .B1(_04730_));
 sg13g2_nand2b_1 _24754_ (.Y(_04732_),
    .B(_03975_),
    .A_N(_03972_));
 sg13g2_o21ai_1 _24755_ (.B1(_04732_),
    .Y(_04733_),
    .A1(net138),
    .A2(net49));
 sg13g2_nor3_1 _24756_ (.A(net90),
    .B(net52),
    .C(_04733_),
    .Y(_04734_));
 sg13g2_nor2_1 _24757_ (.A(_04731_),
    .B(_04734_),
    .Y(_04735_));
 sg13g2_xor2_1 _24758_ (.B(_04679_),
    .A(_04674_),
    .X(_04736_));
 sg13g2_nand2_1 _24759_ (.Y(_04737_),
    .A(_04729_),
    .B(_04735_));
 sg13g2_nand2_1 _24760_ (.Y(_04738_),
    .A(_04736_),
    .B(_04737_));
 sg13g2_o21ai_1 _24761_ (.B1(_04738_),
    .Y(_04739_),
    .A1(_04729_),
    .A2(_04735_));
 sg13g2_buf_1 _24762_ (.A(_04739_),
    .X(_04740_));
 sg13g2_buf_1 _24763_ (.A(net62),
    .X(_04741_));
 sg13g2_nor2_1 _24764_ (.A(net86),
    .B(net56),
    .Y(_04742_));
 sg13g2_nand2_1 _24765_ (.Y(_04743_),
    .A(_04093_),
    .B(_04547_));
 sg13g2_xnor2_1 _24766_ (.Y(_04744_),
    .A(_04742_),
    .B(_04743_));
 sg13g2_nand2b_1 _24767_ (.Y(_04745_),
    .B(_04686_),
    .A_N(_04688_));
 sg13g2_xor2_1 _24768_ (.B(_04745_),
    .A(_04668_),
    .X(_04746_));
 sg13g2_nand2_1 _24769_ (.Y(_04747_),
    .A(_04744_),
    .B(_04746_));
 sg13g2_nor2_1 _24770_ (.A(_04744_),
    .B(_04746_),
    .Y(_04748_));
 sg13g2_a21o_1 _24771_ (.A2(_04747_),
    .A1(_04740_),
    .B1(_04748_),
    .X(_04749_));
 sg13g2_o21ai_1 _24772_ (.B1(_04749_),
    .Y(_04750_),
    .A1(_04634_),
    .A2(_04725_));
 sg13g2_nand2_1 _24773_ (.Y(_04751_),
    .A(_04634_),
    .B(_04725_));
 sg13g2_nand2_1 _24774_ (.Y(_04752_),
    .A(_04750_),
    .B(_04751_));
 sg13g2_nor2b_1 _24775_ (.A(_04740_),
    .B_N(_04744_),
    .Y(_04753_));
 sg13g2_nand2b_1 _24776_ (.Y(_04754_),
    .B(_04740_),
    .A_N(_04744_));
 sg13g2_o21ai_1 _24777_ (.B1(_04754_),
    .Y(_04755_),
    .A1(_04746_),
    .A2(_04753_));
 sg13g2_xor2_1 _24778_ (.B(_04755_),
    .A(_04725_),
    .X(_04756_));
 sg13g2_xnor2_1 _24779_ (.Y(_04757_),
    .A(_04634_),
    .B(_04756_));
 sg13g2_nor4_1 _24780_ (.A(net118),
    .B(net90),
    .C(_04726_),
    .D(net45),
    .Y(_04758_));
 sg13g2_inv_1 _24781_ (.Y(_04759_),
    .A(_04758_));
 sg13g2_nand2_1 _24782_ (.Y(_04760_),
    .A(_04341_),
    .B(_04588_));
 sg13g2_nor2_1 _24783_ (.A(net47),
    .B(_04760_),
    .Y(_04761_));
 sg13g2_a21oi_1 _24784_ (.A1(net178),
    .A2(net54),
    .Y(_04762_),
    .B1(net49));
 sg13g2_xnor2_1 _24785_ (.Y(_04763_),
    .A(_04126_),
    .B(_04762_));
 sg13g2_nand2_1 _24786_ (.Y(_04764_),
    .A(_03973_),
    .B(_04126_));
 sg13g2_o21ai_1 _24787_ (.B1(_04764_),
    .Y(_04765_),
    .A1(net161),
    .A2(net43));
 sg13g2_xnor2_1 _24788_ (.Y(_04766_),
    .A(net43),
    .B(net53));
 sg13g2_nand4_1 _24789_ (.B(_04518_),
    .C(_04343_),
    .A(_03156_),
    .Y(_04767_),
    .D(_04766_));
 sg13g2_buf_1 _24790_ (.A(_04767_),
    .X(_04768_));
 sg13g2_nor2_1 _24791_ (.A(net118),
    .B(net56),
    .Y(_04769_));
 sg13g2_a21oi_1 _24792_ (.A1(net100),
    .A2(net53),
    .Y(_04770_),
    .B1(_04769_));
 sg13g2_or2_1 _24793_ (.X(_04771_),
    .B(_04770_),
    .A(_04768_));
 sg13g2_nor2_1 _24794_ (.A(net138),
    .B(net53),
    .Y(_04772_));
 sg13g2_nor4_1 _24795_ (.A(net160),
    .B(net90),
    .C(net56),
    .D(_04772_),
    .Y(_04773_));
 sg13g2_nand3b_1 _24796_ (.B(_04321_),
    .C(net216),
    .Y(_04774_),
    .A_N(net43));
 sg13g2_nand2b_1 _24797_ (.Y(_04775_),
    .B(_04274_),
    .A_N(_04342_));
 sg13g2_or2_1 _24798_ (.X(_04776_),
    .B(net43),
    .A(_04775_));
 sg13g2_nand3_1 _24799_ (.B(_04775_),
    .C(net43),
    .A(_03744_),
    .Y(_04777_));
 sg13g2_nand3_1 _24800_ (.B(_04776_),
    .C(_04777_),
    .A(_04774_),
    .Y(_04778_));
 sg13g2_nand2_1 _24801_ (.Y(_04779_),
    .A(net161),
    .B(net43));
 sg13g2_a21oi_1 _24802_ (.A1(net216),
    .A2(_04779_),
    .Y(_04780_),
    .B1(_04321_));
 sg13g2_nor4_1 _24803_ (.A(net90),
    .B(_04281_),
    .C(net56),
    .D(_04780_),
    .Y(_04781_));
 sg13g2_a21oi_1 _24804_ (.A1(_04773_),
    .A2(_04778_),
    .Y(_04782_),
    .B1(_04781_));
 sg13g2_nor2_1 _24805_ (.A(_02988_),
    .B(net54),
    .Y(_04783_));
 sg13g2_a21o_1 _24806_ (.A2(net54),
    .A1(_03051_),
    .B1(_04783_),
    .X(_04784_));
 sg13g2_nor3_1 _24807_ (.A(_03081_),
    .B(net44),
    .C(net54),
    .Y(_04785_));
 sg13g2_a21oi_1 _24808_ (.A1(_03051_),
    .A2(net44),
    .Y(_04786_),
    .B1(_04785_));
 sg13g2_nand3b_1 _24809_ (.B(net202),
    .C(_04786_),
    .Y(_04787_),
    .A_N(_04784_));
 sg13g2_xnor2_1 _24810_ (.Y(_04788_),
    .A(net181),
    .B(_04677_));
 sg13g2_o21ai_1 _24811_ (.B1(_04783_),
    .Y(_04789_),
    .A1(net43),
    .A2(_04788_));
 sg13g2_o21ai_1 _24812_ (.B1(_04789_),
    .Y(_04790_),
    .A1(net43),
    .A2(_04787_));
 sg13g2_buf_1 _24813_ (.A(_04790_),
    .X(_04791_));
 sg13g2_a21oi_1 _24814_ (.A1(_04025_),
    .A2(_04027_),
    .Y(_04792_),
    .B1(_04126_));
 sg13g2_nor2_1 _24815_ (.A(net52),
    .B(_04732_),
    .Y(_04793_));
 sg13g2_o21ai_1 _24816_ (.B1(_03744_),
    .Y(_04794_),
    .A1(_04792_),
    .A2(_04793_));
 sg13g2_nand3_1 _24817_ (.B(_04153_),
    .C(_04794_),
    .A(_04362_),
    .Y(_04795_));
 sg13g2_xnor2_1 _24818_ (.Y(_04796_),
    .A(_03974_),
    .B(net52));
 sg13g2_nand3b_1 _24819_ (.B(_04796_),
    .C(_04024_),
    .Y(_04797_),
    .A_N(_03972_));
 sg13g2_nand3_1 _24820_ (.B(_03972_),
    .C(_04033_),
    .A(_04026_),
    .Y(_04798_));
 sg13g2_a21o_1 _24821_ (.A2(_04798_),
    .A1(_04797_),
    .B1(_04636_),
    .X(_04799_));
 sg13g2_nand2_1 _24822_ (.Y(_04800_),
    .A(_03043_),
    .B(net44));
 sg13g2_nand3_1 _24823_ (.B(_04799_),
    .C(_04800_),
    .A(_04795_),
    .Y(_04801_));
 sg13g2_xnor2_1 _24824_ (.Y(_04802_),
    .A(_04675_),
    .B(_04801_));
 sg13g2_xnor2_1 _24825_ (.Y(_04803_),
    .A(_04791_),
    .B(_04802_));
 sg13g2_nand2_1 _24826_ (.Y(_04804_),
    .A(net100),
    .B(net53));
 sg13g2_xnor2_1 _24827_ (.Y(_04805_),
    .A(_04804_),
    .B(_04769_));
 sg13g2_nand2_1 _24828_ (.Y(_04806_),
    .A(_04768_),
    .B(_04805_));
 sg13g2_a22oi_1 _24829_ (.Y(_04807_),
    .B1(_04803_),
    .B2(_04806_),
    .A2(_04782_),
    .A1(_04771_));
 sg13g2_a221oi_1 _24830_ (.B2(_03069_),
    .C1(_04807_),
    .B1(_04765_),
    .A1(net161),
    .Y(_04808_),
    .A2(_04763_));
 sg13g2_a21oi_1 _24831_ (.A1(net139),
    .A2(_04760_),
    .Y(_04809_),
    .B1(net56));
 sg13g2_and2_1 _24832_ (.A(_04727_),
    .B(_04760_),
    .X(_04810_));
 sg13g2_buf_1 _24833_ (.A(_04810_),
    .X(_04811_));
 sg13g2_nand2_1 _24834_ (.Y(_04812_),
    .A(_04800_),
    .B(_04811_));
 sg13g2_and2_1 _24835_ (.A(_04795_),
    .B(_04799_),
    .X(_04813_));
 sg13g2_buf_1 _24836_ (.A(_04813_),
    .X(_04814_));
 sg13g2_mux2_1 _24837_ (.A0(_04809_),
    .A1(_04812_),
    .S(_04814_),
    .X(_04815_));
 sg13g2_nor2_2 _24838_ (.A(_03151_),
    .B(net45),
    .Y(_04816_));
 sg13g2_nor2_1 _24839_ (.A(_04816_),
    .B(_04809_),
    .Y(_04817_));
 sg13g2_a221oi_1 _24840_ (.B2(_04814_),
    .C1(_04791_),
    .B1(_04817_),
    .A1(_04816_),
    .Y(_04818_),
    .A2(_04811_));
 sg13g2_a21o_1 _24841_ (.A2(_04815_),
    .A1(_04791_),
    .B1(_04818_),
    .X(_04819_));
 sg13g2_nor2_1 _24842_ (.A(_04800_),
    .B(_04809_),
    .Y(_04820_));
 sg13g2_a21oi_1 _24843_ (.A1(_04776_),
    .A2(_04777_),
    .Y(_04821_),
    .B1(net160));
 sg13g2_nand2_1 _24844_ (.Y(_04822_),
    .A(net160),
    .B(_04281_));
 sg13g2_nand3_1 _24845_ (.B(_04779_),
    .C(_04822_),
    .A(net216),
    .Y(_04823_));
 sg13g2_nand2b_1 _24846_ (.Y(_04824_),
    .B(_04823_),
    .A_N(_04821_));
 sg13g2_nand3_1 _24847_ (.B(_04518_),
    .C(_04824_),
    .A(net100),
    .Y(_04825_));
 sg13g2_nand2b_1 _24848_ (.Y(_04826_),
    .B(_04811_),
    .A_N(_04814_));
 sg13g2_nor2_1 _24849_ (.A(_04791_),
    .B(_04826_),
    .Y(_04827_));
 sg13g2_a221oi_1 _24850_ (.B2(_04768_),
    .C1(_04827_),
    .B1(_04825_),
    .A1(_04791_),
    .Y(_04828_),
    .A2(_04820_));
 sg13g2_nor2_1 _24851_ (.A(_04770_),
    .B(_04803_),
    .Y(_04829_));
 sg13g2_a21oi_1 _24852_ (.A1(_04819_),
    .A2(_04828_),
    .Y(_04830_),
    .B1(_04829_));
 sg13g2_xnor2_1 _24853_ (.Y(_04831_),
    .A(_04729_),
    .B(_04735_));
 sg13g2_xor2_1 _24854_ (.B(_04831_),
    .A(_04736_),
    .X(_04832_));
 sg13g2_a21oi_1 _24855_ (.A1(net118),
    .A2(net90),
    .Y(_04833_),
    .B1(_04761_));
 sg13g2_a21oi_1 _24856_ (.A1(_03156_),
    .A2(net45),
    .Y(_04834_),
    .B1(_04833_));
 sg13g2_nand2_1 _24857_ (.Y(_04835_),
    .A(net118),
    .B(net47));
 sg13g2_o21ai_1 _24858_ (.B1(net54),
    .Y(_04836_),
    .A1(net90),
    .A2(net47));
 sg13g2_nand2_1 _24859_ (.Y(_04837_),
    .A(_04835_),
    .B(_04836_));
 sg13g2_nor2_2 _24860_ (.A(_04834_),
    .B(_04837_),
    .Y(_04838_));
 sg13g2_nand3_1 _24861_ (.B(_04838_),
    .C(_04816_),
    .A(net56),
    .Y(_04839_));
 sg13g2_nor2_1 _24862_ (.A(net91),
    .B(net56),
    .Y(_04840_));
 sg13g2_nor2_1 _24863_ (.A(_03040_),
    .B(net47),
    .Y(_04841_));
 sg13g2_nand4_1 _24864_ (.B(net53),
    .C(_04453_),
    .A(net45),
    .Y(_04842_),
    .D(_04841_));
 sg13g2_buf_1 _24865_ (.A(_04842_),
    .X(_04843_));
 sg13g2_inv_1 _24866_ (.Y(_04844_),
    .A(_04838_));
 sg13g2_nand3_1 _24867_ (.B(_04843_),
    .C(_04844_),
    .A(_04840_),
    .Y(_04845_));
 sg13g2_nand2b_1 _24868_ (.Y(_04846_),
    .B(net56),
    .A_N(_04843_));
 sg13g2_nand3_1 _24869_ (.B(_04840_),
    .C(_04816_),
    .A(net140),
    .Y(_04847_));
 sg13g2_nand4_1 _24870_ (.B(_04845_),
    .C(_04846_),
    .A(_04839_),
    .Y(_04848_),
    .D(_04847_));
 sg13g2_nand3_1 _24871_ (.B(_04727_),
    .C(_04838_),
    .A(_04716_),
    .Y(_04849_));
 sg13g2_nand3_1 _24872_ (.B(_04675_),
    .C(_04843_),
    .A(_04840_),
    .Y(_04850_));
 sg13g2_nand2_1 _24873_ (.Y(_04851_),
    .A(_04814_),
    .B(_04800_));
 sg13g2_a21oi_1 _24874_ (.A1(_04849_),
    .A2(_04850_),
    .Y(_04852_),
    .B1(_04851_));
 sg13g2_nand3_1 _24875_ (.B(_04838_),
    .C(_04816_),
    .A(net139),
    .Y(_04853_));
 sg13g2_a21oi_1 _24876_ (.A1(_04843_),
    .A2(_04853_),
    .Y(_04854_),
    .B1(net87));
 sg13g2_nand3_1 _24877_ (.B(_04727_),
    .C(_04843_),
    .A(_04840_),
    .Y(_04855_));
 sg13g2_nand3_1 _24878_ (.B(_04675_),
    .C(_04838_),
    .A(_04716_),
    .Y(_04856_));
 sg13g2_a21oi_1 _24879_ (.A1(_04855_),
    .A2(_04856_),
    .Y(_04857_),
    .B1(_04814_));
 sg13g2_nor4_1 _24880_ (.A(_04848_),
    .B(_04852_),
    .C(_04854_),
    .D(_04857_),
    .Y(_04858_));
 sg13g2_xor2_1 _24881_ (.B(_04858_),
    .A(_04832_),
    .X(_04859_));
 sg13g2_o21ai_1 _24882_ (.B1(_04859_),
    .Y(_04860_),
    .A1(_04808_),
    .A2(_04830_));
 sg13g2_nor3_1 _24883_ (.A(_04859_),
    .B(_04808_),
    .C(_04830_),
    .Y(_04861_));
 sg13g2_a21oi_1 _24884_ (.A1(_04761_),
    .A2(_04860_),
    .Y(_04862_),
    .B1(_04861_));
 sg13g2_nor2_1 _24885_ (.A(_04759_),
    .B(_04862_),
    .Y(_04863_));
 sg13g2_xnor2_1 _24886_ (.Y(_04864_),
    .A(_04740_),
    .B(_04744_));
 sg13g2_xnor2_1 _24887_ (.Y(_04865_),
    .A(_04746_),
    .B(_04864_));
 sg13g2_xnor2_1 _24888_ (.Y(_04866_),
    .A(_04727_),
    .B(_04851_));
 sg13g2_o21ai_1 _24889_ (.B1(_04843_),
    .Y(_04867_),
    .A1(_04844_),
    .A2(_04866_));
 sg13g2_nand2_1 _24890_ (.Y(_04868_),
    .A(_04832_),
    .B(_04867_));
 sg13g2_nor2_1 _24891_ (.A(_04865_),
    .B(_04868_),
    .Y(_04869_));
 sg13g2_nand3_1 _24892_ (.B(_04863_),
    .C(_04869_),
    .A(_04757_),
    .Y(_04870_));
 sg13g2_buf_1 _24893_ (.A(_04870_),
    .X(_04871_));
 sg13g2_nor4_2 _24894_ (.A(net118),
    .B(_04695_),
    .C(_04068_),
    .Y(_04872_),
    .D(_04077_));
 sg13g2_xor2_1 _24895_ (.B(_04720_),
    .A(_04711_),
    .X(_04873_));
 sg13g2_a21o_1 _24896_ (.A2(_04702_),
    .A1(_04666_),
    .B1(_04873_),
    .X(_04874_));
 sg13g2_o21ai_1 _24897_ (.B1(_04874_),
    .Y(_04875_),
    .A1(_04666_),
    .A2(_04702_));
 sg13g2_a21oi_1 _24898_ (.A1(net85),
    .A2(_04468_),
    .Y(_04876_),
    .B1(_04475_));
 sg13g2_xnor2_1 _24899_ (.Y(_04877_),
    .A(_04469_),
    .B(_04876_));
 sg13g2_buf_1 _24900_ (.A(_04877_),
    .X(_04878_));
 sg13g2_xor2_1 _24901_ (.B(_04878_),
    .A(_04517_),
    .X(_04879_));
 sg13g2_nor3_1 _24902_ (.A(_04709_),
    .B(_04717_),
    .C(_04710_),
    .Y(_04880_));
 sg13g2_xnor2_1 _24903_ (.Y(_04881_),
    .A(_04715_),
    .B(_04718_));
 sg13g2_o21ai_1 _24904_ (.B1(_04717_),
    .Y(_04882_),
    .A1(_04709_),
    .A2(_04710_));
 sg13g2_o21ai_1 _24905_ (.B1(_04882_),
    .Y(_04883_),
    .A1(_04880_),
    .A2(_04881_));
 sg13g2_buf_1 _24906_ (.A(_04883_),
    .X(_04884_));
 sg13g2_nand2_1 _24907_ (.Y(_04885_),
    .A(_04366_),
    .B(_04714_));
 sg13g2_o21ai_1 _24908_ (.B1(_04885_),
    .Y(_04886_),
    .A1(_03040_),
    .A2(net48));
 sg13g2_nor2_1 _24909_ (.A(net51),
    .B(_04425_),
    .Y(_04887_));
 sg13g2_a22oi_1 _24910_ (.Y(_04888_),
    .B1(_04887_),
    .B2(net44),
    .A2(_04886_),
    .A1(_04041_));
 sg13g2_or2_1 _24911_ (.X(_04889_),
    .B(_04888_),
    .A(net36));
 sg13g2_buf_1 _24912_ (.A(_04889_),
    .X(_04890_));
 sg13g2_and2_1 _24913_ (.A(_04461_),
    .B(_04462_),
    .X(_04891_));
 sg13g2_xor2_1 _24914_ (.B(_04462_),
    .A(_04461_),
    .X(_04892_));
 sg13g2_mux2_1 _24915_ (.A0(_04891_),
    .A1(_04892_),
    .S(_04421_),
    .X(_04893_));
 sg13g2_nor2_1 _24916_ (.A(_04421_),
    .B(_04461_),
    .Y(_04894_));
 sg13g2_a22oi_1 _24917_ (.Y(_04895_),
    .B1(_04894_),
    .B2(_04463_),
    .A2(_04893_),
    .A1(net37));
 sg13g2_buf_1 _24918_ (.A(_04895_),
    .X(_04896_));
 sg13g2_nand2_1 _24919_ (.Y(_04897_),
    .A(_04690_),
    .B(_04692_));
 sg13g2_nand2_1 _24920_ (.Y(_04898_),
    .A(_04691_),
    .B(_04897_));
 sg13g2_o21ai_1 _24921_ (.B1(_04898_),
    .Y(_04899_),
    .A1(_04690_),
    .A2(_04692_));
 sg13g2_buf_1 _24922_ (.A(_04899_),
    .X(_04900_));
 sg13g2_xor2_1 _24923_ (.B(_04900_),
    .A(_04896_),
    .X(_04901_));
 sg13g2_xnor2_1 _24924_ (.Y(_04902_),
    .A(_04890_),
    .B(_04901_));
 sg13g2_a21oi_1 _24925_ (.A1(_04500_),
    .A2(_04039_),
    .Y(_04903_),
    .B1(_04426_));
 sg13g2_nand2_1 _24926_ (.Y(_04904_),
    .A(_04054_),
    .B(_04086_));
 sg13g2_o21ai_1 _24927_ (.B1(_04904_),
    .Y(_04905_),
    .A1(_04054_),
    .A2(_04903_));
 sg13g2_o21ai_1 _24928_ (.B1(net138),
    .Y(_04906_),
    .A1(_04695_),
    .A2(net41));
 sg13g2_nor2_1 _24929_ (.A(_04068_),
    .B(_04906_),
    .Y(_04907_));
 sg13g2_a21oi_2 _24930_ (.B1(_04907_),
    .Y(_04908_),
    .A2(_04905_),
    .A1(_04380_));
 sg13g2_xor2_1 _24931_ (.B(_04908_),
    .A(_04902_),
    .X(_04909_));
 sg13g2_xnor2_1 _24932_ (.Y(_04910_),
    .A(_04884_),
    .B(_04909_));
 sg13g2_xor2_1 _24933_ (.B(_04910_),
    .A(_04879_),
    .X(_04911_));
 sg13g2_xnor2_1 _24934_ (.Y(_04912_),
    .A(_04875_),
    .B(_04911_));
 sg13g2_nand2_1 _24935_ (.Y(_04913_),
    .A(_04668_),
    .B(_04686_));
 sg13g2_nand3b_1 _24936_ (.B(_04913_),
    .C(_04694_),
    .Y(_04914_),
    .A_N(_04688_));
 sg13g2_nor2_1 _24937_ (.A(_04689_),
    .B(_04694_),
    .Y(_04915_));
 sg13g2_a21oi_1 _24938_ (.A1(_04723_),
    .A2(_04914_),
    .Y(_04916_),
    .B1(_04915_));
 sg13g2_xor2_1 _24939_ (.B(_04916_),
    .A(_04912_),
    .X(_04917_));
 sg13g2_xnor2_1 _24940_ (.Y(_04918_),
    .A(_04872_),
    .B(_04917_));
 sg13g2_nor3_2 _24941_ (.A(_04752_),
    .B(_04871_),
    .C(_04918_),
    .Y(_04919_));
 sg13g2_a21o_1 _24942_ (.A2(_04873_),
    .A1(_04666_),
    .B1(_04702_),
    .X(_04920_));
 sg13g2_nand2b_1 _24943_ (.Y(_04921_),
    .B(_04721_),
    .A_N(_04666_));
 sg13g2_a22oi_1 _24944_ (.Y(_04922_),
    .B1(_04920_),
    .B2(_04921_),
    .A2(_04910_),
    .A1(_04879_));
 sg13g2_nor2_1 _24945_ (.A(_04879_),
    .B(_04910_),
    .Y(_04923_));
 sg13g2_or2_1 _24946_ (.X(_04924_),
    .B(_04923_),
    .A(_04922_));
 sg13g2_o21ai_1 _24947_ (.B1(_04896_),
    .Y(_04925_),
    .A1(_04890_),
    .A2(_04900_));
 sg13g2_nand2_1 _24948_ (.Y(_04926_),
    .A(_04890_),
    .B(_04900_));
 sg13g2_nand2_1 _24949_ (.Y(_04927_),
    .A(_04925_),
    .B(_04926_));
 sg13g2_nand2_1 _24950_ (.Y(_04928_),
    .A(net138),
    .B(_04041_));
 sg13g2_a221oi_1 _24951_ (.B2(_04928_),
    .C1(net36),
    .B1(_04502_),
    .A1(_04062_),
    .Y(_04929_),
    .A2(_04588_));
 sg13g2_buf_1 _24952_ (.A(_04929_),
    .X(_04930_));
 sg13g2_nor2b_1 _24953_ (.A(_04421_),
    .B_N(_04461_),
    .Y(_04931_));
 sg13g2_nand2_1 _24954_ (.Y(_04932_),
    .A(_04153_),
    .B(_04493_));
 sg13g2_o21ai_1 _24955_ (.B1(_04932_),
    .Y(_04933_),
    .A1(_04463_),
    .A2(_04931_));
 sg13g2_xnor2_1 _24956_ (.Y(_04934_),
    .A(_04477_),
    .B(_04484_));
 sg13g2_mux2_1 _24957_ (.A0(_04466_),
    .A1(_04933_),
    .S(_04934_),
    .X(_04935_));
 sg13g2_buf_1 _24958_ (.A(_04935_),
    .X(_04936_));
 sg13g2_xnor2_1 _24959_ (.Y(_04937_),
    .A(_04930_),
    .B(_04936_));
 sg13g2_xnor2_1 _24960_ (.Y(_04938_),
    .A(_04927_),
    .B(_04937_));
 sg13g2_o21ai_1 _24961_ (.B1(_04017_),
    .Y(_04939_),
    .A1(net53),
    .A2(_04878_));
 sg13g2_a21oi_1 _24962_ (.A1(net93),
    .A2(_04878_),
    .Y(_04940_),
    .B1(_04741_));
 sg13g2_nor2_1 _24963_ (.A(net53),
    .B(_04741_),
    .Y(_04941_));
 sg13g2_mux2_1 _24964_ (.A0(_04547_),
    .A1(_04941_),
    .S(_04878_),
    .X(_04942_));
 sg13g2_nand2_1 _24965_ (.Y(_04943_),
    .A(_04001_),
    .B(_04942_));
 sg13g2_o21ai_1 _24966_ (.B1(_04943_),
    .Y(_04944_),
    .A1(net54),
    .A2(_04940_));
 sg13g2_a22oi_1 _24967_ (.Y(_04945_),
    .B1(_04944_),
    .B2(_04017_),
    .A2(_04939_),
    .A1(_04546_));
 sg13g2_xor2_1 _24968_ (.B(_04945_),
    .A(_04545_),
    .X(_04946_));
 sg13g2_xnor2_1 _24969_ (.Y(_04947_),
    .A(_04938_),
    .B(_04946_));
 sg13g2_and2_1 _24970_ (.A(_04884_),
    .B(_04902_),
    .X(_04948_));
 sg13g2_buf_1 _24971_ (.A(_04948_),
    .X(_04949_));
 sg13g2_inv_1 _24972_ (.Y(_04950_),
    .A(_04949_));
 sg13g2_nor2_1 _24973_ (.A(_04884_),
    .B(_04902_),
    .Y(_04951_));
 sg13g2_a21oi_1 _24974_ (.A1(_04950_),
    .A2(_04908_),
    .Y(_04952_),
    .B1(_04951_));
 sg13g2_xnor2_1 _24975_ (.Y(_04953_),
    .A(_04947_),
    .B(_04952_));
 sg13g2_nand3_1 _24976_ (.B(_04053_),
    .C(_04588_),
    .A(net35),
    .Y(_04954_));
 sg13g2_buf_1 _24977_ (.A(_04954_),
    .X(_04955_));
 sg13g2_xor2_1 _24978_ (.B(_04955_),
    .A(_04953_),
    .X(_04956_));
 sg13g2_xnor2_1 _24979_ (.Y(_04957_),
    .A(_04924_),
    .B(_04956_));
 sg13g2_nor2_1 _24980_ (.A(_04872_),
    .B(_04912_),
    .Y(_04958_));
 sg13g2_nand2b_1 _24981_ (.Y(_04959_),
    .B(_04723_),
    .A_N(_04694_));
 sg13g2_nor2b_1 _24982_ (.A(_04723_),
    .B_N(_04694_),
    .Y(_04960_));
 sg13g2_a21oi_1 _24983_ (.A1(_04689_),
    .A2(_04959_),
    .Y(_04961_),
    .B1(_04960_));
 sg13g2_nand2_1 _24984_ (.Y(_04962_),
    .A(_04872_),
    .B(_04912_));
 sg13g2_o21ai_1 _24985_ (.B1(_04962_),
    .Y(_04963_),
    .A1(_04958_),
    .A2(_04961_));
 sg13g2_nor2b_1 _24986_ (.A(_04957_),
    .B_N(_04963_),
    .Y(_04964_));
 sg13g2_buf_2 _24987_ (.A(_04964_),
    .X(_04965_));
 sg13g2_nor3_1 _24988_ (.A(_04922_),
    .B(_04955_),
    .C(_04923_),
    .Y(_04966_));
 sg13g2_nand2_1 _24989_ (.Y(_04967_),
    .A(_04955_),
    .B(_04924_));
 sg13g2_o21ai_1 _24990_ (.B1(_04967_),
    .Y(_04968_),
    .A1(_04953_),
    .A2(_04966_));
 sg13g2_buf_2 _24991_ (.A(_04968_),
    .X(_04969_));
 sg13g2_inv_1 _24992_ (.Y(_04970_),
    .A(_04938_));
 sg13g2_nor2_1 _24993_ (.A(_04908_),
    .B(_04951_),
    .Y(_04971_));
 sg13g2_nor3_1 _24994_ (.A(_04949_),
    .B(_04946_),
    .C(_04971_),
    .Y(_04972_));
 sg13g2_o21ai_1 _24995_ (.B1(_04946_),
    .Y(_04973_),
    .A1(_04949_),
    .A2(_04971_));
 sg13g2_o21ai_1 _24996_ (.B1(_04973_),
    .Y(_04974_),
    .A1(_04970_),
    .A2(_04972_));
 sg13g2_buf_1 _24997_ (.A(_04974_),
    .X(_04975_));
 sg13g2_inv_1 _24998_ (.Y(_04976_),
    .A(_04975_));
 sg13g2_nor4_2 _24999_ (.A(net118),
    .B(net90),
    .C(_04048_),
    .Y(_04977_),
    .D(_04101_));
 sg13g2_xor2_1 _25000_ (.B(_04550_),
    .A(_04526_),
    .X(_04978_));
 sg13g2_buf_2 _25001_ (.A(_04978_),
    .X(_04979_));
 sg13g2_nor2b_1 _25002_ (.A(_04930_),
    .B_N(_04936_),
    .Y(_04980_));
 sg13g2_a21oi_1 _25003_ (.A1(_04896_),
    .A2(_04900_),
    .Y(_04981_),
    .B1(_04890_));
 sg13g2_nor2_1 _25004_ (.A(_04896_),
    .B(_04900_),
    .Y(_04982_));
 sg13g2_nor2_1 _25005_ (.A(_04981_),
    .B(_04982_),
    .Y(_04983_));
 sg13g2_nand2b_1 _25006_ (.Y(_04984_),
    .B(_04930_),
    .A_N(_04936_));
 sg13g2_o21ai_1 _25007_ (.B1(_04984_),
    .Y(_04985_),
    .A1(_04980_),
    .A2(_04983_));
 sg13g2_buf_2 _25008_ (.A(_04985_),
    .X(_04986_));
 sg13g2_xnor2_1 _25009_ (.Y(_04987_),
    .A(_04001_),
    .B(_04341_));
 sg13g2_xnor2_1 _25010_ (.Y(_04988_),
    .A(_04545_),
    .B(_04987_));
 sg13g2_and3_1 _25011_ (.X(_04989_),
    .A(_04517_),
    .B(_04988_),
    .C(_04878_));
 sg13g2_buf_2 _25012_ (.A(_04989_),
    .X(_04990_));
 sg13g2_xor2_1 _25013_ (.B(_04498_),
    .A(_04487_),
    .X(_04991_));
 sg13g2_xnor2_1 _25014_ (.Y(_04992_),
    .A(_04504_),
    .B(_04991_));
 sg13g2_buf_8 _25015_ (.A(_04992_),
    .X(_04993_));
 sg13g2_xnor2_1 _25016_ (.Y(_04994_),
    .A(_04990_),
    .B(_04993_));
 sg13g2_xnor2_1 _25017_ (.Y(_04995_),
    .A(_04986_),
    .B(_04994_));
 sg13g2_xor2_1 _25018_ (.B(_04995_),
    .A(_04979_),
    .X(_04996_));
 sg13g2_xnor2_1 _25019_ (.Y(_04997_),
    .A(_04977_),
    .B(_04996_));
 sg13g2_xnor2_1 _25020_ (.Y(_04998_),
    .A(_04976_),
    .B(_04997_));
 sg13g2_buf_2 _25021_ (.A(_04998_),
    .X(_04999_));
 sg13g2_nand2_1 _25022_ (.Y(_05000_),
    .A(_04969_),
    .B(_04999_));
 sg13g2_nor2_1 _25023_ (.A(_04979_),
    .B(_04990_),
    .Y(_05001_));
 sg13g2_nand2b_1 _25024_ (.Y(_05002_),
    .B(_05001_),
    .A_N(_04993_));
 sg13g2_nor2_1 _25025_ (.A(_04979_),
    .B(_04993_),
    .Y(_05003_));
 sg13g2_inv_1 _25026_ (.Y(_05004_),
    .A(_04986_));
 sg13g2_o21ai_1 _25027_ (.B1(_05004_),
    .Y(_05005_),
    .A1(_05001_),
    .A2(_05003_));
 sg13g2_nand4_1 _25028_ (.B(_04986_),
    .C(_04990_),
    .A(_04979_),
    .Y(_05006_),
    .D(_04993_));
 sg13g2_or3_1 _25029_ (.A(_04986_),
    .B(_04990_),
    .C(_04993_),
    .X(_05007_));
 sg13g2_nand4_1 _25030_ (.B(_05005_),
    .C(_05006_),
    .A(_05002_),
    .Y(_05008_),
    .D(_05007_));
 sg13g2_nand2_1 _25031_ (.Y(_05009_),
    .A(_04499_),
    .B(_04505_));
 sg13g2_xor2_1 _25032_ (.B(_04563_),
    .A(_04459_),
    .X(_05010_));
 sg13g2_xnor2_1 _25033_ (.Y(_05011_),
    .A(_05009_),
    .B(_05010_));
 sg13g2_xnor2_1 _25034_ (.Y(_05012_),
    .A(_04551_),
    .B(_05011_));
 sg13g2_xnor2_1 _25035_ (.Y(_05013_),
    .A(net31),
    .B(_05012_));
 sg13g2_xnor2_1 _25036_ (.Y(_05014_),
    .A(_05008_),
    .B(_05013_));
 sg13g2_nand2_1 _25037_ (.Y(_05015_),
    .A(_04977_),
    .B(_04996_));
 sg13g2_nor2_1 _25038_ (.A(_04977_),
    .B(_04996_),
    .Y(_05016_));
 sg13g2_a21oi_1 _25039_ (.A1(_04976_),
    .A2(_05015_),
    .Y(_05017_),
    .B1(_05016_));
 sg13g2_xnor2_1 _25040_ (.Y(_05018_),
    .A(_05014_),
    .B(_05017_));
 sg13g2_a22oi_1 _25041_ (.Y(_05019_),
    .B1(_05000_),
    .B2(_05018_),
    .A2(_04965_),
    .A1(_04919_));
 sg13g2_nor2_1 _25042_ (.A(_04969_),
    .B(_04999_),
    .Y(_05020_));
 sg13g2_or2_1 _25043_ (.X(_05021_),
    .B(_05020_),
    .A(_05018_));
 sg13g2_nor2_1 _25044_ (.A(_04832_),
    .B(_04867_),
    .Y(_05022_));
 sg13g2_a21oi_1 _25045_ (.A1(_04716_),
    .A2(_04868_),
    .Y(_05023_),
    .B1(_05022_));
 sg13g2_inv_1 _25046_ (.Y(_05024_),
    .A(_05023_));
 sg13g2_nor2_1 _25047_ (.A(_04865_),
    .B(_05024_),
    .Y(_05025_));
 sg13g2_o21ai_1 _25048_ (.B1(_04860_),
    .Y(_05026_),
    .A1(_04761_),
    .A2(_04861_));
 sg13g2_a22oi_1 _25049_ (.Y(_05027_),
    .B1(_04759_),
    .B2(_05026_),
    .A2(_05024_),
    .A1(_04865_));
 sg13g2_o21ai_1 _25050_ (.B1(_04757_),
    .Y(_05028_),
    .A1(_05025_),
    .A2(_05027_));
 sg13g2_o21ai_1 _25051_ (.B1(_04863_),
    .Y(_05029_),
    .A1(_04757_),
    .A2(_05025_));
 sg13g2_a22oi_1 _25052_ (.Y(_05030_),
    .B1(_04871_),
    .B2(_04918_),
    .A2(_05029_),
    .A1(_05028_));
 sg13g2_a21oi_2 _25053_ (.B1(_05030_),
    .Y(_05031_),
    .A2(_04751_),
    .A1(_04750_));
 sg13g2_and3_1 _25054_ (.X(_05032_),
    .A(_05028_),
    .B(_05029_),
    .C(_04918_));
 sg13g2_buf_1 _25055_ (.A(_05032_),
    .X(_05033_));
 sg13g2_nor2b_1 _25056_ (.A(_04963_),
    .B_N(_04957_),
    .Y(_05034_));
 sg13g2_or2_1 _25057_ (.X(_05035_),
    .B(_05034_),
    .A(_05033_));
 sg13g2_inv_1 _25058_ (.Y(_05036_),
    .A(_04969_));
 sg13g2_xnor2_1 _25059_ (.Y(_05037_),
    .A(_04975_),
    .B(_04997_));
 sg13g2_inv_1 _25060_ (.Y(_05038_),
    .A(_04957_));
 sg13g2_a221oi_1 _25061_ (.B2(_04963_),
    .C1(_04919_),
    .B1(_05038_),
    .A1(_05036_),
    .Y(_05039_),
    .A2(_05037_));
 sg13g2_o21ai_1 _25062_ (.B1(_05039_),
    .Y(_05040_),
    .A1(_05031_),
    .A2(_05035_));
 sg13g2_nand3b_1 _25063_ (.B(_05021_),
    .C(_05040_),
    .Y(_05041_),
    .A_N(_05019_));
 sg13g2_nand2_1 _25064_ (.Y(_05042_),
    .A(_04979_),
    .B(_04995_));
 sg13g2_nor2_1 _25065_ (.A(net31),
    .B(_05012_),
    .Y(_05043_));
 sg13g2_and2_1 _25066_ (.A(net31),
    .B(_05012_),
    .X(_05044_));
 sg13g2_buf_1 _25067_ (.A(_05044_),
    .X(_05045_));
 sg13g2_a21oi_1 _25068_ (.A1(_04986_),
    .A2(_04993_),
    .Y(_05046_),
    .B1(_04990_));
 sg13g2_nor2_1 _25069_ (.A(_04986_),
    .B(_04993_),
    .Y(_05047_));
 sg13g2_nor2_1 _25070_ (.A(_05046_),
    .B(_05047_),
    .Y(_05048_));
 sg13g2_nor2_1 _25071_ (.A(_05045_),
    .B(_05048_),
    .Y(_05049_));
 sg13g2_or2_1 _25072_ (.X(_05050_),
    .B(_05049_),
    .A(_05043_));
 sg13g2_nand3_1 _25073_ (.B(_04564_),
    .C(_04583_),
    .A(net30),
    .Y(_05051_));
 sg13g2_o21ai_1 _25074_ (.B1(net29),
    .Y(_05052_),
    .A1(net30),
    .A2(_04564_));
 sg13g2_nand3b_1 _25075_ (.B(_05051_),
    .C(_05052_),
    .Y(_05053_),
    .A_N(_04586_));
 sg13g2_xor2_1 _25076_ (.B(_04578_),
    .A(net31),
    .X(_05054_));
 sg13g2_xnor2_1 _25077_ (.Y(_05055_),
    .A(_05053_),
    .B(_05054_));
 sg13g2_buf_1 _25078_ (.A(_05055_),
    .X(_05056_));
 sg13g2_nor2b_1 _25079_ (.A(_05042_),
    .B_N(_05045_),
    .Y(_05057_));
 sg13g2_o21ai_1 _25080_ (.B1(_05048_),
    .Y(_05058_),
    .A1(_05056_),
    .A2(_05057_));
 sg13g2_nand2b_1 _25081_ (.Y(_05059_),
    .B(_05056_),
    .A_N(_05043_));
 sg13g2_a22oi_1 _25082_ (.Y(_05060_),
    .B1(_05058_),
    .B2(_05059_),
    .A2(_05050_),
    .A1(_05042_));
 sg13g2_buf_1 _25083_ (.A(_05060_),
    .X(_05061_));
 sg13g2_nor2_1 _25084_ (.A(_04596_),
    .B(_04597_),
    .Y(_05062_));
 sg13g2_or3_1 _25085_ (.A(_04591_),
    .B(_05062_),
    .C(_04595_),
    .X(_05063_));
 sg13g2_buf_1 _25086_ (.A(_05063_),
    .X(_05064_));
 sg13g2_xnor2_1 _25087_ (.Y(_05065_),
    .A(_04600_),
    .B(_04628_));
 sg13g2_xor2_1 _25088_ (.B(_05065_),
    .A(_05064_),
    .X(_05066_));
 sg13g2_xor2_1 _25089_ (.B(_05066_),
    .A(_05061_),
    .X(_05067_));
 sg13g2_o21ai_1 _25090_ (.B1(_04975_),
    .Y(_05068_),
    .A1(_04977_),
    .A2(_04996_));
 sg13g2_a21oi_1 _25091_ (.A1(_05015_),
    .A2(_05068_),
    .Y(_05069_),
    .B1(_05014_));
 sg13g2_buf_2 _25092_ (.A(_05069_),
    .X(_05070_));
 sg13g2_nand4_1 _25093_ (.B(_04995_),
    .C(_05045_),
    .A(_04979_),
    .Y(_05071_),
    .D(_05048_));
 sg13g2_buf_1 _25094_ (.A(_05071_),
    .X(_05072_));
 sg13g2_a22oi_1 _25095_ (.Y(_05073_),
    .B1(_04590_),
    .B2(_05012_),
    .A2(_04995_),
    .A1(_04979_));
 sg13g2_inv_1 _25096_ (.Y(_05074_),
    .A(_05048_));
 sg13g2_o21ai_1 _25097_ (.B1(_05074_),
    .Y(_05075_),
    .A1(_05043_),
    .A2(_05073_));
 sg13g2_nand2_1 _25098_ (.Y(_05076_),
    .A(_05042_),
    .B(_05043_));
 sg13g2_nand3_1 _25099_ (.B(_05075_),
    .C(_05076_),
    .A(_05072_),
    .Y(_05077_));
 sg13g2_xor2_1 _25100_ (.B(_05077_),
    .A(_05056_),
    .X(_05078_));
 sg13g2_xnor2_1 _25101_ (.Y(_05079_),
    .A(_05070_),
    .B(_05078_));
 sg13g2_nand2b_1 _25102_ (.Y(_05080_),
    .B(_05079_),
    .A_N(_05067_));
 sg13g2_nand2_1 _25103_ (.Y(_05081_),
    .A(_05056_),
    .B(_05070_));
 sg13g2_o21ai_1 _25104_ (.B1(_05066_),
    .Y(_05082_),
    .A1(_05072_),
    .A2(_05081_));
 sg13g2_nand2_1 _25105_ (.Y(_05083_),
    .A(_05075_),
    .B(_05076_));
 sg13g2_nor2_1 _25106_ (.A(_05056_),
    .B(_05070_),
    .Y(_05084_));
 sg13g2_a22oi_1 _25107_ (.Y(_05085_),
    .B1(_05084_),
    .B2(_05072_),
    .A2(_05081_),
    .A1(_05083_));
 sg13g2_nand2_1 _25108_ (.Y(_05086_),
    .A(_05082_),
    .B(_05085_));
 sg13g2_o21ai_1 _25109_ (.B1(_05086_),
    .Y(_05087_),
    .A1(_05041_),
    .A2(_05080_));
 sg13g2_buf_2 _25110_ (.A(_05087_),
    .X(_05088_));
 sg13g2_o21ai_1 _25111_ (.B1(_05088_),
    .Y(_05089_),
    .A1(_04417_),
    .A2(_04632_));
 sg13g2_a21o_1 _25112_ (.A2(_04621_),
    .A1(_04568_),
    .B1(_04620_),
    .X(_05090_));
 sg13g2_a21oi_1 _25113_ (.A1(_04612_),
    .A2(_04614_),
    .Y(_05091_),
    .B1(_04620_));
 sg13g2_nand3_1 _25114_ (.B(_04614_),
    .C(_04621_),
    .A(_04612_),
    .Y(_05092_));
 sg13g2_o21ai_1 _25115_ (.B1(_05092_),
    .Y(_05093_),
    .A1(_04623_),
    .A2(_05091_));
 sg13g2_a22oi_1 _25116_ (.Y(_05094_),
    .B1(_04575_),
    .B2(_05093_),
    .A2(_05090_),
    .A1(_04615_));
 sg13g2_buf_1 _25117_ (.A(_05094_),
    .X(_05095_));
 sg13g2_nor2_1 _25118_ (.A(_05095_),
    .B(_04416_),
    .Y(_05096_));
 sg13g2_nor2_1 _25119_ (.A(_05095_),
    .B(_04403_),
    .Y(_05097_));
 sg13g2_nor2b_1 _25120_ (.A(_04631_),
    .B_N(_05097_),
    .Y(_05098_));
 sg13g2_o21ai_1 _25121_ (.B1(_05088_),
    .Y(_05099_),
    .A1(_05096_),
    .A2(_05098_));
 sg13g2_inv_1 _25122_ (.Y(_05100_),
    .A(_05095_));
 sg13g2_inv_1 _25123_ (.Y(_05101_),
    .A(_04416_));
 sg13g2_nor3_1 _25124_ (.A(_04403_),
    .B(_04631_),
    .C(_04416_),
    .Y(_05102_));
 sg13g2_a221oi_1 _25125_ (.B2(_05101_),
    .C1(_05102_),
    .B1(_05097_),
    .A1(_05100_),
    .Y(_05103_),
    .A2(_04632_));
 sg13g2_nand3_1 _25126_ (.B(_05099_),
    .C(_05103_),
    .A(_05089_),
    .Y(_05104_));
 sg13g2_buf_2 _25127_ (.A(_05104_),
    .X(_05105_));
 sg13g2_o21ai_1 _25128_ (.B1(_04407_),
    .Y(_05106_),
    .A1(_04404_),
    .A2(_04405_));
 sg13g2_nand2_1 _25129_ (.Y(_05107_),
    .A(_04404_),
    .B(_04405_));
 sg13g2_and2_1 _25130_ (.A(_05106_),
    .B(_05107_),
    .X(_05108_));
 sg13g2_buf_1 _25131_ (.A(_05108_),
    .X(_05109_));
 sg13g2_nor2b_1 _25132_ (.A(_04243_),
    .B_N(_04249_),
    .Y(_05110_));
 sg13g2_inv_1 _25133_ (.Y(_05111_),
    .A(_04251_));
 sg13g2_nand2_1 _25134_ (.Y(_05112_),
    .A(_05109_),
    .B(_04249_));
 sg13g2_a221oi_1 _25135_ (.B2(_04242_),
    .C1(_04249_),
    .B1(_04181_),
    .A1(_05106_),
    .Y(_05113_),
    .A2(_05107_));
 sg13g2_a221oi_1 _25136_ (.B2(_05112_),
    .C1(_05113_),
    .B1(_05111_),
    .A1(_05109_),
    .Y(_05114_),
    .A2(_05110_));
 sg13g2_xnor2_1 _25137_ (.Y(_05115_),
    .A(net28),
    .B(_05114_));
 sg13g2_nor2b_1 _25138_ (.A(_04241_),
    .B_N(_04249_),
    .Y(_05116_));
 sg13g2_nand2b_1 _25139_ (.Y(_05117_),
    .B(_04241_),
    .A_N(_04249_));
 sg13g2_nand2b_1 _25140_ (.Y(_05118_),
    .B(_05117_),
    .A_N(_05116_));
 sg13g2_a21o_1 _25141_ (.A2(_04407_),
    .A1(_04404_),
    .B1(_04405_),
    .X(_05119_));
 sg13g2_o21ai_1 _25142_ (.B1(_05119_),
    .Y(_05120_),
    .A1(_04404_),
    .A2(_04407_));
 sg13g2_xor2_1 _25143_ (.B(_05120_),
    .A(_05118_),
    .X(_05121_));
 sg13g2_xnor2_1 _25144_ (.Y(_05122_),
    .A(_04250_),
    .B(_05121_));
 sg13g2_nor2_1 _25145_ (.A(_04410_),
    .B(_04415_),
    .Y(_05123_));
 sg13g2_buf_1 _25146_ (.A(_05123_),
    .X(_05124_));
 sg13g2_xnor2_1 _25147_ (.Y(_05125_),
    .A(_05122_),
    .B(_05124_));
 sg13g2_buf_2 _25148_ (.A(_05125_),
    .X(_05126_));
 sg13g2_and2_1 _25149_ (.A(_05115_),
    .B(_05126_),
    .X(_05127_));
 sg13g2_a21oi_1 _25150_ (.A1(_04181_),
    .A2(_05117_),
    .Y(_05128_),
    .B1(_05116_));
 sg13g2_mux2_1 _25151_ (.A0(_04251_),
    .A1(_05128_),
    .S(net28),
    .X(_05129_));
 sg13g2_nand3b_1 _25152_ (.B(_05124_),
    .C(_05109_),
    .Y(_05130_),
    .A_N(_05129_));
 sg13g2_inv_1 _25153_ (.Y(_05131_),
    .A(_05116_));
 sg13g2_mux2_1 _25154_ (.A0(_05117_),
    .A1(_05131_),
    .S(net28),
    .X(_05132_));
 sg13g2_or3_1 _25155_ (.A(_04259_),
    .B(_04181_),
    .C(_05118_),
    .X(_05133_));
 sg13g2_o21ai_1 _25156_ (.B1(_05133_),
    .Y(_05134_),
    .A1(_04250_),
    .A2(_05132_));
 sg13g2_o21ai_1 _25157_ (.B1(_05134_),
    .Y(_05135_),
    .A1(_05109_),
    .A2(_05124_));
 sg13g2_and2_1 _25158_ (.A(_05130_),
    .B(_05135_),
    .X(_05136_));
 sg13g2_inv_1 _25159_ (.Y(_05137_),
    .A(_05136_));
 sg13g2_a21oi_1 _25160_ (.A1(_05105_),
    .A2(_05127_),
    .Y(_05138_),
    .B1(_05137_));
 sg13g2_xnor2_1 _25161_ (.Y(_05139_),
    .A(_04262_),
    .B(_05138_));
 sg13g2_buf_1 _25162_ (.A(net303),
    .X(_05140_));
 sg13g2_xnor2_1 _25163_ (.Y(_05141_),
    .A(_04969_),
    .B(_04999_));
 sg13g2_nor4_1 _25164_ (.A(_05031_),
    .B(_05033_),
    .C(_05141_),
    .D(_05034_),
    .Y(_05142_));
 sg13g2_or3_1 _25165_ (.A(_04752_),
    .B(_04871_),
    .C(_04918_),
    .X(_05143_));
 sg13g2_buf_1 _25166_ (.A(_05143_),
    .X(_05144_));
 sg13g2_o21ai_1 _25167_ (.B1(_05037_),
    .Y(_05145_),
    .A1(_05036_),
    .A2(_04919_));
 sg13g2_o21ai_1 _25168_ (.B1(_05145_),
    .Y(_05146_),
    .A1(_04969_),
    .A2(_05144_));
 sg13g2_o21ai_1 _25169_ (.B1(_05018_),
    .Y(_05147_),
    .A1(_05142_),
    .A2(_05146_));
 sg13g2_inv_1 _25170_ (.Y(_05148_),
    .A(_05070_));
 sg13g2_xor2_1 _25171_ (.B(_05017_),
    .A(_05014_),
    .X(_05149_));
 sg13g2_a21oi_1 _25172_ (.A1(_05141_),
    .A2(_05144_),
    .Y(_05150_),
    .B1(_05149_));
 sg13g2_nor3_1 _25173_ (.A(_04969_),
    .B(_04999_),
    .C(_05144_),
    .Y(_05151_));
 sg13g2_o21ai_1 _25174_ (.B1(_04965_),
    .Y(_05152_),
    .A1(_05150_),
    .A2(_05151_));
 sg13g2_nand3_1 _25175_ (.B(_05148_),
    .C(_05152_),
    .A(_05147_),
    .Y(_05153_));
 sg13g2_and2_1 _25176_ (.A(_05070_),
    .B(_04965_),
    .X(_05154_));
 sg13g2_o21ai_1 _25177_ (.B1(_05154_),
    .Y(_05155_),
    .A1(_05150_),
    .A2(_05151_));
 sg13g2_xor2_1 _25178_ (.B(_04403_),
    .A(_05095_),
    .X(_05156_));
 sg13g2_nor2b_1 _25179_ (.A(_05156_),
    .B_N(_04631_),
    .Y(_05157_));
 sg13g2_or2_1 _25180_ (.X(_05158_),
    .B(_05157_),
    .A(_05067_));
 sg13g2_a21oi_1 _25181_ (.A1(_05078_),
    .A2(_05155_),
    .Y(_05159_),
    .B1(_05158_));
 sg13g2_nor3_1 _25182_ (.A(_04600_),
    .B(_04628_),
    .C(_04610_),
    .Y(_05160_));
 sg13g2_nand2_1 _25183_ (.Y(_05161_),
    .A(_04600_),
    .B(_04628_));
 sg13g2_nand3b_1 _25184_ (.B(_04628_),
    .C(_04610_),
    .Y(_05162_),
    .A_N(_04600_));
 sg13g2_mux2_1 _25185_ (.A0(_05161_),
    .A1(_05162_),
    .S(_05064_),
    .X(_05163_));
 sg13g2_and2_1 _25186_ (.A(_05156_),
    .B(_05163_),
    .X(_05164_));
 sg13g2_nand2b_1 _25187_ (.Y(_05165_),
    .B(_04631_),
    .A_N(_05061_));
 sg13g2_a22oi_1 _25188_ (.Y(_05166_),
    .B1(_05164_),
    .B2(_05165_),
    .A2(_05160_),
    .A1(_05061_));
 sg13g2_inv_1 _25189_ (.Y(_05167_),
    .A(_05166_));
 sg13g2_a21o_1 _25190_ (.A2(_05159_),
    .A1(_05153_),
    .B1(_05167_),
    .X(_05168_));
 sg13g2_buf_1 _25191_ (.A(_05168_),
    .X(_05169_));
 sg13g2_nor2_1 _25192_ (.A(_04397_),
    .B(_04412_),
    .Y(_05170_));
 sg13g2_and2_1 _25193_ (.A(_04397_),
    .B(_04414_),
    .X(_05171_));
 sg13g2_o21ai_1 _25194_ (.B1(_04412_),
    .Y(_05172_),
    .A1(_04397_),
    .A2(_04414_));
 sg13g2_mux2_1 _25195_ (.A0(_05171_),
    .A1(_05172_),
    .S(_05095_),
    .X(_05173_));
 sg13g2_nor2_1 _25196_ (.A(_05170_),
    .B(_05173_),
    .Y(_05174_));
 sg13g2_xnor2_1 _25197_ (.Y(_05175_),
    .A(_04410_),
    .B(_05174_));
 sg13g2_nand2_1 _25198_ (.Y(_05176_),
    .A(_05175_),
    .B(_05126_));
 sg13g2_inv_1 _25199_ (.Y(_05177_),
    .A(_05176_));
 sg13g2_nand2b_1 _25200_ (.Y(_05178_),
    .B(_04410_),
    .A_N(_04414_));
 sg13g2_nor2b_1 _25201_ (.A(_04410_),
    .B_N(_04412_),
    .Y(_05179_));
 sg13g2_a21o_1 _25202_ (.A2(_05178_),
    .A1(_04397_),
    .B1(_05179_),
    .X(_05180_));
 sg13g2_a21oi_1 _25203_ (.A1(_05100_),
    .A2(_05180_),
    .Y(_05181_),
    .B1(_05124_));
 sg13g2_or2_1 _25204_ (.X(_05182_),
    .B(_05181_),
    .A(_05122_));
 sg13g2_buf_1 _25205_ (.A(_05182_),
    .X(_05183_));
 sg13g2_inv_1 _25206_ (.Y(_05184_),
    .A(_05183_));
 sg13g2_a21oi_1 _25207_ (.A1(_05169_),
    .A2(_05177_),
    .Y(_05185_),
    .B1(_05184_));
 sg13g2_xnor2_1 _25208_ (.Y(_05186_),
    .A(_05115_),
    .B(_05185_));
 sg13g2_nor2_1 _25209_ (.A(_05140_),
    .B(_05186_),
    .Y(_05187_));
 sg13g2_a21o_1 _25210_ (.A2(_05139_),
    .A1(_02409_),
    .B1(_05187_),
    .X(_05188_));
 sg13g2_buf_1 _25211_ (.A(net296),
    .X(_05189_));
 sg13g2_nor2b_1 _25212_ (.A(_04255_),
    .B_N(_04119_),
    .Y(_05190_));
 sg13g2_a22oi_1 _25213_ (.Y(_05191_),
    .B1(_04112_),
    .B2(net102),
    .A2(_03995_),
    .A1(_04113_));
 sg13g2_o21ai_1 _25214_ (.B1(_04044_),
    .Y(_05192_),
    .A1(_03999_),
    .A2(net32));
 sg13g2_o21ai_1 _25215_ (.B1(_05192_),
    .Y(_05193_),
    .A1(net103),
    .A2(_05191_));
 sg13g2_and3_1 _25216_ (.X(_05194_),
    .A(net241),
    .B(_04111_),
    .C(_05193_));
 sg13g2_nor3_1 _25217_ (.A(net254),
    .B(_04099_),
    .C(_04108_),
    .Y(_05195_));
 sg13g2_xor2_1 _25218_ (.B(_05195_),
    .A(_05194_),
    .X(_05196_));
 sg13g2_xnor2_1 _25219_ (.Y(_05197_),
    .A(_05190_),
    .B(_05196_));
 sg13g2_nor2_1 _25220_ (.A(_05122_),
    .B(_05124_),
    .Y(_05198_));
 sg13g2_and2_1 _25221_ (.A(_05122_),
    .B(_05124_),
    .X(_05199_));
 sg13g2_o21ai_1 _25222_ (.B1(_05175_),
    .Y(_05200_),
    .A1(_05198_),
    .A2(_05199_));
 sg13g2_nand2_1 _25223_ (.Y(_05201_),
    .A(_05183_),
    .B(_05200_));
 sg13g2_a21o_1 _25224_ (.A2(_04175_),
    .A1(_04119_),
    .B1(_04176_),
    .X(_05202_));
 sg13g2_buf_1 _25225_ (.A(_05202_),
    .X(_05203_));
 sg13g2_or2_1 _25226_ (.X(_05204_),
    .B(_05112_),
    .A(_04243_));
 sg13g2_o21ai_1 _25227_ (.B1(_05112_),
    .Y(_05205_),
    .A1(_05113_),
    .A2(_05111_));
 sg13g2_nand3_1 _25228_ (.B(_05204_),
    .C(_05205_),
    .A(_05203_),
    .Y(_05206_));
 sg13g2_nor4_1 _25229_ (.A(_04250_),
    .B(_04241_),
    .C(_05112_),
    .D(_05203_),
    .Y(_05207_));
 sg13g2_or2_1 _25230_ (.X(_05208_),
    .B(_04251_),
    .A(_04249_));
 sg13g2_nand2b_1 _25231_ (.Y(_05209_),
    .B(_04252_),
    .A_N(_05109_));
 sg13g2_a221oi_1 _25232_ (.B2(_05209_),
    .C1(_04177_),
    .B1(_05208_),
    .A1(_04181_),
    .Y(_05210_),
    .A2(_04242_));
 sg13g2_nor3_1 _25233_ (.A(net28),
    .B(_05207_),
    .C(_05210_),
    .Y(_05211_));
 sg13g2_a21oi_2 _25234_ (.B1(_05211_),
    .Y(_05212_),
    .A2(_05206_),
    .A1(net28));
 sg13g2_nand3_1 _25235_ (.B(_05201_),
    .C(_05212_),
    .A(_05197_),
    .Y(_05213_));
 sg13g2_nand2_1 _25236_ (.Y(_05214_),
    .A(_05166_),
    .B(_05183_));
 sg13g2_a21oi_1 _25237_ (.A1(_05153_),
    .A2(_05159_),
    .Y(_05215_),
    .B1(_05214_));
 sg13g2_nand2_1 _25238_ (.Y(_05216_),
    .A(_05109_),
    .B(_05208_));
 sg13g2_a21oi_1 _25239_ (.A1(_04252_),
    .A2(_05216_),
    .Y(_05217_),
    .B1(net28));
 sg13g2_a21oi_1 _25240_ (.A1(net28),
    .A2(_05112_),
    .Y(_05218_),
    .B1(_04243_));
 sg13g2_o21ai_1 _25241_ (.B1(_05203_),
    .Y(_05219_),
    .A1(_05217_),
    .A2(_05218_));
 sg13g2_nand2b_1 _25242_ (.Y(_05220_),
    .B(_05197_),
    .A_N(_05219_));
 sg13g2_o21ai_1 _25243_ (.B1(_05220_),
    .Y(_05221_),
    .A1(_05213_),
    .A2(_05215_));
 sg13g2_o21ai_1 _25244_ (.B1(_05212_),
    .Y(_05222_),
    .A1(_05184_),
    .A2(_05177_));
 sg13g2_nor2b_1 _25245_ (.A(_05197_),
    .B_N(_05219_),
    .Y(_05223_));
 sg13g2_o21ai_1 _25246_ (.B1(_05223_),
    .Y(_05224_),
    .A1(_05215_),
    .A2(_05222_));
 sg13g2_nand2b_1 _25247_ (.Y(_05225_),
    .B(_05224_),
    .A_N(_05221_));
 sg13g2_buf_1 _25248_ (.A(_05225_),
    .X(_05226_));
 sg13g2_xnor2_1 _25249_ (.Y(_05227_),
    .A(_05126_),
    .B(_05105_));
 sg13g2_nand2_1 _25250_ (.Y(_05228_),
    .A(net296),
    .B(_05227_));
 sg13g2_o21ai_1 _25251_ (.B1(_05228_),
    .Y(_05229_),
    .A1(net290),
    .A2(_05226_));
 sg13g2_buf_1 _25252_ (.A(net324),
    .X(_05230_));
 sg13g2_buf_1 _25253_ (.A(net315),
    .X(_05231_));
 sg13g2_mux2_1 _25254_ (.A0(_05188_),
    .A1(_05229_),
    .S(net310),
    .X(_05232_));
 sg13g2_buf_1 _25255_ (.A(_05232_),
    .X(_05233_));
 sg13g2_buf_1 _25256_ (.A(net297),
    .X(_05234_));
 sg13g2_xor2_1 _25257_ (.B(_05169_),
    .A(_05175_),
    .X(_05235_));
 sg13g2_xnor2_1 _25258_ (.Y(_05236_),
    .A(_05041_),
    .B(_05079_));
 sg13g2_inv_1 _25259_ (.Y(_05237_),
    .A(_05236_));
 sg13g2_nand2_1 _25260_ (.Y(_05238_),
    .A(_05237_),
    .B(_02409_));
 sg13g2_o21ai_1 _25261_ (.B1(_05238_),
    .Y(_05239_),
    .A1(net296),
    .A2(_05235_));
 sg13g2_xor2_1 _25262_ (.B(_04631_),
    .A(_05156_),
    .X(_05240_));
 sg13g2_xor2_1 _25263_ (.B(_05240_),
    .A(_05088_),
    .X(_05241_));
 sg13g2_nor2_1 _25264_ (.A(_05070_),
    .B(_05021_),
    .Y(_05242_));
 sg13g2_inv_1 _25265_ (.Y(_05243_),
    .A(_05078_));
 sg13g2_a21oi_1 _25266_ (.A1(_05070_),
    .A2(_05020_),
    .Y(_05244_),
    .B1(_05243_));
 sg13g2_inv_1 _25267_ (.Y(_05245_),
    .A(_05031_));
 sg13g2_nor3_1 _25268_ (.A(_05033_),
    .B(_05141_),
    .C(_05034_),
    .Y(_05246_));
 sg13g2_xnor2_1 _25269_ (.Y(_05247_),
    .A(_05036_),
    .B(_04999_));
 sg13g2_a21o_1 _25270_ (.A2(_04965_),
    .A1(_05247_),
    .B1(_04919_),
    .X(_05248_));
 sg13g2_nand2b_1 _25271_ (.Y(_05249_),
    .B(_05141_),
    .A_N(_04965_));
 sg13g2_nand2_1 _25272_ (.Y(_05250_),
    .A(_05149_),
    .B(_05078_));
 sg13g2_a221oi_1 _25273_ (.B2(_05249_),
    .C1(_05250_),
    .B1(_05248_),
    .A1(_05245_),
    .Y(_05251_),
    .A2(_05246_));
 sg13g2_or2_1 _25274_ (.X(_05252_),
    .B(_05020_),
    .A(_05070_));
 sg13g2_nand2_1 _25275_ (.Y(_05253_),
    .A(_05149_),
    .B(_05148_));
 sg13g2_a221oi_1 _25276_ (.B2(_05253_),
    .C1(_05142_),
    .B1(_05252_),
    .A1(_05248_),
    .Y(_05254_),
    .A2(_05249_));
 sg13g2_nor4_2 _25277_ (.A(_05242_),
    .B(_05244_),
    .C(_05251_),
    .Y(_05255_),
    .D(_05254_));
 sg13g2_xnor2_1 _25278_ (.Y(_05256_),
    .A(_05067_),
    .B(_05255_));
 sg13g2_nor2_1 _25279_ (.A(net303),
    .B(_05256_),
    .Y(_05257_));
 sg13g2_a21o_1 _25280_ (.A2(_05241_),
    .A1(net296),
    .B1(_05257_),
    .X(_05258_));
 sg13g2_mux2_1 _25281_ (.A0(_05239_),
    .A1(_05258_),
    .S(net316),
    .X(_05259_));
 sg13g2_nand2_1 _25282_ (.Y(_05260_),
    .A(net289),
    .B(_05259_));
 sg13g2_inv_1 _25283_ (.Y(_05261_),
    .A(_05260_));
 sg13g2_a21oi_1 _25284_ (.A1(net298),
    .A2(_05233_),
    .Y(_05262_),
    .B1(_05261_));
 sg13g2_nor2_1 _25285_ (.A(_04105_),
    .B(_04107_),
    .Y(_05263_));
 sg13g2_nand2_1 _25286_ (.Y(_05264_),
    .A(net96),
    .B(_04443_));
 sg13g2_nand3_1 _25287_ (.B(_04044_),
    .C(_05264_),
    .A(_04218_),
    .Y(_05265_));
 sg13g2_nand2b_1 _25288_ (.Y(_05266_),
    .B(_02807_),
    .A_N(_05265_));
 sg13g2_o21ai_1 _25289_ (.B1(_05266_),
    .Y(_05267_),
    .A1(_02807_),
    .A2(_05263_));
 sg13g2_nor2_1 _25290_ (.A(_05263_),
    .B(_05265_),
    .Y(_05268_));
 sg13g2_a21oi_1 _25291_ (.A1(net230),
    .A2(_05267_),
    .Y(_05269_),
    .B1(_05268_));
 sg13g2_a21oi_1 _25292_ (.A1(_05194_),
    .A2(_05195_),
    .Y(_05270_),
    .B1(_05269_));
 sg13g2_buf_2 _25293_ (.A(_05270_),
    .X(_05271_));
 sg13g2_nor2b_1 _25294_ (.A(_05197_),
    .B_N(_05212_),
    .Y(_05272_));
 sg13g2_nor2b_1 _25295_ (.A(_05271_),
    .B_N(_05272_),
    .Y(_05273_));
 sg13g2_nor2_1 _25296_ (.A(_05067_),
    .B(_05157_),
    .Y(_05274_));
 sg13g2_a21oi_1 _25297_ (.A1(_05274_),
    .A2(_05255_),
    .Y(_05275_),
    .B1(_05167_));
 sg13g2_o21ai_1 _25298_ (.B1(_05183_),
    .Y(_05276_),
    .A1(_05176_),
    .A2(_05275_));
 sg13g2_nand2_1 _25299_ (.Y(_05277_),
    .A(_05273_),
    .B(_05276_));
 sg13g2_buf_1 _25300_ (.A(_05277_),
    .X(_05278_));
 sg13g2_o21ai_1 _25301_ (.B1(_04218_),
    .Y(_05279_),
    .A1(net290),
    .A2(net27));
 sg13g2_nand2_1 _25302_ (.Y(_05280_),
    .A(_05190_),
    .B(_05196_));
 sg13g2_o21ai_1 _25303_ (.B1(_05280_),
    .Y(_05281_),
    .A1(_04262_),
    .A2(_05136_));
 sg13g2_o21ai_1 _25304_ (.B1(_05281_),
    .Y(_05282_),
    .A1(_05190_),
    .A2(_05196_));
 sg13g2_buf_1 _25305_ (.A(_05282_),
    .X(_05283_));
 sg13g2_nand2b_1 _25306_ (.Y(_05284_),
    .B(_05283_),
    .A_N(_05271_));
 sg13g2_and2_1 _25307_ (.A(_05126_),
    .B(_05272_),
    .X(_05285_));
 sg13g2_buf_1 _25308_ (.A(_05285_),
    .X(_05286_));
 sg13g2_nand2_1 _25309_ (.Y(_05287_),
    .A(_05271_),
    .B(_05286_));
 sg13g2_mux2_1 _25310_ (.A0(_05284_),
    .A1(_05287_),
    .S(_05105_),
    .X(_05288_));
 sg13g2_inv_1 _25311_ (.Y(_05289_),
    .A(_05283_));
 sg13g2_nor2_1 _25312_ (.A(_05284_),
    .B(_05286_),
    .Y(_05290_));
 sg13g2_a21oi_1 _25313_ (.A1(_05271_),
    .A2(_05289_),
    .Y(_05291_),
    .B1(_05290_));
 sg13g2_nand2_2 _25314_ (.Y(_05292_),
    .A(net296),
    .B(_02569_));
 sg13g2_a21oi_1 _25315_ (.A1(_05288_),
    .A2(_05291_),
    .Y(_05293_),
    .B1(_05292_));
 sg13g2_a21oi_1 _25316_ (.A1(net316),
    .A2(_05279_),
    .Y(_05294_),
    .B1(_05293_));
 sg13g2_nor3_1 _25317_ (.A(net299),
    .B(net298),
    .C(_05294_),
    .Y(_05295_));
 sg13g2_a21o_1 _25318_ (.A2(_05262_),
    .A1(net299),
    .B1(_05295_),
    .X(_05296_));
 sg13g2_xnor2_1 _25319_ (.Y(_05297_),
    .A(_05149_),
    .B(_05020_));
 sg13g2_o21ai_1 _25320_ (.B1(_05144_),
    .Y(_05298_),
    .A1(_05031_),
    .A2(_05035_));
 sg13g2_a21o_1 _25321_ (.A2(_05298_),
    .A1(_05247_),
    .B1(_04965_),
    .X(_05299_));
 sg13g2_o21ai_1 _25322_ (.B1(_05299_),
    .Y(_05300_),
    .A1(_05247_),
    .A2(_04919_));
 sg13g2_xnor2_1 _25323_ (.Y(_05301_),
    .A(_05297_),
    .B(_05300_));
 sg13g2_nor2_1 _25324_ (.A(net305),
    .B(_02569_),
    .Y(_05302_));
 sg13g2_a22oi_1 _25325_ (.Y(_05303_),
    .B1(_05301_),
    .B2(_05302_),
    .A2(_05236_),
    .A1(_02538_));
 sg13g2_nand3_1 _25326_ (.B(net241),
    .C(_05303_),
    .A(net297),
    .Y(_05304_));
 sg13g2_nor2_1 _25327_ (.A(net304),
    .B(_05304_),
    .Y(_05305_));
 sg13g2_buf_1 _25328_ (.A(_02660_),
    .X(_05306_));
 sg13g2_buf_1 _25329_ (.A(_02377_),
    .X(_05307_));
 sg13g2_a21oi_1 _25330_ (.A1(_05105_),
    .A2(_05286_),
    .Y(_05308_),
    .B1(_05289_));
 sg13g2_xnor2_1 _25331_ (.Y(_05309_),
    .A(_05271_),
    .B(_05308_));
 sg13g2_nand2_1 _25332_ (.Y(_05310_),
    .A(net303),
    .B(_04100_));
 sg13g2_nor2_1 _25333_ (.A(_05310_),
    .B(_05186_),
    .Y(_05311_));
 sg13g2_a21oi_1 _25334_ (.A1(net295),
    .A2(_05309_),
    .Y(_05312_),
    .B1(_05311_));
 sg13g2_nor4_1 _25335_ (.A(net309),
    .B(net299),
    .C(_02373_),
    .D(_05312_),
    .Y(_05313_));
 sg13g2_a21oi_1 _25336_ (.A1(_02382_),
    .A2(net27),
    .Y(_05314_),
    .B1(_05292_));
 sg13g2_xor2_1 _25337_ (.B(_05105_),
    .A(_05126_),
    .X(_05315_));
 sg13g2_nand2_1 _25338_ (.Y(_05316_),
    .A(net305),
    .B(_05241_));
 sg13g2_nand2b_1 _25339_ (.Y(_05317_),
    .B(_02409_),
    .A_N(_05256_));
 sg13g2_nand2b_1 _25340_ (.Y(_05318_),
    .B(net241),
    .A_N(_05235_));
 sg13g2_mux4_1 _25341_ (.S0(net316),
    .A0(_05315_),
    .A1(_05316_),
    .A2(_05317_),
    .A3(_05318_),
    .S1(_05189_),
    .X(_05319_));
 sg13g2_mux2_1 _25342_ (.A0(_05314_),
    .A1(_05319_),
    .S(_02367_),
    .X(_05320_));
 sg13g2_nor2_1 _25343_ (.A(net289),
    .B(_05320_),
    .Y(_05321_));
 sg13g2_nand2_1 _25344_ (.Y(_05322_),
    .A(net290),
    .B(_05226_));
 sg13g2_o21ai_1 _25345_ (.B1(_05322_),
    .Y(_05323_),
    .A1(net290),
    .A2(_05139_));
 sg13g2_nor2_1 _25346_ (.A(_02524_),
    .B(_05323_),
    .Y(_05324_));
 sg13g2_or4_1 _25347_ (.A(_05305_),
    .B(_05313_),
    .C(_05321_),
    .D(_05324_),
    .X(_05325_));
 sg13g2_a21oi_1 _25348_ (.A1(net296),
    .A2(_05318_),
    .Y(_05326_),
    .B1(net316));
 sg13g2_nand2_1 _25349_ (.Y(_05327_),
    .A(_05139_),
    .B(_05326_));
 sg13g2_nand2_1 _25350_ (.Y(_05328_),
    .A(_02377_),
    .B(_02660_));
 sg13g2_nor2_1 _25351_ (.A(_05315_),
    .B(_05328_),
    .Y(_05329_));
 sg13g2_a221oi_1 _25352_ (.B2(net296),
    .C1(_05329_),
    .B1(_05326_),
    .A1(net316),
    .Y(_05330_),
    .A2(_05311_));
 sg13g2_and2_1 _25353_ (.A(_05327_),
    .B(_05330_),
    .X(_05331_));
 sg13g2_buf_1 _25354_ (.A(_05331_),
    .X(_05332_));
 sg13g2_nor2_2 _25355_ (.A(net304),
    .B(net289),
    .Y(_05333_));
 sg13g2_nand2_1 _25356_ (.Y(_05334_),
    .A(net295),
    .B(_05309_));
 sg13g2_a21oi_1 _25357_ (.A1(net290),
    .A2(net27),
    .Y(_05335_),
    .B1(net310));
 sg13g2_nand2_1 _25358_ (.Y(_05336_),
    .A(_05184_),
    .B(_05212_));
 sg13g2_a21oi_1 _25359_ (.A1(_05223_),
    .A2(_05336_),
    .Y(_05337_),
    .B1(_05221_));
 sg13g2_and3_1 _25360_ (.X(_05338_),
    .A(_05169_),
    .B(_05177_),
    .C(_05272_));
 sg13g2_nor3_1 _25361_ (.A(_05292_),
    .B(_05337_),
    .C(_05338_),
    .Y(_05339_));
 sg13g2_a21o_1 _25362_ (.A2(_05335_),
    .A1(_05334_),
    .B1(_05339_),
    .X(_05340_));
 sg13g2_nor2_2 _25363_ (.A(net299),
    .B(_02372_),
    .Y(_05341_));
 sg13g2_nor2_1 _25364_ (.A(net330),
    .B(_02364_),
    .Y(_05342_));
 sg13g2_nand2b_1 _25365_ (.Y(_05343_),
    .B(net403),
    .A_N(_02260_));
 sg13g2_nor2_1 _25366_ (.A(_05310_),
    .B(_05256_),
    .Y(_05344_));
 sg13g2_a21oi_1 _25367_ (.A1(net305),
    .A2(_05237_),
    .Y(_05345_),
    .B1(_05344_));
 sg13g2_xnor2_1 _25368_ (.Y(_05346_),
    .A(_05088_),
    .B(_05240_));
 sg13g2_nor2_1 _25369_ (.A(_05140_),
    .B(_05346_),
    .Y(_05347_));
 sg13g2_nor3_1 _25370_ (.A(net305),
    .B(_02407_),
    .C(_05301_),
    .Y(_05348_));
 sg13g2_o21ai_1 _25371_ (.B1(_05230_),
    .Y(_05349_),
    .A1(_05347_),
    .A2(_05348_));
 sg13g2_o21ai_1 _25372_ (.B1(_05349_),
    .Y(_05350_),
    .A1(net315),
    .A2(_05345_));
 sg13g2_buf_1 _25373_ (.A(_05350_),
    .X(_05351_));
 sg13g2_a21oi_1 _25374_ (.A1(_05342_),
    .A2(_05343_),
    .Y(_05352_),
    .B1(_05351_));
 sg13g2_a221oi_1 _25375_ (.B2(_05341_),
    .C1(_05352_),
    .B1(_05340_),
    .A1(_05332_),
    .Y(_05353_),
    .A2(_05333_));
 sg13g2_buf_1 _25376_ (.A(_05353_),
    .X(_05354_));
 sg13g2_or2_1 _25377_ (.X(_05355_),
    .B(_02364_),
    .A(net330));
 sg13g2_mux4_1 _25378_ (.S0(_05230_),
    .A0(_05235_),
    .A1(_05186_),
    .A2(_05315_),
    .A3(_05346_),
    .S1(_05189_),
    .X(_05356_));
 sg13g2_nand2_1 _25379_ (.Y(_05357_),
    .A(_02409_),
    .B(_05139_));
 sg13g2_a21oi_1 _25380_ (.A1(net295),
    .A2(net27),
    .Y(_05358_),
    .B1(net316));
 sg13g2_nand2_1 _25381_ (.Y(_05359_),
    .A(_05271_),
    .B(_05283_));
 sg13g2_nor2_1 _25382_ (.A(_05286_),
    .B(_05359_),
    .Y(_05360_));
 sg13g2_nor2_1 _25383_ (.A(_05271_),
    .B(_05283_),
    .Y(_05361_));
 sg13g2_o21ai_1 _25384_ (.B1(net303),
    .Y(_05362_),
    .A1(_05360_),
    .A2(_05361_));
 sg13g2_o21ai_1 _25385_ (.B1(_05362_),
    .Y(_05363_),
    .A1(net296),
    .A2(_05226_));
 sg13g2_nand3_1 _25386_ (.B(_05126_),
    .C(_05273_),
    .A(_02518_),
    .Y(_05364_));
 sg13g2_nand3_1 _25387_ (.B(_05271_),
    .C(_05283_),
    .A(_02518_),
    .Y(_05365_));
 sg13g2_nor2b_1 _25388_ (.A(_05105_),
    .B_N(_05365_),
    .Y(_05366_));
 sg13g2_a21oi_1 _25389_ (.A1(_05105_),
    .A2(_05364_),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_nor3_1 _25390_ (.A(net315),
    .B(_05363_),
    .C(_05367_),
    .Y(_05368_));
 sg13g2_a21o_1 _25391_ (.A2(_05358_),
    .A1(_05357_),
    .B1(_05368_),
    .X(_05369_));
 sg13g2_buf_1 _25392_ (.A(_05369_),
    .X(_05370_));
 sg13g2_nor2b_1 _25393_ (.A(_05343_),
    .B_N(_05356_),
    .Y(_05371_));
 sg13g2_a221oi_1 _25394_ (.B2(_05333_),
    .C1(_05371_),
    .B1(_05370_),
    .A1(_05355_),
    .Y(_05372_),
    .A2(_05356_));
 sg13g2_nand3_1 _25395_ (.B(_05354_),
    .C(_05372_),
    .A(_05325_),
    .Y(_05373_));
 sg13g2_nand3_1 _25396_ (.B(net465),
    .C(net453),
    .A(_02318_),
    .Y(_05374_));
 sg13g2_o21ai_1 _25397_ (.B1(net325),
    .Y(_05375_),
    .A1(_02324_),
    .A2(_05374_));
 sg13g2_buf_1 _25398_ (.A(_05375_),
    .X(_05376_));
 sg13g2_nand2b_1 _25399_ (.Y(_05377_),
    .B(_05307_),
    .A_N(_05186_));
 sg13g2_and2_1 _25400_ (.A(net315),
    .B(_05377_),
    .X(_05378_));
 sg13g2_a21o_1 _25401_ (.A2(_05378_),
    .A1(_05357_),
    .B1(_05368_),
    .X(_05379_));
 sg13g2_buf_1 _25402_ (.A(_05379_),
    .X(_05380_));
 sg13g2_nand2b_1 _25403_ (.Y(_05381_),
    .B(net295),
    .A_N(_05235_));
 sg13g2_o21ai_1 _25404_ (.B1(_05381_),
    .Y(_05382_),
    .A1(net295),
    .A2(_05315_));
 sg13g2_nor2_1 _25405_ (.A(net305),
    .B(_05241_),
    .Y(_05383_));
 sg13g2_a21oi_1 _25406_ (.A1(_05307_),
    .A2(_05256_),
    .Y(_05384_),
    .B1(_05383_));
 sg13g2_mux2_1 _25407_ (.A0(_05382_),
    .A1(_05384_),
    .S(_05231_),
    .X(_05385_));
 sg13g2_nand2_1 _25408_ (.Y(_05386_),
    .A(net305),
    .B(_05301_));
 sg13g2_o21ai_1 _25409_ (.B1(_05386_),
    .Y(_05387_),
    .A1(net305),
    .A2(_05237_));
 sg13g2_a21o_1 _25410_ (.A2(_05387_),
    .A1(net316),
    .B1(net230),
    .X(_05388_));
 sg13g2_nor3_1 _25411_ (.A(_02514_),
    .B(_02370_),
    .C(net27),
    .Y(_05389_));
 sg13g2_a21oi_1 _25412_ (.A1(_02469_),
    .A2(_05388_),
    .Y(_05390_),
    .B1(_05389_));
 sg13g2_o21ai_1 _25413_ (.B1(_05390_),
    .Y(_05391_),
    .A1(_02643_),
    .A2(_05385_));
 sg13g2_a21o_1 _25414_ (.A2(_05380_),
    .A1(_02459_),
    .B1(_05391_),
    .X(_05392_));
 sg13g2_buf_1 _25415_ (.A(_05392_),
    .X(_05393_));
 sg13g2_nand2_1 _25416_ (.Y(_05394_),
    .A(_02367_),
    .B(_02372_));
 sg13g2_nor2_1 _25417_ (.A(net290),
    .B(net315),
    .Y(_05395_));
 sg13g2_a22oi_1 _25418_ (.Y(_05396_),
    .B1(_05395_),
    .B2(_05139_),
    .A2(_05309_),
    .A1(_02538_));
 sg13g2_nor2b_1 _25419_ (.A(_05226_),
    .B_N(_05302_),
    .Y(_05397_));
 sg13g2_a21oi_1 _25420_ (.A1(net315),
    .A2(_05311_),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nand2_1 _25421_ (.Y(_05399_),
    .A(_05396_),
    .B(_05398_));
 sg13g2_nand2_1 _25422_ (.Y(_05400_),
    .A(net289),
    .B(_05320_));
 sg13g2_o21ai_1 _25423_ (.B1(_05400_),
    .Y(_05401_),
    .A1(_05394_),
    .A2(_05399_));
 sg13g2_or2_1 _25424_ (.X(_05402_),
    .B(_05401_),
    .A(_05393_));
 sg13g2_nor4_1 _25425_ (.A(_05296_),
    .B(_05373_),
    .C(_05376_),
    .D(_05402_),
    .Y(_05403_));
 sg13g2_nand2_1 _25426_ (.Y(_05404_),
    .A(net241),
    .B(_05303_));
 sg13g2_and4_1 _25427_ (.A(_02260_),
    .B(_02373_),
    .C(_05396_),
    .D(_05398_),
    .X(_05405_));
 sg13g2_a221oi_1 _25428_ (.B2(_05404_),
    .C1(_05405_),
    .B1(_05333_),
    .A1(_05341_),
    .Y(_05406_),
    .A2(_05319_));
 sg13g2_nor2_1 _25429_ (.A(_02409_),
    .B(_05257_),
    .Y(_05407_));
 sg13g2_nor2_1 _25430_ (.A(net230),
    .B(_05301_),
    .Y(_05408_));
 sg13g2_a221oi_1 _25431_ (.B2(net295),
    .C1(net315),
    .B1(_05408_),
    .A1(_05237_),
    .Y(_05409_),
    .A2(_02409_));
 sg13g2_a21oi_1 _25432_ (.A1(net315),
    .A2(_05407_),
    .Y(_05410_),
    .B1(_05409_));
 sg13g2_a21oi_1 _25433_ (.A1(net289),
    .A2(_05410_),
    .Y(_05411_),
    .B1(net299));
 sg13g2_o21ai_1 _25434_ (.B1(_05411_),
    .Y(_05412_),
    .A1(net289),
    .A2(_05356_));
 sg13g2_o21ai_1 _25435_ (.B1(net304),
    .Y(_05413_),
    .A1(_05234_),
    .A2(_05319_));
 sg13g2_nand2b_1 _25436_ (.Y(_05414_),
    .B(_05351_),
    .A_N(_05304_));
 sg13g2_nand2b_1 _25437_ (.Y(_05415_),
    .B(_05414_),
    .A_N(_05413_));
 sg13g2_and2_1 _25438_ (.A(_05412_),
    .B(_05415_),
    .X(_05416_));
 sg13g2_nand2_1 _25439_ (.Y(_05417_),
    .A(net290),
    .B(net27));
 sg13g2_and3_1 _25440_ (.X(_05418_),
    .A(net309),
    .B(_02630_),
    .C(_05417_));
 sg13g2_nand2_1 _25441_ (.Y(_05419_),
    .A(_02630_),
    .B(_05339_));
 sg13g2_o21ai_1 _25442_ (.B1(_05419_),
    .Y(_05420_),
    .A1(_05351_),
    .A2(_05394_));
 sg13g2_a221oi_1 _25443_ (.B2(_05334_),
    .C1(_05420_),
    .B1(_05418_),
    .A1(_05341_),
    .Y(_05421_),
    .A2(_05332_));
 sg13g2_a21oi_1 _25444_ (.A1(_02630_),
    .A2(_05332_),
    .Y(_05422_),
    .B1(_05376_));
 sg13g2_nand4_1 _25445_ (.B(_05416_),
    .C(_05421_),
    .A(_05406_),
    .Y(_05423_),
    .D(_05422_));
 sg13g2_buf_1 _25446_ (.A(_05423_),
    .X(_05424_));
 sg13g2_nand2_1 _25447_ (.Y(_05425_),
    .A(net304),
    .B(_05260_));
 sg13g2_nor2_1 _25448_ (.A(_02370_),
    .B(_05408_),
    .Y(_05426_));
 sg13g2_a22oi_1 _25449_ (.Y(_05427_),
    .B1(_05333_),
    .B2(_05426_),
    .A2(_05260_),
    .A1(_05341_));
 sg13g2_o21ai_1 _25450_ (.B1(_05427_),
    .Y(_05428_),
    .A1(_05233_),
    .A2(_05425_));
 sg13g2_nand3_1 _25451_ (.B(net298),
    .C(_05370_),
    .A(_02260_),
    .Y(_05429_));
 sg13g2_inv_1 _25452_ (.Y(_05430_),
    .A(_05410_));
 sg13g2_a22oi_1 _25453_ (.Y(_05431_),
    .B1(_05430_),
    .B2(_05333_),
    .A2(_05356_),
    .A1(_05341_));
 sg13g2_nand3b_1 _25454_ (.B(_05429_),
    .C(_05431_),
    .Y(_05432_),
    .A_N(_05428_));
 sg13g2_buf_1 _25455_ (.A(_05432_),
    .X(_05433_));
 sg13g2_mux2_1 _25456_ (.A0(_05233_),
    .A1(_05294_),
    .S(net298),
    .X(_05434_));
 sg13g2_nor2_1 _25457_ (.A(net298),
    .B(_05426_),
    .Y(_05435_));
 sg13g2_a21oi_1 _25458_ (.A1(net298),
    .A2(_05259_),
    .Y(_05436_),
    .B1(_05435_));
 sg13g2_nand2_1 _25459_ (.Y(_05437_),
    .A(net299),
    .B(_05436_));
 sg13g2_o21ai_1 _25460_ (.B1(_05437_),
    .Y(_05438_),
    .A1(net299),
    .A2(_05434_));
 sg13g2_nor3_1 _25461_ (.A(_05424_),
    .B(_05433_),
    .C(_05438_),
    .Y(_05439_));
 sg13g2_a21oi_1 _25462_ (.A1(net241),
    .A2(net27),
    .Y(_05440_),
    .B1(_05292_));
 sg13g2_nor2b_1 _25463_ (.A(_05440_),
    .B_N(_05294_),
    .Y(_05441_));
 sg13g2_a21oi_1 _25464_ (.A1(_05292_),
    .A2(_05328_),
    .Y(_05442_),
    .B1(_04218_));
 sg13g2_nor2_1 _25465_ (.A(net289),
    .B(_05442_),
    .Y(_05443_));
 sg13g2_a21oi_1 _25466_ (.A1(_05334_),
    .A2(_05335_),
    .Y(_05444_),
    .B1(_05339_));
 sg13g2_and4_1 _25467_ (.A(net289),
    .B(_05444_),
    .C(_05399_),
    .D(_05441_),
    .X(_05445_));
 sg13g2_nor2b_1 _25468_ (.A(_05370_),
    .B_N(_05233_),
    .Y(_05446_));
 sg13g2_a221oi_1 _25469_ (.B2(_05446_),
    .C1(net304),
    .B1(_05445_),
    .A1(_05441_),
    .Y(_05447_),
    .A2(_05443_));
 sg13g2_o21ai_1 _25470_ (.B1(_05447_),
    .Y(_05448_),
    .A1(_05424_),
    .A2(_05433_));
 sg13g2_a22oi_1 _25471_ (.Y(_05449_),
    .B1(_05448_),
    .B2(net241),
    .A2(_05439_),
    .A1(_05403_));
 sg13g2_nand2_1 _25472_ (.Y(_05450_),
    .A(_02254_),
    .B(_05449_));
 sg13g2_inv_1 _25473_ (.Y(_05451_),
    .A(_08644_));
 sg13g2_buf_1 _25474_ (.A(_05451_),
    .X(_05452_));
 sg13g2_a21oi_1 _25475_ (.A1(net325),
    .A2(_05393_),
    .Y(_05453_),
    .B1(net689));
 sg13g2_buf_1 _25476_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-11] ),
    .X(_05454_));
 sg13g2_o21ai_1 _25477_ (.B1(net608),
    .Y(_05455_),
    .A1(net724),
    .A2(_05454_));
 sg13g2_a21oi_1 _25478_ (.A1(_05450_),
    .A2(_05453_),
    .Y(_01598_),
    .B1(_05455_));
 sg13g2_buf_1 _25479_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-1] ),
    .X(_05456_));
 sg13g2_nand2_1 _25480_ (.Y(_05457_),
    .A(_05452_),
    .B(_05456_));
 sg13g2_nor3_1 _25481_ (.A(net309),
    .B(_05363_),
    .C(_05367_),
    .Y(_05458_));
 sg13g2_a21o_1 _25482_ (.A2(_05279_),
    .A1(net309),
    .B1(_05458_),
    .X(_05459_));
 sg13g2_a21oi_1 _25483_ (.A1(net317),
    .A2(_05459_),
    .Y(_05460_),
    .B1(net230));
 sg13g2_o21ai_1 _25484_ (.B1(net325),
    .Y(_05461_),
    .A1(_02437_),
    .A2(_05460_));
 sg13g2_nand2_1 _25485_ (.Y(_05462_),
    .A(net788),
    .B(_05461_));
 sg13g2_nand2_1 _25486_ (.Y(_05463_),
    .A(_08644_),
    .B(_02254_));
 sg13g2_nor2_1 _25487_ (.A(_05449_),
    .B(_05463_),
    .Y(_05464_));
 sg13g2_buf_1 _25488_ (.A(_05464_),
    .X(_05465_));
 sg13g2_inv_1 _25489_ (.Y(_05466_),
    .A(_05428_));
 sg13g2_a221oi_1 _25490_ (.B2(_05466_),
    .C1(net635),
    .B1(net26),
    .A1(_05457_),
    .Y(_01599_),
    .A2(_05462_));
 sg13g2_nor2_1 _25491_ (.A(net689),
    .B(net331),
    .Y(_05467_));
 sg13g2_buf_2 _25492_ (.A(_05467_),
    .X(_05468_));
 sg13g2_a22oi_1 _25493_ (.Y(_05469_),
    .B1(_05309_),
    .B2(net295),
    .A2(net27),
    .A1(_02409_));
 sg13g2_a21o_1 _25494_ (.A2(_05469_),
    .A1(_02596_),
    .B1(net230),
    .X(_05470_));
 sg13g2_nand2_1 _25495_ (.Y(_05471_),
    .A(net318),
    .B(_05470_));
 sg13g2_buf_1 _25496_ (.A(_08645_),
    .X(_05472_));
 sg13g2_buf_1 _25497_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[0] ),
    .X(_05473_));
 sg13g2_o21ai_1 _25498_ (.B1(net610),
    .Y(_05474_),
    .A1(_05472_),
    .A2(_05473_));
 sg13g2_a221oi_1 _25499_ (.B2(_05471_),
    .C1(_05474_),
    .B1(_05468_),
    .A1(_05406_),
    .Y(_01600_),
    .A2(net26));
 sg13g2_nand2_1 _25500_ (.Y(_05475_),
    .A(_05429_),
    .B(_05431_));
 sg13g2_inv_1 _25501_ (.Y(_05476_),
    .A(_05475_));
 sg13g2_buf_1 _25502_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[1] ),
    .X(_05477_));
 sg13g2_nand2_1 _25503_ (.Y(_05478_),
    .A(_05452_),
    .B(_05477_));
 sg13g2_o21ai_1 _25504_ (.B1(_03998_),
    .Y(_05479_),
    .A1(net290),
    .A2(_05278_));
 sg13g2_a21oi_1 _25505_ (.A1(_02596_),
    .A2(_05479_),
    .Y(_05480_),
    .B1(net230));
 sg13g2_o21ai_1 _25506_ (.B1(net325),
    .Y(_05481_),
    .A1(_02437_),
    .A2(_05480_));
 sg13g2_nand2_1 _25507_ (.Y(_05482_),
    .A(net688),
    .B(_05481_));
 sg13g2_a221oi_1 _25508_ (.B2(_05482_),
    .C1(_11527_),
    .B1(_05478_),
    .A1(_05476_),
    .Y(_01601_),
    .A2(net26));
 sg13g2_or2_1 _25509_ (.X(_05483_),
    .B(_05433_),
    .A(_05424_));
 sg13g2_a22oi_1 _25510_ (.Y(_05484_),
    .B1(_05403_),
    .B2(_05439_),
    .A2(_05376_),
    .A1(net241));
 sg13g2_a21oi_1 _25511_ (.A1(_05483_),
    .A2(_05447_),
    .Y(_05485_),
    .B1(_05484_));
 sg13g2_buf_1 _25512_ (.A(_05485_),
    .X(_05486_));
 sg13g2_and2_1 _25513_ (.A(net788),
    .B(_05421_),
    .X(_05487_));
 sg13g2_buf_1 _25514_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[2] ),
    .X(_05488_));
 sg13g2_nor2_1 _25515_ (.A(_08411_),
    .B(_05468_),
    .Y(_05489_));
 sg13g2_buf_2 _25516_ (.A(_05489_),
    .X(_05490_));
 sg13g2_o21ai_1 _25517_ (.B1(_05490_),
    .Y(_05491_),
    .A1(net724),
    .A2(_05488_));
 sg13g2_a21oi_1 _25518_ (.A1(net25),
    .A2(_05487_),
    .Y(_01602_),
    .B1(_05491_));
 sg13g2_nor2_1 _25519_ (.A(net689),
    .B(_05438_),
    .Y(_05492_));
 sg13g2_buf_1 _25520_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[3] ),
    .X(_05493_));
 sg13g2_o21ai_1 _25521_ (.B1(_05490_),
    .Y(_05494_),
    .A1(net724),
    .A2(_05493_));
 sg13g2_a21oi_1 _25522_ (.A1(net25),
    .A2(_05492_),
    .Y(_01603_),
    .B1(_05494_));
 sg13g2_and2_1 _25523_ (.A(net788),
    .B(_05325_),
    .X(_05495_));
 sg13g2_buf_1 _25524_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[4] ),
    .X(_05496_));
 sg13g2_o21ai_1 _25525_ (.B1(_05490_),
    .Y(_05497_),
    .A1(net724),
    .A2(_05496_));
 sg13g2_a21oi_1 _25526_ (.A1(net25),
    .A2(_05495_),
    .Y(_01604_),
    .B1(_05497_));
 sg13g2_nor2_1 _25527_ (.A(net689),
    .B(_05393_),
    .Y(_05498_));
 sg13g2_buf_1 _25528_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[5] ),
    .X(_05499_));
 sg13g2_o21ai_1 _25529_ (.B1(_05490_),
    .Y(_05500_),
    .A1(net724),
    .A2(_05499_));
 sg13g2_a21oi_1 _25530_ (.A1(_05486_),
    .A2(_05498_),
    .Y(_01605_),
    .B1(_05500_));
 sg13g2_and2_1 _25531_ (.A(net788),
    .B(_05354_),
    .X(_05501_));
 sg13g2_buf_1 _25532_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[6] ),
    .X(_05502_));
 sg13g2_o21ai_1 _25533_ (.B1(_05490_),
    .Y(_05503_),
    .A1(net724),
    .A2(_05502_));
 sg13g2_a21oi_1 _25534_ (.A1(net25),
    .A2(_05501_),
    .Y(_01606_),
    .B1(_05503_));
 sg13g2_nor2_1 _25535_ (.A(net689),
    .B(_05296_),
    .Y(_05504_));
 sg13g2_buf_1 _25536_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[7] ),
    .X(_05505_));
 sg13g2_o21ai_1 _25537_ (.B1(_05490_),
    .Y(_05506_),
    .A1(_08646_),
    .A2(_05505_));
 sg13g2_a21oi_1 _25538_ (.A1(net25),
    .A2(_05504_),
    .Y(_01607_),
    .B1(_05506_));
 sg13g2_nor2_1 _25539_ (.A(net689),
    .B(_05401_),
    .Y(_05507_));
 sg13g2_buf_1 _25540_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[8] ),
    .X(_05508_));
 sg13g2_o21ai_1 _25541_ (.B1(_05490_),
    .Y(_05509_),
    .A1(_08646_),
    .A2(_05508_));
 sg13g2_a21oi_1 _25542_ (.A1(net25),
    .A2(_05507_),
    .Y(_01608_),
    .B1(_05509_));
 sg13g2_o21ai_1 _25543_ (.B1(net788),
    .Y(_05510_),
    .A1(_05354_),
    .A2(_05376_));
 sg13g2_inv_1 _25544_ (.Y(_05511_),
    .A(_05510_));
 sg13g2_buf_1 _25545_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-10] ),
    .X(_05512_));
 sg13g2_o21ai_1 _25546_ (.B1(net608),
    .Y(_05513_),
    .A1(net724),
    .A2(_05512_));
 sg13g2_a21oi_1 _25547_ (.A1(_05450_),
    .A2(_05511_),
    .Y(_01609_),
    .B1(_05513_));
 sg13g2_and2_1 _25548_ (.A(net788),
    .B(_05372_),
    .X(_05514_));
 sg13g2_buf_1 _25549_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[9] ),
    .X(_05515_));
 sg13g2_o21ai_1 _25550_ (.B1(_05490_),
    .Y(_05516_),
    .A1(net688),
    .A2(_05515_));
 sg13g2_a21oi_1 _25551_ (.A1(_05486_),
    .A2(_05514_),
    .Y(_01610_),
    .B1(_05516_));
 sg13g2_nor2b_1 _25552_ (.A(_05342_),
    .B_N(_05332_),
    .Y(_05517_));
 sg13g2_a21oi_1 _25553_ (.A1(_02381_),
    .A2(_05340_),
    .Y(_05518_),
    .B1(_05517_));
 sg13g2_or3_1 _25554_ (.A(_05449_),
    .B(_05463_),
    .C(_05518_),
    .X(_05519_));
 sg13g2_buf_1 _25555_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[10] ),
    .X(_05520_));
 sg13g2_nand2_1 _25556_ (.Y(_05521_),
    .A(net689),
    .B(_05520_));
 sg13g2_a21oi_1 _25557_ (.A1(_05519_),
    .A2(_05521_),
    .Y(_01611_),
    .B1(net562));
 sg13g2_nand2_1 _25558_ (.Y(_05522_),
    .A(_08644_),
    .B(net325));
 sg13g2_and2_1 _25559_ (.A(net310),
    .B(_05382_),
    .X(_05523_));
 sg13g2_a21oi_1 _25560_ (.A1(net309),
    .A2(_05188_),
    .Y(_05524_),
    .B1(_05523_));
 sg13g2_o21ai_1 _25561_ (.B1(net310),
    .Y(_05525_),
    .A1(net230),
    .A2(_05387_));
 sg13g2_o21ai_1 _25562_ (.B1(_05525_),
    .Y(_05526_),
    .A1(_05231_),
    .A2(_05384_));
 sg13g2_a22oi_1 _25563_ (.Y(_05527_),
    .B1(_05526_),
    .B2(net360),
    .A2(_05524_),
    .A1(net312));
 sg13g2_o21ai_1 _25564_ (.B1(_05527_),
    .Y(_05528_),
    .A1(net318),
    .A2(_05460_));
 sg13g2_nor2_1 _25565_ (.A(_05522_),
    .B(_05528_),
    .Y(_05529_));
 sg13g2_buf_1 _25566_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-9] ),
    .X(_05530_));
 sg13g2_o21ai_1 _25567_ (.B1(_09043_),
    .Y(_05531_),
    .A1(net688),
    .A2(_05530_));
 sg13g2_nor3_1 _25568_ (.A(net26),
    .B(_05529_),
    .C(_05531_),
    .Y(_01612_));
 sg13g2_a21oi_1 _25569_ (.A1(_02630_),
    .A2(_05404_),
    .Y(_05532_),
    .B1(_05463_));
 sg13g2_o21ai_1 _25570_ (.B1(_05316_),
    .Y(_05533_),
    .A1(_05235_),
    .A2(_05310_));
 sg13g2_nand2_1 _25571_ (.Y(_05534_),
    .A(net310),
    .B(_05345_));
 sg13g2_o21ai_1 _25572_ (.B1(_05534_),
    .Y(_05535_),
    .A1(net310),
    .A2(_05533_));
 sg13g2_a21oi_1 _25573_ (.A1(net360),
    .A2(_05535_),
    .Y(_05536_),
    .B1(_05522_));
 sg13g2_a21o_1 _25574_ (.A2(_05227_),
    .A1(net295),
    .B1(_05311_),
    .X(_05537_));
 sg13g2_inv_1 _25575_ (.Y(_05538_),
    .A(_05537_));
 sg13g2_and2_1 _25576_ (.A(net309),
    .B(_05323_),
    .X(_05539_));
 sg13g2_a21oi_1 _25577_ (.A1(net310),
    .A2(_05538_),
    .Y(_05540_),
    .B1(_05539_));
 sg13g2_inv_1 _25578_ (.Y(_05541_),
    .A(_05540_));
 sg13g2_a22oi_1 _25579_ (.Y(_05542_),
    .B1(_05541_),
    .B2(net312),
    .A2(_05470_),
    .A1(_02437_));
 sg13g2_buf_1 _25580_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-8] ),
    .X(_05543_));
 sg13g2_o21ai_1 _25581_ (.B1(net610),
    .Y(_05544_),
    .A1(_05472_),
    .A2(_05543_));
 sg13g2_a221oi_1 _25582_ (.B2(_05542_),
    .C1(_05544_),
    .B1(_05536_),
    .A1(net25),
    .Y(_01613_),
    .A2(_05532_));
 sg13g2_nor2_1 _25583_ (.A(_02479_),
    .B(_05480_),
    .Y(_05545_));
 sg13g2_o21ai_1 _25584_ (.B1(_05468_),
    .Y(_05546_),
    .A1(_02355_),
    .A2(_05385_));
 sg13g2_nor2_1 _25585_ (.A(_05545_),
    .B(_05546_),
    .Y(_05547_));
 sg13g2_nand2_1 _25586_ (.Y(_05548_),
    .A(net312),
    .B(_05380_));
 sg13g2_a21oi_1 _25587_ (.A1(_02630_),
    .A2(_05430_),
    .Y(_05549_),
    .B1(_05463_));
 sg13g2_buf_1 _25588_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-7] ),
    .X(_05550_));
 sg13g2_o21ai_1 _25589_ (.B1(net610),
    .Y(_05551_),
    .A1(net688),
    .A2(_05550_));
 sg13g2_a221oi_1 _25590_ (.B2(net25),
    .C1(_05551_),
    .B1(_05549_),
    .A1(_05547_),
    .Y(_01614_),
    .A2(_05548_));
 sg13g2_nand2_1 _25591_ (.Y(_05552_),
    .A(net309),
    .B(_05538_));
 sg13g2_o21ai_1 _25592_ (.B1(_05552_),
    .Y(_05553_),
    .A1(net309),
    .A2(_05533_));
 sg13g2_a21oi_1 _25593_ (.A1(net360),
    .A2(_05553_),
    .Y(_05554_),
    .B1(_05522_));
 sg13g2_mux2_1 _25594_ (.A0(_05323_),
    .A1(_05469_),
    .S(_05306_),
    .X(_05555_));
 sg13g2_nand2_1 _25595_ (.Y(_05556_),
    .A(_02422_),
    .B(_05555_));
 sg13g2_or3_1 _25596_ (.A(net299),
    .B(_05234_),
    .C(_05351_),
    .X(_05557_));
 sg13g2_buf_1 _25597_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-6] ),
    .X(_05558_));
 sg13g2_o21ai_1 _25598_ (.B1(net610),
    .Y(_05559_),
    .A1(net688),
    .A2(_05558_));
 sg13g2_a221oi_1 _25599_ (.B2(net26),
    .C1(_05559_),
    .B1(_05557_),
    .A1(_05554_),
    .Y(_01615_),
    .A2(_05556_));
 sg13g2_a22oi_1 _25600_ (.Y(_05560_),
    .B1(_05524_),
    .B2(net360),
    .A2(_05459_),
    .A1(_02422_));
 sg13g2_nand2_1 _25601_ (.Y(_05561_),
    .A(net304),
    .B(_05436_));
 sg13g2_buf_1 _25602_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-5] ),
    .X(_05562_));
 sg13g2_o21ai_1 _25603_ (.B1(net610),
    .Y(_05563_),
    .A1(net688),
    .A2(_05562_));
 sg13g2_a221oi_1 _25604_ (.B2(net26),
    .C1(_05563_),
    .B1(_05561_),
    .A1(_05468_),
    .Y(_01616_),
    .A2(_05560_));
 sg13g2_nor2_1 _25605_ (.A(_05306_),
    .B(_02643_),
    .Y(_05564_));
 sg13g2_a21oi_1 _25606_ (.A1(_05564_),
    .A2(_05469_),
    .Y(_05565_),
    .B1(_05522_));
 sg13g2_nand2_1 _25607_ (.Y(_05566_),
    .A(_02469_),
    .B(_05541_));
 sg13g2_nand2b_1 _25608_ (.Y(_05567_),
    .B(_05304_),
    .A_N(_05413_));
 sg13g2_buf_1 _25609_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-4] ),
    .X(_05568_));
 sg13g2_o21ai_1 _25610_ (.B1(net610),
    .Y(_05569_),
    .A1(net688),
    .A2(_05568_));
 sg13g2_a221oi_1 _25611_ (.B2(_05465_),
    .C1(_05569_),
    .B1(_05567_),
    .A1(_05565_),
    .Y(_01617_),
    .A2(_05566_));
 sg13g2_nand2_1 _25612_ (.Y(_05570_),
    .A(net317),
    .B(_05380_));
 sg13g2_nand3b_1 _25613_ (.B(net310),
    .C(_05279_),
    .Y(_05571_),
    .A_N(_02565_));
 sg13g2_a21o_1 _25614_ (.A2(_05571_),
    .A1(_05570_),
    .B1(_02437_),
    .X(_05572_));
 sg13g2_buf_1 _25615_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-3] ),
    .X(_05573_));
 sg13g2_o21ai_1 _25616_ (.B1(_08641_),
    .Y(_05574_),
    .A1(net688),
    .A2(_05573_));
 sg13g2_a221oi_1 _25617_ (.B2(_05572_),
    .C1(_05574_),
    .B1(_05468_),
    .A1(_05412_),
    .Y(_01618_),
    .A2(net26));
 sg13g2_nor2_1 _25618_ (.A(net298),
    .B(_05351_),
    .Y(_05575_));
 sg13g2_a21oi_1 _25619_ (.A1(net298),
    .A2(_05332_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_nand2b_1 _25620_ (.Y(_05577_),
    .B(net304),
    .A_N(_05576_));
 sg13g2_a21oi_1 _25621_ (.A1(_02565_),
    .A2(_05555_),
    .Y(_05578_),
    .B1(net230));
 sg13g2_or2_1 _25622_ (.X(_05579_),
    .B(_05578_),
    .A(_02437_));
 sg13g2_buf_1 _25623_ (.A(\rbzero.wall_tracer.rcp_fsm.o_data[-2] ),
    .X(_05580_));
 sg13g2_o21ai_1 _25624_ (.B1(_08641_),
    .Y(_05581_),
    .A1(_08645_),
    .A2(_05580_));
 sg13g2_a221oi_1 _25625_ (.B2(_05468_),
    .C1(_05581_),
    .B1(_05579_),
    .A1(net26),
    .Y(_01619_),
    .A2(_05577_));
 sg13g2_and2_1 _25626_ (.A(net832),
    .B(_08643_),
    .X(_05582_));
 sg13g2_buf_1 _25627_ (.A(_05582_),
    .X(_05583_));
 sg13g2_buf_1 _25628_ (.A(_05583_),
    .X(_05584_));
 sg13g2_inv_1 _25629_ (.Y(_05585_),
    .A(_08643_));
 sg13g2_o21ai_1 _25630_ (.B1(net788),
    .Y(_05586_),
    .A1(net832),
    .A2(_05585_));
 sg13g2_a221oi_1 _25631_ (.B2(_08434_),
    .C1(_11527_),
    .B1(_05586_),
    .A1(net689),
    .Y(_01620_),
    .A2(_05584_));
 sg13g2_nand2_1 _25632_ (.Y(_05587_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-11] ),
    .B(net623));
 sg13g2_nand2_1 _25633_ (.Y(_05588_),
    .A(net806),
    .B(net681));
 sg13g2_a21oi_1 _25634_ (.A1(_05587_),
    .A2(_05588_),
    .Y(_01621_),
    .B1(net562));
 sg13g2_nand2_1 _25635_ (.Y(_05589_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-1] ),
    .B(net623));
 sg13g2_nand2_1 _25636_ (.Y(_05590_),
    .A(_02139_),
    .B(net681));
 sg13g2_a21oi_1 _25637_ (.A1(_05589_),
    .A2(_05590_),
    .Y(_01622_),
    .B1(net562));
 sg13g2_nand2_1 _25638_ (.Y(_05591_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[0] ),
    .B(net623));
 sg13g2_nand2_1 _25639_ (.Y(_05592_),
    .A(_02140_),
    .B(net681));
 sg13g2_a21oi_1 _25640_ (.A1(_05591_),
    .A2(_05592_),
    .Y(_01623_),
    .B1(net562));
 sg13g2_nand2_1 _25641_ (.Y(_05593_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[1] ),
    .B(net623));
 sg13g2_nand2_1 _25642_ (.Y(_05594_),
    .A(net733),
    .B(net681));
 sg13g2_a21oi_1 _25643_ (.A1(_05593_),
    .A2(_05594_),
    .Y(_01624_),
    .B1(_01989_));
 sg13g2_nand2_1 _25644_ (.Y(_05595_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[2] ),
    .B(net623));
 sg13g2_nand2_1 _25645_ (.Y(_05596_),
    .A(_02144_),
    .B(_08692_));
 sg13g2_a21oi_1 _25646_ (.A1(_05595_),
    .A2(_05596_),
    .Y(_01625_),
    .B1(_01989_));
 sg13g2_nand2_1 _25647_ (.Y(_05597_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[3] ),
    .B(net623));
 sg13g2_nand2_1 _25648_ (.Y(_05598_),
    .A(net805),
    .B(net681));
 sg13g2_buf_1 _25649_ (.A(_11764_),
    .X(_05599_));
 sg13g2_a21oi_1 _25650_ (.A1(_05597_),
    .A2(_05598_),
    .Y(_01626_),
    .B1(net560));
 sg13g2_nand2_1 _25651_ (.Y(_05600_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[4] ),
    .B(net623));
 sg13g2_nand2_1 _25652_ (.Y(_05601_),
    .A(_02195_),
    .B(net681));
 sg13g2_a21oi_1 _25653_ (.A1(_05600_),
    .A2(_05601_),
    .Y(_01627_),
    .B1(net560));
 sg13g2_nand2_1 _25654_ (.Y(_05602_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[5] ),
    .B(_05584_));
 sg13g2_nand2_1 _25655_ (.Y(_05603_),
    .A(net732),
    .B(net681));
 sg13g2_a21oi_1 _25656_ (.A1(_05602_),
    .A2(_05603_),
    .Y(_01628_),
    .B1(net560));
 sg13g2_nand2_1 _25657_ (.Y(_05604_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[6] ),
    .B(net623));
 sg13g2_nand2_1 _25658_ (.Y(_05605_),
    .A(net802),
    .B(net681));
 sg13g2_a21oi_1 _25659_ (.A1(_05604_),
    .A2(_05605_),
    .Y(_01629_),
    .B1(net560));
 sg13g2_buf_1 _25660_ (.A(_05583_),
    .X(_05606_));
 sg13g2_nand2_1 _25661_ (.Y(_05607_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[7] ),
    .B(net622));
 sg13g2_buf_1 _25662_ (.A(_08691_),
    .X(_05608_));
 sg13g2_nand2_1 _25663_ (.Y(_05609_),
    .A(_02219_),
    .B(net621));
 sg13g2_a21oi_1 _25664_ (.A1(_05607_),
    .A2(_05609_),
    .Y(_01630_),
    .B1(_05599_));
 sg13g2_nand2_1 _25665_ (.Y(_05610_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[8] ),
    .B(net622));
 sg13g2_nand2_1 _25666_ (.Y(_05611_),
    .A(_02220_),
    .B(net621));
 sg13g2_a21oi_1 _25667_ (.A1(_05610_),
    .A2(_05611_),
    .Y(_01631_),
    .B1(net560));
 sg13g2_nand2_1 _25668_ (.Y(_05612_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-10] ),
    .B(net622));
 sg13g2_nand2_1 _25669_ (.Y(_05613_),
    .A(_02014_),
    .B(net621));
 sg13g2_a21oi_1 _25670_ (.A1(_05612_),
    .A2(_05613_),
    .Y(_01632_),
    .B1(net560));
 sg13g2_nand2_1 _25671_ (.Y(_05614_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[9] ),
    .B(net622));
 sg13g2_nand2_1 _25672_ (.Y(_05615_),
    .A(_02236_),
    .B(net621));
 sg13g2_a21oi_1 _25673_ (.A1(_05614_),
    .A2(_05615_),
    .Y(_01633_),
    .B1(_05599_));
 sg13g2_nand2_1 _25674_ (.Y(_05616_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[10] ),
    .B(_05606_));
 sg13g2_nand2_1 _25675_ (.Y(_05617_),
    .A(net561),
    .B(_05608_));
 sg13g2_a21oi_1 _25676_ (.A1(_05616_),
    .A2(_05617_),
    .Y(_01634_),
    .B1(net560));
 sg13g2_nand2_1 _25677_ (.Y(_05618_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-9] ),
    .B(_05606_));
 sg13g2_nand2_1 _25678_ (.Y(_05619_),
    .A(_02015_),
    .B(_05608_));
 sg13g2_a21oi_1 _25679_ (.A1(_05618_),
    .A2(_05619_),
    .Y(_01635_),
    .B1(net560));
 sg13g2_nand2_1 _25680_ (.Y(_05620_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-8] ),
    .B(net622));
 sg13g2_nand2_1 _25681_ (.Y(_05621_),
    .A(_02016_),
    .B(net621));
 sg13g2_buf_1 _25682_ (.A(_11764_),
    .X(_05622_));
 sg13g2_a21oi_1 _25683_ (.A1(_05620_),
    .A2(_05621_),
    .Y(_01636_),
    .B1(net559));
 sg13g2_nand2_1 _25684_ (.Y(_05623_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-7] ),
    .B(net622));
 sg13g2_nand2_1 _25685_ (.Y(_05624_),
    .A(_02064_),
    .B(net621));
 sg13g2_a21oi_1 _25686_ (.A1(_05623_),
    .A2(_05624_),
    .Y(_01637_),
    .B1(net559));
 sg13g2_nand2_1 _25687_ (.Y(_05625_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-6] ),
    .B(net622));
 sg13g2_nand2_1 _25688_ (.Y(_05626_),
    .A(_02035_),
    .B(net621));
 sg13g2_a21oi_1 _25689_ (.A1(_05625_),
    .A2(_05626_),
    .Y(_01638_),
    .B1(net559));
 sg13g2_nand2_1 _25690_ (.Y(_05627_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-5] ),
    .B(net622));
 sg13g2_nand2_1 _25691_ (.Y(_05628_),
    .A(_02021_),
    .B(net621));
 sg13g2_a21oi_1 _25692_ (.A1(_05627_),
    .A2(_05628_),
    .Y(_01639_),
    .B1(net559));
 sg13g2_nand2_1 _25693_ (.Y(_05629_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-4] ),
    .B(_05583_));
 sg13g2_nand2_1 _25694_ (.Y(_05630_),
    .A(net807),
    .B(_08691_));
 sg13g2_a21oi_1 _25695_ (.A1(_05629_),
    .A2(_05630_),
    .Y(_01640_),
    .B1(net559));
 sg13g2_nand2_1 _25696_ (.Y(_05631_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-3] ),
    .B(_05583_));
 sg13g2_nand2_1 _25697_ (.Y(_05632_),
    .A(net737),
    .B(_08691_));
 sg13g2_a21oi_1 _25698_ (.A1(_05631_),
    .A2(_05632_),
    .Y(_01641_),
    .B1(net559));
 sg13g2_nand2_1 _25699_ (.Y(_05633_),
    .A(\rbzero.wall_tracer.rcp_fsm.i_data[-2] ),
    .B(_05583_));
 sg13g2_nand2_1 _25700_ (.Y(_05634_),
    .A(_02009_),
    .B(_08691_));
 sg13g2_a21oi_1 _25701_ (.A1(_05633_),
    .A2(_05634_),
    .Y(_01642_),
    .B1(net559));
 sg13g2_o21ai_1 _25702_ (.B1(_08422_),
    .Y(_05635_),
    .A1(_08423_),
    .A2(net832));
 sg13g2_nor3_1 _25703_ (.A(_08431_),
    .B(\rbzero.wall_tracer.state[0] ),
    .C(_08669_),
    .Y(_05636_));
 sg13g2_a21o_1 _25704_ (.A2(_05635_),
    .A1(_08431_),
    .B1(_05636_),
    .X(_05637_));
 sg13g2_buf_1 _25705_ (.A(_05637_),
    .X(_05638_));
 sg13g2_buf_1 _25706_ (.A(_05638_),
    .X(_05639_));
 sg13g2_a22oi_1 _25707_ (.Y(_05640_),
    .B1(_09115_),
    .B2(net799),
    .A2(_08669_),
    .A1(_11846_));
 sg13g2_nor2_1 _25708_ (.A(_08431_),
    .B(_08669_),
    .Y(_05641_));
 sg13g2_buf_1 _25709_ (.A(_05641_),
    .X(_05642_));
 sg13g2_nand2_1 _25710_ (.Y(_05643_),
    .A(_08781_),
    .B(_05642_));
 sg13g2_a21oi_1 _25711_ (.A1(_05640_),
    .A2(_05643_),
    .Y(_05644_),
    .B1(_05638_));
 sg13g2_a21oi_1 _25712_ (.A1(\rbzero.wall_tracer.rcp_fsm.i_data[-11] ),
    .A2(net558),
    .Y(_05645_),
    .B1(_05644_));
 sg13g2_nor2_1 _25713_ (.A(net634),
    .B(_05645_),
    .Y(_01643_));
 sg13g2_buf_1 _25714_ (.A(_08669_),
    .X(_05646_));
 sg13g2_a221oi_1 _25715_ (.B2(net727),
    .C1(net558),
    .B1(_11570_),
    .A1(_08533_),
    .Y(_05647_),
    .A2(net731));
 sg13g2_buf_1 _25716_ (.A(_05642_),
    .X(_05648_));
 sg13g2_nand2_1 _25717_ (.Y(_05649_),
    .A(_11400_),
    .B(net620));
 sg13g2_a21oi_1 _25718_ (.A1(_08431_),
    .A2(_05635_),
    .Y(_05650_),
    .B1(_05636_));
 sg13g2_buf_1 _25719_ (.A(_05650_),
    .X(_05651_));
 sg13g2_buf_1 _25720_ (.A(_05651_),
    .X(_05652_));
 sg13g2_o21ai_1 _25721_ (.B1(net608),
    .Y(_05653_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-1] ),
    .A2(net557));
 sg13g2_a21oi_1 _25722_ (.A1(_05647_),
    .A2(_05649_),
    .Y(_01644_),
    .B1(_05653_));
 sg13g2_a221oi_1 _25723_ (.B2(_08433_),
    .C1(net558),
    .B1(_11849_),
    .A1(_08532_),
    .Y(_05654_),
    .A2(net731));
 sg13g2_nand2_1 _25724_ (.Y(_05655_),
    .A(_11850_),
    .B(_05648_));
 sg13g2_o21ai_1 _25725_ (.B1(_09078_),
    .Y(_05656_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[0] ),
    .A2(net557));
 sg13g2_a21oi_1 _25726_ (.A1(_05654_),
    .A2(_05655_),
    .Y(_01645_),
    .B1(_05656_));
 sg13g2_nor2b_1 _25727_ (.A(_12098_),
    .B_N(net799),
    .Y(_05657_));
 sg13g2_a21oi_1 _25728_ (.A1(_08538_),
    .A2(_08669_),
    .Y(_05658_),
    .B1(_05638_));
 sg13g2_nor2b_1 _25729_ (.A(_05657_),
    .B_N(_05658_),
    .Y(_05659_));
 sg13g2_nand2_1 _25730_ (.Y(_05660_),
    .A(_12100_),
    .B(_05648_));
 sg13g2_o21ai_1 _25731_ (.B1(_09078_),
    .Y(_05661_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[1] ),
    .A2(net557));
 sg13g2_a21oi_1 _25732_ (.A1(_05659_),
    .A2(_05660_),
    .Y(_01646_),
    .B1(_05661_));
 sg13g2_nand2_1 _25733_ (.Y(_05662_),
    .A(net727),
    .B(_12599_));
 sg13g2_a221oi_1 _25734_ (.B2(net620),
    .C1(_05638_),
    .B1(_12602_),
    .A1(_08537_),
    .Y(_05663_),
    .A2(_05646_));
 sg13g2_buf_1 _25735_ (.A(_08640_),
    .X(_05664_));
 sg13g2_o21ai_1 _25736_ (.B1(net556),
    .Y(_05665_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[2] ),
    .A2(net557));
 sg13g2_a21oi_1 _25737_ (.A1(_05662_),
    .A2(_05663_),
    .Y(_01647_),
    .B1(_05665_));
 sg13g2_a221oi_1 _25738_ (.B2(_12696_),
    .C1(_05638_),
    .B1(_05642_),
    .A1(net799),
    .Y(_05666_),
    .A2(_12693_));
 sg13g2_buf_2 _25739_ (.A(_05666_),
    .X(_05667_));
 sg13g2_nand2_1 _25740_ (.Y(_05668_),
    .A(_08536_),
    .B(net784));
 sg13g2_o21ai_1 _25741_ (.B1(net556),
    .Y(_05669_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[3] ),
    .A2(net557));
 sg13g2_a21oi_1 _25742_ (.A1(_05667_),
    .A2(_05668_),
    .Y(_01648_),
    .B1(_05669_));
 sg13g2_nand2_1 _25743_ (.Y(_05670_),
    .A(_08535_),
    .B(net784));
 sg13g2_o21ai_1 _25744_ (.B1(net556),
    .Y(_05671_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[4] ),
    .A2(net557));
 sg13g2_a21oi_1 _25745_ (.A1(_05667_),
    .A2(_05670_),
    .Y(_01649_),
    .B1(_05671_));
 sg13g2_nand2_1 _25746_ (.Y(_05672_),
    .A(_08547_),
    .B(net784));
 sg13g2_o21ai_1 _25747_ (.B1(net556),
    .Y(_05673_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[5] ),
    .A2(net557));
 sg13g2_a21oi_1 _25748_ (.A1(_05667_),
    .A2(_05672_),
    .Y(_01650_),
    .B1(_05673_));
 sg13g2_nand2_1 _25749_ (.Y(_05674_),
    .A(_08546_),
    .B(net784));
 sg13g2_o21ai_1 _25750_ (.B1(net556),
    .Y(_05675_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[6] ),
    .A2(_05652_));
 sg13g2_a21oi_1 _25751_ (.A1(_05667_),
    .A2(_05674_),
    .Y(_01651_),
    .B1(_05675_));
 sg13g2_nand2_1 _25752_ (.Y(_05676_),
    .A(_08545_),
    .B(net784));
 sg13g2_o21ai_1 _25753_ (.B1(net556),
    .Y(_05677_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[7] ),
    .A2(_05652_));
 sg13g2_a21oi_1 _25754_ (.A1(_05667_),
    .A2(_05676_),
    .Y(_01652_),
    .B1(_05677_));
 sg13g2_nand2_1 _25755_ (.Y(_05678_),
    .A(_08542_),
    .B(_08670_));
 sg13g2_buf_1 _25756_ (.A(_05651_),
    .X(_05679_));
 sg13g2_o21ai_1 _25757_ (.B1(_05664_),
    .Y(_05680_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[8] ),
    .A2(net555));
 sg13g2_a21oi_1 _25758_ (.A1(_05667_),
    .A2(_05678_),
    .Y(_01653_),
    .B1(_05680_));
 sg13g2_a22oi_1 _25759_ (.Y(_05681_),
    .B1(_09118_),
    .B2(net799),
    .A2(_08669_),
    .A1(_11796_));
 sg13g2_nand2_1 _25760_ (.Y(_05682_),
    .A(_08784_),
    .B(_05642_));
 sg13g2_a21oi_1 _25761_ (.A1(_05681_),
    .A2(_05682_),
    .Y(_05683_),
    .B1(_05638_));
 sg13g2_a21oi_1 _25762_ (.A1(\rbzero.wall_tracer.rcp_fsm.i_data[-10] ),
    .A2(net558),
    .Y(_05684_),
    .B1(_05683_));
 sg13g2_nor2_1 _25763_ (.A(_11690_),
    .B(_05684_),
    .Y(_01654_));
 sg13g2_nand2_1 _25764_ (.Y(_05685_),
    .A(_08543_),
    .B(_08670_));
 sg13g2_o21ai_1 _25765_ (.B1(_05664_),
    .Y(_05686_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[9] ),
    .A2(_05679_));
 sg13g2_a21oi_1 _25766_ (.A1(_05667_),
    .A2(_05685_),
    .Y(_01655_),
    .B1(_05686_));
 sg13g2_nand2_1 _25767_ (.Y(_05687_),
    .A(_08481_),
    .B(net784));
 sg13g2_o21ai_1 _25768_ (.B1(net556),
    .Y(_05688_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[10] ),
    .A2(_05679_));
 sg13g2_a21oi_1 _25769_ (.A1(_05667_),
    .A2(_05687_),
    .Y(_01656_),
    .B1(_05688_));
 sg13g2_nor2b_1 _25770_ (.A(_11423_),
    .B_N(_05642_),
    .Y(_05689_));
 sg13g2_a221oi_1 _25771_ (.B2(net799),
    .C1(_05689_),
    .B1(_11599_),
    .A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .Y(_05690_),
    .A2(net731));
 sg13g2_o21ai_1 _25772_ (.B1(net556),
    .Y(_05691_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-9] ),
    .A2(net555));
 sg13g2_a21oi_1 _25773_ (.A1(net557),
    .A2(_05690_),
    .Y(_01657_),
    .B1(_05691_));
 sg13g2_a21oi_1 _25774_ (.A1(\rbzero.wall_tracer.visualWallDist[-8] ),
    .A2(net731),
    .Y(_05692_),
    .B1(net558));
 sg13g2_inv_1 _25775_ (.Y(_05693_),
    .A(_11422_));
 sg13g2_a22oi_1 _25776_ (.Y(_05694_),
    .B1(net620),
    .B2(_05693_),
    .A2(_11598_),
    .A1(net727));
 sg13g2_o21ai_1 _25777_ (.B1(_09043_),
    .Y(_05695_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-8] ),
    .A2(net555));
 sg13g2_a21oi_1 _25778_ (.A1(_05692_),
    .A2(_05694_),
    .Y(_01658_),
    .B1(_05695_));
 sg13g2_nand2b_1 _25779_ (.Y(_05696_),
    .B(net727),
    .A_N(_11595_));
 sg13g2_a221oi_1 _25780_ (.B2(_05642_),
    .C1(_05638_),
    .B1(_11916_),
    .A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .Y(_05697_),
    .A2(_08669_));
 sg13g2_o21ai_1 _25781_ (.B1(net609),
    .Y(_05698_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-7] ),
    .A2(net555));
 sg13g2_a21oi_1 _25782_ (.A1(_05696_),
    .A2(_05697_),
    .Y(_01659_),
    .B1(_05698_));
 sg13g2_a21oi_1 _25783_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_05646_),
    .Y(_05699_),
    .B1(_05639_));
 sg13g2_a22oi_1 _25784_ (.Y(_05700_),
    .B1(net620),
    .B2(_11416_),
    .A2(_11592_),
    .A1(net727));
 sg13g2_o21ai_1 _25785_ (.B1(net609),
    .Y(_05701_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-6] ),
    .A2(net555));
 sg13g2_a21oi_1 _25786_ (.A1(_05699_),
    .A2(_05700_),
    .Y(_01660_),
    .B1(_05701_));
 sg13g2_a21oi_1 _25787_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(net731),
    .Y(_05702_),
    .B1(_05639_));
 sg13g2_a22oi_1 _25788_ (.Y(_05703_),
    .B1(net620),
    .B2(_11413_),
    .A2(_11589_),
    .A1(net727));
 sg13g2_o21ai_1 _25789_ (.B1(net609),
    .Y(_05704_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-5] ),
    .A2(net555));
 sg13g2_a21oi_1 _25790_ (.A1(_05702_),
    .A2(_05703_),
    .Y(_01661_),
    .B1(_05704_));
 sg13g2_a21oi_1 _25791_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(net731),
    .Y(_05705_),
    .B1(net558));
 sg13g2_a22oi_1 _25792_ (.Y(_05706_),
    .B1(net620),
    .B2(_11410_),
    .A2(_11587_),
    .A1(net727));
 sg13g2_o21ai_1 _25793_ (.B1(net609),
    .Y(_05707_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-4] ),
    .A2(net555));
 sg13g2_a21oi_1 _25794_ (.A1(_05705_),
    .A2(_05706_),
    .Y(_01662_),
    .B1(_05707_));
 sg13g2_a221oi_1 _25795_ (.B2(net727),
    .C1(net558),
    .B1(_11785_),
    .A1(_08541_),
    .Y(_05708_),
    .A2(net731));
 sg13g2_nand2b_1 _25796_ (.Y(_05709_),
    .B(net620),
    .A_N(_11405_));
 sg13g2_o21ai_1 _25797_ (.B1(net609),
    .Y(_05710_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-3] ),
    .A2(net555));
 sg13g2_a21oi_1 _25798_ (.A1(_05708_),
    .A2(_05709_),
    .Y(_01663_),
    .B1(_05710_));
 sg13g2_a221oi_1 _25799_ (.B2(net799),
    .C1(net558),
    .B1(_11581_),
    .A1(_08540_),
    .Y(_05711_),
    .A2(net731));
 sg13g2_nand2b_1 _25800_ (.Y(_05712_),
    .B(net620),
    .A_N(_11402_));
 sg13g2_o21ai_1 _25801_ (.B1(net609),
    .Y(_05713_),
    .A1(\rbzero.wall_tracer.rcp_fsm.i_data[-2] ),
    .A2(_05651_));
 sg13g2_a21oi_1 _25802_ (.A1(_05711_),
    .A2(_05712_),
    .Y(_01664_),
    .B1(_05713_));
 sg13g2_nor2_1 _25803_ (.A(\rbzero.wall_tracer.state[0] ),
    .B(net784),
    .Y(_05714_));
 sg13g2_nor2_1 _25804_ (.A(net685),
    .B(net611),
    .Y(_05715_));
 sg13g2_buf_1 _25805_ (.A(_05715_),
    .X(_05716_));
 sg13g2_nor2_1 _25806_ (.A(_08434_),
    .B(net832),
    .Y(_05717_));
 sg13g2_mux2_1 _25807_ (.A0(net832),
    .A1(_05717_),
    .S(_08432_),
    .X(_05718_));
 sg13g2_nand2_1 _25808_ (.Y(_05719_),
    .A(_05716_),
    .B(_05718_));
 sg13g2_a21oi_1 _25809_ (.A1(_05714_),
    .A2(_05719_),
    .Y(_01665_),
    .B1(net559));
 sg13g2_buf_1 _25810_ (.A(_11325_),
    .X(_05720_));
 sg13g2_buf_1 _25811_ (.A(_11322_),
    .X(_05721_));
 sg13g2_buf_1 _25812_ (.A(_05721_),
    .X(_05722_));
 sg13g2_nor2_1 _25813_ (.A(net73),
    .B(_11325_),
    .Y(_05723_));
 sg13g2_a21oi_1 _25814_ (.A1(net573),
    .A2(_05720_),
    .Y(_05724_),
    .B1(_05723_));
 sg13g2_nor2_1 _25815_ (.A(net634),
    .B(_05724_),
    .Y(_01666_));
 sg13g2_nand2_1 _25816_ (.Y(_05725_),
    .A(_05454_),
    .B(net492));
 sg13g2_nand2_1 _25817_ (.Y(_05726_),
    .A(net685),
    .B(_08425_));
 sg13g2_buf_1 _25818_ (.A(_05726_),
    .X(_05727_));
 sg13g2_buf_1 _25819_ (.A(net516),
    .X(_05728_));
 sg13g2_nand2_1 _25820_ (.Y(_05729_),
    .A(\rbzero.wall_tracer.size_full[-11] ),
    .B(net496));
 sg13g2_a21oi_1 _25821_ (.A1(_05725_),
    .A2(_05729_),
    .Y(_01667_),
    .B1(_05622_));
 sg13g2_nand2_1 _25822_ (.Y(_05730_),
    .A(_05456_),
    .B(net492));
 sg13g2_nand2_1 _25823_ (.Y(_05731_),
    .A(_11752_),
    .B(net496));
 sg13g2_a21oi_1 _25824_ (.A1(_05730_),
    .A2(_05731_),
    .Y(_01668_),
    .B1(_05622_));
 sg13g2_nand2_1 _25825_ (.Y(_05732_),
    .A(_05473_),
    .B(_08429_));
 sg13g2_nand2_1 _25826_ (.Y(_05733_),
    .A(_11756_),
    .B(_05728_));
 sg13g2_buf_1 _25827_ (.A(_08746_),
    .X(_05734_));
 sg13g2_buf_1 _25828_ (.A(_05734_),
    .X(_05735_));
 sg13g2_a21oi_1 _25829_ (.A1(_05732_),
    .A2(_05733_),
    .Y(_01669_),
    .B1(net554));
 sg13g2_nand2_1 _25830_ (.Y(_05736_),
    .A(_05477_),
    .B(net492));
 sg13g2_nand2_1 _25831_ (.Y(_05737_),
    .A(_11760_),
    .B(_05728_));
 sg13g2_a21oi_1 _25832_ (.A1(_05736_),
    .A2(_05737_),
    .Y(_01670_),
    .B1(net554));
 sg13g2_nand2_1 _25833_ (.Y(_05738_),
    .A(_05488_),
    .B(net492));
 sg13g2_buf_1 _25834_ (.A(_05727_),
    .X(_05739_));
 sg13g2_nand2_1 _25835_ (.Y(_05740_),
    .A(_11727_),
    .B(net495));
 sg13g2_a21oi_1 _25836_ (.A1(_05738_),
    .A2(_05740_),
    .Y(_01671_),
    .B1(net554));
 sg13g2_nand2_1 _25837_ (.Y(_05741_),
    .A(_05493_),
    .B(net492));
 sg13g2_nand2_1 _25838_ (.Y(_05742_),
    .A(_12701_),
    .B(net495));
 sg13g2_a21oi_1 _25839_ (.A1(_05741_),
    .A2(_05742_),
    .Y(_01672_),
    .B1(net554));
 sg13g2_nand2_1 _25840_ (.Y(_05743_),
    .A(_05496_),
    .B(net492));
 sg13g2_nand2_1 _25841_ (.Y(_05744_),
    .A(_12797_),
    .B(net495));
 sg13g2_a21oi_1 _25842_ (.A1(_05743_),
    .A2(_05744_),
    .Y(_01673_),
    .B1(net554));
 sg13g2_nand2_1 _25843_ (.Y(_05745_),
    .A(_05499_),
    .B(net492));
 sg13g2_nand2_1 _25844_ (.Y(_05746_),
    .A(_12911_),
    .B(net495));
 sg13g2_a21oi_1 _25845_ (.A1(_05745_),
    .A2(_05746_),
    .Y(_01674_),
    .B1(net554));
 sg13g2_nand2_1 _25846_ (.Y(_05747_),
    .A(_05502_),
    .B(_08429_));
 sg13g2_nand2_1 _25847_ (.Y(_05748_),
    .A(_13033_),
    .B(net495));
 sg13g2_a21oi_1 _25848_ (.A1(_05747_),
    .A2(_05748_),
    .Y(_01675_),
    .B1(net554));
 sg13g2_buf_1 _25849_ (.A(_08427_),
    .X(_05749_));
 sg13g2_nand2_1 _25850_ (.Y(_05750_),
    .A(_05505_),
    .B(net494));
 sg13g2_nand2_1 _25851_ (.Y(_05751_),
    .A(_13182_),
    .B(net495));
 sg13g2_a21oi_1 _25852_ (.A1(_05750_),
    .A2(_05751_),
    .Y(_01676_),
    .B1(_05735_));
 sg13g2_nand2_1 _25853_ (.Y(_05752_),
    .A(_05508_),
    .B(net494));
 sg13g2_nand2_1 _25854_ (.Y(_05753_),
    .A(_13320_),
    .B(net495));
 sg13g2_a21oi_1 _25855_ (.A1(_05752_),
    .A2(_05753_),
    .Y(_01677_),
    .B1(_05735_));
 sg13g2_nand2_1 _25856_ (.Y(_05754_),
    .A(_05512_),
    .B(net494));
 sg13g2_nand2_1 _25857_ (.Y(_05755_),
    .A(\rbzero.wall_tracer.size_full[-10] ),
    .B(net495));
 sg13g2_a21oi_1 _25858_ (.A1(_05754_),
    .A2(_05755_),
    .Y(_01678_),
    .B1(net554));
 sg13g2_nand2_1 _25859_ (.Y(_05756_),
    .A(_05515_),
    .B(_05749_));
 sg13g2_nand2_1 _25860_ (.Y(_05757_),
    .A(\rbzero.wall_tracer.size_full[9] ),
    .B(_05739_));
 sg13g2_buf_1 _25861_ (.A(_05734_),
    .X(_05758_));
 sg13g2_a21oi_1 _25862_ (.A1(_05756_),
    .A2(_05757_),
    .Y(_01679_),
    .B1(_05758_));
 sg13g2_nand2_1 _25863_ (.Y(_05759_),
    .A(_05520_),
    .B(_05749_));
 sg13g2_nand2_1 _25864_ (.Y(_05760_),
    .A(\rbzero.wall_tracer.size_full[10] ),
    .B(_05739_));
 sg13g2_a21oi_1 _25865_ (.A1(_05759_),
    .A2(_05760_),
    .Y(_01680_),
    .B1(_05758_));
 sg13g2_nand2_1 _25866_ (.Y(_05761_),
    .A(_05530_),
    .B(net494));
 sg13g2_nand2_1 _25867_ (.Y(_05762_),
    .A(\rbzero.wall_tracer.size_full[-9] ),
    .B(_05727_));
 sg13g2_a21oi_1 _25868_ (.A1(_05761_),
    .A2(_05762_),
    .Y(_01681_),
    .B1(net553));
 sg13g2_nand2_1 _25869_ (.Y(_05763_),
    .A(_05543_),
    .B(net494));
 sg13g2_nand2_1 _25870_ (.Y(_05764_),
    .A(\rbzero.wall_tracer.size[0] ),
    .B(net516));
 sg13g2_a21oi_1 _25871_ (.A1(_05763_),
    .A2(_05764_),
    .Y(_01682_),
    .B1(net553));
 sg13g2_nand2_1 _25872_ (.Y(_05765_),
    .A(_05550_),
    .B(net494));
 sg13g2_nand2_1 _25873_ (.Y(_05766_),
    .A(\rbzero.wall_tracer.size[1] ),
    .B(net516));
 sg13g2_a21oi_1 _25874_ (.A1(_05765_),
    .A2(_05766_),
    .Y(_01683_),
    .B1(net553));
 sg13g2_nand2_1 _25875_ (.Y(_05767_),
    .A(_05558_),
    .B(net494));
 sg13g2_nand2_1 _25876_ (.Y(_05768_),
    .A(\rbzero.wall_tracer.size[2] ),
    .B(net516));
 sg13g2_a21oi_1 _25877_ (.A1(_05767_),
    .A2(_05768_),
    .Y(_01684_),
    .B1(net553));
 sg13g2_nand2_1 _25878_ (.Y(_05769_),
    .A(_05562_),
    .B(net494));
 sg13g2_nand2_1 _25879_ (.Y(_05770_),
    .A(\rbzero.wall_tracer.size[3] ),
    .B(net516));
 sg13g2_a21oi_1 _25880_ (.A1(_05769_),
    .A2(_05770_),
    .Y(_01685_),
    .B1(net553));
 sg13g2_nand2_1 _25881_ (.Y(_05771_),
    .A(_05568_),
    .B(net512));
 sg13g2_nand2_1 _25882_ (.Y(_05772_),
    .A(\rbzero.wall_tracer.size[4] ),
    .B(net516));
 sg13g2_a21oi_1 _25883_ (.A1(_05771_),
    .A2(_05772_),
    .Y(_01686_),
    .B1(net553));
 sg13g2_nand2_1 _25884_ (.Y(_05773_),
    .A(_05573_),
    .B(_08428_));
 sg13g2_nand2_1 _25885_ (.Y(_05774_),
    .A(\rbzero.wall_tracer.size[5] ),
    .B(net516));
 sg13g2_a21oi_1 _25886_ (.A1(_05773_),
    .A2(_05774_),
    .Y(_01687_),
    .B1(net553));
 sg13g2_nand2_1 _25887_ (.Y(_05775_),
    .A(_05580_),
    .B(_08428_));
 sg13g2_nand2_1 _25888_ (.Y(_05776_),
    .A(_11748_),
    .B(net516));
 sg13g2_a21oi_1 _25889_ (.A1(_05775_),
    .A2(_05776_),
    .Y(_01688_),
    .B1(net553));
 sg13g2_nand2_1 _25890_ (.Y(_05777_),
    .A(_05454_),
    .B(net546));
 sg13g2_nand2_1 _25891_ (.Y(_05778_),
    .A(net799),
    .B(_08425_));
 sg13g2_buf_1 _25892_ (.A(_05778_),
    .X(_05779_));
 sg13g2_buf_1 _25893_ (.A(_05779_),
    .X(_05780_));
 sg13g2_nand2_1 _25894_ (.Y(_05781_),
    .A(_12013_),
    .B(net515));
 sg13g2_buf_1 _25895_ (.A(_05734_),
    .X(_05782_));
 sg13g2_a21oi_1 _25896_ (.A1(_05777_),
    .A2(_05781_),
    .Y(_01689_),
    .B1(net552));
 sg13g2_nand2_1 _25897_ (.Y(_05783_),
    .A(_05456_),
    .B(_08635_));
 sg13g2_nand2_1 _25898_ (.Y(_05784_),
    .A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(net515));
 sg13g2_a21oi_1 _25899_ (.A1(_05783_),
    .A2(_05784_),
    .Y(_01690_),
    .B1(net552));
 sg13g2_nand2_1 _25900_ (.Y(_05785_),
    .A(_05473_),
    .B(_08635_));
 sg13g2_buf_1 _25901_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_05786_));
 sg13g2_nand2_1 _25902_ (.Y(_05787_),
    .A(_05786_),
    .B(net515));
 sg13g2_a21oi_1 _25903_ (.A1(_05785_),
    .A2(_05787_),
    .Y(_01691_),
    .B1(net552));
 sg13g2_nand2_1 _25904_ (.Y(_05788_),
    .A(_05477_),
    .B(net546));
 sg13g2_buf_1 _25905_ (.A(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_05789_));
 sg13g2_nand2_1 _25906_ (.Y(_05790_),
    .A(_05789_),
    .B(net515));
 sg13g2_a21oi_1 _25907_ (.A1(_05788_),
    .A2(_05790_),
    .Y(_01692_),
    .B1(net552));
 sg13g2_nand2_1 _25908_ (.Y(_05791_),
    .A(_05488_),
    .B(net546));
 sg13g2_buf_1 _25909_ (.A(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_05792_));
 sg13g2_nand2_1 _25910_ (.Y(_05793_),
    .A(_05792_),
    .B(net515));
 sg13g2_a21oi_1 _25911_ (.A1(_05791_),
    .A2(_05793_),
    .Y(_01693_),
    .B1(net552));
 sg13g2_nand2_1 _25912_ (.Y(_05794_),
    .A(_05493_),
    .B(net546));
 sg13g2_buf_1 _25913_ (.A(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_05795_));
 sg13g2_nand2_1 _25914_ (.Y(_05796_),
    .A(_05795_),
    .B(net515));
 sg13g2_a21oi_1 _25915_ (.A1(_05794_),
    .A2(_05796_),
    .Y(_01694_),
    .B1(net552));
 sg13g2_nand2_1 _25916_ (.Y(_05797_),
    .A(_05496_),
    .B(net546));
 sg13g2_buf_1 _25917_ (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_05798_));
 sg13g2_nand2_1 _25918_ (.Y(_05799_),
    .A(_05798_),
    .B(net515));
 sg13g2_a21oi_1 _25919_ (.A1(_05797_),
    .A2(_05799_),
    .Y(_01695_),
    .B1(net552));
 sg13g2_nand2_1 _25920_ (.Y(_05800_),
    .A(_05499_),
    .B(net546));
 sg13g2_buf_1 _25921_ (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_05801_));
 sg13g2_nand2_1 _25922_ (.Y(_05802_),
    .A(_05801_),
    .B(net515));
 sg13g2_a21oi_1 _25923_ (.A1(_05800_),
    .A2(_05802_),
    .Y(_01696_),
    .B1(net552));
 sg13g2_nand2_1 _25924_ (.Y(_05803_),
    .A(_05502_),
    .B(net546));
 sg13g2_buf_1 _25925_ (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .X(_05804_));
 sg13g2_nand2_1 _25926_ (.Y(_05805_),
    .A(_05804_),
    .B(_05780_));
 sg13g2_a21oi_1 _25927_ (.A1(_05803_),
    .A2(_05805_),
    .Y(_01697_),
    .B1(_05782_));
 sg13g2_buf_1 _25928_ (.A(_08634_),
    .X(_05806_));
 sg13g2_nand2_1 _25929_ (.Y(_05807_),
    .A(_05505_),
    .B(net514));
 sg13g2_buf_1 _25930_ (.A(\rbzero.wall_tracer.stepDistX[7] ),
    .X(_05808_));
 sg13g2_nand2_1 _25931_ (.Y(_05809_),
    .A(_05808_),
    .B(_05780_));
 sg13g2_a21oi_1 _25932_ (.A1(_05807_),
    .A2(_05809_),
    .Y(_01698_),
    .B1(_05782_));
 sg13g2_nand2_1 _25933_ (.Y(_05810_),
    .A(_05508_),
    .B(net514));
 sg13g2_buf_1 _25934_ (.A(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_05811_));
 sg13g2_buf_1 _25935_ (.A(_05779_),
    .X(_05812_));
 sg13g2_nand2_1 _25936_ (.Y(_05813_),
    .A(_05811_),
    .B(_05812_));
 sg13g2_buf_1 _25937_ (.A(_05734_),
    .X(_05814_));
 sg13g2_a21oi_1 _25938_ (.A1(_05810_),
    .A2(_05813_),
    .Y(_01699_),
    .B1(_05814_));
 sg13g2_nand2_1 _25939_ (.Y(_05815_),
    .A(_05512_),
    .B(net514));
 sg13g2_nand2_1 _25940_ (.Y(_05816_),
    .A(_12023_),
    .B(net513));
 sg13g2_a21oi_1 _25941_ (.A1(_05815_),
    .A2(_05816_),
    .Y(_01700_),
    .B1(net551));
 sg13g2_nand2_1 _25942_ (.Y(_05817_),
    .A(_05515_),
    .B(_05806_));
 sg13g2_buf_1 _25943_ (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_05818_));
 sg13g2_nand2_1 _25944_ (.Y(_05819_),
    .A(_05818_),
    .B(net513));
 sg13g2_a21oi_1 _25945_ (.A1(_05817_),
    .A2(_05819_),
    .Y(_01701_),
    .B1(_05814_));
 sg13g2_nand2_1 _25946_ (.Y(_05820_),
    .A(_05520_),
    .B(_05806_));
 sg13g2_nand2_1 _25947_ (.Y(_05821_),
    .A(\rbzero.wall_tracer.stepDistX[10] ),
    .B(_05812_));
 sg13g2_a21oi_1 _25948_ (.A1(_05820_),
    .A2(_05821_),
    .Y(_01702_),
    .B1(net551));
 sg13g2_nand2_1 _25949_ (.Y(_05822_),
    .A(_05530_),
    .B(net514));
 sg13g2_buf_1 _25950_ (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_05823_));
 sg13g2_nand2_1 _25951_ (.Y(_05824_),
    .A(_05823_),
    .B(net513));
 sg13g2_a21oi_1 _25952_ (.A1(_05822_),
    .A2(_05824_),
    .Y(_01703_),
    .B1(net551));
 sg13g2_nand2_1 _25953_ (.Y(_05825_),
    .A(_05543_),
    .B(net514));
 sg13g2_buf_1 _25954_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_05826_));
 sg13g2_nand2_1 _25955_ (.Y(_05827_),
    .A(_05826_),
    .B(net513));
 sg13g2_a21oi_1 _25956_ (.A1(_05825_),
    .A2(_05827_),
    .Y(_01704_),
    .B1(net551));
 sg13g2_nand2_1 _25957_ (.Y(_05828_),
    .A(_05550_),
    .B(net514));
 sg13g2_nand2_1 _25958_ (.Y(_05829_),
    .A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(net513));
 sg13g2_a21oi_1 _25959_ (.A1(_05828_),
    .A2(_05829_),
    .Y(_01705_),
    .B1(net551));
 sg13g2_nand2_1 _25960_ (.Y(_05830_),
    .A(_05558_),
    .B(net514));
 sg13g2_buf_1 _25961_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_05831_));
 sg13g2_nand2_1 _25962_ (.Y(_05832_),
    .A(_05831_),
    .B(net513));
 sg13g2_a21oi_1 _25963_ (.A1(_05830_),
    .A2(_05832_),
    .Y(_01706_),
    .B1(net551));
 sg13g2_nand2_1 _25964_ (.Y(_05833_),
    .A(_05562_),
    .B(net514));
 sg13g2_nand2_1 _25965_ (.Y(_05834_),
    .A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(net513));
 sg13g2_a21oi_1 _25966_ (.A1(_05833_),
    .A2(_05834_),
    .Y(_01707_),
    .B1(net551));
 sg13g2_nand2_1 _25967_ (.Y(_05835_),
    .A(_05568_),
    .B(_08634_));
 sg13g2_buf_1 _25968_ (.A(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_05836_));
 sg13g2_nand2_1 _25969_ (.Y(_05837_),
    .A(_05836_),
    .B(net513));
 sg13g2_a21oi_1 _25970_ (.A1(_05835_),
    .A2(_05837_),
    .Y(_01708_),
    .B1(net551));
 sg13g2_nand2_1 _25971_ (.Y(_05838_),
    .A(_05573_),
    .B(_08634_));
 sg13g2_buf_1 _25972_ (.A(\rbzero.wall_tracer.stepDistX[-3] ),
    .X(_05839_));
 sg13g2_nand2_1 _25973_ (.Y(_05840_),
    .A(_05839_),
    .B(_05779_));
 sg13g2_buf_1 _25974_ (.A(_05734_),
    .X(_05841_));
 sg13g2_a21oi_1 _25975_ (.A1(_05838_),
    .A2(_05840_),
    .Y(_01709_),
    .B1(net550));
 sg13g2_nand2_1 _25976_ (.Y(_05842_),
    .A(_05580_),
    .B(_08634_));
 sg13g2_buf_1 _25977_ (.A(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_05843_));
 sg13g2_nand2_1 _25978_ (.Y(_05844_),
    .A(_05843_),
    .B(_05779_));
 sg13g2_a21oi_1 _25979_ (.A1(_05842_),
    .A2(_05844_),
    .Y(_01710_),
    .B1(net550));
 sg13g2_nand2_1 _25980_ (.Y(_05845_),
    .A(_05454_),
    .B(net491));
 sg13g2_nand2_1 _25981_ (.Y(_05846_),
    .A(net611),
    .B(_08425_));
 sg13g2_buf_1 _25982_ (.A(_05846_),
    .X(_05847_));
 sg13g2_buf_1 _25983_ (.A(_05847_),
    .X(_05848_));
 sg13g2_nand2_1 _25984_ (.Y(_05849_),
    .A(_12018_),
    .B(net476));
 sg13g2_a21oi_1 _25985_ (.A1(_05845_),
    .A2(_05849_),
    .Y(_01711_),
    .B1(net550));
 sg13g2_nand2_1 _25986_ (.Y(_05850_),
    .A(_05456_),
    .B(net491));
 sg13g2_nand2_1 _25987_ (.Y(_05851_),
    .A(\rbzero.wall_tracer.stepDistY[-1] ),
    .B(net476));
 sg13g2_a21oi_1 _25988_ (.A1(_05850_),
    .A2(_05851_),
    .Y(_01712_),
    .B1(net550));
 sg13g2_nand2_1 _25989_ (.Y(_05852_),
    .A(_05473_),
    .B(net491));
 sg13g2_buf_1 _25990_ (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_05853_));
 sg13g2_nand2_1 _25991_ (.Y(_05854_),
    .A(_05853_),
    .B(net476));
 sg13g2_a21oi_1 _25992_ (.A1(_05852_),
    .A2(_05854_),
    .Y(_01713_),
    .B1(net550));
 sg13g2_nand2_1 _25993_ (.Y(_05855_),
    .A(_05477_),
    .B(net491));
 sg13g2_buf_1 _25994_ (.A(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_05856_));
 sg13g2_nand2_1 _25995_ (.Y(_05857_),
    .A(_05856_),
    .B(net476));
 sg13g2_a21oi_1 _25996_ (.A1(_05855_),
    .A2(_05857_),
    .Y(_01714_),
    .B1(net550));
 sg13g2_nand2_1 _25997_ (.Y(_05858_),
    .A(_05488_),
    .B(net491));
 sg13g2_buf_1 _25998_ (.A(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_05859_));
 sg13g2_nand2_1 _25999_ (.Y(_05860_),
    .A(_05859_),
    .B(net476));
 sg13g2_a21oi_1 _26000_ (.A1(_05858_),
    .A2(_05860_),
    .Y(_01715_),
    .B1(net550));
 sg13g2_nand2_1 _26001_ (.Y(_05861_),
    .A(_05493_),
    .B(net491));
 sg13g2_buf_1 _26002_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_05862_));
 sg13g2_nand2_1 _26003_ (.Y(_05863_),
    .A(_05862_),
    .B(net476));
 sg13g2_a21oi_1 _26004_ (.A1(_05861_),
    .A2(_05863_),
    .Y(_01716_),
    .B1(net550));
 sg13g2_nand2_1 _26005_ (.Y(_05864_),
    .A(_05496_),
    .B(net491));
 sg13g2_buf_1 _26006_ (.A(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_05865_));
 sg13g2_nand2_1 _26007_ (.Y(_05866_),
    .A(_05865_),
    .B(net476));
 sg13g2_a21oi_1 _26008_ (.A1(_05864_),
    .A2(_05866_),
    .Y(_01717_),
    .B1(_05841_));
 sg13g2_nand2_1 _26009_ (.Y(_05867_),
    .A(_05499_),
    .B(_08450_));
 sg13g2_buf_1 _26010_ (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_05868_));
 sg13g2_nand2_1 _26011_ (.Y(_05869_),
    .A(_05868_),
    .B(net476));
 sg13g2_a21oi_1 _26012_ (.A1(_05867_),
    .A2(_05869_),
    .Y(_01718_),
    .B1(_05841_));
 sg13g2_nand2_1 _26013_ (.Y(_05870_),
    .A(_05502_),
    .B(_08450_));
 sg13g2_buf_1 _26014_ (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_05871_));
 sg13g2_nand2_1 _26015_ (.Y(_05872_),
    .A(_05871_),
    .B(_05848_));
 sg13g2_buf_1 _26016_ (.A(_05734_),
    .X(_05873_));
 sg13g2_a21oi_1 _26017_ (.A1(_05870_),
    .A2(_05872_),
    .Y(_01719_),
    .B1(net549));
 sg13g2_buf_1 _26018_ (.A(_08449_),
    .X(_05874_));
 sg13g2_nand2_1 _26019_ (.Y(_05875_),
    .A(_05505_),
    .B(net475));
 sg13g2_buf_1 _26020_ (.A(\rbzero.wall_tracer.stepDistY[7] ),
    .X(_05876_));
 sg13g2_nand2_1 _26021_ (.Y(_05877_),
    .A(_05876_),
    .B(_05848_));
 sg13g2_a21oi_1 _26022_ (.A1(_05875_),
    .A2(_05877_),
    .Y(_01720_),
    .B1(net549));
 sg13g2_nand2_1 _26023_ (.Y(_05878_),
    .A(_05508_),
    .B(net475));
 sg13g2_buf_1 _26024_ (.A(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_05879_));
 sg13g2_buf_1 _26025_ (.A(_05847_),
    .X(_05880_));
 sg13g2_nand2_1 _26026_ (.Y(_05881_),
    .A(_05879_),
    .B(_05880_));
 sg13g2_a21oi_1 _26027_ (.A1(_05878_),
    .A2(_05881_),
    .Y(_01721_),
    .B1(_05873_));
 sg13g2_nand2_1 _26028_ (.Y(_05882_),
    .A(_05512_),
    .B(net475));
 sg13g2_nand2_1 _26029_ (.Y(_05883_),
    .A(_12029_),
    .B(net474));
 sg13g2_a21oi_1 _26030_ (.A1(_05882_),
    .A2(_05883_),
    .Y(_01722_),
    .B1(net549));
 sg13g2_nand2_1 _26031_ (.Y(_05884_),
    .A(_05515_),
    .B(_05874_));
 sg13g2_buf_1 _26032_ (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_05885_));
 sg13g2_nand2_1 _26033_ (.Y(_05886_),
    .A(_05885_),
    .B(net474));
 sg13g2_a21oi_1 _26034_ (.A1(_05884_),
    .A2(_05886_),
    .Y(_01723_),
    .B1(net549));
 sg13g2_nand2_1 _26035_ (.Y(_05887_),
    .A(_05520_),
    .B(_05874_));
 sg13g2_nand2_1 _26036_ (.Y(_05888_),
    .A(\rbzero.wall_tracer.stepDistY[10] ),
    .B(_05880_));
 sg13g2_a21oi_1 _26037_ (.A1(_05887_),
    .A2(_05888_),
    .Y(_01724_),
    .B1(_05873_));
 sg13g2_nand2_1 _26038_ (.Y(_05889_),
    .A(_05530_),
    .B(net475));
 sg13g2_buf_1 _26039_ (.A(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_05890_));
 sg13g2_nand2_1 _26040_ (.Y(_05891_),
    .A(_05890_),
    .B(net474));
 sg13g2_a21oi_1 _26041_ (.A1(_05889_),
    .A2(_05891_),
    .Y(_01725_),
    .B1(net549));
 sg13g2_nand2_1 _26042_ (.Y(_05892_),
    .A(_05543_),
    .B(net475));
 sg13g2_buf_1 _26043_ (.A(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_05893_));
 sg13g2_nand2_1 _26044_ (.Y(_05894_),
    .A(_05893_),
    .B(net474));
 sg13g2_a21oi_1 _26045_ (.A1(_05892_),
    .A2(_05894_),
    .Y(_01726_),
    .B1(net549));
 sg13g2_nand2_1 _26046_ (.Y(_05895_),
    .A(_05550_),
    .B(net475));
 sg13g2_nand2_1 _26047_ (.Y(_05896_),
    .A(\rbzero.wall_tracer.stepDistY[-7] ),
    .B(net474));
 sg13g2_a21oi_1 _26048_ (.A1(_05895_),
    .A2(_05896_),
    .Y(_01727_),
    .B1(net549));
 sg13g2_nand2_1 _26049_ (.Y(_05897_),
    .A(_05558_),
    .B(net475));
 sg13g2_buf_1 _26050_ (.A(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_05898_));
 sg13g2_nand2_1 _26051_ (.Y(_05899_),
    .A(_05898_),
    .B(net474));
 sg13g2_a21oi_1 _26052_ (.A1(_05897_),
    .A2(_05899_),
    .Y(_01728_),
    .B1(net549));
 sg13g2_nand2_1 _26053_ (.Y(_05900_),
    .A(_05562_),
    .B(net475));
 sg13g2_nand2_1 _26054_ (.Y(_05901_),
    .A(\rbzero.wall_tracer.stepDistY[-5] ),
    .B(net474));
 sg13g2_buf_1 _26055_ (.A(_05734_),
    .X(_05902_));
 sg13g2_a21oi_1 _26056_ (.A1(_05900_),
    .A2(_05901_),
    .Y(_01729_),
    .B1(net548));
 sg13g2_nand2_1 _26057_ (.Y(_05903_),
    .A(_05568_),
    .B(_08449_));
 sg13g2_buf_1 _26058_ (.A(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_05904_));
 sg13g2_nand2_1 _26059_ (.Y(_05905_),
    .A(_05904_),
    .B(net474));
 sg13g2_a21oi_1 _26060_ (.A1(_05903_),
    .A2(_05905_),
    .Y(_01730_),
    .B1(net548));
 sg13g2_nand2_1 _26061_ (.Y(_05906_),
    .A(_05573_),
    .B(_08449_));
 sg13g2_buf_1 _26062_ (.A(\rbzero.wall_tracer.stepDistY[-3] ),
    .X(_05907_));
 sg13g2_nand2_1 _26063_ (.Y(_05908_),
    .A(_05907_),
    .B(_05847_));
 sg13g2_a21oi_1 _26064_ (.A1(_05906_),
    .A2(_05908_),
    .Y(_01731_),
    .B1(_05902_));
 sg13g2_nand2_1 _26065_ (.Y(_05909_),
    .A(_05580_),
    .B(_08449_));
 sg13g2_buf_1 _26066_ (.A(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_05910_));
 sg13g2_nand2_1 _26067_ (.Y(_05911_),
    .A(_05910_),
    .B(_05847_));
 sg13g2_a21oi_1 _26068_ (.A1(_05909_),
    .A2(_05911_),
    .Y(_01732_),
    .B1(_05902_));
 sg13g2_nand2_1 _26069_ (.Y(_05912_),
    .A(\rbzero.wall_tracer.texu[0] ),
    .B(net496));
 sg13g2_o21ai_1 _26070_ (.B1(_12657_),
    .Y(_05913_),
    .A1(_12560_),
    .A2(_12658_));
 sg13g2_nor2_1 _26071_ (.A(_12659_),
    .B(_05913_),
    .Y(_05914_));
 sg13g2_a21oi_1 _26072_ (.A1(_12656_),
    .A2(_12659_),
    .Y(_05915_),
    .B1(_05914_));
 sg13g2_nand2_1 _26073_ (.Y(_05916_),
    .A(_09820_),
    .B(net633));
 sg13g2_o21ai_1 _26074_ (.B1(_05916_),
    .Y(_05917_),
    .A1(_11889_),
    .A2(net633));
 sg13g2_nor2_1 _26075_ (.A(_05915_),
    .B(_05917_),
    .Y(_05918_));
 sg13g2_nand2b_1 _26076_ (.Y(_05919_),
    .B(net633),
    .A_N(_00443_));
 sg13g2_o21ai_1 _26077_ (.B1(_05919_),
    .Y(_05920_),
    .A1(net633),
    .A2(_00442_));
 sg13g2_o21ai_1 _26078_ (.B1(_05920_),
    .Y(_05921_),
    .A1(_12777_),
    .A2(_05918_));
 sg13g2_nand2_1 _26079_ (.Y(_05922_),
    .A(_12777_),
    .B(_05918_));
 sg13g2_nand2_1 _26080_ (.Y(_05923_),
    .A(_05921_),
    .B(_05922_));
 sg13g2_nand2b_1 _26081_ (.Y(_05924_),
    .B(net633),
    .A_N(_00437_));
 sg13g2_o21ai_1 _26082_ (.B1(_05924_),
    .Y(_05925_),
    .A1(net633),
    .A2(_00436_));
 sg13g2_a21o_1 _26083_ (.A2(_05923_),
    .A1(_12890_),
    .B1(_05925_),
    .X(_05926_));
 sg13g2_o21ai_1 _26084_ (.B1(_05926_),
    .Y(_05927_),
    .A1(_12890_),
    .A2(_05923_));
 sg13g2_buf_1 _26085_ (.A(_05927_),
    .X(_05928_));
 sg13g2_nor2_1 _26086_ (.A(net573),
    .B(net302),
    .Y(_05929_));
 sg13g2_a21oi_1 _26087_ (.A1(net573),
    .A2(_11638_),
    .Y(_05930_),
    .B1(_05929_));
 sg13g2_buf_2 _26088_ (.A(_05930_),
    .X(_05931_));
 sg13g2_mux2_1 _26089_ (.A0(_00430_),
    .A1(_00431_),
    .S(net633),
    .X(_05932_));
 sg13g2_xnor2_1 _26090_ (.Y(_05933_),
    .A(_05931_),
    .B(_05932_));
 sg13g2_xnor2_1 _26091_ (.Y(_05934_),
    .A(_13013_),
    .B(_05933_));
 sg13g2_xnor2_1 _26092_ (.Y(_05935_),
    .A(_05928_),
    .B(_05934_));
 sg13g2_nand2_1 _26093_ (.Y(_05936_),
    .A(net512),
    .B(_05935_));
 sg13g2_a21oi_1 _26094_ (.A1(_05912_),
    .A2(_05936_),
    .Y(_01733_),
    .B1(net548));
 sg13g2_nand2_1 _26095_ (.Y(_05937_),
    .A(\rbzero.wall_tracer.texu[1] ),
    .B(net496));
 sg13g2_a21oi_1 _26096_ (.A1(_13013_),
    .A2(_05928_),
    .Y(_05938_),
    .B1(_05932_));
 sg13g2_nor2_1 _26097_ (.A(_13013_),
    .B(_05928_),
    .Y(_05939_));
 sg13g2_nor2_1 _26098_ (.A(_05938_),
    .B(_05939_),
    .Y(_05940_));
 sg13g2_mux2_1 _26099_ (.A0(_00424_),
    .A1(_00425_),
    .S(net573),
    .X(_05941_));
 sg13g2_xor2_1 _26100_ (.B(_05941_),
    .A(_05931_),
    .X(_05942_));
 sg13g2_xnor2_1 _26101_ (.Y(_05943_),
    .A(_13142_),
    .B(_05942_));
 sg13g2_xnor2_1 _26102_ (.Y(_05944_),
    .A(_05940_),
    .B(_05943_));
 sg13g2_nand2_1 _26103_ (.Y(_05945_),
    .A(net512),
    .B(_05944_));
 sg13g2_a21oi_1 _26104_ (.A1(_05937_),
    .A2(_05945_),
    .Y(_01734_),
    .B1(net548));
 sg13g2_nand2_1 _26105_ (.Y(_05946_),
    .A(\rbzero.wall_tracer.texu[2] ),
    .B(net496));
 sg13g2_inv_1 _26106_ (.Y(_05947_),
    .A(_05940_));
 sg13g2_inv_1 _26107_ (.Y(_05948_),
    .A(_13142_));
 sg13g2_a21oi_1 _26108_ (.A1(_05948_),
    .A2(_05940_),
    .Y(_05949_),
    .B1(_05941_));
 sg13g2_a21oi_1 _26109_ (.A1(_13142_),
    .A2(_05947_),
    .Y(_05950_),
    .B1(_05949_));
 sg13g2_mux2_1 _26110_ (.A0(_00418_),
    .A1(_00419_),
    .S(net573),
    .X(_05951_));
 sg13g2_buf_1 _26111_ (.A(_05951_),
    .X(_05952_));
 sg13g2_xor2_1 _26112_ (.B(_05952_),
    .A(_05931_),
    .X(_05953_));
 sg13g2_xnor2_1 _26113_ (.Y(_05954_),
    .A(_13282_),
    .B(_05953_));
 sg13g2_xnor2_1 _26114_ (.Y(_05955_),
    .A(_05950_),
    .B(_05954_));
 sg13g2_nand2_1 _26115_ (.Y(_05956_),
    .A(net512),
    .B(_05955_));
 sg13g2_a21oi_1 _26116_ (.A1(_05946_),
    .A2(_05956_),
    .Y(_01735_),
    .B1(net548));
 sg13g2_nand2_1 _26117_ (.Y(_05957_),
    .A(\rbzero.wall_tracer.texu[3] ),
    .B(net496));
 sg13g2_nand2_1 _26118_ (.Y(_05958_),
    .A(_05950_),
    .B(_05952_));
 sg13g2_nor2_1 _26119_ (.A(_05950_),
    .B(_05952_),
    .Y(_05959_));
 sg13g2_a21oi_2 _26120_ (.B1(_05959_),
    .Y(_05960_),
    .A2(_05958_),
    .A1(_13282_));
 sg13g2_mux2_1 _26121_ (.A0(_00412_),
    .A1(_00413_),
    .S(net573),
    .X(_05961_));
 sg13g2_xnor2_1 _26122_ (.Y(_05962_),
    .A(_05931_),
    .B(_05961_));
 sg13g2_xnor2_1 _26123_ (.Y(_05963_),
    .A(_13422_),
    .B(_05962_));
 sg13g2_xnor2_1 _26124_ (.Y(_05964_),
    .A(_05960_),
    .B(_05963_));
 sg13g2_nand2_1 _26125_ (.Y(_05965_),
    .A(net512),
    .B(_05964_));
 sg13g2_a21oi_1 _26126_ (.A1(_05957_),
    .A2(_05965_),
    .Y(_01736_),
    .B1(net548));
 sg13g2_nand2_1 _26127_ (.Y(_05966_),
    .A(\rbzero.wall_tracer.texu[4] ),
    .B(net496));
 sg13g2_a21o_1 _26128_ (.A2(_05960_),
    .A1(_13422_),
    .B1(_05961_),
    .X(_05967_));
 sg13g2_o21ai_1 _26129_ (.B1(_05967_),
    .Y(_05968_),
    .A1(_13422_),
    .A2(_05960_));
 sg13g2_buf_1 _26130_ (.A(_05968_),
    .X(_05969_));
 sg13g2_mux2_1 _26131_ (.A0(_00407_),
    .A1(_00408_),
    .S(_11713_),
    .X(_05970_));
 sg13g2_xnor2_1 _26132_ (.Y(_05971_),
    .A(_05931_),
    .B(_05970_));
 sg13g2_xnor2_1 _26133_ (.Y(_05972_),
    .A(_13559_),
    .B(_05971_));
 sg13g2_xnor2_1 _26134_ (.Y(_05973_),
    .A(_05969_),
    .B(_05972_));
 sg13g2_nand2_1 _26135_ (.Y(_05974_),
    .A(net512),
    .B(_05973_));
 sg13g2_a21oi_1 _26136_ (.A1(_05966_),
    .A2(_05974_),
    .Y(_01737_),
    .B1(net548));
 sg13g2_nand2_1 _26137_ (.Y(_05975_),
    .A(\rbzero.wall_tracer.texu[5] ),
    .B(net496));
 sg13g2_mux2_1 _26138_ (.A0(_00401_),
    .A1(_00402_),
    .S(_11713_),
    .X(_05976_));
 sg13g2_xnor2_1 _26139_ (.Y(_05977_),
    .A(_05931_),
    .B(_05976_));
 sg13g2_xnor2_1 _26140_ (.Y(_05978_),
    .A(_13724_),
    .B(_05977_));
 sg13g2_nor2_1 _26141_ (.A(_13559_),
    .B(_05969_),
    .Y(_05979_));
 sg13g2_nand2_1 _26142_ (.Y(_05980_),
    .A(_13559_),
    .B(_05969_));
 sg13g2_o21ai_1 _26143_ (.B1(_05980_),
    .Y(_05981_),
    .A1(_05970_),
    .A2(_05979_));
 sg13g2_xnor2_1 _26144_ (.Y(_05982_),
    .A(_05978_),
    .B(_05981_));
 sg13g2_nand2_1 _26145_ (.Y(_05983_),
    .A(net512),
    .B(_05982_));
 sg13g2_a21oi_1 _26146_ (.A1(_05975_),
    .A2(_05983_),
    .Y(_01738_),
    .B1(net548));
 sg13g2_and2_1 _26147_ (.A(_12348_),
    .B(_12558_),
    .X(_05984_));
 sg13g2_nor2_1 _26148_ (.A(_12348_),
    .B(_12558_),
    .Y(_05985_));
 sg13g2_or3_1 _26149_ (.A(_08480_),
    .B(_05984_),
    .C(_05985_),
    .X(_05986_));
 sg13g2_or2_1 _26150_ (.X(_05987_),
    .B(_05986_),
    .A(net68));
 sg13g2_buf_1 _26151_ (.A(net69),
    .X(_05988_));
 sg13g2_nand2_1 _26152_ (.Y(_05989_),
    .A(_12013_),
    .B(_11472_));
 sg13g2_nand2b_1 _26153_ (.Y(_05990_),
    .B(_11267_),
    .A_N(_12013_));
 sg13g2_o21ai_1 _26154_ (.B1(_05990_),
    .Y(_05991_),
    .A1(_11267_),
    .A2(_05989_));
 sg13g2_buf_1 _26155_ (.A(net700),
    .X(_05992_));
 sg13g2_a22oi_1 _26156_ (.Y(_05993_),
    .B1(_05991_),
    .B2(net619),
    .A2(net61),
    .A1(_11267_));
 sg13g2_buf_1 _26157_ (.A(_08675_),
    .X(_05994_));
 sg13g2_a21oi_1 _26158_ (.A1(_05987_),
    .A2(_05993_),
    .Y(_01739_),
    .B1(net618));
 sg13g2_nor2_1 _26159_ (.A(_08479_),
    .B(_11341_),
    .Y(_05995_));
 sg13g2_buf_2 _26160_ (.A(_05995_),
    .X(_05996_));
 sg13g2_buf_1 _26161_ (.A(_05996_),
    .X(_05997_));
 sg13g2_nand2_1 _26162_ (.Y(_05998_),
    .A(_13724_),
    .B(net60));
 sg13g2_inv_1 _26163_ (.Y(_05999_),
    .A(\rbzero.wall_tracer.stepDistX[-1] ));
 sg13g2_inv_1 _26164_ (.Y(_06000_),
    .A(\rbzero.wall_tracer.stepDistX[-5] ));
 sg13g2_inv_1 _26165_ (.Y(_06001_),
    .A(\rbzero.wall_tracer.stepDistX[-7] ));
 sg13g2_inv_1 _26166_ (.Y(_06002_),
    .A(_05823_));
 sg13g2_a21oi_1 _26167_ (.A1(_11267_),
    .A2(_12013_),
    .Y(_06003_),
    .B1(_12023_));
 sg13g2_nand3_1 _26168_ (.B(_12013_),
    .C(_12023_),
    .A(_11267_),
    .Y(_06004_));
 sg13g2_o21ai_1 _26169_ (.B1(_06004_),
    .Y(_06005_),
    .A1(_11266_),
    .A2(_06003_));
 sg13g2_a21oi_1 _26170_ (.A1(_11262_),
    .A2(_05823_),
    .Y(_06006_),
    .B1(_06005_));
 sg13g2_a21oi_2 _26171_ (.B1(_06006_),
    .Y(_06007_),
    .A2(_06002_),
    .A1(_11263_));
 sg13g2_a21o_1 _26172_ (.A2(_06007_),
    .A1(_05826_),
    .B1(_11261_),
    .X(_06008_));
 sg13g2_o21ai_1 _26173_ (.B1(_06008_),
    .Y(_06009_),
    .A1(_05826_),
    .A2(_06007_));
 sg13g2_buf_1 _26174_ (.A(_06009_),
    .X(_06010_));
 sg13g2_a21o_1 _26175_ (.A2(_06010_),
    .A1(_06001_),
    .B1(_11259_),
    .X(_06011_));
 sg13g2_o21ai_1 _26176_ (.B1(_06011_),
    .Y(_06012_),
    .A1(_06001_),
    .A2(_06010_));
 sg13g2_buf_1 _26177_ (.A(_06012_),
    .X(_06013_));
 sg13g2_a21o_1 _26178_ (.A2(_06013_),
    .A1(_05831_),
    .B1(_11256_),
    .X(_06014_));
 sg13g2_o21ai_1 _26179_ (.B1(_06014_),
    .Y(_06015_),
    .A1(_05831_),
    .A2(_06013_));
 sg13g2_buf_1 _26180_ (.A(_06015_),
    .X(_06016_));
 sg13g2_a21o_1 _26181_ (.A2(_06016_),
    .A1(_06000_),
    .B1(_11253_),
    .X(_06017_));
 sg13g2_o21ai_1 _26182_ (.B1(_06017_),
    .Y(_06018_),
    .A1(_06000_),
    .A2(_06016_));
 sg13g2_buf_1 _26183_ (.A(_06018_),
    .X(_06019_));
 sg13g2_nor2_1 _26184_ (.A(_05836_),
    .B(_06019_),
    .Y(_06020_));
 sg13g2_a21oi_1 _26185_ (.A1(_05836_),
    .A2(_06019_),
    .Y(_06021_),
    .B1(_11249_));
 sg13g2_nor2_1 _26186_ (.A(_06020_),
    .B(_06021_),
    .Y(_06022_));
 sg13g2_nor2_1 _26187_ (.A(_05839_),
    .B(_06022_),
    .Y(_06023_));
 sg13g2_a21oi_1 _26188_ (.A1(_05839_),
    .A2(_06022_),
    .Y(_06024_),
    .B1(_11247_));
 sg13g2_nor2_1 _26189_ (.A(_06023_),
    .B(_06024_),
    .Y(_06025_));
 sg13g2_a21o_1 _26190_ (.A2(_06025_),
    .A1(_05843_),
    .B1(_11243_),
    .X(_06026_));
 sg13g2_o21ai_1 _26191_ (.B1(_06026_),
    .Y(_06027_),
    .A1(_05843_),
    .A2(_06025_));
 sg13g2_buf_1 _26192_ (.A(_06027_),
    .X(_06028_));
 sg13g2_xnor2_1 _26193_ (.Y(_06029_),
    .A(_05999_),
    .B(_06028_));
 sg13g2_nor3_1 _26194_ (.A(_11291_),
    .B(net71),
    .C(_06029_),
    .Y(_06030_));
 sg13g2_a21o_1 _26195_ (.A2(_06029_),
    .A1(_11291_),
    .B1(_06030_),
    .X(_06031_));
 sg13g2_a22oi_1 _26196_ (.Y(_06032_),
    .B1(_06031_),
    .B2(net619),
    .A2(net61),
    .A1(_11291_));
 sg13g2_a21oi_1 _26197_ (.A1(_05998_),
    .A2(_06032_),
    .Y(_01740_),
    .B1(net618));
 sg13g2_nand2_1 _26198_ (.Y(_06033_),
    .A(_13880_),
    .B(net60));
 sg13g2_inv_1 _26199_ (.Y(_06034_),
    .A(_06028_));
 sg13g2_a21oi_1 _26200_ (.A1(\rbzero.wall_tracer.stepDistX[-1] ),
    .A2(_06034_),
    .Y(_06035_),
    .B1(_11291_));
 sg13g2_a21oi_1 _26201_ (.A1(_05999_),
    .A2(_06028_),
    .Y(_06036_),
    .B1(_06035_));
 sg13g2_xnor2_1 _26202_ (.Y(_06037_),
    .A(_05786_),
    .B(_06036_));
 sg13g2_nor3_1 _26203_ (.A(_11239_),
    .B(net71),
    .C(_06037_),
    .Y(_06038_));
 sg13g2_a21o_1 _26204_ (.A2(_06037_),
    .A1(_11239_),
    .B1(_06038_),
    .X(_06039_));
 sg13g2_a22oi_1 _26205_ (.Y(_06040_),
    .B1(_06039_),
    .B2(net619),
    .A2(net61),
    .A1(_11239_));
 sg13g2_a21oi_1 _26206_ (.A1(_06033_),
    .A2(_06040_),
    .Y(_01741_),
    .B1(net618));
 sg13g2_nand2b_1 _26207_ (.Y(_06041_),
    .B(_05996_),
    .A_N(_14050_));
 sg13g2_nor2_1 _26208_ (.A(_05786_),
    .B(_06036_),
    .Y(_06042_));
 sg13g2_a21oi_1 _26209_ (.A1(_05786_),
    .A2(_06036_),
    .Y(_06043_),
    .B1(_11239_));
 sg13g2_nor2_1 _26210_ (.A(_06042_),
    .B(_06043_),
    .Y(_06044_));
 sg13g2_xnor2_1 _26211_ (.Y(_06045_),
    .A(_05789_),
    .B(_06044_));
 sg13g2_nor3_1 _26212_ (.A(_11237_),
    .B(net71),
    .C(_06045_),
    .Y(_06046_));
 sg13g2_a21o_1 _26213_ (.A2(_06045_),
    .A1(_11237_),
    .B1(_06046_),
    .X(_06047_));
 sg13g2_a22oi_1 _26214_ (.Y(_06048_),
    .B1(_06047_),
    .B2(net619),
    .A2(net61),
    .A1(_11237_));
 sg13g2_a21oi_1 _26215_ (.A1(_06041_),
    .A2(_06048_),
    .Y(_01742_),
    .B1(net618));
 sg13g2_nand2_1 _26216_ (.Y(_06049_),
    .A(_01905_),
    .B(_05997_));
 sg13g2_nor2_1 _26217_ (.A(_05789_),
    .B(_06044_),
    .Y(_06050_));
 sg13g2_a21oi_1 _26218_ (.A1(_05789_),
    .A2(_06044_),
    .Y(_06051_),
    .B1(_11237_));
 sg13g2_nor2_1 _26219_ (.A(_06050_),
    .B(_06051_),
    .Y(_06052_));
 sg13g2_xnor2_1 _26220_ (.Y(_06053_),
    .A(_05792_),
    .B(_06052_));
 sg13g2_nor3_1 _26221_ (.A(_11233_),
    .B(net71),
    .C(_06053_),
    .Y(_06054_));
 sg13g2_a21o_1 _26222_ (.A2(_06053_),
    .A1(_11233_),
    .B1(_06054_),
    .X(_06055_));
 sg13g2_a22oi_1 _26223_ (.Y(_06056_),
    .B1(_06055_),
    .B2(net619),
    .A2(net61),
    .A1(_11233_));
 sg13g2_a21oi_1 _26224_ (.A1(_06049_),
    .A2(_06056_),
    .Y(_01743_),
    .B1(net618));
 sg13g2_nor2_1 _26225_ (.A(_05792_),
    .B(_06052_),
    .Y(_06057_));
 sg13g2_a21oi_1 _26226_ (.A1(_05792_),
    .A2(_06052_),
    .Y(_06058_),
    .B1(_11233_));
 sg13g2_nor2_1 _26227_ (.A(_06057_),
    .B(_06058_),
    .Y(_06059_));
 sg13g2_xnor2_1 _26228_ (.Y(_06060_),
    .A(_05795_),
    .B(_06059_));
 sg13g2_nor3_1 _26229_ (.A(_11231_),
    .B(net72),
    .C(_06060_),
    .Y(_06061_));
 sg13g2_a21o_1 _26230_ (.A2(_06060_),
    .A1(_11231_),
    .B1(_06061_),
    .X(_06062_));
 sg13g2_o21ai_1 _26231_ (.B1(_01903_),
    .Y(_06063_),
    .A1(_14055_),
    .A2(_01902_));
 sg13g2_buf_1 _26232_ (.A(_06063_),
    .X(_06064_));
 sg13g2_or2_1 _26233_ (.X(_06065_),
    .B(_01895_),
    .A(_01888_));
 sg13g2_inv_1 _26234_ (.Y(_06066_),
    .A(_14060_));
 sg13g2_o21ai_1 _26235_ (.B1(_01885_),
    .Y(_06067_),
    .A1(_06066_),
    .A2(_01896_));
 sg13g2_nand2_1 _26236_ (.Y(_06068_),
    .A(_06066_),
    .B(_01896_));
 sg13g2_a21oi_1 _26237_ (.A1(_14080_),
    .A2(_14091_),
    .Y(_06069_),
    .B1(_14090_));
 sg13g2_a21oi_2 _26238_ (.B1(_01830_),
    .Y(_06070_),
    .A2(_01831_),
    .A1(_14104_));
 sg13g2_nor2_1 _26239_ (.A(_14074_),
    .B(_14078_),
    .Y(_06071_));
 sg13g2_nand2_1 _26240_ (.Y(_06072_),
    .A(_14074_),
    .B(_14078_));
 sg13g2_o21ai_1 _26241_ (.B1(_06072_),
    .Y(_06073_),
    .A1(_14069_),
    .A2(_06071_));
 sg13g2_inv_1 _26242_ (.Y(_06074_),
    .A(_14064_));
 sg13g2_a22oi_1 _26243_ (.Y(_06075_),
    .B1(_06074_),
    .B2(_14065_),
    .A2(net174),
    .A1(net210));
 sg13g2_a21oi_2 _26244_ (.B1(_06075_),
    .Y(_06076_),
    .A2(_14066_),
    .A1(_14064_));
 sg13g2_nor2_1 _26245_ (.A(_01821_),
    .B(_01822_),
    .Y(_06077_));
 sg13g2_nor2_1 _26246_ (.A(_01820_),
    .B(_06077_),
    .Y(_06078_));
 sg13g2_a21oi_1 _26247_ (.A1(_01821_),
    .A2(_01822_),
    .Y(_06079_),
    .B1(_06078_));
 sg13g2_buf_2 _26248_ (.A(_06079_),
    .X(_06080_));
 sg13g2_xnor2_1 _26249_ (.Y(_06081_),
    .A(_06076_),
    .B(_06080_));
 sg13g2_nor2_1 _26250_ (.A(net262),
    .B(net206),
    .Y(_06082_));
 sg13g2_nand2_1 _26251_ (.Y(_06083_),
    .A(net237),
    .B(_13903_));
 sg13g2_xor2_1 _26252_ (.B(_06083_),
    .A(_06082_),
    .X(_06084_));
 sg13g2_nand2_1 _26253_ (.Y(_06085_),
    .A(net205),
    .B(net257));
 sg13g2_buf_2 _26254_ (.A(_06085_),
    .X(_06086_));
 sg13g2_inv_1 _26255_ (.Y(_06087_),
    .A(_06086_));
 sg13g2_xnor2_1 _26256_ (.Y(_06088_),
    .A(_06084_),
    .B(_06087_));
 sg13g2_xnor2_1 _26257_ (.Y(_06089_),
    .A(_06081_),
    .B(_06088_));
 sg13g2_buf_1 _26258_ (.A(_13910_),
    .X(_06090_));
 sg13g2_nand3_1 _26259_ (.B(net520),
    .C(_13023_),
    .A(net235),
    .Y(_06091_));
 sg13g2_nand2b_1 _26260_ (.Y(_06092_),
    .B(_06091_),
    .A_N(_14087_));
 sg13g2_xnor2_1 _26261_ (.Y(_06093_),
    .A(net505),
    .B(_06092_));
 sg13g2_and2_1 _26262_ (.A(net212),
    .B(_06093_),
    .X(_06094_));
 sg13g2_buf_1 _26263_ (.A(_06094_),
    .X(_06095_));
 sg13g2_xnor2_1 _26264_ (.Y(_06096_),
    .A(_06089_),
    .B(_06095_));
 sg13g2_xnor2_1 _26265_ (.Y(_06097_),
    .A(_06073_),
    .B(_06096_));
 sg13g2_xnor2_1 _26266_ (.Y(_06098_),
    .A(_06070_),
    .B(_06097_));
 sg13g2_xnor2_1 _26267_ (.Y(_06099_),
    .A(_06069_),
    .B(_06098_));
 sg13g2_a21o_1 _26268_ (.A2(_01824_),
    .A1(_01816_),
    .B1(_01819_),
    .X(_06100_));
 sg13g2_o21ai_1 _26269_ (.B1(_06100_),
    .Y(_06101_),
    .A1(_01816_),
    .A2(_01824_));
 sg13g2_nand2b_1 _26270_ (.Y(_06102_),
    .B(_01814_),
    .A_N(_01811_));
 sg13g2_a21oi_1 _26271_ (.A1(net256),
    .A2(net500),
    .Y(_06103_),
    .B1(_01814_));
 sg13g2_a21oi_1 _26272_ (.A1(_01813_),
    .A2(_06102_),
    .Y(_06104_),
    .B1(_06103_));
 sg13g2_nand2_1 _26273_ (.Y(_06105_),
    .A(net236),
    .B(net172));
 sg13g2_nand2_1 _26274_ (.Y(_06106_),
    .A(_13789_),
    .B(net255));
 sg13g2_nand2_1 _26275_ (.Y(_06107_),
    .A(net234),
    .B(_13951_));
 sg13g2_xnor2_1 _26276_ (.Y(_06108_),
    .A(_06106_),
    .B(_06107_));
 sg13g2_xnor2_1 _26277_ (.Y(_06109_),
    .A(_06105_),
    .B(_06108_));
 sg13g2_nor2b_1 _26278_ (.A(net208),
    .B_N(net233),
    .Y(_06110_));
 sg13g2_nand2_1 _26279_ (.Y(_06111_),
    .A(net232),
    .B(net173));
 sg13g2_nand2_1 _26280_ (.Y(_06112_),
    .A(net204),
    .B(_13506_));
 sg13g2_xnor2_1 _26281_ (.Y(_06113_),
    .A(_06111_),
    .B(_06112_));
 sg13g2_xnor2_1 _26282_ (.Y(_06114_),
    .A(_06110_),
    .B(_06113_));
 sg13g2_xnor2_1 _26283_ (.Y(_06115_),
    .A(_06109_),
    .B(_06114_));
 sg13g2_xnor2_1 _26284_ (.Y(_06116_),
    .A(_06104_),
    .B(_06115_));
 sg13g2_a21o_1 _26285_ (.A2(_01853_),
    .A1(_01849_),
    .B1(_01845_),
    .X(_06117_));
 sg13g2_o21ai_1 _26286_ (.B1(_06117_),
    .Y(_06118_),
    .A1(_01849_),
    .A2(_01853_));
 sg13g2_buf_1 _26287_ (.A(_06118_),
    .X(_06119_));
 sg13g2_xor2_1 _26288_ (.B(_06119_),
    .A(_06116_),
    .X(_06120_));
 sg13g2_xnor2_1 _26289_ (.Y(_06121_),
    .A(_06101_),
    .B(_06120_));
 sg13g2_and2_1 _26290_ (.A(net256),
    .B(net499),
    .X(_06122_));
 sg13g2_buf_1 _26291_ (.A(_06122_),
    .X(_06123_));
 sg13g2_nand2_1 _26292_ (.Y(_06124_),
    .A(net300),
    .B(net501));
 sg13g2_buf_1 _26293_ (.A(_12928_),
    .X(_06125_));
 sg13g2_nand2_1 _26294_ (.Y(_06126_),
    .A(net284),
    .B(net498));
 sg13g2_xnor2_1 _26295_ (.Y(_06127_),
    .A(_06124_),
    .B(_06126_));
 sg13g2_xnor2_1 _26296_ (.Y(_06128_),
    .A(_06123_),
    .B(_06127_));
 sg13g2_a22oi_1 _26297_ (.Y(_06129_),
    .B1(_01838_),
    .B2(_01843_),
    .A2(net501),
    .A1(net288));
 sg13g2_nor2_1 _26298_ (.A(_01838_),
    .B(_01843_),
    .Y(_06130_));
 sg13g2_nor2_1 _26299_ (.A(_06129_),
    .B(_06130_),
    .Y(_06131_));
 sg13g2_nand3_1 _26300_ (.B(net479),
    .C(_01856_),
    .A(net319),
    .Y(_06132_));
 sg13g2_buf_1 _26301_ (.A(net479),
    .X(_06133_));
 sg13g2_a21oi_1 _26302_ (.A1(net319),
    .A2(net469),
    .Y(_06134_),
    .B1(_01856_));
 sg13g2_a21oi_1 _26303_ (.A1(_01857_),
    .A2(_06132_),
    .Y(_06135_),
    .B1(_06134_));
 sg13g2_xnor2_1 _26304_ (.Y(_06136_),
    .A(_06131_),
    .B(_06135_));
 sg13g2_xnor2_1 _26305_ (.Y(_06137_),
    .A(_06128_),
    .B(_06136_));
 sg13g2_nand2_1 _26306_ (.Y(_06138_),
    .A(_01866_),
    .B(_01869_));
 sg13g2_o21ai_1 _26307_ (.B1(_01860_),
    .Y(_06139_),
    .A1(_01866_),
    .A2(_01869_));
 sg13g2_nand2_1 _26308_ (.Y(_06140_),
    .A(_06138_),
    .B(_06139_));
 sg13g2_a21oi_2 _26309_ (.B1(_13387_),
    .Y(_06141_),
    .A2(_11823_),
    .A1(_11816_));
 sg13g2_nand2_1 _26310_ (.Y(_06142_),
    .A(net319),
    .B(net478));
 sg13g2_nand2_1 _26311_ (.Y(_06143_),
    .A(net301),
    .B(net479));
 sg13g2_xnor2_1 _26312_ (.Y(_06144_),
    .A(_06142_),
    .B(_06143_));
 sg13g2_xor2_1 _26313_ (.B(_06144_),
    .A(_06141_),
    .X(_06145_));
 sg13g2_nor2_1 _26314_ (.A(_12069_),
    .B(_13633_),
    .Y(_06146_));
 sg13g2_nor2_1 _26315_ (.A(net362),
    .B(net517),
    .Y(_06147_));
 sg13g2_and2_1 _26316_ (.A(_12362_),
    .B(net477),
    .X(_06148_));
 sg13g2_buf_1 _26317_ (.A(_06148_),
    .X(_06149_));
 sg13g2_xnor2_1 _26318_ (.Y(_06150_),
    .A(_06147_),
    .B(_06149_));
 sg13g2_xnor2_1 _26319_ (.Y(_06151_),
    .A(_06146_),
    .B(_06150_));
 sg13g2_a22oi_1 _26320_ (.Y(_06152_),
    .B1(_01861_),
    .B2(_01862_),
    .A2(net477),
    .A1(net362));
 sg13g2_nor2_1 _26321_ (.A(_01861_),
    .B(_01862_),
    .Y(_06153_));
 sg13g2_nor2_1 _26322_ (.A(_06152_),
    .B(_06153_),
    .Y(_06154_));
 sg13g2_nor2_1 _26323_ (.A(_06151_),
    .B(_06154_),
    .Y(_06155_));
 sg13g2_nand2_1 _26324_ (.Y(_06156_),
    .A(_06151_),
    .B(_06154_));
 sg13g2_nand2b_1 _26325_ (.Y(_06157_),
    .B(_06156_),
    .A_N(_06155_));
 sg13g2_xor2_1 _26326_ (.B(_06157_),
    .A(_06145_),
    .X(_06158_));
 sg13g2_xnor2_1 _26327_ (.Y(_06159_),
    .A(_06140_),
    .B(_06158_));
 sg13g2_xnor2_1 _26328_ (.Y(_06160_),
    .A(_06137_),
    .B(_06159_));
 sg13g2_o21ai_1 _26329_ (.B1(_01855_),
    .Y(_06161_),
    .A1(_01871_),
    .A2(_01873_));
 sg13g2_nand2_1 _26330_ (.Y(_06162_),
    .A(_01871_),
    .B(_01873_));
 sg13g2_nand2_2 _26331_ (.Y(_06163_),
    .A(_06161_),
    .B(_06162_));
 sg13g2_xor2_1 _26332_ (.B(_06163_),
    .A(_06160_),
    .X(_06164_));
 sg13g2_xnor2_1 _26333_ (.Y(_06165_),
    .A(_06121_),
    .B(_06164_));
 sg13g2_nor3_1 _26334_ (.A(_01875_),
    .B(_01835_),
    .C(_01836_),
    .Y(_06166_));
 sg13g2_a21o_1 _26335_ (.A2(_01876_),
    .A1(_01833_),
    .B1(_06166_),
    .X(_06167_));
 sg13g2_buf_1 _26336_ (.A(_06167_),
    .X(_06168_));
 sg13g2_xnor2_1 _26337_ (.Y(_06169_),
    .A(_06165_),
    .B(_06168_));
 sg13g2_xnor2_1 _26338_ (.Y(_06170_),
    .A(_06099_),
    .B(_06169_));
 sg13g2_a21oi_1 _26339_ (.A1(_01879_),
    .A2(_01883_),
    .Y(_06171_),
    .B1(_14101_));
 sg13g2_nor2_1 _26340_ (.A(_01879_),
    .B(_01883_),
    .Y(_06172_));
 sg13g2_nor2_1 _26341_ (.A(_06171_),
    .B(_06172_),
    .Y(_06173_));
 sg13g2_o21ai_1 _26342_ (.B1(_14099_),
    .Y(_06174_),
    .A1(_14063_),
    .A2(_14098_));
 sg13g2_nand3_1 _26343_ (.B(net206),
    .C(_14086_),
    .A(_13748_),
    .Y(_06175_));
 sg13g2_nand3b_1 _26344_ (.B(_06175_),
    .C(_12363_),
    .Y(_06176_),
    .A_N(_14087_));
 sg13g2_a21o_1 _26345_ (.A2(_06176_),
    .A1(_06091_),
    .B1(net231),
    .X(_06177_));
 sg13g2_xor2_1 _26346_ (.B(_06177_),
    .A(_06174_),
    .X(_06178_));
 sg13g2_xnor2_1 _26347_ (.Y(_06179_),
    .A(_06173_),
    .B(_06178_));
 sg13g2_xnor2_1 _26348_ (.Y(_06180_),
    .A(_06170_),
    .B(_06179_));
 sg13g2_nand3_1 _26349_ (.B(_06068_),
    .C(_06180_),
    .A(_06067_),
    .Y(_06181_));
 sg13g2_a21o_1 _26350_ (.A2(_06068_),
    .A1(_06067_),
    .B1(_06180_),
    .X(_06182_));
 sg13g2_nand2_1 _26351_ (.Y(_06183_),
    .A(_06181_),
    .B(_06182_));
 sg13g2_xor2_1 _26352_ (.B(_06183_),
    .A(_06065_),
    .X(_06184_));
 sg13g2_nand2_1 _26353_ (.Y(_06185_),
    .A(_01898_),
    .B(_01899_));
 sg13g2_nor2_1 _26354_ (.A(_01898_),
    .B(_01899_),
    .Y(_06186_));
 sg13g2_a21oi_1 _26355_ (.A1(_14037_),
    .A2(_06185_),
    .Y(_06187_),
    .B1(_06186_));
 sg13g2_and2_1 _26356_ (.A(_06184_),
    .B(_06187_),
    .X(_06188_));
 sg13g2_buf_1 _26357_ (.A(_06188_),
    .X(_06189_));
 sg13g2_or2_1 _26358_ (.X(_06190_),
    .B(_06187_),
    .A(_06184_));
 sg13g2_buf_1 _26359_ (.A(_06190_),
    .X(_06191_));
 sg13g2_nand2b_1 _26360_ (.Y(_06192_),
    .B(_06191_),
    .A_N(_06189_));
 sg13g2_xor2_1 _26361_ (.B(_06192_),
    .A(_06064_),
    .X(_06193_));
 sg13g2_nor3_1 _26362_ (.A(net700),
    .B(_11343_),
    .C(_06193_),
    .Y(_06194_));
 sg13g2_a221oi_1 _26363_ (.B2(_11471_),
    .C1(_06194_),
    .B1(_06062_),
    .A1(_11231_),
    .Y(_06195_),
    .A2(net68));
 sg13g2_nor2_1 _26364_ (.A(_11690_),
    .B(_06195_),
    .Y(_01744_));
 sg13g2_nor2_1 _26365_ (.A(_05795_),
    .B(_06059_),
    .Y(_06196_));
 sg13g2_a21oi_1 _26366_ (.A1(_05795_),
    .A2(_06059_),
    .Y(_06197_),
    .B1(_11231_));
 sg13g2_nor2_1 _26367_ (.A(_06196_),
    .B(_06197_),
    .Y(_06198_));
 sg13g2_xnor2_1 _26368_ (.Y(_06199_),
    .A(_05798_),
    .B(_06198_));
 sg13g2_nor3_1 _26369_ (.A(_11228_),
    .B(_11342_),
    .C(_06199_),
    .Y(_06200_));
 sg13g2_a21o_1 _26370_ (.A2(_06199_),
    .A1(_11228_),
    .B1(_06200_),
    .X(_06201_));
 sg13g2_a21oi_1 _26371_ (.A1(_06064_),
    .A2(_06191_),
    .Y(_06202_),
    .B1(_06189_));
 sg13g2_inv_1 _26372_ (.Y(_06203_),
    .A(_06178_));
 sg13g2_inv_1 _26373_ (.Y(_06204_),
    .A(_06173_));
 sg13g2_o21ai_1 _26374_ (.B1(_06170_),
    .Y(_06205_),
    .A1(_06204_),
    .A2(_06178_));
 sg13g2_o21ai_1 _26375_ (.B1(_06205_),
    .Y(_06206_),
    .A1(_06173_),
    .A2(_06203_));
 sg13g2_buf_1 _26376_ (.A(_06206_),
    .X(_06207_));
 sg13g2_nor2_1 _26377_ (.A(_06174_),
    .B(_06177_),
    .Y(_06208_));
 sg13g2_nand2_1 _26378_ (.Y(_06209_),
    .A(_06116_),
    .B(_06119_));
 sg13g2_o21ai_1 _26379_ (.B1(_06101_),
    .Y(_06210_),
    .A1(_06116_),
    .A2(_06119_));
 sg13g2_nand2_1 _26380_ (.Y(_06211_),
    .A(_06209_),
    .B(_06210_));
 sg13g2_mux2_1 _26381_ (.A0(_06086_),
    .A1(_06084_),
    .S(_06080_),
    .X(_06212_));
 sg13g2_mux2_1 _26382_ (.A0(_06084_),
    .A1(_06087_),
    .S(_06080_),
    .X(_06213_));
 sg13g2_mux2_1 _26383_ (.A0(_06212_),
    .A1(_06213_),
    .S(_06076_),
    .X(_06214_));
 sg13g2_nand2_1 _26384_ (.Y(_06215_),
    .A(net212),
    .B(_06093_));
 sg13g2_buf_2 _26385_ (.A(_06215_),
    .X(_06216_));
 sg13g2_nor2_1 _26386_ (.A(_06083_),
    .B(_06086_),
    .Y(_06217_));
 sg13g2_nand2_1 _26387_ (.Y(_06218_),
    .A(_06083_),
    .B(_06086_));
 sg13g2_o21ai_1 _26388_ (.B1(_06218_),
    .Y(_06219_),
    .A1(_06082_),
    .A2(_06217_));
 sg13g2_buf_1 _26389_ (.A(_06219_),
    .X(_06220_));
 sg13g2_nand2_1 _26390_ (.Y(_06221_),
    .A(_06111_),
    .B(_06112_));
 sg13g2_nor2_1 _26391_ (.A(_06111_),
    .B(_06112_),
    .Y(_06222_));
 sg13g2_a21oi_1 _26392_ (.A1(_06110_),
    .A2(_06221_),
    .Y(_06223_),
    .B1(_06222_));
 sg13g2_xnor2_1 _26393_ (.Y(_06224_),
    .A(_06220_),
    .B(_06223_));
 sg13g2_nand2_1 _26394_ (.Y(_06225_),
    .A(net237),
    .B(net150));
 sg13g2_nor2_1 _26395_ (.A(net262),
    .B(_13676_),
    .Y(_06226_));
 sg13g2_xnor2_1 _26396_ (.Y(_06227_),
    .A(_06225_),
    .B(_06226_));
 sg13g2_xnor2_1 _26397_ (.Y(_06228_),
    .A(_06224_),
    .B(_06227_));
 sg13g2_xnor2_1 _26398_ (.Y(_06229_),
    .A(_06216_),
    .B(_06228_));
 sg13g2_xnor2_1 _26399_ (.Y(_06230_),
    .A(_06214_),
    .B(_06229_));
 sg13g2_inv_1 _26400_ (.Y(_06231_),
    .A(_06089_));
 sg13g2_buf_1 _26401_ (.A(_06095_),
    .X(_06232_));
 sg13g2_a21oi_1 _26402_ (.A1(_06089_),
    .A2(net89),
    .Y(_06233_),
    .B1(_06073_));
 sg13g2_a21oi_1 _26403_ (.A1(_06231_),
    .A2(_06216_),
    .Y(_06234_),
    .B1(_06233_));
 sg13g2_xnor2_1 _26404_ (.Y(_06235_),
    .A(_06230_),
    .B(_06234_));
 sg13g2_xor2_1 _26405_ (.B(_06235_),
    .A(_06211_),
    .X(_06236_));
 sg13g2_inv_1 _26406_ (.Y(_06237_),
    .A(_06114_));
 sg13g2_nand2_1 _26407_ (.Y(_06238_),
    .A(_06109_),
    .B(_06237_));
 sg13g2_nor2_1 _26408_ (.A(_06109_),
    .B(_06237_),
    .Y(_06239_));
 sg13g2_a21oi_1 _26409_ (.A1(_06104_),
    .A2(_06238_),
    .Y(_06240_),
    .B1(_06239_));
 sg13g2_a21o_1 _26410_ (.A2(_06107_),
    .A1(_06105_),
    .B1(_06106_),
    .X(_06241_));
 sg13g2_o21ai_1 _26411_ (.B1(_06241_),
    .Y(_06242_),
    .A1(_06105_),
    .A2(_06107_));
 sg13g2_nand2_1 _26412_ (.Y(_06243_),
    .A(net233),
    .B(net149));
 sg13g2_and2_1 _26413_ (.A(net232),
    .B(_13506_),
    .X(_06244_));
 sg13g2_buf_1 _26414_ (.A(_06244_),
    .X(_06245_));
 sg13g2_nor2b_1 _26415_ (.A(net208),
    .B_N(net204),
    .Y(_06246_));
 sg13g2_xnor2_1 _26416_ (.Y(_06247_),
    .A(_06245_),
    .B(_06246_));
 sg13g2_xnor2_1 _26417_ (.Y(_06248_),
    .A(_06243_),
    .B(_06247_));
 sg13g2_nand2_1 _26418_ (.Y(_06249_),
    .A(net236),
    .B(net173));
 sg13g2_nor2_1 _26419_ (.A(_12630_),
    .B(net258),
    .Y(_06250_));
 sg13g2_nand2_1 _26420_ (.Y(_06251_),
    .A(_13791_),
    .B(net172));
 sg13g2_xor2_1 _26421_ (.B(_06251_),
    .A(_06250_),
    .X(_06252_));
 sg13g2_xnor2_1 _26422_ (.Y(_06253_),
    .A(_06249_),
    .B(_06252_));
 sg13g2_xnor2_1 _26423_ (.Y(_06254_),
    .A(_06248_),
    .B(_06253_));
 sg13g2_xnor2_1 _26424_ (.Y(_06255_),
    .A(_06242_),
    .B(_06254_));
 sg13g2_a21oi_1 _26425_ (.A1(_06128_),
    .A2(_06135_),
    .Y(_06256_),
    .B1(_06131_));
 sg13g2_nor2_1 _26426_ (.A(_06128_),
    .B(_06135_),
    .Y(_06257_));
 sg13g2_nor2_1 _26427_ (.A(_06256_),
    .B(_06257_),
    .Y(_06258_));
 sg13g2_xor2_1 _26428_ (.B(_06258_),
    .A(_06255_),
    .X(_06259_));
 sg13g2_xnor2_1 _26429_ (.Y(_06260_),
    .A(_06240_),
    .B(_06259_));
 sg13g2_nand2_1 _26430_ (.Y(_06261_),
    .A(_01812_),
    .B(net499));
 sg13g2_nand2_1 _26431_ (.Y(_06262_),
    .A(net284),
    .B(net501));
 sg13g2_nand2_1 _26432_ (.Y(_06263_),
    .A(net256),
    .B(_01841_));
 sg13g2_xnor2_1 _26433_ (.Y(_06264_),
    .A(_06262_),
    .B(_06263_));
 sg13g2_xnor2_1 _26434_ (.Y(_06265_),
    .A(_06261_),
    .B(_06264_));
 sg13g2_nand3_1 _26435_ (.B(net469),
    .C(_06141_),
    .A(net301),
    .Y(_06266_));
 sg13g2_nor2b_1 _26436_ (.A(_06141_),
    .B_N(_06143_),
    .Y(_06267_));
 sg13g2_a21oi_2 _26437_ (.B1(_06267_),
    .Y(_06268_),
    .A2(_06266_),
    .A1(_06142_));
 sg13g2_nor2b_1 _26438_ (.A(_06123_),
    .B_N(_06126_),
    .Y(_06269_));
 sg13g2_nand3_1 _26439_ (.B(net498),
    .C(_06123_),
    .A(net284),
    .Y(_06270_));
 sg13g2_o21ai_1 _26440_ (.B1(_06270_),
    .Y(_06271_),
    .A1(_06124_),
    .A2(_06269_));
 sg13g2_buf_1 _26441_ (.A(_06271_),
    .X(_06272_));
 sg13g2_xnor2_1 _26442_ (.Y(_06273_),
    .A(_06268_),
    .B(_06272_));
 sg13g2_xnor2_1 _26443_ (.Y(_06274_),
    .A(_06265_),
    .B(_06273_));
 sg13g2_and2_1 _26444_ (.A(net300),
    .B(net482),
    .X(_06275_));
 sg13g2_buf_1 _26445_ (.A(_06275_),
    .X(_06276_));
 sg13g2_nand2_1 _26446_ (.Y(_06277_),
    .A(net301),
    .B(net478));
 sg13g2_nand2_1 _26447_ (.Y(_06278_),
    .A(_01839_),
    .B(_13391_));
 sg13g2_xnor2_1 _26448_ (.Y(_06279_),
    .A(_06277_),
    .B(_06278_));
 sg13g2_xnor2_1 _26449_ (.Y(_06280_),
    .A(_06276_),
    .B(_06279_));
 sg13g2_nor2_1 _26450_ (.A(_12197_),
    .B(_13633_),
    .Y(_06281_));
 sg13g2_nor2_1 _26451_ (.A(_12362_),
    .B(net517),
    .Y(_06282_));
 sg13g2_and2_1 _26452_ (.A(_12739_),
    .B(net477),
    .X(_06283_));
 sg13g2_buf_1 _26453_ (.A(_06283_),
    .X(_06284_));
 sg13g2_xnor2_1 _26454_ (.Y(_06285_),
    .A(_06282_),
    .B(_06284_));
 sg13g2_xnor2_1 _26455_ (.Y(_06286_),
    .A(_06281_),
    .B(_06285_));
 sg13g2_a21oi_1 _26456_ (.A1(_06146_),
    .A2(_06149_),
    .Y(_06287_),
    .B1(_06147_));
 sg13g2_nor2_1 _26457_ (.A(_06146_),
    .B(_06149_),
    .Y(_06288_));
 sg13g2_nor2_1 _26458_ (.A(_06287_),
    .B(_06288_),
    .Y(_06289_));
 sg13g2_xnor2_1 _26459_ (.Y(_06290_),
    .A(_06286_),
    .B(_06289_));
 sg13g2_xnor2_1 _26460_ (.Y(_06291_),
    .A(_06280_),
    .B(_06290_));
 sg13g2_o21ai_1 _26461_ (.B1(_06156_),
    .Y(_06292_),
    .A1(_06145_),
    .A2(_06155_));
 sg13g2_buf_1 _26462_ (.A(_06292_),
    .X(_06293_));
 sg13g2_xor2_1 _26463_ (.B(_06293_),
    .A(_06291_),
    .X(_06294_));
 sg13g2_xnor2_1 _26464_ (.Y(_06295_),
    .A(_06274_),
    .B(_06294_));
 sg13g2_a21o_1 _26465_ (.A2(_06158_),
    .A1(_06140_),
    .B1(_06137_),
    .X(_06296_));
 sg13g2_o21ai_1 _26466_ (.B1(_06296_),
    .Y(_06297_),
    .A1(_06140_),
    .A2(_06158_));
 sg13g2_buf_1 _26467_ (.A(_06297_),
    .X(_06298_));
 sg13g2_xnor2_1 _26468_ (.Y(_06299_),
    .A(_06295_),
    .B(_06298_));
 sg13g2_xnor2_1 _26469_ (.Y(_06300_),
    .A(_06260_),
    .B(_06299_));
 sg13g2_o21ai_1 _26470_ (.B1(_06121_),
    .Y(_06301_),
    .A1(_06160_),
    .A2(_06163_));
 sg13g2_inv_1 _26471_ (.Y(_06302_),
    .A(_06301_));
 sg13g2_a21oi_2 _26472_ (.B1(_06302_),
    .Y(_06303_),
    .A2(_06163_),
    .A1(_06160_));
 sg13g2_xor2_1 _26473_ (.B(_06303_),
    .A(_06300_),
    .X(_06304_));
 sg13g2_xnor2_1 _26474_ (.Y(_06305_),
    .A(_06236_),
    .B(_06304_));
 sg13g2_nor2_1 _26475_ (.A(_06165_),
    .B(_06168_),
    .Y(_06306_));
 sg13g2_nand2_1 _26476_ (.Y(_06307_),
    .A(_06165_),
    .B(_06168_));
 sg13g2_o21ai_1 _26477_ (.B1(_06307_),
    .Y(_06308_),
    .A1(_06099_),
    .A2(_06306_));
 sg13g2_buf_1 _26478_ (.A(_06308_),
    .X(_06309_));
 sg13g2_a21oi_1 _26479_ (.A1(_06070_),
    .A2(_06097_),
    .Y(_06310_),
    .B1(_06069_));
 sg13g2_nor2_1 _26480_ (.A(_06070_),
    .B(_06097_),
    .Y(_06311_));
 sg13g2_nor2_1 _26481_ (.A(_06310_),
    .B(_06311_),
    .Y(_06312_));
 sg13g2_o21ai_1 _26482_ (.B1(net521),
    .Y(_06313_),
    .A1(_12199_),
    .A2(_12403_));
 sg13g2_nand2_1 _26483_ (.Y(_06314_),
    .A(net235),
    .B(_06313_));
 sg13g2_nand2_1 _26484_ (.Y(_06315_),
    .A(net505),
    .B(_14086_));
 sg13g2_a21oi_1 _26485_ (.A1(_06314_),
    .A2(_06315_),
    .Y(_06316_),
    .B1(net231));
 sg13g2_buf_1 _26486_ (.A(_06316_),
    .X(_06317_));
 sg13g2_xnor2_1 _26487_ (.Y(_06318_),
    .A(_06312_),
    .B(net136));
 sg13g2_xor2_1 _26488_ (.B(_06318_),
    .A(_06309_),
    .X(_06319_));
 sg13g2_xnor2_1 _26489_ (.Y(_06320_),
    .A(_06305_),
    .B(_06319_));
 sg13g2_xor2_1 _26490_ (.B(_06320_),
    .A(_06208_),
    .X(_06321_));
 sg13g2_xnor2_1 _26491_ (.Y(_06322_),
    .A(_06207_),
    .B(_06321_));
 sg13g2_nand2_1 _26492_ (.Y(_06323_),
    .A(_06065_),
    .B(_06182_));
 sg13g2_nand2_1 _26493_ (.Y(_06324_),
    .A(_06181_),
    .B(_06323_));
 sg13g2_xnor2_1 _26494_ (.Y(_06325_),
    .A(_06322_),
    .B(_06324_));
 sg13g2_xnor2_1 _26495_ (.Y(_06326_),
    .A(_06202_),
    .B(_06325_));
 sg13g2_nor3_1 _26496_ (.A(net700),
    .B(net69),
    .C(_06326_),
    .Y(_06327_));
 sg13g2_a221oi_1 _26497_ (.B2(_11471_),
    .C1(_06327_),
    .B1(_06201_),
    .A1(_11228_),
    .Y(_06328_),
    .A2(net68));
 sg13g2_nor2_1 _26498_ (.A(net682),
    .B(_06328_),
    .Y(_01745_));
 sg13g2_or2_1 _26499_ (.X(_06329_),
    .B(_06324_),
    .A(_06322_));
 sg13g2_o21ai_1 _26500_ (.B1(_06191_),
    .Y(_06330_),
    .A1(_06064_),
    .A2(_06189_));
 sg13g2_and2_1 _26501_ (.A(_06322_),
    .B(_06324_),
    .X(_06331_));
 sg13g2_a21oi_1 _26502_ (.A1(_06329_),
    .A2(_06330_),
    .Y(_06332_),
    .B1(_06331_));
 sg13g2_nand2_1 _26503_ (.Y(_06333_),
    .A(_06309_),
    .B(_06318_));
 sg13g2_o21ai_1 _26504_ (.B1(_06305_),
    .Y(_06334_),
    .A1(_06309_),
    .A2(_06318_));
 sg13g2_nand2_1 _26505_ (.Y(_06335_),
    .A(_06333_),
    .B(_06334_));
 sg13g2_a21o_1 _26506_ (.A2(_06315_),
    .A1(_06314_),
    .B1(net231),
    .X(_06336_));
 sg13g2_buf_2 _26507_ (.A(_06336_),
    .X(_06337_));
 sg13g2_nor3_1 _26508_ (.A(_06310_),
    .B(_06311_),
    .C(_06337_),
    .Y(_06338_));
 sg13g2_nand2_1 _26509_ (.Y(_06339_),
    .A(_06300_),
    .B(_06303_));
 sg13g2_nor2_1 _26510_ (.A(_06300_),
    .B(_06303_),
    .Y(_06340_));
 sg13g2_a21oi_1 _26511_ (.A1(_06236_),
    .A2(_06339_),
    .Y(_06341_),
    .B1(_06340_));
 sg13g2_nor2_1 _26512_ (.A(_06084_),
    .B(_06086_),
    .Y(_06342_));
 sg13g2_o21ai_1 _26513_ (.B1(_06342_),
    .Y(_06343_),
    .A1(_06216_),
    .A2(_06228_));
 sg13g2_nand2_1 _26514_ (.Y(_06344_),
    .A(_06095_),
    .B(_06228_));
 sg13g2_nand3_1 _26515_ (.B(_06086_),
    .C(_06344_),
    .A(_06084_),
    .Y(_06345_));
 sg13g2_a22oi_1 _26516_ (.Y(_06346_),
    .B1(_06343_),
    .B2(_06345_),
    .A2(_06080_),
    .A1(_06076_));
 sg13g2_nor2_1 _26517_ (.A(_06076_),
    .B(_06080_),
    .Y(_06347_));
 sg13g2_nor2_1 _26518_ (.A(_06216_),
    .B(_06347_),
    .Y(_06348_));
 sg13g2_xnor2_1 _26519_ (.Y(_06349_),
    .A(_06086_),
    .B(_06228_));
 sg13g2_nand2_1 _26520_ (.Y(_06350_),
    .A(_06216_),
    .B(_06347_));
 sg13g2_o21ai_1 _26521_ (.B1(_06350_),
    .Y(_06351_),
    .A1(_06348_),
    .A2(_06349_));
 sg13g2_nor2_1 _26522_ (.A(_06346_),
    .B(_06351_),
    .Y(_06352_));
 sg13g2_xnor2_1 _26523_ (.Y(_06353_),
    .A(net205),
    .B(net262));
 sg13g2_nand2_1 _26524_ (.Y(_06354_),
    .A(net212),
    .B(_06353_));
 sg13g2_xnor2_1 _26525_ (.Y(_06355_),
    .A(_06225_),
    .B(_06354_));
 sg13g2_a21oi_1 _26526_ (.A1(_06220_),
    .A2(_06223_),
    .Y(_06356_),
    .B1(_06355_));
 sg13g2_nor2_1 _26527_ (.A(_06220_),
    .B(_06223_),
    .Y(_06357_));
 sg13g2_nor2_1 _26528_ (.A(_06356_),
    .B(_06357_),
    .Y(_06358_));
 sg13g2_nand2_1 _26529_ (.Y(_06359_),
    .A(_06245_),
    .B(_06246_));
 sg13g2_nand2_1 _26530_ (.Y(_06360_),
    .A(_06243_),
    .B(_06359_));
 sg13g2_o21ai_1 _26531_ (.B1(_06360_),
    .Y(_06361_),
    .A1(_06245_),
    .A2(_06246_));
 sg13g2_buf_1 _26532_ (.A(_06361_),
    .X(_06362_));
 sg13g2_o21ai_1 _26533_ (.B1(net210),
    .Y(_06363_),
    .A1(_13920_),
    .A2(_13904_));
 sg13g2_o21ai_1 _26534_ (.B1(_06363_),
    .Y(_06364_),
    .A1(net279),
    .A2(_13913_));
 sg13g2_xnor2_1 _26535_ (.Y(_06365_),
    .A(_12071_),
    .B(_06353_));
 sg13g2_and2_1 _26536_ (.A(_13910_),
    .B(_06365_),
    .X(_06366_));
 sg13g2_buf_2 _26537_ (.A(_06366_),
    .X(_06367_));
 sg13g2_nand2_1 _26538_ (.Y(_06368_),
    .A(net205),
    .B(net237));
 sg13g2_o21ai_1 _26539_ (.B1(_13049_),
    .Y(_06369_),
    .A1(_13920_),
    .A2(net237));
 sg13g2_a21oi_1 _26540_ (.A1(_06368_),
    .A2(_06369_),
    .Y(_06370_),
    .B1(_13676_));
 sg13g2_buf_1 _26541_ (.A(_06370_),
    .X(_06371_));
 sg13g2_nor2_1 _26542_ (.A(_06367_),
    .B(net117),
    .Y(_06372_));
 sg13g2_a21oi_1 _26543_ (.A1(net237),
    .A2(_06364_),
    .Y(_06373_),
    .B1(_06372_));
 sg13g2_xnor2_1 _26544_ (.Y(_06374_),
    .A(_06362_),
    .B(_06373_));
 sg13g2_xnor2_1 _26545_ (.Y(_06375_),
    .A(_06095_),
    .B(_06374_));
 sg13g2_xnor2_1 _26546_ (.Y(_06376_),
    .A(_06358_),
    .B(_06375_));
 sg13g2_nand2_1 _26547_ (.Y(_06377_),
    .A(_06255_),
    .B(_06258_));
 sg13g2_nor2_1 _26548_ (.A(_06255_),
    .B(_06258_),
    .Y(_06378_));
 sg13g2_a21oi_2 _26549_ (.B1(_06378_),
    .Y(_06379_),
    .A2(_06377_),
    .A1(_06240_));
 sg13g2_xnor2_1 _26550_ (.Y(_06380_),
    .A(_06376_),
    .B(_06379_));
 sg13g2_xnor2_1 _26551_ (.Y(_06381_),
    .A(_06352_),
    .B(_06380_));
 sg13g2_nor2_1 _26552_ (.A(_06248_),
    .B(_06253_),
    .Y(_06382_));
 sg13g2_nor2_1 _26553_ (.A(_06242_),
    .B(_06382_),
    .Y(_06383_));
 sg13g2_a21oi_1 _26554_ (.A1(_06248_),
    .A2(_06253_),
    .Y(_06384_),
    .B1(_06383_));
 sg13g2_nand2_1 _26555_ (.Y(_06385_),
    .A(_06249_),
    .B(_06251_));
 sg13g2_nand2_1 _26556_ (.Y(_06386_),
    .A(_06250_),
    .B(_06385_));
 sg13g2_o21ai_1 _26557_ (.B1(_06386_),
    .Y(_06387_),
    .A1(_06249_),
    .A2(_06251_));
 sg13g2_nand2_1 _26558_ (.Y(_06388_),
    .A(net233),
    .B(net150));
 sg13g2_and2_1 _26559_ (.A(net232),
    .B(_13664_),
    .X(_06389_));
 sg13g2_buf_1 _26560_ (.A(_06389_),
    .X(_06390_));
 sg13g2_nand2_1 _26561_ (.Y(_06391_),
    .A(_14071_),
    .B(net149));
 sg13g2_xor2_1 _26562_ (.B(_06391_),
    .A(_06390_),
    .X(_06392_));
 sg13g2_xnor2_1 _26563_ (.Y(_06393_),
    .A(_06388_),
    .B(_06392_));
 sg13g2_nor2_1 _26564_ (.A(_12153_),
    .B(net207),
    .Y(_06394_));
 sg13g2_nand2_1 _26565_ (.Y(_06395_),
    .A(net500),
    .B(net172));
 sg13g2_nand2_1 _26566_ (.Y(_06396_),
    .A(_13791_),
    .B(net173));
 sg13g2_xor2_1 _26567_ (.B(_06396_),
    .A(_06395_),
    .X(_06397_));
 sg13g2_xnor2_1 _26568_ (.Y(_06398_),
    .A(_06394_),
    .B(_06397_));
 sg13g2_xnor2_1 _26569_ (.Y(_06399_),
    .A(_06393_),
    .B(_06398_));
 sg13g2_xnor2_1 _26570_ (.Y(_06400_),
    .A(_06387_),
    .B(_06399_));
 sg13g2_nor2_1 _26571_ (.A(_06268_),
    .B(_06272_),
    .Y(_06401_));
 sg13g2_nor2_1 _26572_ (.A(_06265_),
    .B(_06401_),
    .Y(_06402_));
 sg13g2_a21oi_2 _26573_ (.B1(_06402_),
    .Y(_06403_),
    .A2(_06272_),
    .A1(_06268_));
 sg13g2_xnor2_1 _26574_ (.Y(_06404_),
    .A(_06400_),
    .B(_06403_));
 sg13g2_xnor2_1 _26575_ (.Y(_06405_),
    .A(_06384_),
    .B(_06404_));
 sg13g2_nand2_1 _26576_ (.Y(_06406_),
    .A(_06261_),
    .B(_06263_));
 sg13g2_o21ai_1 _26577_ (.B1(_06262_),
    .Y(_06407_),
    .A1(_06261_),
    .A2(_06263_));
 sg13g2_and2_1 _26578_ (.A(_06406_),
    .B(_06407_),
    .X(_06408_));
 sg13g2_nand2_1 _26579_ (.Y(_06409_),
    .A(net256),
    .B(net501));
 sg13g2_and2_1 _26580_ (.A(_01812_),
    .B(_01841_),
    .X(_06410_));
 sg13g2_buf_1 _26581_ (.A(_06410_),
    .X(_06411_));
 sg13g2_nor2_1 _26582_ (.A(net503),
    .B(net258),
    .Y(_06412_));
 sg13g2_xor2_1 _26583_ (.B(_06412_),
    .A(_06411_),
    .X(_06413_));
 sg13g2_xnor2_1 _26584_ (.Y(_06414_),
    .A(_06409_),
    .B(_06413_));
 sg13g2_nor2b_1 _26585_ (.A(_06276_),
    .B_N(_06278_),
    .Y(_06415_));
 sg13g2_nand3_1 _26586_ (.B(net469),
    .C(_06276_),
    .A(_01839_),
    .Y(_06416_));
 sg13g2_o21ai_1 _26587_ (.B1(_06416_),
    .Y(_06417_),
    .A1(_06277_),
    .A2(_06415_));
 sg13g2_or2_1 _26588_ (.X(_06418_),
    .B(_06417_),
    .A(_06414_));
 sg13g2_nand2_1 _26589_ (.Y(_06419_),
    .A(_06414_),
    .B(_06417_));
 sg13g2_nand2_1 _26590_ (.Y(_06420_),
    .A(_06418_),
    .B(_06419_));
 sg13g2_xnor2_1 _26591_ (.Y(_06421_),
    .A(_06408_),
    .B(_06420_));
 sg13g2_and2_1 _26592_ (.A(_06125_),
    .B(net482),
    .X(_06422_));
 sg13g2_buf_1 _26593_ (.A(_06422_),
    .X(_06423_));
 sg13g2_nand2_1 _26594_ (.Y(_06424_),
    .A(net288),
    .B(net478));
 sg13g2_and2_1 _26595_ (.A(net300),
    .B(_13391_),
    .X(_06425_));
 sg13g2_buf_1 _26596_ (.A(_06425_),
    .X(_06426_));
 sg13g2_xor2_1 _26597_ (.B(_06426_),
    .A(_06424_),
    .X(_06427_));
 sg13g2_xnor2_1 _26598_ (.Y(_06428_),
    .A(_06423_),
    .B(_06427_));
 sg13g2_nand2_1 _26599_ (.Y(_06429_),
    .A(net301),
    .B(net480));
 sg13g2_nor2_1 _26600_ (.A(_12739_),
    .B(net517),
    .Y(_06430_));
 sg13g2_and2_1 _26601_ (.A(_13216_),
    .B(net477),
    .X(_06431_));
 sg13g2_buf_1 _26602_ (.A(_06431_),
    .X(_06432_));
 sg13g2_xor2_1 _26603_ (.B(_06432_),
    .A(_06430_),
    .X(_06433_));
 sg13g2_xnor2_1 _26604_ (.Y(_06434_),
    .A(_06429_),
    .B(_06433_));
 sg13g2_a21oi_1 _26605_ (.A1(_06281_),
    .A2(_06284_),
    .Y(_06435_),
    .B1(_06282_));
 sg13g2_nor2_1 _26606_ (.A(_06281_),
    .B(_06284_),
    .Y(_06436_));
 sg13g2_nor2_1 _26607_ (.A(_06435_),
    .B(_06436_),
    .Y(_06437_));
 sg13g2_xnor2_1 _26608_ (.Y(_06438_),
    .A(_06434_),
    .B(_06437_));
 sg13g2_xnor2_1 _26609_ (.Y(_06439_),
    .A(_06428_),
    .B(_06438_));
 sg13g2_nor2_1 _26610_ (.A(_06286_),
    .B(_06289_),
    .Y(_06440_));
 sg13g2_a21oi_1 _26611_ (.A1(_06286_),
    .A2(_06289_),
    .Y(_06441_),
    .B1(_06280_));
 sg13g2_nor2_1 _26612_ (.A(_06440_),
    .B(_06441_),
    .Y(_06442_));
 sg13g2_xnor2_1 _26613_ (.Y(_06443_),
    .A(_06439_),
    .B(_06442_));
 sg13g2_xnor2_1 _26614_ (.Y(_06444_),
    .A(_06421_),
    .B(_06443_));
 sg13g2_nand2_1 _26615_ (.Y(_06445_),
    .A(_06291_),
    .B(_06293_));
 sg13g2_nor2_1 _26616_ (.A(_06291_),
    .B(_06293_),
    .Y(_06446_));
 sg13g2_a21oi_1 _26617_ (.A1(_06274_),
    .A2(_06445_),
    .Y(_06447_),
    .B1(_06446_));
 sg13g2_nor2_1 _26618_ (.A(_06444_),
    .B(_06447_),
    .Y(_06448_));
 sg13g2_nand2_1 _26619_ (.Y(_06449_),
    .A(_06444_),
    .B(_06447_));
 sg13g2_nor2b_1 _26620_ (.A(_06448_),
    .B_N(_06449_),
    .Y(_06450_));
 sg13g2_xnor2_1 _26621_ (.Y(_06451_),
    .A(_06405_),
    .B(_06450_));
 sg13g2_inv_1 _26622_ (.Y(_06452_),
    .A(_06295_));
 sg13g2_nand2_1 _26623_ (.Y(_06453_),
    .A(_06452_),
    .B(_06298_));
 sg13g2_nor2_1 _26624_ (.A(_06452_),
    .B(_06298_),
    .Y(_06454_));
 sg13g2_a21oi_1 _26625_ (.A1(_06260_),
    .A2(_06453_),
    .Y(_06455_),
    .B1(_06454_));
 sg13g2_xor2_1 _26626_ (.B(_06455_),
    .A(_06451_),
    .X(_06456_));
 sg13g2_xnor2_1 _26627_ (.Y(_06457_),
    .A(_06381_),
    .B(_06456_));
 sg13g2_nand2_1 _26628_ (.Y(_06458_),
    .A(_06230_),
    .B(_06234_));
 sg13g2_nor2_1 _26629_ (.A(_06230_),
    .B(_06234_),
    .Y(_06459_));
 sg13g2_a21oi_1 _26630_ (.A1(_06211_),
    .A2(_06458_),
    .Y(_06460_),
    .B1(_06459_));
 sg13g2_xnor2_1 _26631_ (.Y(_06461_),
    .A(net136),
    .B(_06460_));
 sg13g2_xnor2_1 _26632_ (.Y(_06462_),
    .A(_06457_),
    .B(_06461_));
 sg13g2_xnor2_1 _26633_ (.Y(_06463_),
    .A(_06341_),
    .B(_06462_));
 sg13g2_xnor2_1 _26634_ (.Y(_06464_),
    .A(_06338_),
    .B(_06463_));
 sg13g2_xnor2_1 _26635_ (.Y(_06465_),
    .A(_06335_),
    .B(_06464_));
 sg13g2_o21ai_1 _26636_ (.B1(_06208_),
    .Y(_06466_),
    .A1(_06207_),
    .A2(_06320_));
 sg13g2_nand2_1 _26637_ (.Y(_06467_),
    .A(_06207_),
    .B(_06320_));
 sg13g2_nand2_1 _26638_ (.Y(_06468_),
    .A(_06466_),
    .B(_06467_));
 sg13g2_xnor2_1 _26639_ (.Y(_06469_),
    .A(_06465_),
    .B(_06468_));
 sg13g2_xnor2_1 _26640_ (.Y(_06470_),
    .A(_06332_),
    .B(_06469_));
 sg13g2_nand2_1 _26641_ (.Y(_06471_),
    .A(net60),
    .B(_06470_));
 sg13g2_nor2_1 _26642_ (.A(_05798_),
    .B(_06198_),
    .Y(_06472_));
 sg13g2_a21oi_1 _26643_ (.A1(_05798_),
    .A2(_06198_),
    .Y(_06473_),
    .B1(_11228_));
 sg13g2_nor2_1 _26644_ (.A(_06472_),
    .B(_06473_),
    .Y(_06474_));
 sg13g2_xnor2_1 _26645_ (.Y(_06475_),
    .A(_05801_),
    .B(_06474_));
 sg13g2_nor3_1 _26646_ (.A(_11227_),
    .B(net71),
    .C(_06475_),
    .Y(_06476_));
 sg13g2_a21o_1 _26647_ (.A2(_06475_),
    .A1(_11227_),
    .B1(_06476_),
    .X(_06477_));
 sg13g2_a22oi_1 _26648_ (.Y(_06478_),
    .B1(_06477_),
    .B2(net619),
    .A2(net61),
    .A1(_11227_));
 sg13g2_a21oi_1 _26649_ (.A1(_06471_),
    .A2(_06478_),
    .Y(_01746_),
    .B1(net618));
 sg13g2_nor2_1 _26650_ (.A(_06465_),
    .B(_06468_),
    .Y(_06479_));
 sg13g2_o21ai_1 _26651_ (.B1(_06329_),
    .Y(_06480_),
    .A1(_06202_),
    .A2(_06331_));
 sg13g2_nor2b_1 _26652_ (.A(_06479_),
    .B_N(_06480_),
    .Y(_06481_));
 sg13g2_nand2_1 _26653_ (.Y(_06482_),
    .A(_06465_),
    .B(_06468_));
 sg13g2_nor2b_1 _26654_ (.A(_06481_),
    .B_N(_06482_),
    .Y(_06483_));
 sg13g2_nor2_1 _26655_ (.A(_06335_),
    .B(_06463_),
    .Y(_06484_));
 sg13g2_nand2_1 _26656_ (.Y(_06485_),
    .A(_06335_),
    .B(_06463_));
 sg13g2_o21ai_1 _26657_ (.B1(_06485_),
    .Y(_06486_),
    .A1(_06338_),
    .A2(_06484_));
 sg13g2_buf_1 _26658_ (.A(_06486_),
    .X(_06487_));
 sg13g2_a21o_1 _26659_ (.A2(_06461_),
    .A1(_06457_),
    .B1(_06341_),
    .X(_06488_));
 sg13g2_o21ai_1 _26660_ (.B1(_06488_),
    .Y(_06489_),
    .A1(_06457_),
    .A2(_06461_));
 sg13g2_buf_1 _26661_ (.A(_06489_),
    .X(_06490_));
 sg13g2_and2_1 _26662_ (.A(net136),
    .B(_06460_),
    .X(_06491_));
 sg13g2_nand2b_1 _26663_ (.Y(_06492_),
    .B(_06451_),
    .A_N(_06455_));
 sg13g2_nor2b_1 _26664_ (.A(_06451_),
    .B_N(_06455_),
    .Y(_06493_));
 sg13g2_a21oi_2 _26665_ (.B1(_06493_),
    .Y(_06494_),
    .A2(_06492_),
    .A1(_06381_));
 sg13g2_inv_1 _26666_ (.Y(_06495_),
    .A(_06379_));
 sg13g2_inv_1 _26667_ (.Y(_06496_),
    .A(_06376_));
 sg13g2_o21ai_1 _26668_ (.B1(_06352_),
    .Y(_06497_),
    .A1(_06496_),
    .A2(_06379_));
 sg13g2_o21ai_1 _26669_ (.B1(_06497_),
    .Y(_06498_),
    .A1(_06376_),
    .A2(_06495_));
 sg13g2_buf_1 _26670_ (.A(_06498_),
    .X(_06499_));
 sg13g2_inv_1 _26671_ (.Y(_06500_),
    .A(_06358_));
 sg13g2_a21oi_1 _26672_ (.A1(_06500_),
    .A2(_06374_),
    .Y(_06501_),
    .B1(net89));
 sg13g2_nor2_1 _26673_ (.A(_06500_),
    .B(_06374_),
    .Y(_06502_));
 sg13g2_nor2_1 _26674_ (.A(_06501_),
    .B(_06502_),
    .Y(_06503_));
 sg13g2_inv_1 _26675_ (.Y(_06504_),
    .A(_06400_));
 sg13g2_nand2_1 _26676_ (.Y(_06505_),
    .A(_06504_),
    .B(_06403_));
 sg13g2_nor2_1 _26677_ (.A(_06504_),
    .B(_06403_),
    .Y(_06506_));
 sg13g2_a21oi_2 _26678_ (.B1(_06506_),
    .Y(_06507_),
    .A2(_06505_),
    .A1(_06384_));
 sg13g2_nand2_1 _26679_ (.Y(_06508_),
    .A(_06362_),
    .B(_06368_));
 sg13g2_nand3_1 _26680_ (.B(net206),
    .C(_06353_),
    .A(_13160_),
    .Y(_06509_));
 sg13g2_nor2_1 _26681_ (.A(net205),
    .B(_13160_),
    .Y(_06510_));
 sg13g2_o21ai_1 _26682_ (.B1(_12388_),
    .Y(_06511_),
    .A1(_06362_),
    .A2(_06510_));
 sg13g2_and4_1 _26683_ (.A(net212),
    .B(_06508_),
    .C(_06509_),
    .D(_06511_),
    .X(_06512_));
 sg13g2_nand3_1 _26684_ (.B(net149),
    .C(_06390_),
    .A(net204),
    .Y(_06513_));
 sg13g2_nor2b_1 _26685_ (.A(_06390_),
    .B_N(_06391_),
    .Y(_06514_));
 sg13g2_a21oi_1 _26686_ (.A1(_06388_),
    .A2(_06513_),
    .Y(_06515_),
    .B1(_06514_));
 sg13g2_buf_2 _26687_ (.A(_06515_),
    .X(_06516_));
 sg13g2_xnor2_1 _26688_ (.Y(_06517_),
    .A(_06512_),
    .B(_06516_));
 sg13g2_xnor2_1 _26689_ (.Y(_06518_),
    .A(_06507_),
    .B(_06517_));
 sg13g2_xnor2_1 _26690_ (.Y(_06519_),
    .A(_06503_),
    .B(_06518_));
 sg13g2_buf_1 _26691_ (.A(net172),
    .X(_06520_));
 sg13g2_nand3_1 _26692_ (.B(net135),
    .C(_06394_),
    .A(net500),
    .Y(_06521_));
 sg13g2_a21oi_1 _26693_ (.A1(_13789_),
    .A2(net135),
    .Y(_06522_),
    .B1(_06394_));
 sg13g2_a21oi_1 _26694_ (.A1(_06396_),
    .A2(_06521_),
    .Y(_06523_),
    .B1(_06522_));
 sg13g2_nand2_1 _26695_ (.Y(_06524_),
    .A(net233),
    .B(net212));
 sg13g2_nand2_1 _26696_ (.Y(_06525_),
    .A(net232),
    .B(net149));
 sg13g2_nand2_1 _26697_ (.Y(_06526_),
    .A(net204),
    .B(net150));
 sg13g2_xnor2_1 _26698_ (.Y(_06527_),
    .A(_06525_),
    .B(_06526_));
 sg13g2_xnor2_1 _26699_ (.Y(_06528_),
    .A(_06524_),
    .B(_06527_));
 sg13g2_nor2_1 _26700_ (.A(_12153_),
    .B(net208),
    .Y(_06529_));
 sg13g2_nand2_1 _26701_ (.Y(_06530_),
    .A(net500),
    .B(net173));
 sg13g2_nor2_1 _26702_ (.A(_12238_),
    .B(net207),
    .Y(_06531_));
 sg13g2_xnor2_1 _26703_ (.Y(_06532_),
    .A(_06530_),
    .B(_06531_));
 sg13g2_xnor2_1 _26704_ (.Y(_06533_),
    .A(_06529_),
    .B(_06532_));
 sg13g2_xnor2_1 _26705_ (.Y(_06534_),
    .A(_06528_),
    .B(_06533_));
 sg13g2_xnor2_1 _26706_ (.Y(_06535_),
    .A(_06523_),
    .B(_06534_));
 sg13g2_nand2_1 _26707_ (.Y(_06536_),
    .A(_06408_),
    .B(_06418_));
 sg13g2_nor2_1 _26708_ (.A(_06393_),
    .B(_06398_),
    .Y(_06537_));
 sg13g2_nand2_1 _26709_ (.Y(_06538_),
    .A(_06393_),
    .B(_06398_));
 sg13g2_o21ai_1 _26710_ (.B1(_06538_),
    .Y(_06539_),
    .A1(_06387_),
    .A2(_06537_));
 sg13g2_a21oi_1 _26711_ (.A1(_06419_),
    .A2(_06536_),
    .Y(_06540_),
    .B1(_06539_));
 sg13g2_nand3_1 _26712_ (.B(_06539_),
    .C(_06536_),
    .A(_06419_),
    .Y(_06541_));
 sg13g2_nor2b_1 _26713_ (.A(_06540_),
    .B_N(_06541_),
    .Y(_06542_));
 sg13g2_xnor2_1 _26714_ (.Y(_06543_),
    .A(_06535_),
    .B(_06542_));
 sg13g2_nor2_1 _26715_ (.A(_06411_),
    .B(_06412_),
    .Y(_06544_));
 sg13g2_nand2_1 _26716_ (.Y(_06545_),
    .A(_06411_),
    .B(_06412_));
 sg13g2_o21ai_1 _26717_ (.B1(_06545_),
    .Y(_06546_),
    .A1(_06409_),
    .A2(_06544_));
 sg13g2_nand2_1 _26718_ (.Y(_06547_),
    .A(net255),
    .B(net501));
 sg13g2_nor2_1 _26719_ (.A(_13179_),
    .B(_12729_),
    .Y(_06548_));
 sg13g2_nand2_1 _26720_ (.Y(_06549_),
    .A(net499),
    .B(net172));
 sg13g2_xnor2_1 _26721_ (.Y(_06550_),
    .A(_06548_),
    .B(_06549_));
 sg13g2_xnor2_1 _26722_ (.Y(_06551_),
    .A(_06547_),
    .B(_06550_));
 sg13g2_a22oi_1 _26723_ (.Y(_06552_),
    .B1(_06423_),
    .B2(_06426_),
    .A2(net478),
    .A1(net288));
 sg13g2_nor2_1 _26724_ (.A(_06423_),
    .B(_06426_),
    .Y(_06553_));
 sg13g2_nor2_1 _26725_ (.A(_06552_),
    .B(_06553_),
    .Y(_06554_));
 sg13g2_xnor2_1 _26726_ (.Y(_06555_),
    .A(_06551_),
    .B(_06554_));
 sg13g2_xnor2_1 _26727_ (.Y(_06556_),
    .A(_06546_),
    .B(_06555_));
 sg13g2_and2_1 _26728_ (.A(net256),
    .B(net482),
    .X(_06557_));
 sg13g2_buf_1 _26729_ (.A(_06557_),
    .X(_06558_));
 sg13g2_nand2_1 _26730_ (.Y(_06559_),
    .A(net300),
    .B(net478));
 sg13g2_nand2_1 _26731_ (.Y(_06560_),
    .A(net284),
    .B(net469));
 sg13g2_xnor2_1 _26732_ (.Y(_06561_),
    .A(_06559_),
    .B(_06560_));
 sg13g2_xnor2_1 _26733_ (.Y(_06562_),
    .A(_06558_),
    .B(_06561_));
 sg13g2_nand2_1 _26734_ (.Y(_06563_),
    .A(net288),
    .B(net480));
 sg13g2_or2_1 _26735_ (.X(_06564_),
    .B(net517),
    .A(_13216_));
 sg13g2_buf_1 _26736_ (.A(_06564_),
    .X(_06565_));
 sg13g2_nand2_1 _26737_ (.Y(_06566_),
    .A(_13221_),
    .B(net477));
 sg13g2_xor2_1 _26738_ (.B(_06566_),
    .A(_06565_),
    .X(_06567_));
 sg13g2_xor2_1 _26739_ (.B(_06567_),
    .A(_06563_),
    .X(_06568_));
 sg13g2_nor2_1 _26740_ (.A(_06430_),
    .B(_06432_),
    .Y(_06569_));
 sg13g2_nor2_1 _26741_ (.A(_06429_),
    .B(_06569_),
    .Y(_06570_));
 sg13g2_a21oi_1 _26742_ (.A1(_06430_),
    .A2(_06432_),
    .Y(_06571_),
    .B1(_06570_));
 sg13g2_nand2_1 _26743_ (.Y(_06572_),
    .A(_06568_),
    .B(_06571_));
 sg13g2_or2_1 _26744_ (.X(_06573_),
    .B(_06571_),
    .A(_06568_));
 sg13g2_nand2_1 _26745_ (.Y(_06574_),
    .A(_06572_),
    .B(_06573_));
 sg13g2_xnor2_1 _26746_ (.Y(_06575_),
    .A(_06562_),
    .B(_06574_));
 sg13g2_nor2_1 _26747_ (.A(_06434_),
    .B(_06437_),
    .Y(_06576_));
 sg13g2_a21oi_1 _26748_ (.A1(_06434_),
    .A2(_06437_),
    .Y(_06577_),
    .B1(_06428_));
 sg13g2_nor2_1 _26749_ (.A(_06576_),
    .B(_06577_),
    .Y(_06578_));
 sg13g2_xnor2_1 _26750_ (.Y(_06579_),
    .A(_06575_),
    .B(_06578_));
 sg13g2_xnor2_1 _26751_ (.Y(_06580_),
    .A(_06556_),
    .B(_06579_));
 sg13g2_nand2_1 _26752_ (.Y(_06581_),
    .A(_06439_),
    .B(_06442_));
 sg13g2_o21ai_1 _26753_ (.B1(_06421_),
    .Y(_06582_),
    .A1(_06439_),
    .A2(_06442_));
 sg13g2_nand2_1 _26754_ (.Y(_06583_),
    .A(_06581_),
    .B(_06582_));
 sg13g2_xor2_1 _26755_ (.B(_06583_),
    .A(_06580_),
    .X(_06584_));
 sg13g2_xnor2_1 _26756_ (.Y(_06585_),
    .A(_06543_),
    .B(_06584_));
 sg13g2_a21oi_2 _26757_ (.B1(_06448_),
    .Y(_06586_),
    .A2(_06449_),
    .A1(_06405_));
 sg13g2_xnor2_1 _26758_ (.Y(_06587_),
    .A(_06585_),
    .B(_06586_));
 sg13g2_xnor2_1 _26759_ (.Y(_06588_),
    .A(_06519_),
    .B(_06587_));
 sg13g2_nand2_1 _26760_ (.Y(_06589_),
    .A(net212),
    .B(_06365_));
 sg13g2_buf_1 _26761_ (.A(_06589_),
    .X(_06590_));
 sg13g2_xnor2_1 _26762_ (.Y(_06591_),
    .A(_06590_),
    .B(net117));
 sg13g2_xnor2_1 _26763_ (.Y(_06592_),
    .A(net89),
    .B(_06591_));
 sg13g2_buf_1 _26764_ (.A(_06592_),
    .X(_06593_));
 sg13g2_xnor2_1 _26765_ (.Y(_06594_),
    .A(net136),
    .B(net82));
 sg13g2_xor2_1 _26766_ (.B(_06594_),
    .A(_06588_),
    .X(_06595_));
 sg13g2_xnor2_1 _26767_ (.Y(_06596_),
    .A(_06499_),
    .B(_06595_));
 sg13g2_xnor2_1 _26768_ (.Y(_06597_),
    .A(_06494_),
    .B(_06596_));
 sg13g2_xor2_1 _26769_ (.B(_06597_),
    .A(_06491_),
    .X(_06598_));
 sg13g2_xnor2_1 _26770_ (.Y(_06599_),
    .A(_06490_),
    .B(_06598_));
 sg13g2_xnor2_1 _26771_ (.Y(_06600_),
    .A(_06487_),
    .B(_06599_));
 sg13g2_xnor2_1 _26772_ (.Y(_06601_),
    .A(_06483_),
    .B(_06600_));
 sg13g2_nand2b_1 _26773_ (.Y(_06602_),
    .B(_05996_),
    .A_N(_06601_));
 sg13g2_nor2_1 _26774_ (.A(_05801_),
    .B(_06474_),
    .Y(_06603_));
 sg13g2_a21oi_1 _26775_ (.A1(_05801_),
    .A2(_06474_),
    .Y(_06604_),
    .B1(_11227_));
 sg13g2_nor2_1 _26776_ (.A(_06603_),
    .B(_06604_),
    .Y(_06605_));
 sg13g2_xnor2_1 _26777_ (.Y(_06606_),
    .A(_05804_),
    .B(_06605_));
 sg13g2_nor3_1 _26778_ (.A(_11224_),
    .B(net71),
    .C(_06606_),
    .Y(_06607_));
 sg13g2_a21o_1 _26779_ (.A2(_06606_),
    .A1(_11224_),
    .B1(_06607_),
    .X(_06608_));
 sg13g2_a22oi_1 _26780_ (.Y(_06609_),
    .B1(_06608_),
    .B2(net619),
    .A2(net61),
    .A1(_11224_));
 sg13g2_a21oi_1 _26781_ (.A1(_06602_),
    .A2(_06609_),
    .Y(_01747_),
    .B1(net618));
 sg13g2_o21ai_1 _26782_ (.B1(_06482_),
    .Y(_06610_),
    .A1(_06487_),
    .A2(_06599_));
 sg13g2_nand2_1 _26783_ (.Y(_06611_),
    .A(_06487_),
    .B(_06599_));
 sg13g2_o21ai_1 _26784_ (.B1(_06611_),
    .Y(_06612_),
    .A1(_06481_),
    .A2(_06610_));
 sg13g2_buf_1 _26785_ (.A(_06612_),
    .X(_06613_));
 sg13g2_a21oi_1 _26786_ (.A1(_06490_),
    .A2(_06597_),
    .Y(_06614_),
    .B1(_06491_));
 sg13g2_nor2_1 _26787_ (.A(_06490_),
    .B(_06597_),
    .Y(_06615_));
 sg13g2_nor2_1 _26788_ (.A(_06614_),
    .B(_06615_),
    .Y(_06616_));
 sg13g2_buf_1 _26789_ (.A(_06616_),
    .X(_06617_));
 sg13g2_xnor2_1 _26790_ (.Y(_06618_),
    .A(_06337_),
    .B(_06499_));
 sg13g2_xnor2_1 _26791_ (.Y(_06619_),
    .A(_06588_),
    .B(net82));
 sg13g2_o21ai_1 _26792_ (.B1(_06619_),
    .Y(_06620_),
    .A1(_06494_),
    .A2(_06618_));
 sg13g2_nand2_1 _26793_ (.Y(_06621_),
    .A(_06494_),
    .B(_06618_));
 sg13g2_nand2_1 _26794_ (.Y(_06622_),
    .A(_06620_),
    .B(_06621_));
 sg13g2_and2_1 _26795_ (.A(net136),
    .B(_06499_),
    .X(_06623_));
 sg13g2_buf_1 _26796_ (.A(_06623_),
    .X(_06624_));
 sg13g2_inv_1 _26797_ (.Y(_06625_),
    .A(_06624_));
 sg13g2_nor2_1 _26798_ (.A(_06585_),
    .B(_06586_),
    .Y(_06626_));
 sg13g2_xor2_1 _26799_ (.B(net82),
    .A(_06519_),
    .X(_06627_));
 sg13g2_nand2_1 _26800_ (.Y(_06628_),
    .A(_06585_),
    .B(_06586_));
 sg13g2_o21ai_1 _26801_ (.B1(_06628_),
    .Y(_06629_),
    .A1(_06626_),
    .A2(_06627_));
 sg13g2_xnor2_1 _26802_ (.Y(_06630_),
    .A(_06517_),
    .B(net82));
 sg13g2_nand2_1 _26803_ (.Y(_06631_),
    .A(_06507_),
    .B(_06630_));
 sg13g2_nand2b_1 _26804_ (.Y(_06632_),
    .B(_06630_),
    .A_N(_06503_));
 sg13g2_nand2b_1 _26805_ (.Y(_06633_),
    .B(_06507_),
    .A_N(_06503_));
 sg13g2_and3_1 _26806_ (.X(_06634_),
    .A(_06631_),
    .B(_06632_),
    .C(_06633_));
 sg13g2_buf_1 _26807_ (.A(_06634_),
    .X(_06635_));
 sg13g2_xor2_1 _26808_ (.B(_06591_),
    .A(_06516_),
    .X(_06636_));
 sg13g2_nand2_1 _26809_ (.Y(_06637_),
    .A(net89),
    .B(_06636_));
 sg13g2_o21ai_1 _26810_ (.B1(_06512_),
    .Y(_06638_),
    .A1(net89),
    .A2(_06636_));
 sg13g2_and2_1 _26811_ (.A(_06637_),
    .B(_06638_),
    .X(_06639_));
 sg13g2_buf_1 _26812_ (.A(_06639_),
    .X(_06640_));
 sg13g2_o21ai_1 _26813_ (.B1(_06524_),
    .Y(_06641_),
    .A1(_06525_),
    .A2(_06526_));
 sg13g2_nand2_1 _26814_ (.Y(_06642_),
    .A(_06525_),
    .B(_06526_));
 sg13g2_and2_1 _26815_ (.A(_06641_),
    .B(_06642_),
    .X(_06643_));
 sg13g2_buf_1 _26816_ (.A(_06643_),
    .X(_06644_));
 sg13g2_inv_1 _26817_ (.Y(_06645_),
    .A(_06368_));
 sg13g2_o21ai_1 _26818_ (.B1(_13049_),
    .Y(_06646_),
    .A1(_06645_),
    .A2(_06516_));
 sg13g2_nand2b_1 _26819_ (.Y(_06647_),
    .B(_06516_),
    .A_N(_06510_));
 sg13g2_a21oi_1 _26820_ (.A1(_06646_),
    .A2(_06647_),
    .Y(_06648_),
    .B1(net231));
 sg13g2_xnor2_1 _26821_ (.Y(_06649_),
    .A(net84),
    .B(_06648_));
 sg13g2_a21o_1 _26822_ (.A2(_06541_),
    .A1(_06535_),
    .B1(_06540_),
    .X(_06650_));
 sg13g2_buf_1 _26823_ (.A(_06650_),
    .X(_06651_));
 sg13g2_xor2_1 _26824_ (.B(_06651_),
    .A(_06649_),
    .X(_06652_));
 sg13g2_xnor2_1 _26825_ (.Y(_06653_),
    .A(_06640_),
    .B(_06652_));
 sg13g2_nor2_1 _26826_ (.A(_06529_),
    .B(_06531_),
    .Y(_06654_));
 sg13g2_nand2_1 _26827_ (.Y(_06655_),
    .A(_06529_),
    .B(_06531_));
 sg13g2_o21ai_1 _26828_ (.B1(_06655_),
    .Y(_06656_),
    .A1(_06530_),
    .A2(_06654_));
 sg13g2_nand2_1 _26829_ (.Y(_06657_),
    .A(net232),
    .B(net150));
 sg13g2_xnor2_1 _26830_ (.Y(_06658_),
    .A(_14071_),
    .B(_13947_));
 sg13g2_nor2_1 _26831_ (.A(_01891_),
    .B(_06658_),
    .Y(_06659_));
 sg13g2_xnor2_1 _26832_ (.Y(_06660_),
    .A(_06657_),
    .B(_06659_));
 sg13g2_nand2_1 _26833_ (.Y(_06661_),
    .A(net236),
    .B(net149));
 sg13g2_nor2_1 _26834_ (.A(_12630_),
    .B(_13758_),
    .Y(_06662_));
 sg13g2_nand2_1 _26835_ (.Y(_06663_),
    .A(net234),
    .B(_13664_));
 sg13g2_xor2_1 _26836_ (.B(_06663_),
    .A(_06662_),
    .X(_06664_));
 sg13g2_xnor2_1 _26837_ (.Y(_06665_),
    .A(_06661_),
    .B(_06664_));
 sg13g2_xnor2_1 _26838_ (.Y(_06666_),
    .A(_06660_),
    .B(_06665_));
 sg13g2_xnor2_1 _26839_ (.Y(_06667_),
    .A(_06656_),
    .B(_06666_));
 sg13g2_nor2_1 _26840_ (.A(_06528_),
    .B(_06533_),
    .Y(_06668_));
 sg13g2_nand2_1 _26841_ (.Y(_06669_),
    .A(_06528_),
    .B(_06533_));
 sg13g2_o21ai_1 _26842_ (.B1(_06669_),
    .Y(_06670_),
    .A1(_06523_),
    .A2(_06668_));
 sg13g2_buf_1 _26843_ (.A(_06670_),
    .X(_06671_));
 sg13g2_nand2_1 _26844_ (.Y(_06672_),
    .A(_06551_),
    .B(_06554_));
 sg13g2_o21ai_1 _26845_ (.B1(_06546_),
    .Y(_06673_),
    .A1(_06551_),
    .A2(_06554_));
 sg13g2_nand2_2 _26846_ (.Y(_06674_),
    .A(_06672_),
    .B(_06673_));
 sg13g2_xnor2_1 _26847_ (.Y(_06675_),
    .A(_06671_),
    .B(_06674_));
 sg13g2_xnor2_1 _26848_ (.Y(_06676_),
    .A(_06667_),
    .B(_06675_));
 sg13g2_nand2_1 _26849_ (.Y(_06677_),
    .A(net499),
    .B(_13948_));
 sg13g2_nand2_1 _26850_ (.Y(_06678_),
    .A(net498),
    .B(_13954_));
 sg13g2_nor2_1 _26851_ (.A(net258),
    .B(_12979_),
    .Y(_06679_));
 sg13g2_xnor2_1 _26852_ (.Y(_06680_),
    .A(_06678_),
    .B(_06679_));
 sg13g2_xnor2_1 _26853_ (.Y(_06681_),
    .A(_06677_),
    .B(_06680_));
 sg13g2_a21oi_1 _26854_ (.A1(net499),
    .A2(net135),
    .Y(_06682_),
    .B1(_06548_));
 sg13g2_nand3_1 _26855_ (.B(net135),
    .C(_06548_),
    .A(_13807_),
    .Y(_06683_));
 sg13g2_o21ai_1 _26856_ (.B1(_06683_),
    .Y(_06684_),
    .A1(_06547_),
    .A2(_06682_));
 sg13g2_nor2b_1 _26857_ (.A(_06558_),
    .B_N(_06560_),
    .Y(_06685_));
 sg13g2_nand3_1 _26858_ (.B(net469),
    .C(_06558_),
    .A(net284),
    .Y(_06686_));
 sg13g2_o21ai_1 _26859_ (.B1(_06686_),
    .Y(_06687_),
    .A1(_06559_),
    .A2(_06685_));
 sg13g2_buf_1 _26860_ (.A(_06687_),
    .X(_06688_));
 sg13g2_xnor2_1 _26861_ (.Y(_06689_),
    .A(_06684_),
    .B(_06688_));
 sg13g2_xnor2_1 _26862_ (.Y(_06690_),
    .A(_06681_),
    .B(_06689_));
 sg13g2_nand2_1 _26863_ (.Y(_06691_),
    .A(net255),
    .B(_12987_));
 sg13g2_nand2_1 _26864_ (.Y(_06692_),
    .A(_06125_),
    .B(net478));
 sg13g2_nand2_1 _26865_ (.Y(_06693_),
    .A(net256),
    .B(net469));
 sg13g2_xnor2_1 _26866_ (.Y(_06694_),
    .A(_06692_),
    .B(_06693_));
 sg13g2_xnor2_1 _26867_ (.Y(_06695_),
    .A(_06691_),
    .B(_06694_));
 sg13g2_nand2_1 _26868_ (.Y(_06696_),
    .A(net300),
    .B(net480));
 sg13g2_or2_1 _26869_ (.X(_06697_),
    .B(_13712_),
    .A(_13221_));
 sg13g2_nand2_1 _26870_ (.Y(_06698_),
    .A(net288),
    .B(net477));
 sg13g2_xor2_1 _26871_ (.B(_06698_),
    .A(_06697_),
    .X(_06699_));
 sg13g2_xnor2_1 _26872_ (.Y(_06700_),
    .A(_06696_),
    .B(_06699_));
 sg13g2_a21o_1 _26873_ (.A2(_06565_),
    .A1(_06563_),
    .B1(_06566_),
    .X(_06701_));
 sg13g2_o21ai_1 _26874_ (.B1(_06701_),
    .Y(_06702_),
    .A1(_06563_),
    .A2(_06565_));
 sg13g2_nor2_1 _26875_ (.A(_06700_),
    .B(_06702_),
    .Y(_06703_));
 sg13g2_nand2_1 _26876_ (.Y(_06704_),
    .A(_06700_),
    .B(_06702_));
 sg13g2_nand2b_1 _26877_ (.Y(_06705_),
    .B(_06704_),
    .A_N(_06703_));
 sg13g2_xor2_1 _26878_ (.B(_06705_),
    .A(_06695_),
    .X(_06706_));
 sg13g2_nand2_1 _26879_ (.Y(_06707_),
    .A(_06562_),
    .B(_06572_));
 sg13g2_nand2_1 _26880_ (.Y(_06708_),
    .A(_06573_),
    .B(_06707_));
 sg13g2_xnor2_1 _26881_ (.Y(_06709_),
    .A(_06706_),
    .B(_06708_));
 sg13g2_xnor2_1 _26882_ (.Y(_06710_),
    .A(_06690_),
    .B(_06709_));
 sg13g2_nand2_1 _26883_ (.Y(_06711_),
    .A(_06575_),
    .B(_06578_));
 sg13g2_o21ai_1 _26884_ (.B1(_06556_),
    .Y(_06712_),
    .A1(_06575_),
    .A2(_06578_));
 sg13g2_nand2_1 _26885_ (.Y(_06713_),
    .A(_06711_),
    .B(_06712_));
 sg13g2_xor2_1 _26886_ (.B(_06713_),
    .A(_06710_),
    .X(_06714_));
 sg13g2_xnor2_1 _26887_ (.Y(_06715_),
    .A(_06676_),
    .B(_06714_));
 sg13g2_nand2_1 _26888_ (.Y(_06716_),
    .A(_06580_),
    .B(_06583_));
 sg13g2_nor2_1 _26889_ (.A(_06580_),
    .B(_06583_),
    .Y(_06717_));
 sg13g2_a21oi_1 _26890_ (.A1(_06543_),
    .A2(_06716_),
    .Y(_06718_),
    .B1(_06717_));
 sg13g2_xnor2_1 _26891_ (.Y(_06719_),
    .A(_06715_),
    .B(_06718_));
 sg13g2_xnor2_1 _26892_ (.Y(_06720_),
    .A(_06653_),
    .B(_06719_));
 sg13g2_xor2_1 _26893_ (.B(_06720_),
    .A(_06594_),
    .X(_06721_));
 sg13g2_xnor2_1 _26894_ (.Y(_06722_),
    .A(_06635_),
    .B(_06721_));
 sg13g2_xnor2_1 _26895_ (.Y(_06723_),
    .A(_06629_),
    .B(_06722_));
 sg13g2_xnor2_1 _26896_ (.Y(_06724_),
    .A(_06625_),
    .B(_06723_));
 sg13g2_xnor2_1 _26897_ (.Y(_06725_),
    .A(_06622_),
    .B(_06724_));
 sg13g2_xnor2_1 _26898_ (.Y(_06726_),
    .A(_06617_),
    .B(_06725_));
 sg13g2_xnor2_1 _26899_ (.Y(_06727_),
    .A(_06613_),
    .B(_06726_));
 sg13g2_nand2_1 _26900_ (.Y(_06728_),
    .A(net60),
    .B(_06727_));
 sg13g2_nor2_1 _26901_ (.A(_05804_),
    .B(_06605_),
    .Y(_06729_));
 sg13g2_a21oi_1 _26902_ (.A1(_05804_),
    .A2(_06605_),
    .Y(_06730_),
    .B1(_11224_));
 sg13g2_nor2_1 _26903_ (.A(_06729_),
    .B(_06730_),
    .Y(_06731_));
 sg13g2_xnor2_1 _26904_ (.Y(_06732_),
    .A(_05808_),
    .B(_06731_));
 sg13g2_nor3_1 _26905_ (.A(_11311_),
    .B(_11345_),
    .C(_06732_),
    .Y(_06733_));
 sg13g2_a21o_1 _26906_ (.A2(_06732_),
    .A1(_11311_),
    .B1(_06733_),
    .X(_06734_));
 sg13g2_a22oi_1 _26907_ (.Y(_06735_),
    .B1(_06734_),
    .B2(_05992_),
    .A2(_05988_),
    .A1(_11311_));
 sg13g2_a21oi_1 _26908_ (.A1(_06728_),
    .A2(_06735_),
    .Y(_01748_),
    .B1(net618));
 sg13g2_xnor2_1 _26909_ (.Y(_06736_),
    .A(_06593_),
    .B(_06720_));
 sg13g2_xnor2_1 _26910_ (.Y(_06737_),
    .A(_06337_),
    .B(_06635_));
 sg13g2_a21o_1 _26911_ (.A2(_06737_),
    .A1(_06736_),
    .B1(_06629_),
    .X(_06738_));
 sg13g2_o21ai_1 _26912_ (.B1(_06738_),
    .Y(_06739_),
    .A1(_06736_),
    .A2(_06737_));
 sg13g2_buf_1 _26913_ (.A(_06739_),
    .X(_06740_));
 sg13g2_nand2_1 _26914_ (.Y(_06741_),
    .A(net136),
    .B(_06635_));
 sg13g2_inv_1 _26915_ (.Y(_06742_),
    .A(_06718_));
 sg13g2_nor2_1 _26916_ (.A(_06715_),
    .B(_06742_),
    .Y(_06743_));
 sg13g2_xnor2_1 _26917_ (.Y(_06744_),
    .A(net82),
    .B(_06653_));
 sg13g2_a21oi_1 _26918_ (.A1(_06715_),
    .A2(_06742_),
    .Y(_06745_),
    .B1(_06744_));
 sg13g2_nor2_1 _26919_ (.A(_06743_),
    .B(_06745_),
    .Y(_06746_));
 sg13g2_inv_1 _26920_ (.Y(_06747_),
    .A(_06651_));
 sg13g2_inv_1 _26921_ (.Y(_06748_),
    .A(_06640_));
 sg13g2_xor2_1 _26922_ (.B(_06649_),
    .A(net82),
    .X(_06749_));
 sg13g2_a21oi_1 _26923_ (.A1(_06748_),
    .A2(_06651_),
    .Y(_06750_),
    .B1(_06749_));
 sg13g2_a21oi_2 _26924_ (.B1(_06750_),
    .Y(_06751_),
    .A2(_06747_),
    .A1(_06640_));
 sg13g2_a21oi_1 _26925_ (.A1(_06367_),
    .A2(net117),
    .Y(_06752_),
    .B1(net89));
 sg13g2_nand2b_1 _26926_ (.Y(_06753_),
    .B(_06516_),
    .A_N(net84));
 sg13g2_inv_1 _26927_ (.Y(_06754_),
    .A(net117));
 sg13g2_nor2b_1 _26928_ (.A(_06516_),
    .B_N(net84),
    .Y(_06755_));
 sg13g2_nor2_1 _26929_ (.A(_06367_),
    .B(_06644_),
    .Y(_06756_));
 sg13g2_a21oi_1 _26930_ (.A1(_06367_),
    .A2(_06755_),
    .Y(_06757_),
    .B1(_06756_));
 sg13g2_nor3_1 _26931_ (.A(net89),
    .B(_06590_),
    .C(net84),
    .Y(_06758_));
 sg13g2_a21oi_1 _26932_ (.A1(_06590_),
    .A2(_06755_),
    .Y(_06759_),
    .B1(_06758_));
 sg13g2_and2_1 _26933_ (.A(net117),
    .B(_06759_),
    .X(_06760_));
 sg13g2_a21oi_1 _26934_ (.A1(_06754_),
    .A2(_06757_),
    .Y(_06761_),
    .B1(_06760_));
 sg13g2_a21o_1 _26935_ (.A2(_06753_),
    .A1(_06752_),
    .B1(_06761_),
    .X(_06762_));
 sg13g2_buf_1 _26936_ (.A(_06762_),
    .X(_06763_));
 sg13g2_inv_1 _26937_ (.Y(_06764_),
    .A(_06671_));
 sg13g2_inv_1 _26938_ (.Y(_06765_),
    .A(_06674_));
 sg13g2_a21oi_1 _26939_ (.A1(_06671_),
    .A2(_06765_),
    .Y(_06766_),
    .B1(_06667_));
 sg13g2_a21oi_2 _26940_ (.B1(_06766_),
    .Y(_06767_),
    .A2(_06674_),
    .A1(_06764_));
 sg13g2_inv_1 _26941_ (.Y(_06768_),
    .A(_06657_));
 sg13g2_o21ai_1 _26942_ (.B1(_13947_),
    .Y(_06769_),
    .A1(net204),
    .A2(_06768_));
 sg13g2_nand2_1 _26943_ (.Y(_06770_),
    .A(net204),
    .B(_06768_));
 sg13g2_a21oi_1 _26944_ (.A1(_06769_),
    .A2(_06770_),
    .Y(_06771_),
    .B1(net231));
 sg13g2_buf_1 _26945_ (.A(_06771_),
    .X(_06772_));
 sg13g2_a21oi_1 _26946_ (.A1(_06367_),
    .A2(net84),
    .Y(_06773_),
    .B1(net117));
 sg13g2_nor2_1 _26947_ (.A(_06756_),
    .B(_06773_),
    .Y(_06774_));
 sg13g2_xnor2_1 _26948_ (.Y(_06775_),
    .A(net81),
    .B(_06774_));
 sg13g2_xnor2_1 _26949_ (.Y(_06776_),
    .A(_06767_),
    .B(_06775_));
 sg13g2_xnor2_1 _26950_ (.Y(_06777_),
    .A(_06763_),
    .B(_06776_));
 sg13g2_nand2_1 _26951_ (.Y(_06778_),
    .A(_06661_),
    .B(_06663_));
 sg13g2_nand2_1 _26952_ (.Y(_06779_),
    .A(_06662_),
    .B(_06778_));
 sg13g2_o21ai_1 _26953_ (.B1(_06779_),
    .Y(_06780_),
    .A1(_06661_),
    .A2(_06663_));
 sg13g2_xnor2_1 _26954_ (.Y(_06781_),
    .A(net232),
    .B(_06658_));
 sg13g2_nand2_1 _26955_ (.Y(_06782_),
    .A(net212),
    .B(_06781_));
 sg13g2_nand2_1 _26956_ (.Y(_06783_),
    .A(net236),
    .B(net150));
 sg13g2_nor2_1 _26957_ (.A(_12630_),
    .B(_13191_),
    .Y(_06784_));
 sg13g2_inv_1 _26958_ (.Y(_06785_),
    .A(_06784_));
 sg13g2_nand2_1 _26959_ (.Y(_06786_),
    .A(net234),
    .B(net149));
 sg13g2_xnor2_1 _26960_ (.Y(_06787_),
    .A(_06785_),
    .B(_06786_));
 sg13g2_xnor2_1 _26961_ (.Y(_06788_),
    .A(_06783_),
    .B(_06787_));
 sg13g2_xnor2_1 _26962_ (.Y(_06789_),
    .A(_06782_),
    .B(_06788_));
 sg13g2_xnor2_1 _26963_ (.Y(_06790_),
    .A(_06780_),
    .B(_06789_));
 sg13g2_inv_1 _26964_ (.Y(_06791_),
    .A(_06660_));
 sg13g2_nor2_1 _26965_ (.A(_06791_),
    .B(_06665_),
    .Y(_06792_));
 sg13g2_nand2_1 _26966_ (.Y(_06793_),
    .A(_06791_),
    .B(_06665_));
 sg13g2_o21ai_1 _26967_ (.B1(_06793_),
    .Y(_06794_),
    .A1(_06656_),
    .A2(_06792_));
 sg13g2_nor2_1 _26968_ (.A(_06681_),
    .B(_06688_),
    .Y(_06795_));
 sg13g2_a21oi_1 _26969_ (.A1(_06681_),
    .A2(_06688_),
    .Y(_06796_),
    .B1(_06684_));
 sg13g2_nor3_1 _26970_ (.A(_06794_),
    .B(_06795_),
    .C(_06796_),
    .Y(_06797_));
 sg13g2_o21ai_1 _26971_ (.B1(_06794_),
    .Y(_06798_),
    .A1(_06795_),
    .A2(_06796_));
 sg13g2_nor2b_1 _26972_ (.A(_06797_),
    .B_N(_06798_),
    .Y(_06799_));
 sg13g2_xnor2_1 _26973_ (.Y(_06800_),
    .A(_06790_),
    .B(_06799_));
 sg13g2_nor2_1 _26974_ (.A(net503),
    .B(net207),
    .Y(_06801_));
 sg13g2_nand2_1 _26975_ (.Y(_06802_),
    .A(_06520_),
    .B(_13368_));
 sg13g2_nand2_1 _26976_ (.Y(_06803_),
    .A(net498),
    .B(net173));
 sg13g2_xnor2_1 _26977_ (.Y(_06804_),
    .A(_06802_),
    .B(_06803_));
 sg13g2_xnor2_1 _26978_ (.Y(_06805_),
    .A(_06801_),
    .B(_06804_));
 sg13g2_a21oi_1 _26979_ (.A1(net498),
    .A2(_13954_),
    .Y(_06806_),
    .B1(_06679_));
 sg13g2_nand3_1 _26980_ (.B(_06520_),
    .C(_06679_),
    .A(net498),
    .Y(_06807_));
 sg13g2_o21ai_1 _26981_ (.B1(_06807_),
    .Y(_06808_),
    .A1(_06677_),
    .A2(_06806_));
 sg13g2_buf_1 _26982_ (.A(_06808_),
    .X(_06809_));
 sg13g2_nand2_1 _26983_ (.Y(_06810_),
    .A(_06691_),
    .B(_06693_));
 sg13g2_o21ai_1 _26984_ (.B1(_06692_),
    .Y(_06811_),
    .A1(_06691_),
    .A2(_06693_));
 sg13g2_and2_1 _26985_ (.A(_06810_),
    .B(_06811_),
    .X(_06812_));
 sg13g2_buf_1 _26986_ (.A(_06812_),
    .X(_06813_));
 sg13g2_xnor2_1 _26987_ (.Y(_06814_),
    .A(_06809_),
    .B(_06813_));
 sg13g2_xnor2_1 _26988_ (.Y(_06815_),
    .A(_06805_),
    .B(_06814_));
 sg13g2_nand2_1 _26989_ (.Y(_06816_),
    .A(_01810_),
    .B(_01846_));
 sg13g2_nand2_1 _26990_ (.Y(_06817_),
    .A(net255),
    .B(net469));
 sg13g2_nor2_1 _26991_ (.A(net258),
    .B(_13387_),
    .Y(_06818_));
 sg13g2_xnor2_1 _26992_ (.Y(_06819_),
    .A(_06817_),
    .B(_06818_));
 sg13g2_xnor2_1 _26993_ (.Y(_06820_),
    .A(_06816_),
    .B(_06819_));
 sg13g2_nand2_1 _26994_ (.Y(_06821_),
    .A(net284),
    .B(_13384_));
 sg13g2_or2_1 _26995_ (.X(_06822_),
    .B(_13712_),
    .A(net288));
 sg13g2_buf_1 _26996_ (.A(_06822_),
    .X(_06823_));
 sg13g2_nand2_1 _26997_ (.Y(_06824_),
    .A(_13788_),
    .B(_01863_));
 sg13g2_xor2_1 _26998_ (.B(_06824_),
    .A(_06823_),
    .X(_06825_));
 sg13g2_xnor2_1 _26999_ (.Y(_06826_),
    .A(_06821_),
    .B(_06825_));
 sg13g2_and2_1 _27000_ (.A(_06696_),
    .B(_06698_),
    .X(_06827_));
 sg13g2_or2_1 _27001_ (.X(_06828_),
    .B(_06698_),
    .A(_06696_));
 sg13g2_o21ai_1 _27002_ (.B1(_06828_),
    .Y(_06829_),
    .A1(_06697_),
    .A2(_06827_));
 sg13g2_buf_1 _27003_ (.A(_06829_),
    .X(_06830_));
 sg13g2_xnor2_1 _27004_ (.Y(_06831_),
    .A(_06826_),
    .B(_06830_));
 sg13g2_xnor2_1 _27005_ (.Y(_06832_),
    .A(_06820_),
    .B(_06831_));
 sg13g2_o21ai_1 _27006_ (.B1(_06704_),
    .Y(_06833_),
    .A1(_06695_),
    .A2(_06703_));
 sg13g2_buf_1 _27007_ (.A(_06833_),
    .X(_06834_));
 sg13g2_xnor2_1 _27008_ (.Y(_06835_),
    .A(_06832_),
    .B(_06834_));
 sg13g2_xnor2_1 _27009_ (.Y(_06836_),
    .A(_06815_),
    .B(_06835_));
 sg13g2_nand2_1 _27010_ (.Y(_06837_),
    .A(_06706_),
    .B(_06708_));
 sg13g2_o21ai_1 _27011_ (.B1(_06690_),
    .Y(_06838_),
    .A1(_06706_),
    .A2(_06708_));
 sg13g2_nand2_1 _27012_ (.Y(_06839_),
    .A(_06837_),
    .B(_06838_));
 sg13g2_xor2_1 _27013_ (.B(_06839_),
    .A(_06836_),
    .X(_06840_));
 sg13g2_xnor2_1 _27014_ (.Y(_06841_),
    .A(_06800_),
    .B(_06840_));
 sg13g2_nor2_1 _27015_ (.A(_06710_),
    .B(_06713_),
    .Y(_06842_));
 sg13g2_a21oi_1 _27016_ (.A1(_06710_),
    .A2(_06713_),
    .Y(_06843_),
    .B1(_06676_));
 sg13g2_nor2_2 _27017_ (.A(_06842_),
    .B(_06843_),
    .Y(_06844_));
 sg13g2_xnor2_1 _27018_ (.Y(_06845_),
    .A(_06841_),
    .B(_06844_));
 sg13g2_xnor2_1 _27019_ (.Y(_06846_),
    .A(_06777_),
    .B(_06845_));
 sg13g2_xnor2_1 _27020_ (.Y(_06847_),
    .A(_06594_),
    .B(_06846_));
 sg13g2_xnor2_1 _27021_ (.Y(_06848_),
    .A(_06751_),
    .B(_06847_));
 sg13g2_xnor2_1 _27022_ (.Y(_06849_),
    .A(_06746_),
    .B(_06848_));
 sg13g2_xnor2_1 _27023_ (.Y(_06850_),
    .A(_06741_),
    .B(_06849_));
 sg13g2_xnor2_1 _27024_ (.Y(_06851_),
    .A(_06740_),
    .B(_06850_));
 sg13g2_buf_1 _27025_ (.A(_06851_),
    .X(_06852_));
 sg13g2_nand2_1 _27026_ (.Y(_06853_),
    .A(_06622_),
    .B(_06723_));
 sg13g2_buf_1 _27027_ (.A(_06853_),
    .X(_06854_));
 sg13g2_inv_1 _27028_ (.Y(_06855_),
    .A(_06854_));
 sg13g2_nor2_1 _27029_ (.A(_06622_),
    .B(_06723_),
    .Y(_06856_));
 sg13g2_buf_1 _27030_ (.A(_06856_),
    .X(_06857_));
 sg13g2_o21ai_1 _27031_ (.B1(_06854_),
    .Y(_06858_),
    .A1(_06625_),
    .A2(_06857_));
 sg13g2_a221oi_1 _27032_ (.B2(_06617_),
    .C1(_06613_),
    .B1(_06858_),
    .A1(_06624_),
    .Y(_06859_),
    .A2(_06855_));
 sg13g2_a21oi_1 _27033_ (.A1(_06625_),
    .A2(_06854_),
    .Y(_06860_),
    .B1(_06857_));
 sg13g2_nor2_1 _27034_ (.A(_06617_),
    .B(_06860_),
    .Y(_06861_));
 sg13g2_a21oi_1 _27035_ (.A1(_06625_),
    .A2(_06857_),
    .Y(_06862_),
    .B1(_06861_));
 sg13g2_and2_1 _27036_ (.A(_06613_),
    .B(_06862_),
    .X(_06863_));
 sg13g2_nor2_1 _27037_ (.A(_06617_),
    .B(_06624_),
    .Y(_06864_));
 sg13g2_nand2_1 _27038_ (.Y(_06865_),
    .A(_06617_),
    .B(_06624_));
 sg13g2_nor2_1 _27039_ (.A(_06854_),
    .B(_06865_),
    .Y(_06866_));
 sg13g2_a21oi_1 _27040_ (.A1(_06857_),
    .A2(_06864_),
    .Y(_06867_),
    .B1(_06866_));
 sg13g2_o21ai_1 _27041_ (.B1(_06867_),
    .Y(_06868_),
    .A1(_06859_),
    .A2(_06863_));
 sg13g2_xor2_1 _27042_ (.B(_06868_),
    .A(_06852_),
    .X(_06869_));
 sg13g2_nand2_1 _27043_ (.Y(_06870_),
    .A(_05997_),
    .B(_06869_));
 sg13g2_nor2_1 _27044_ (.A(_05808_),
    .B(_06731_),
    .Y(_06871_));
 sg13g2_a21oi_1 _27045_ (.A1(_05808_),
    .A2(_06731_),
    .Y(_06872_),
    .B1(_11311_));
 sg13g2_nor2_1 _27046_ (.A(_06871_),
    .B(_06872_),
    .Y(_06873_));
 sg13g2_xnor2_1 _27047_ (.Y(_06874_),
    .A(_05811_),
    .B(_06873_));
 sg13g2_nor3_1 _27048_ (.A(_11219_),
    .B(_11345_),
    .C(_06874_),
    .Y(_06875_));
 sg13g2_a21o_1 _27049_ (.A2(_06874_),
    .A1(_11219_),
    .B1(_06875_),
    .X(_06876_));
 sg13g2_a22oi_1 _27050_ (.Y(_06877_),
    .B1(_06876_),
    .B2(net619),
    .A2(net61),
    .A1(_11219_));
 sg13g2_a21oi_1 _27051_ (.A1(_06870_),
    .A2(_06877_),
    .Y(_01749_),
    .B1(_05994_));
 sg13g2_xor2_1 _27052_ (.B(_12559_),
    .A(_12301_),
    .X(_06878_));
 sg13g2_xnor2_1 _27053_ (.Y(_06879_),
    .A(_05984_),
    .B(_06878_));
 sg13g2_nand2_1 _27054_ (.Y(_06880_),
    .A(net638),
    .B(_06879_));
 sg13g2_nand2_1 _27055_ (.Y(_06881_),
    .A(_11267_),
    .B(_12013_));
 sg13g2_xor2_1 _27056_ (.B(_12023_),
    .A(\rbzero.wall_tracer.trackDistX[-10] ),
    .X(_06882_));
 sg13g2_xnor2_1 _27057_ (.Y(_06883_),
    .A(_06881_),
    .B(_06882_));
 sg13g2_a21oi_1 _27058_ (.A1(net700),
    .A2(_06883_),
    .Y(_06884_),
    .B1(_11346_));
 sg13g2_a221oi_1 _27059_ (.B2(_06884_),
    .C1(net635),
    .B1(_06880_),
    .A1(_11266_),
    .Y(_01750_),
    .A2(_11344_));
 sg13g2_a21o_1 _27060_ (.A2(_06865_),
    .A1(_06613_),
    .B1(_06864_),
    .X(_06885_));
 sg13g2_o21ai_1 _27061_ (.B1(_06885_),
    .Y(_06886_),
    .A1(_06852_),
    .A2(_06857_));
 sg13g2_or2_1 _27062_ (.X(_06887_),
    .B(_06864_),
    .A(_06852_));
 sg13g2_nand3_1 _27063_ (.B(_06854_),
    .C(_06887_),
    .A(_06613_),
    .Y(_06888_));
 sg13g2_nand3_1 _27064_ (.B(_06854_),
    .C(_06865_),
    .A(_06852_),
    .Y(_06889_));
 sg13g2_nand2_1 _27065_ (.Y(_06890_),
    .A(_06852_),
    .B(_06857_));
 sg13g2_and4_1 _27066_ (.A(_06886_),
    .B(_06888_),
    .C(_06889_),
    .D(_06890_),
    .X(_06891_));
 sg13g2_xnor2_1 _27067_ (.Y(_06892_),
    .A(net82),
    .B(_06846_));
 sg13g2_xnor2_1 _27068_ (.Y(_06893_),
    .A(net136),
    .B(_06751_));
 sg13g2_a21o_1 _27069_ (.A2(_06893_),
    .A1(_06892_),
    .B1(_06746_),
    .X(_06894_));
 sg13g2_o21ai_1 _27070_ (.B1(_06894_),
    .Y(_06895_),
    .A1(_06892_),
    .A2(_06893_));
 sg13g2_inv_1 _27071_ (.Y(_06896_),
    .A(_06895_));
 sg13g2_nand2_1 _27072_ (.Y(_06897_),
    .A(net136),
    .B(_06751_));
 sg13g2_nor2_1 _27073_ (.A(_06841_),
    .B(_06844_),
    .Y(_06898_));
 sg13g2_xnor2_1 _27074_ (.Y(_06899_),
    .A(_06593_),
    .B(_06777_));
 sg13g2_nor2_1 _27075_ (.A(_06898_),
    .B(_06899_),
    .Y(_06900_));
 sg13g2_a21oi_2 _27076_ (.B1(_06900_),
    .Y(_06901_),
    .A2(_06844_),
    .A1(_06841_));
 sg13g2_nand2b_1 _27077_ (.Y(_06902_),
    .B(net84),
    .A_N(net81));
 sg13g2_nor2_1 _27078_ (.A(_06590_),
    .B(net81),
    .Y(_06903_));
 sg13g2_nand2_1 _27079_ (.Y(_06904_),
    .A(_06590_),
    .B(net81));
 sg13g2_nor2_1 _27080_ (.A(net84),
    .B(_06904_),
    .Y(_06905_));
 sg13g2_a21oi_1 _27081_ (.A1(_06216_),
    .A2(_06903_),
    .Y(_06906_),
    .B1(_06905_));
 sg13g2_nand3b_1 _27082_ (.B(net81),
    .C(_06367_),
    .Y(_06907_),
    .A_N(net84));
 sg13g2_o21ai_1 _27083_ (.B1(_06907_),
    .Y(_06908_),
    .A1(_06367_),
    .A2(_06772_));
 sg13g2_nor2_1 _27084_ (.A(_06371_),
    .B(_06908_),
    .Y(_06909_));
 sg13g2_a21oi_1 _27085_ (.A1(net117),
    .A2(_06906_),
    .Y(_06910_),
    .B1(_06909_));
 sg13g2_a21o_1 _27086_ (.A2(_06902_),
    .A1(_06752_),
    .B1(_06910_),
    .X(_06911_));
 sg13g2_buf_1 _27087_ (.A(_06911_),
    .X(_06912_));
 sg13g2_o21ai_1 _27088_ (.B1(net204),
    .Y(_06913_),
    .A1(net233),
    .A2(_13950_));
 sg13g2_nand2_1 _27089_ (.Y(_06914_),
    .A(net233),
    .B(_13950_));
 sg13g2_a21o_1 _27090_ (.A2(_06914_),
    .A1(_06913_),
    .B1(_01891_),
    .X(_06915_));
 sg13g2_buf_1 _27091_ (.A(_06915_),
    .X(_06916_));
 sg13g2_xnor2_1 _27092_ (.Y(_06917_),
    .A(_06232_),
    .B(_06916_));
 sg13g2_a21o_1 _27093_ (.A2(net81),
    .A1(_06368_),
    .B1(_12388_),
    .X(_06918_));
 sg13g2_or2_1 _27094_ (.X(_06919_),
    .B(net81),
    .A(_06510_));
 sg13g2_a21oi_1 _27095_ (.A1(_06918_),
    .A2(_06919_),
    .Y(_06920_),
    .B1(net231));
 sg13g2_xnor2_1 _27096_ (.Y(_06921_),
    .A(_06917_),
    .B(_06920_));
 sg13g2_a21o_1 _27097_ (.A2(_06813_),
    .A1(_06809_),
    .B1(_06805_),
    .X(_06922_));
 sg13g2_o21ai_1 _27098_ (.B1(_06922_),
    .Y(_06923_),
    .A1(_06809_),
    .A2(_06813_));
 sg13g2_inv_1 _27099_ (.Y(_06924_),
    .A(_06783_));
 sg13g2_a22oi_1 _27100_ (.Y(_06925_),
    .B1(_06924_),
    .B2(_06784_),
    .A2(net149),
    .A1(net234));
 sg13g2_a21oi_1 _27101_ (.A1(_06783_),
    .A2(_06785_),
    .Y(_06926_),
    .B1(_06925_));
 sg13g2_nand2_1 _27102_ (.Y(_06927_),
    .A(_13351_),
    .B(net212));
 sg13g2_nand2_1 _27103_ (.Y(_06928_),
    .A(net500),
    .B(_01890_));
 sg13g2_nand2_1 _27104_ (.Y(_06929_),
    .A(net234),
    .B(net150));
 sg13g2_xnor2_1 _27105_ (.Y(_06930_),
    .A(_06928_),
    .B(_06929_));
 sg13g2_xnor2_1 _27106_ (.Y(_06931_),
    .A(_06927_),
    .B(_06930_));
 sg13g2_nand2b_1 _27107_ (.Y(_06932_),
    .B(_06931_),
    .A_N(_06782_));
 sg13g2_a21o_1 _27108_ (.A2(_06781_),
    .A1(_06090_),
    .B1(_06931_),
    .X(_06933_));
 sg13g2_and2_1 _27109_ (.A(_06932_),
    .B(_06933_),
    .X(_06934_));
 sg13g2_xnor2_1 _27110_ (.Y(_06935_),
    .A(_06926_),
    .B(_06934_));
 sg13g2_nor2_1 _27111_ (.A(_06782_),
    .B(_06788_),
    .Y(_06936_));
 sg13g2_nand2_1 _27112_ (.Y(_06937_),
    .A(_06782_),
    .B(_06788_));
 sg13g2_o21ai_1 _27113_ (.B1(_06937_),
    .Y(_06938_),
    .A1(_06780_),
    .A2(_06936_));
 sg13g2_xor2_1 _27114_ (.B(_06938_),
    .A(_06935_),
    .X(_06939_));
 sg13g2_xnor2_1 _27115_ (.Y(_06940_),
    .A(_06923_),
    .B(_06939_));
 sg13g2_a21o_1 _27116_ (.A2(_06834_),
    .A1(_06832_),
    .B1(_06815_),
    .X(_06941_));
 sg13g2_o21ai_1 _27117_ (.B1(_06941_),
    .Y(_06942_),
    .A1(_06832_),
    .A2(_06834_));
 sg13g2_xnor2_1 _27118_ (.Y(_06943_),
    .A(_06940_),
    .B(_06942_));
 sg13g2_nor2_1 _27119_ (.A(_12732_),
    .B(net208),
    .Y(_06944_));
 sg13g2_nand2_1 _27120_ (.Y(_06945_),
    .A(net501),
    .B(_13948_));
 sg13g2_nor2_1 _27121_ (.A(_12729_),
    .B(_13758_),
    .Y(_06946_));
 sg13g2_xor2_1 _27122_ (.B(_06946_),
    .A(_06945_),
    .X(_06947_));
 sg13g2_xnor2_1 _27123_ (.Y(_06948_),
    .A(_06944_),
    .B(_06947_));
 sg13g2_nand2_1 _27124_ (.Y(_06949_),
    .A(_06802_),
    .B(_06803_));
 sg13g2_nand2_1 _27125_ (.Y(_06950_),
    .A(_06801_),
    .B(_06949_));
 sg13g2_o21ai_1 _27126_ (.B1(_06950_),
    .Y(_06951_),
    .A1(_06802_),
    .A2(_06803_));
 sg13g2_buf_1 _27127_ (.A(_06951_),
    .X(_06952_));
 sg13g2_a21oi_1 _27128_ (.A1(net255),
    .A2(_06133_),
    .Y(_06953_),
    .B1(_06818_));
 sg13g2_nand2b_1 _27129_ (.Y(_06954_),
    .B(_06818_),
    .A_N(_06817_));
 sg13g2_o21ai_1 _27130_ (.B1(_06954_),
    .Y(_06955_),
    .A1(_06816_),
    .A2(_06953_));
 sg13g2_buf_1 _27131_ (.A(_06955_),
    .X(_06956_));
 sg13g2_xnor2_1 _27132_ (.Y(_06957_),
    .A(_06952_),
    .B(_06956_));
 sg13g2_xnor2_1 _27133_ (.Y(_06958_),
    .A(_06948_),
    .B(_06957_));
 sg13g2_nand2_1 _27134_ (.Y(_06959_),
    .A(net255),
    .B(_01846_));
 sg13g2_nand2_1 _27135_ (.Y(_06960_),
    .A(net135),
    .B(_12987_));
 sg13g2_nor2b_1 _27136_ (.A(net258),
    .B_N(_06133_),
    .Y(_06961_));
 sg13g2_xor2_1 _27137_ (.B(_06961_),
    .A(_06960_),
    .X(_06962_));
 sg13g2_xnor2_1 _27138_ (.Y(_06963_),
    .A(_06959_),
    .B(_06962_));
 sg13g2_nand2_1 _27139_ (.Y(_06964_),
    .A(_01810_),
    .B(_13384_));
 sg13g2_nor2_1 _27140_ (.A(_13788_),
    .B(net517),
    .Y(_06965_));
 sg13g2_nand2_1 _27141_ (.Y(_06966_),
    .A(net284),
    .B(_01863_));
 sg13g2_xnor2_1 _27142_ (.Y(_06967_),
    .A(_06965_),
    .B(_06966_));
 sg13g2_xnor2_1 _27143_ (.Y(_06968_),
    .A(_06964_),
    .B(_06967_));
 sg13g2_a21o_1 _27144_ (.A2(_06823_),
    .A1(_06821_),
    .B1(_06824_),
    .X(_06969_));
 sg13g2_o21ai_1 _27145_ (.B1(_06969_),
    .Y(_06970_),
    .A1(_06821_),
    .A2(_06823_));
 sg13g2_buf_1 _27146_ (.A(_06970_),
    .X(_06971_));
 sg13g2_xor2_1 _27147_ (.B(_06971_),
    .A(_06968_),
    .X(_06972_));
 sg13g2_xnor2_1 _27148_ (.Y(_06973_),
    .A(_06963_),
    .B(_06972_));
 sg13g2_buf_1 _27149_ (.A(_06973_),
    .X(_06974_));
 sg13g2_a21o_1 _27150_ (.A2(_06830_),
    .A1(_06826_),
    .B1(_06820_),
    .X(_06975_));
 sg13g2_o21ai_1 _27151_ (.B1(_06975_),
    .Y(_06976_),
    .A1(_06826_),
    .A2(_06830_));
 sg13g2_buf_1 _27152_ (.A(_06976_),
    .X(_06977_));
 sg13g2_xnor2_1 _27153_ (.Y(_06978_),
    .A(_06974_),
    .B(_06977_));
 sg13g2_xnor2_1 _27154_ (.Y(_06979_),
    .A(_06958_),
    .B(_06978_));
 sg13g2_xnor2_1 _27155_ (.Y(_06980_),
    .A(_06943_),
    .B(_06979_));
 sg13g2_xnor2_1 _27156_ (.Y(_06981_),
    .A(_06921_),
    .B(_06980_));
 sg13g2_xnor2_1 _27157_ (.Y(_06982_),
    .A(_06912_),
    .B(_06981_));
 sg13g2_nand2_1 _27158_ (.Y(_06983_),
    .A(_06836_),
    .B(_06839_));
 sg13g2_nand2_1 _27159_ (.Y(_06984_),
    .A(_06800_),
    .B(_06983_));
 sg13g2_o21ai_1 _27160_ (.B1(_06984_),
    .Y(_06985_),
    .A1(_06836_),
    .A2(_06839_));
 sg13g2_buf_1 _27161_ (.A(_06985_),
    .X(_06986_));
 sg13g2_a21oi_1 _27162_ (.A1(_06790_),
    .A2(_06798_),
    .Y(_06987_),
    .B1(_06797_));
 sg13g2_xor2_1 _27163_ (.B(_06987_),
    .A(_06986_),
    .X(_06988_));
 sg13g2_xnor2_1 _27164_ (.Y(_06989_),
    .A(_06982_),
    .B(_06988_));
 sg13g2_xnor2_1 _27165_ (.Y(_06990_),
    .A(net82),
    .B(_06775_));
 sg13g2_o21ai_1 _27166_ (.B1(_06990_),
    .Y(_06991_),
    .A1(_06763_),
    .A2(_06767_));
 sg13g2_nand2_1 _27167_ (.Y(_06992_),
    .A(_06763_),
    .B(_06767_));
 sg13g2_nand2_2 _27168_ (.Y(_06993_),
    .A(_06991_),
    .B(_06992_));
 sg13g2_xor2_1 _27169_ (.B(_06993_),
    .A(_06989_),
    .X(_06994_));
 sg13g2_xnor2_1 _27170_ (.Y(_06995_),
    .A(_06901_),
    .B(_06994_));
 sg13g2_xnor2_1 _27171_ (.Y(_06996_),
    .A(_06337_),
    .B(_06995_));
 sg13g2_xor2_1 _27172_ (.B(_06996_),
    .A(_06897_),
    .X(_06997_));
 sg13g2_xnor2_1 _27173_ (.Y(_06998_),
    .A(_06896_),
    .B(_06997_));
 sg13g2_a21o_1 _27174_ (.A2(_06849_),
    .A1(_06740_),
    .B1(_06741_),
    .X(_06999_));
 sg13g2_o21ai_1 _27175_ (.B1(_06999_),
    .Y(_07000_),
    .A1(_06740_),
    .A2(_06849_));
 sg13g2_buf_1 _27176_ (.A(_07000_),
    .X(_07001_));
 sg13g2_xnor2_1 _27177_ (.Y(_07002_),
    .A(_06998_),
    .B(_07001_));
 sg13g2_xnor2_1 _27178_ (.Y(_07003_),
    .A(_06891_),
    .B(_07002_));
 sg13g2_nand2_1 _27179_ (.Y(_07004_),
    .A(net60),
    .B(_07003_));
 sg13g2_a21o_1 _27180_ (.A2(_06873_),
    .A1(_05811_),
    .B1(_11219_),
    .X(_07005_));
 sg13g2_o21ai_1 _27181_ (.B1(_07005_),
    .Y(_07006_),
    .A1(_05811_),
    .A2(_06873_));
 sg13g2_xnor2_1 _27182_ (.Y(_07007_),
    .A(_05818_),
    .B(_07006_));
 sg13g2_nand3_1 _27183_ (.B(_11472_),
    .C(_07007_),
    .A(_11217_),
    .Y(_07008_));
 sg13g2_o21ai_1 _27184_ (.B1(_07008_),
    .Y(_07009_),
    .A1(_11217_),
    .A2(_07007_));
 sg13g2_a22oi_1 _27185_ (.Y(_07010_),
    .B1(_07009_),
    .B2(_05992_),
    .A2(_05988_),
    .A1(_11216_));
 sg13g2_a21oi_1 _27186_ (.A1(_07004_),
    .A2(_07010_),
    .Y(_01751_),
    .B1(_05994_));
 sg13g2_inv_1 _27187_ (.Y(_07011_),
    .A(_06989_));
 sg13g2_nand2_1 _27188_ (.Y(_07012_),
    .A(_07011_),
    .B(_06993_));
 sg13g2_nand2_1 _27189_ (.Y(_07013_),
    .A(_06901_),
    .B(_07012_));
 sg13g2_nor3_1 _27190_ (.A(_06337_),
    .B(_07011_),
    .C(_06993_),
    .Y(_07014_));
 sg13g2_or2_1 _27191_ (.X(_07015_),
    .B(_07014_),
    .A(_06901_));
 sg13g2_o21ai_1 _27192_ (.B1(_06901_),
    .Y(_07016_),
    .A1(_07011_),
    .A2(_06993_));
 sg13g2_a21oi_1 _27193_ (.A1(_07012_),
    .A2(_07016_),
    .Y(_07017_),
    .B1(_06317_));
 sg13g2_a21oi_1 _27194_ (.A1(_07013_),
    .A2(_07015_),
    .Y(_07018_),
    .B1(_07017_));
 sg13g2_and2_1 _27195_ (.A(_06940_),
    .B(_06942_),
    .X(_07019_));
 sg13g2_buf_1 _27196_ (.A(_07019_),
    .X(_07020_));
 sg13g2_nand2_1 _27197_ (.Y(_07021_),
    .A(_06977_),
    .B(_07020_));
 sg13g2_or2_1 _27198_ (.X(_07022_),
    .B(_07021_),
    .A(_06974_));
 sg13g2_or2_1 _27199_ (.X(_07023_),
    .B(_06942_),
    .A(_06940_));
 sg13g2_buf_1 _27200_ (.A(_07023_),
    .X(_07024_));
 sg13g2_nor2_1 _27201_ (.A(_06977_),
    .B(_07024_),
    .Y(_07025_));
 sg13g2_o21ai_1 _27202_ (.B1(_07025_),
    .Y(_07026_),
    .A1(_06958_),
    .A2(_06974_));
 sg13g2_o21ai_1 _27203_ (.B1(_07024_),
    .Y(_07027_),
    .A1(_06977_),
    .A2(_07020_));
 sg13g2_nand3_1 _27204_ (.B(_06974_),
    .C(_07027_),
    .A(_06958_),
    .Y(_07028_));
 sg13g2_a21oi_1 _27205_ (.A1(_06977_),
    .A2(_07024_),
    .Y(_07029_),
    .B1(_07020_));
 sg13g2_o21ai_1 _27206_ (.B1(_07021_),
    .Y(_07030_),
    .A1(_06974_),
    .A2(_07029_));
 sg13g2_nand2b_1 _27207_ (.Y(_07031_),
    .B(_07030_),
    .A_N(_06958_));
 sg13g2_nand4_1 _27208_ (.B(_07026_),
    .C(_07028_),
    .A(_07022_),
    .Y(_07032_),
    .D(_07031_));
 sg13g2_a21oi_1 _27209_ (.A1(_06590_),
    .A2(net81),
    .Y(_07033_),
    .B1(_06916_));
 sg13g2_o21ai_1 _27210_ (.B1(_07033_),
    .Y(_07034_),
    .A1(net117),
    .A2(_06903_));
 sg13g2_a22oi_1 _27211_ (.Y(_07035_),
    .B1(_07034_),
    .B2(net89),
    .A2(_06916_),
    .A1(_06372_));
 sg13g2_mux2_1 _27212_ (.A0(_06932_),
    .A1(_06933_),
    .S(_06926_),
    .X(_07036_));
 sg13g2_a21o_1 _27213_ (.A2(_06956_),
    .A1(_06952_),
    .B1(_06948_),
    .X(_07037_));
 sg13g2_o21ai_1 _27214_ (.B1(_07037_),
    .Y(_07038_),
    .A1(_06952_),
    .A2(_06956_));
 sg13g2_xnor2_1 _27215_ (.Y(_07039_),
    .A(_07036_),
    .B(_07038_));
 sg13g2_xnor2_1 _27216_ (.Y(_07040_),
    .A(_07035_),
    .B(_07039_));
 sg13g2_nor2_1 _27217_ (.A(_12630_),
    .B(net206),
    .Y(_07041_));
 sg13g2_nand2_1 _27218_ (.Y(_07042_),
    .A(net255),
    .B(net480));
 sg13g2_xor2_1 _27219_ (.B(_07042_),
    .A(_07041_),
    .X(_07043_));
 sg13g2_nand2b_1 _27220_ (.Y(_07044_),
    .B(_06927_),
    .A_N(_06928_));
 sg13g2_nand4_1 _27221_ (.B(_06090_),
    .C(_06928_),
    .A(net236),
    .Y(_07045_),
    .D(_06929_));
 sg13g2_o21ai_1 _27222_ (.B1(_07045_),
    .Y(_07046_),
    .A1(_06929_),
    .A2(_07044_));
 sg13g2_xnor2_1 _27223_ (.Y(_07047_),
    .A(_07043_),
    .B(_07046_));
 sg13g2_a21oi_1 _27224_ (.A1(net135),
    .A2(net482),
    .Y(_07048_),
    .B1(_06961_));
 sg13g2_nand3_1 _27225_ (.B(net482),
    .C(_06961_),
    .A(net135),
    .Y(_07049_));
 sg13g2_o21ai_1 _27226_ (.B1(_07049_),
    .Y(_07050_),
    .A1(_06959_),
    .A2(_07048_));
 sg13g2_o21ai_1 _27227_ (.B1(_06945_),
    .Y(_07051_),
    .A1(_12729_),
    .A2(net207));
 sg13g2_nor2b_1 _27228_ (.A(_06945_),
    .B_N(_06946_),
    .Y(_07052_));
 sg13g2_a21oi_1 _27229_ (.A1(_06944_),
    .A2(_07051_),
    .Y(_07053_),
    .B1(_07052_));
 sg13g2_xor2_1 _27230_ (.B(_07053_),
    .A(_07050_),
    .X(_07054_));
 sg13g2_xnor2_1 _27231_ (.Y(_07055_),
    .A(_07047_),
    .B(_07054_));
 sg13g2_nand2_1 _27232_ (.Y(_07056_),
    .A(_13951_),
    .B(net478));
 sg13g2_nor2_1 _27233_ (.A(_12729_),
    .B(net208),
    .Y(_07057_));
 sg13g2_xnor2_1 _27234_ (.Y(_07058_),
    .A(_07056_),
    .B(_07057_));
 sg13g2_nand2_1 _27235_ (.Y(_07059_),
    .A(_06964_),
    .B(_06966_));
 sg13g2_nor2_1 _27236_ (.A(_06964_),
    .B(_06966_),
    .Y(_07060_));
 sg13g2_a21oi_1 _27237_ (.A1(_06965_),
    .A2(_07059_),
    .Y(_07061_),
    .B1(_07060_));
 sg13g2_xnor2_1 _27238_ (.Y(_07062_),
    .A(_07058_),
    .B(_07061_));
 sg13g2_xnor2_1 _27239_ (.Y(_07063_),
    .A(_06232_),
    .B(_07062_));
 sg13g2_nor2_1 _27240_ (.A(_12238_),
    .B(net231),
    .Y(_07064_));
 sg13g2_nor2_1 _27241_ (.A(_12979_),
    .B(net207),
    .Y(_07065_));
 sg13g2_xor2_1 _27242_ (.B(_07065_),
    .A(_07064_),
    .X(_07066_));
 sg13g2_nand2_1 _27243_ (.Y(_07067_),
    .A(net135),
    .B(net469));
 sg13g2_nand2_1 _27244_ (.Y(_07068_),
    .A(net173),
    .B(net482));
 sg13g2_xnor2_1 _27245_ (.Y(_07069_),
    .A(_07067_),
    .B(_07068_));
 sg13g2_xnor2_1 _27246_ (.Y(_07070_),
    .A(_07066_),
    .B(_07069_));
 sg13g2_nor2_1 _27247_ (.A(net284),
    .B(net517),
    .Y(_07071_));
 sg13g2_nand2_1 _27248_ (.Y(_07072_),
    .A(net256),
    .B(net477));
 sg13g2_xnor2_1 _27249_ (.Y(_07073_),
    .A(_07071_),
    .B(_07072_));
 sg13g2_nand2_1 _27250_ (.Y(_07074_),
    .A(net499),
    .B(net149));
 sg13g2_xnor2_1 _27251_ (.Y(_07075_),
    .A(_07073_),
    .B(_07074_));
 sg13g2_xnor2_1 _27252_ (.Y(_07076_),
    .A(_06337_),
    .B(_07075_));
 sg13g2_xnor2_1 _27253_ (.Y(_07077_),
    .A(_07070_),
    .B(_07076_));
 sg13g2_xnor2_1 _27254_ (.Y(_07078_),
    .A(_07063_),
    .B(_07077_));
 sg13g2_nor2_1 _27255_ (.A(_06968_),
    .B(_06971_),
    .Y(_07079_));
 sg13g2_nor2_1 _27256_ (.A(_06963_),
    .B(_07079_),
    .Y(_07080_));
 sg13g2_a21oi_1 _27257_ (.A1(_06968_),
    .A2(_06971_),
    .Y(_07081_),
    .B1(_07080_));
 sg13g2_xnor2_1 _27258_ (.Y(_07082_),
    .A(_07078_),
    .B(_07081_));
 sg13g2_xnor2_1 _27259_ (.Y(_07083_),
    .A(_07055_),
    .B(_07082_));
 sg13g2_xnor2_1 _27260_ (.Y(_07084_),
    .A(_07040_),
    .B(_07083_));
 sg13g2_nor2b_1 _27261_ (.A(_06935_),
    .B_N(_06938_),
    .Y(_07085_));
 sg13g2_nand2b_1 _27262_ (.Y(_07086_),
    .B(_06935_),
    .A_N(_06938_));
 sg13g2_o21ai_1 _27263_ (.B1(_07086_),
    .Y(_07087_),
    .A1(_06923_),
    .A2(_07085_));
 sg13g2_xnor2_1 _27264_ (.Y(_07088_),
    .A(_07084_),
    .B(_07087_));
 sg13g2_xnor2_1 _27265_ (.Y(_07089_),
    .A(_07032_),
    .B(_07088_));
 sg13g2_and2_1 _27266_ (.A(_06980_),
    .B(_06987_),
    .X(_07090_));
 sg13g2_buf_1 _27267_ (.A(_07090_),
    .X(_07091_));
 sg13g2_and2_1 _27268_ (.A(_06921_),
    .B(_07091_),
    .X(_07092_));
 sg13g2_nor2_1 _27269_ (.A(_06980_),
    .B(_06987_),
    .Y(_07093_));
 sg13g2_nor2b_1 _27270_ (.A(_07093_),
    .B_N(_06921_),
    .Y(_07094_));
 sg13g2_o21ai_1 _27271_ (.B1(_06986_),
    .Y(_07095_),
    .A1(_07091_),
    .A2(_07094_));
 sg13g2_nand2b_1 _27272_ (.Y(_07096_),
    .B(_07095_),
    .A_N(_07092_));
 sg13g2_nand2b_1 _27273_ (.Y(_07097_),
    .B(_07093_),
    .A_N(_06921_));
 sg13g2_a21oi_1 _27274_ (.A1(_06912_),
    .A2(_06986_),
    .Y(_07098_),
    .B1(_07097_));
 sg13g2_nor2_1 _27275_ (.A(_06921_),
    .B(_07091_),
    .Y(_07099_));
 sg13g2_nor2_1 _27276_ (.A(_06912_),
    .B(_06986_),
    .Y(_07100_));
 sg13g2_o21ai_1 _27277_ (.B1(_07100_),
    .Y(_07101_),
    .A1(_07093_),
    .A2(_07099_));
 sg13g2_nand2b_1 _27278_ (.Y(_07102_),
    .B(_07101_),
    .A_N(_07098_));
 sg13g2_a221oi_1 _27279_ (.B2(_06912_),
    .C1(_07102_),
    .B1(_07096_),
    .A1(_06986_),
    .Y(_07103_),
    .A2(_07092_));
 sg13g2_xnor2_1 _27280_ (.Y(_07104_),
    .A(_07089_),
    .B(_07103_));
 sg13g2_xnor2_1 _27281_ (.Y(_07105_),
    .A(_07018_),
    .B(_07104_));
 sg13g2_inv_1 _27282_ (.Y(_07106_),
    .A(_06996_));
 sg13g2_a21oi_1 _27283_ (.A1(_06896_),
    .A2(_06996_),
    .Y(_07107_),
    .B1(_06897_));
 sg13g2_a21oi_1 _27284_ (.A1(_06895_),
    .A2(_07106_),
    .Y(_07108_),
    .B1(_07107_));
 sg13g2_xnor2_1 _27285_ (.Y(_07109_),
    .A(_07105_),
    .B(_07108_));
 sg13g2_a21o_1 _27286_ (.A2(_07001_),
    .A1(_06998_),
    .B1(_06891_),
    .X(_07110_));
 sg13g2_o21ai_1 _27287_ (.B1(_07110_),
    .Y(_07111_),
    .A1(_06998_),
    .A2(_07001_));
 sg13g2_xnor2_1 _27288_ (.Y(_07112_),
    .A(_07109_),
    .B(_07111_));
 sg13g2_nand2_1 _27289_ (.Y(_07113_),
    .A(_11353_),
    .B(_07112_));
 sg13g2_xnor2_1 _27290_ (.Y(_07114_),
    .A(_11212_),
    .B(\rbzero.wall_tracer.stepDistX[10] ));
 sg13g2_nor2_1 _27291_ (.A(_11216_),
    .B(_05818_),
    .Y(_07115_));
 sg13g2_nand2_1 _27292_ (.Y(_07116_),
    .A(_11216_),
    .B(_05818_));
 sg13g2_o21ai_1 _27293_ (.B1(_07116_),
    .Y(_07117_),
    .A1(_07006_),
    .A2(_07115_));
 sg13g2_xnor2_1 _27294_ (.Y(_07118_),
    .A(_07114_),
    .B(_07117_));
 sg13g2_a21oi_1 _27295_ (.A1(net700),
    .A2(_07118_),
    .Y(_07119_),
    .B1(_11346_));
 sg13g2_a221oi_1 _27296_ (.B2(_07119_),
    .C1(net635),
    .B1(_07113_),
    .A1(_11213_),
    .Y(_01752_),
    .A2(_11344_));
 sg13g2_nand2b_1 _27297_ (.Y(_07120_),
    .B(_05996_),
    .A_N(_05915_));
 sg13g2_xnor2_1 _27298_ (.Y(_07121_),
    .A(_05823_),
    .B(_06005_));
 sg13g2_nor3_1 _27299_ (.A(_11262_),
    .B(net71),
    .C(_07121_),
    .Y(_07122_));
 sg13g2_a21o_1 _27300_ (.A2(_07121_),
    .A1(_11262_),
    .B1(_07122_),
    .X(_07123_));
 sg13g2_buf_1 _27301_ (.A(_11470_),
    .X(_07124_));
 sg13g2_a22oi_1 _27302_ (.Y(_07125_),
    .B1(_07123_),
    .B2(_07124_),
    .A2(net63),
    .A1(_11262_));
 sg13g2_buf_1 _27303_ (.A(_08675_),
    .X(_07126_));
 sg13g2_a21oi_1 _27304_ (.A1(_07120_),
    .A2(_07125_),
    .Y(_01753_),
    .B1(_07126_));
 sg13g2_nand2_1 _27305_ (.Y(_07127_),
    .A(_12777_),
    .B(net60));
 sg13g2_xnor2_1 _27306_ (.Y(_07128_),
    .A(_05826_),
    .B(_06007_));
 sg13g2_nor3_1 _27307_ (.A(_11261_),
    .B(net72),
    .C(_07128_),
    .Y(_07129_));
 sg13g2_a21o_1 _27308_ (.A2(_07128_),
    .A1(_11261_),
    .B1(_07129_),
    .X(_07130_));
 sg13g2_a22oi_1 _27309_ (.Y(_07131_),
    .B1(_07130_),
    .B2(net617),
    .A2(net63),
    .A1(_11261_));
 sg13g2_a21oi_1 _27310_ (.A1(_07127_),
    .A2(_07131_),
    .Y(_01754_),
    .B1(net616));
 sg13g2_nand2_1 _27311_ (.Y(_07132_),
    .A(_12890_),
    .B(net60));
 sg13g2_xnor2_1 _27312_ (.Y(_07133_),
    .A(_06001_),
    .B(_06010_));
 sg13g2_nor3_1 _27313_ (.A(_11258_),
    .B(net72),
    .C(_07133_),
    .Y(_07134_));
 sg13g2_a21o_1 _27314_ (.A2(_07133_),
    .A1(_11258_),
    .B1(_07134_),
    .X(_07135_));
 sg13g2_a22oi_1 _27315_ (.Y(_07136_),
    .B1(_07135_),
    .B2(net617),
    .A2(net63),
    .A1(_11258_));
 sg13g2_a21oi_1 _27316_ (.A1(_07132_),
    .A2(_07136_),
    .Y(_01755_),
    .B1(net616));
 sg13g2_nand2b_1 _27317_ (.Y(_07137_),
    .B(_05996_),
    .A_N(_13013_));
 sg13g2_xnor2_1 _27318_ (.Y(_07138_),
    .A(_05831_),
    .B(_06013_));
 sg13g2_nor3_1 _27319_ (.A(_11256_),
    .B(net72),
    .C(_07138_),
    .Y(_07139_));
 sg13g2_a21o_1 _27320_ (.A2(_07138_),
    .A1(_11256_),
    .B1(_07139_),
    .X(_07140_));
 sg13g2_a22oi_1 _27321_ (.Y(_07141_),
    .B1(_07140_),
    .B2(net617),
    .A2(net63),
    .A1(_11256_));
 sg13g2_a21oi_1 _27322_ (.A1(_07137_),
    .A2(_07141_),
    .Y(_01756_),
    .B1(net616));
 sg13g2_nand2_1 _27323_ (.Y(_07142_),
    .A(_13142_),
    .B(net60));
 sg13g2_xnor2_1 _27324_ (.Y(_07143_),
    .A(_06000_),
    .B(_06016_));
 sg13g2_nor3_1 _27325_ (.A(_11252_),
    .B(net72),
    .C(_07143_),
    .Y(_07144_));
 sg13g2_a21o_1 _27326_ (.A2(_07143_),
    .A1(_11252_),
    .B1(_07144_),
    .X(_07145_));
 sg13g2_a22oi_1 _27327_ (.Y(_07146_),
    .B1(_07145_),
    .B2(net617),
    .A2(net63),
    .A1(_11252_));
 sg13g2_a21oi_1 _27328_ (.A1(_07142_),
    .A2(_07146_),
    .Y(_01757_),
    .B1(net616));
 sg13g2_nand2_1 _27329_ (.Y(_07147_),
    .A(_13282_),
    .B(_05996_));
 sg13g2_xnor2_1 _27330_ (.Y(_07148_),
    .A(_05836_),
    .B(_06019_));
 sg13g2_nor3_1 _27331_ (.A(_11249_),
    .B(net72),
    .C(_07148_),
    .Y(_07149_));
 sg13g2_a21o_1 _27332_ (.A2(_07148_),
    .A1(_11249_),
    .B1(_07149_),
    .X(_07150_));
 sg13g2_a22oi_1 _27333_ (.Y(_07151_),
    .B1(_07150_),
    .B2(net617),
    .A2(net63),
    .A1(_11249_));
 sg13g2_a21oi_1 _27334_ (.A1(_07147_),
    .A2(_07151_),
    .Y(_01758_),
    .B1(net616));
 sg13g2_nand2b_1 _27335_ (.Y(_07152_),
    .B(_05996_),
    .A_N(_13422_));
 sg13g2_xnor2_1 _27336_ (.Y(_07153_),
    .A(_05839_),
    .B(_06022_));
 sg13g2_nor3_1 _27337_ (.A(_11247_),
    .B(net72),
    .C(_07153_),
    .Y(_07154_));
 sg13g2_a21o_1 _27338_ (.A2(_07153_),
    .A1(_11247_),
    .B1(_07154_),
    .X(_07155_));
 sg13g2_a22oi_1 _27339_ (.Y(_07156_),
    .B1(_07155_),
    .B2(net617),
    .A2(_11478_),
    .A1(_11247_));
 sg13g2_a21oi_1 _27340_ (.A1(_07152_),
    .A2(_07156_),
    .Y(_01759_),
    .B1(net616));
 sg13g2_nand2_1 _27341_ (.Y(_07157_),
    .A(_13559_),
    .B(_05996_));
 sg13g2_xnor2_1 _27342_ (.Y(_07158_),
    .A(_05843_),
    .B(_06025_));
 sg13g2_nor3_1 _27343_ (.A(_11243_),
    .B(net72),
    .C(_07158_),
    .Y(_07159_));
 sg13g2_a21o_1 _27344_ (.A2(_07158_),
    .A1(_11243_),
    .B1(_07159_),
    .X(_07160_));
 sg13g2_a22oi_1 _27345_ (.Y(_07161_),
    .B1(_07160_),
    .B2(net617),
    .A2(_11478_),
    .A1(_11243_));
 sg13g2_a21oi_1 _27346_ (.A1(_07157_),
    .A2(_07161_),
    .Y(_01760_),
    .B1(net616));
 sg13g2_nand2_1 _27347_ (.Y(_07162_),
    .A(net697),
    .B(_08479_));
 sg13g2_a21oi_1 _27348_ (.A1(_08674_),
    .A2(_07162_),
    .Y(_07163_),
    .B1(_11331_));
 sg13g2_a21o_1 _27349_ (.A2(_11334_),
    .A1(_08629_),
    .B1(_11323_),
    .X(_07164_));
 sg13g2_nand3_1 _27350_ (.B(_07163_),
    .C(_07164_),
    .A(_11528_),
    .Y(_07165_));
 sg13g2_buf_1 _27351_ (.A(_07165_),
    .X(_07166_));
 sg13g2_buf_1 _27352_ (.A(net70),
    .X(_07167_));
 sg13g2_or2_1 _27353_ (.X(_07168_),
    .B(_07167_),
    .A(_05986_));
 sg13g2_buf_1 _27354_ (.A(net66),
    .X(_07169_));
 sg13g2_nand2b_1 _27355_ (.Y(_07170_),
    .B(_12018_),
    .A_N(_11268_));
 sg13g2_nand2b_1 _27356_ (.Y(_07171_),
    .B(_11268_),
    .A_N(_12018_));
 sg13g2_o21ai_1 _27357_ (.B1(_07171_),
    .Y(_07172_),
    .A1(_07167_),
    .A2(_07170_));
 sg13g2_a22oi_1 _27358_ (.Y(_07173_),
    .B1(_07172_),
    .B2(_07124_),
    .A2(net59),
    .A1(_11268_));
 sg13g2_a21oi_1 _27359_ (.A1(_07168_),
    .A2(_07173_),
    .Y(_01761_),
    .B1(net616));
 sg13g2_nor2_1 _27360_ (.A(_08479_),
    .B(net70),
    .Y(_07174_));
 sg13g2_buf_1 _27361_ (.A(_07174_),
    .X(_07175_));
 sg13g2_buf_1 _27362_ (.A(net58),
    .X(_07176_));
 sg13g2_nand2_1 _27363_ (.Y(_07177_),
    .A(_13724_),
    .B(net55));
 sg13g2_inv_1 _27364_ (.Y(_07178_),
    .A(\rbzero.wall_tracer.stepDistY[-1] ));
 sg13g2_inv_1 _27365_ (.Y(_07179_),
    .A(\rbzero.wall_tracer.stepDistY[-5] ));
 sg13g2_inv_1 _27366_ (.Y(_07180_),
    .A(\rbzero.wall_tracer.stepDistY[-7] ));
 sg13g2_inv_1 _27367_ (.Y(_07181_),
    .A(_05890_));
 sg13g2_inv_1 _27368_ (.Y(_07182_),
    .A(\rbzero.wall_tracer.trackDistY[-10] ));
 sg13g2_a21oi_1 _27369_ (.A1(_11268_),
    .A2(_12018_),
    .Y(_07183_),
    .B1(_12029_));
 sg13g2_nand3_1 _27370_ (.B(_12018_),
    .C(_12029_),
    .A(_11268_),
    .Y(_07184_));
 sg13g2_o21ai_1 _27371_ (.B1(_07184_),
    .Y(_07185_),
    .A1(_07182_),
    .A2(_07183_));
 sg13g2_a21oi_1 _27372_ (.A1(_11264_),
    .A2(_05890_),
    .Y(_07186_),
    .B1(_07185_));
 sg13g2_a21oi_2 _27373_ (.B1(_07186_),
    .Y(_07187_),
    .A2(_07181_),
    .A1(_11265_));
 sg13g2_a21o_1 _27374_ (.A2(_07187_),
    .A1(_05893_),
    .B1(_11274_),
    .X(_07188_));
 sg13g2_o21ai_1 _27375_ (.B1(_07188_),
    .Y(_07189_),
    .A1(_05893_),
    .A2(_07187_));
 sg13g2_buf_1 _27376_ (.A(_07189_),
    .X(_07190_));
 sg13g2_a21o_1 _27377_ (.A2(_07190_),
    .A1(_07180_),
    .B1(_11260_),
    .X(_07191_));
 sg13g2_o21ai_1 _27378_ (.B1(_07191_),
    .Y(_07192_),
    .A1(_07180_),
    .A2(_07190_));
 sg13g2_buf_1 _27379_ (.A(_07192_),
    .X(_07193_));
 sg13g2_a21o_1 _27380_ (.A2(_07193_),
    .A1(_05898_),
    .B1(_11279_),
    .X(_07194_));
 sg13g2_o21ai_1 _27381_ (.B1(_07194_),
    .Y(_07195_),
    .A1(_05898_),
    .A2(_07193_));
 sg13g2_buf_1 _27382_ (.A(_07195_),
    .X(_07196_));
 sg13g2_a21o_1 _27383_ (.A2(_07196_),
    .A1(_07179_),
    .B1(_11255_),
    .X(_07197_));
 sg13g2_o21ai_1 _27384_ (.B1(_07197_),
    .Y(_07198_),
    .A1(_07179_),
    .A2(_07196_));
 sg13g2_buf_1 _27385_ (.A(_07198_),
    .X(_07199_));
 sg13g2_nor2_1 _27386_ (.A(_05904_),
    .B(_07199_),
    .Y(_07200_));
 sg13g2_a21oi_1 _27387_ (.A1(_05904_),
    .A2(_07199_),
    .Y(_07201_),
    .B1(_11248_));
 sg13g2_nor2_1 _27388_ (.A(_07200_),
    .B(_07201_),
    .Y(_07202_));
 sg13g2_nor2_1 _27389_ (.A(_05907_),
    .B(_07202_),
    .Y(_07203_));
 sg13g2_a21oi_1 _27390_ (.A1(_05907_),
    .A2(_07202_),
    .Y(_07204_),
    .B1(_11246_));
 sg13g2_nor2_1 _27391_ (.A(_07203_),
    .B(_07204_),
    .Y(_07205_));
 sg13g2_a21o_1 _27392_ (.A2(_07205_),
    .A1(_05910_),
    .B1(_11244_),
    .X(_07206_));
 sg13g2_o21ai_1 _27393_ (.B1(_07206_),
    .Y(_07207_),
    .A1(_05910_),
    .A2(_07205_));
 sg13g2_buf_1 _27394_ (.A(_07207_),
    .X(_07208_));
 sg13g2_xnor2_1 _27395_ (.Y(_07209_),
    .A(_07178_),
    .B(_07208_));
 sg13g2_nor3_1 _27396_ (.A(_11242_),
    .B(net66),
    .C(_07209_),
    .Y(_07210_));
 sg13g2_a21o_1 _27397_ (.A2(_07209_),
    .A1(_11242_),
    .B1(_07210_),
    .X(_07211_));
 sg13g2_a22oi_1 _27398_ (.Y(_07212_),
    .B1(_07211_),
    .B2(net617),
    .A2(net59),
    .A1(_11242_));
 sg13g2_a21oi_1 _27399_ (.A1(_07177_),
    .A2(_07212_),
    .Y(_01762_),
    .B1(_07126_));
 sg13g2_nand2_1 _27400_ (.Y(_07213_),
    .A(_13880_),
    .B(net55));
 sg13g2_inv_1 _27401_ (.Y(_07214_),
    .A(_07208_));
 sg13g2_a21oi_1 _27402_ (.A1(\rbzero.wall_tracer.stepDistY[-1] ),
    .A2(_07214_),
    .Y(_07215_),
    .B1(_11242_));
 sg13g2_a21oi_1 _27403_ (.A1(_07178_),
    .A2(_07208_),
    .Y(_07216_),
    .B1(_07215_));
 sg13g2_xnor2_1 _27404_ (.Y(_07217_),
    .A(_05853_),
    .B(_07216_));
 sg13g2_buf_1 _27405_ (.A(net70),
    .X(_07218_));
 sg13g2_nor3_1 _27406_ (.A(_11238_),
    .B(net65),
    .C(_07217_),
    .Y(_07219_));
 sg13g2_a21o_1 _27407_ (.A2(_07217_),
    .A1(_11238_),
    .B1(_07219_),
    .X(_07220_));
 sg13g2_buf_1 _27408_ (.A(_11470_),
    .X(_07221_));
 sg13g2_a22oi_1 _27409_ (.Y(_07222_),
    .B1(_07220_),
    .B2(net615),
    .A2(net59),
    .A1(_11238_));
 sg13g2_buf_1 _27410_ (.A(_08675_),
    .X(_07223_));
 sg13g2_a21oi_1 _27411_ (.A1(_07213_),
    .A2(_07222_),
    .Y(_01763_),
    .B1(net614));
 sg13g2_nand2b_1 _27412_ (.Y(_07224_),
    .B(_07175_),
    .A_N(_14050_));
 sg13g2_nor2_1 _27413_ (.A(_05853_),
    .B(_07216_),
    .Y(_07225_));
 sg13g2_a21oi_1 _27414_ (.A1(_05853_),
    .A2(_07216_),
    .Y(_07226_),
    .B1(_11238_));
 sg13g2_nor2_1 _27415_ (.A(_07225_),
    .B(_07226_),
    .Y(_07227_));
 sg13g2_xnor2_1 _27416_ (.Y(_07228_),
    .A(_05856_),
    .B(_07227_));
 sg13g2_nor3_1 _27417_ (.A(_11236_),
    .B(net65),
    .C(_07228_),
    .Y(_07229_));
 sg13g2_a21o_1 _27418_ (.A2(_07228_),
    .A1(_11236_),
    .B1(_07229_),
    .X(_07230_));
 sg13g2_a22oi_1 _27419_ (.Y(_07231_),
    .B1(_07230_),
    .B2(_07221_),
    .A2(net59),
    .A1(_11236_));
 sg13g2_a21oi_1 _27420_ (.A1(_07224_),
    .A2(_07231_),
    .Y(_01764_),
    .B1(net614));
 sg13g2_nand2_1 _27421_ (.Y(_07232_),
    .A(_01905_),
    .B(_07176_));
 sg13g2_nor2_1 _27422_ (.A(_05856_),
    .B(_07227_),
    .Y(_07233_));
 sg13g2_a21oi_1 _27423_ (.A1(_05856_),
    .A2(_07227_),
    .Y(_07234_),
    .B1(_11236_));
 sg13g2_nor2_1 _27424_ (.A(_07233_),
    .B(_07234_),
    .Y(_07235_));
 sg13g2_xnor2_1 _27425_ (.Y(_07236_),
    .A(_05859_),
    .B(_07235_));
 sg13g2_nor3_1 _27426_ (.A(_11234_),
    .B(_07218_),
    .C(_07236_),
    .Y(_07237_));
 sg13g2_a21o_1 _27427_ (.A2(_07236_),
    .A1(_11234_),
    .B1(_07237_),
    .X(_07238_));
 sg13g2_a22oi_1 _27428_ (.Y(_07239_),
    .B1(_07238_),
    .B2(_07221_),
    .A2(net59),
    .A1(_11234_));
 sg13g2_a21oi_1 _27429_ (.A1(_07232_),
    .A2(_07239_),
    .Y(_01765_),
    .B1(net614));
 sg13g2_nand2b_1 _27430_ (.Y(_07240_),
    .B(net58),
    .A_N(_06193_));
 sg13g2_nor2_1 _27431_ (.A(_05859_),
    .B(_07235_),
    .Y(_07241_));
 sg13g2_a21oi_1 _27432_ (.A1(_05859_),
    .A2(_07235_),
    .Y(_07242_),
    .B1(_11234_));
 sg13g2_nor2_1 _27433_ (.A(_07241_),
    .B(_07242_),
    .Y(_07243_));
 sg13g2_xnor2_1 _27434_ (.Y(_07244_),
    .A(_05862_),
    .B(_07243_));
 sg13g2_nor3_1 _27435_ (.A(_11232_),
    .B(net65),
    .C(_07244_),
    .Y(_07245_));
 sg13g2_a21o_1 _27436_ (.A2(_07244_),
    .A1(_11232_),
    .B1(_07245_),
    .X(_07246_));
 sg13g2_a22oi_1 _27437_ (.Y(_07247_),
    .B1(_07246_),
    .B2(net615),
    .A2(net59),
    .A1(_11232_));
 sg13g2_a21oi_1 _27438_ (.A1(_07240_),
    .A2(_07247_),
    .Y(_01766_),
    .B1(net614));
 sg13g2_nand2b_1 _27439_ (.Y(_07248_),
    .B(net58),
    .A_N(_06326_));
 sg13g2_buf_1 _27440_ (.A(net66),
    .X(_07249_));
 sg13g2_nor2_1 _27441_ (.A(_05862_),
    .B(_07243_),
    .Y(_07250_));
 sg13g2_a21oi_1 _27442_ (.A1(_05862_),
    .A2(_07243_),
    .Y(_07251_),
    .B1(_11232_));
 sg13g2_nor2_1 _27443_ (.A(_07250_),
    .B(_07251_),
    .Y(_07252_));
 sg13g2_xnor2_1 _27444_ (.Y(_07253_),
    .A(_05865_),
    .B(_07252_));
 sg13g2_nor3_1 _27445_ (.A(_11229_),
    .B(net65),
    .C(_07253_),
    .Y(_07254_));
 sg13g2_a21o_1 _27446_ (.A2(_07253_),
    .A1(_11229_),
    .B1(_07254_),
    .X(_07255_));
 sg13g2_a22oi_1 _27447_ (.Y(_07256_),
    .B1(_07255_),
    .B2(net615),
    .A2(net57),
    .A1(_11229_));
 sg13g2_a21oi_1 _27448_ (.A1(_07248_),
    .A2(_07256_),
    .Y(_01767_),
    .B1(_07223_));
 sg13g2_nand2_1 _27449_ (.Y(_07257_),
    .A(_06470_),
    .B(net55));
 sg13g2_nor2_1 _27450_ (.A(_05865_),
    .B(_07252_),
    .Y(_07258_));
 sg13g2_a21oi_1 _27451_ (.A1(_05865_),
    .A2(_07252_),
    .Y(_07259_),
    .B1(_11229_));
 sg13g2_nor2_1 _27452_ (.A(_07258_),
    .B(_07259_),
    .Y(_07260_));
 sg13g2_xnor2_1 _27453_ (.Y(_07261_),
    .A(_05868_),
    .B(_07260_));
 sg13g2_nor3_1 _27454_ (.A(_11226_),
    .B(net65),
    .C(_07261_),
    .Y(_07262_));
 sg13g2_a21o_1 _27455_ (.A2(_07261_),
    .A1(_11226_),
    .B1(_07262_),
    .X(_07263_));
 sg13g2_a22oi_1 _27456_ (.Y(_07264_),
    .B1(_07263_),
    .B2(net615),
    .A2(net57),
    .A1(_11226_));
 sg13g2_a21oi_1 _27457_ (.A1(_07257_),
    .A2(_07264_),
    .Y(_01768_),
    .B1(net614));
 sg13g2_nand2b_1 _27458_ (.Y(_07265_),
    .B(net58),
    .A_N(_06601_));
 sg13g2_nor2_1 _27459_ (.A(_05868_),
    .B(_07260_),
    .Y(_07266_));
 sg13g2_a21oi_1 _27460_ (.A1(_05868_),
    .A2(_07260_),
    .Y(_07267_),
    .B1(_11226_));
 sg13g2_nor2_1 _27461_ (.A(_07266_),
    .B(_07267_),
    .Y(_07268_));
 sg13g2_xnor2_1 _27462_ (.Y(_07269_),
    .A(_05871_),
    .B(_07268_));
 sg13g2_nor3_1 _27463_ (.A(_11222_),
    .B(net65),
    .C(_07269_),
    .Y(_07270_));
 sg13g2_a21o_1 _27464_ (.A2(_07269_),
    .A1(_11222_),
    .B1(_07270_),
    .X(_07271_));
 sg13g2_a22oi_1 _27465_ (.Y(_07272_),
    .B1(_07271_),
    .B2(net615),
    .A2(net57),
    .A1(_11222_));
 sg13g2_a21oi_1 _27466_ (.A1(_07265_),
    .A2(_07272_),
    .Y(_01769_),
    .B1(net614));
 sg13g2_nand2_1 _27467_ (.Y(_07273_),
    .A(_06727_),
    .B(_07176_));
 sg13g2_nor2_1 _27468_ (.A(_05871_),
    .B(_07268_),
    .Y(_07274_));
 sg13g2_a21oi_1 _27469_ (.A1(_05871_),
    .A2(_07268_),
    .Y(_07275_),
    .B1(_11222_));
 sg13g2_nor2_1 _27470_ (.A(_07274_),
    .B(_07275_),
    .Y(_07276_));
 sg13g2_xnor2_1 _27471_ (.Y(_07277_),
    .A(_05876_),
    .B(_07276_));
 sg13g2_nor3_1 _27472_ (.A(_11221_),
    .B(net65),
    .C(_07277_),
    .Y(_07278_));
 sg13g2_a21o_1 _27473_ (.A2(_07277_),
    .A1(_11221_),
    .B1(_07278_),
    .X(_07279_));
 sg13g2_a22oi_1 _27474_ (.Y(_07280_),
    .B1(_07279_),
    .B2(net615),
    .A2(_07249_),
    .A1(_11221_));
 sg13g2_a21oi_1 _27475_ (.A1(_07273_),
    .A2(_07280_),
    .Y(_01770_),
    .B1(net614));
 sg13g2_nand2_1 _27476_ (.Y(_07281_),
    .A(_06869_),
    .B(net55));
 sg13g2_nor2_1 _27477_ (.A(_05876_),
    .B(_07276_),
    .Y(_07282_));
 sg13g2_a21oi_1 _27478_ (.A1(_05876_),
    .A2(_07276_),
    .Y(_07283_),
    .B1(_11221_));
 sg13g2_nor2_1 _27479_ (.A(_07282_),
    .B(_07283_),
    .Y(_07284_));
 sg13g2_xnor2_1 _27480_ (.Y(_07285_),
    .A(_05879_),
    .B(_07284_));
 sg13g2_nor3_1 _27481_ (.A(_11218_),
    .B(_07218_),
    .C(_07285_),
    .Y(_07286_));
 sg13g2_a21o_1 _27482_ (.A2(_07285_),
    .A1(_11218_),
    .B1(_07286_),
    .X(_07287_));
 sg13g2_a22oi_1 _27483_ (.Y(_07288_),
    .B1(_07287_),
    .B2(net615),
    .A2(_07249_),
    .A1(_11218_));
 sg13g2_a21oi_1 _27484_ (.A1(_07281_),
    .A2(_07288_),
    .Y(_01771_),
    .B1(_07223_));
 sg13g2_nand2_1 _27485_ (.Y(_07289_),
    .A(_11268_),
    .B(_12018_));
 sg13g2_xor2_1 _27486_ (.B(_12029_),
    .A(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_07290_));
 sg13g2_xnor2_1 _27487_ (.Y(_07291_),
    .A(_07289_),
    .B(_07290_));
 sg13g2_a21oi_1 _27488_ (.A1(_11486_),
    .A2(_07291_),
    .Y(_07292_),
    .B1(net66));
 sg13g2_a221oi_1 _27489_ (.B2(_06880_),
    .C1(net635),
    .B1(_07292_),
    .A1(_07182_),
    .Y(_01772_),
    .A2(net59));
 sg13g2_a21o_1 _27490_ (.A2(_07284_),
    .A1(_05879_),
    .B1(_11218_),
    .X(_07293_));
 sg13g2_o21ai_1 _27491_ (.B1(_07293_),
    .Y(_07294_),
    .A1(_05879_),
    .A2(_07284_));
 sg13g2_xnor2_1 _27492_ (.Y(_07295_),
    .A(_11317_),
    .B(_05885_));
 sg13g2_xnor2_1 _27493_ (.Y(_07296_),
    .A(_07294_),
    .B(_07295_));
 sg13g2_nand2_1 _27494_ (.Y(_07297_),
    .A(_11347_),
    .B(_07003_));
 sg13g2_o21ai_1 _27495_ (.B1(_07297_),
    .Y(_07298_),
    .A1(_11353_),
    .A2(_07296_));
 sg13g2_nand2b_1 _27496_ (.Y(_07299_),
    .B(_07298_),
    .A_N(_07169_));
 sg13g2_nand2_1 _27497_ (.Y(_07300_),
    .A(_11317_),
    .B(net59));
 sg13g2_a21oi_1 _27498_ (.A1(_07299_),
    .A2(_07300_),
    .Y(_01773_),
    .B1(net614));
 sg13g2_xnor2_1 _27499_ (.Y(_07301_),
    .A(_11214_),
    .B(\rbzero.wall_tracer.stepDistY[10] ));
 sg13g2_nor2_1 _27500_ (.A(_11317_),
    .B(_05885_),
    .Y(_07302_));
 sg13g2_nand2_1 _27501_ (.Y(_07303_),
    .A(_11317_),
    .B(_05885_));
 sg13g2_o21ai_1 _27502_ (.B1(_07303_),
    .Y(_07304_),
    .A1(_07294_),
    .A2(_07302_));
 sg13g2_xnor2_1 _27503_ (.Y(_07305_),
    .A(_07301_),
    .B(_07304_));
 sg13g2_a21oi_1 _27504_ (.A1(_11486_),
    .A2(_07305_),
    .Y(_07306_),
    .B1(net66));
 sg13g2_a221oi_1 _27505_ (.B2(_07113_),
    .C1(net635),
    .B1(_07306_),
    .A1(_11215_),
    .Y(_01774_),
    .A2(_07169_));
 sg13g2_nand2b_1 _27506_ (.Y(_07307_),
    .B(net58),
    .A_N(_05915_));
 sg13g2_xnor2_1 _27507_ (.Y(_07308_),
    .A(_05890_),
    .B(_07185_));
 sg13g2_nor3_1 _27508_ (.A(_11264_),
    .B(net65),
    .C(_07308_),
    .Y(_07309_));
 sg13g2_a21o_1 _27509_ (.A2(_07308_),
    .A1(_11264_),
    .B1(_07309_),
    .X(_07310_));
 sg13g2_a22oi_1 _27510_ (.Y(_07311_),
    .B1(_07310_),
    .B2(net615),
    .A2(net57),
    .A1(_11264_));
 sg13g2_buf_1 _27511_ (.A(_08675_),
    .X(_07312_));
 sg13g2_a21oi_1 _27512_ (.A1(_07307_),
    .A2(_07311_),
    .Y(_01775_),
    .B1(net613));
 sg13g2_nand2_1 _27513_ (.Y(_07313_),
    .A(_12777_),
    .B(net55));
 sg13g2_xnor2_1 _27514_ (.Y(_07314_),
    .A(_05893_),
    .B(_07187_));
 sg13g2_nor3_1 _27515_ (.A(_11274_),
    .B(net70),
    .C(_07314_),
    .Y(_07315_));
 sg13g2_a21o_1 _27516_ (.A2(_07314_),
    .A1(_11274_),
    .B1(_07315_),
    .X(_07316_));
 sg13g2_a22oi_1 _27517_ (.Y(_07317_),
    .B1(_07316_),
    .B2(net637),
    .A2(net57),
    .A1(_11274_));
 sg13g2_a21oi_1 _27518_ (.A1(_07313_),
    .A2(_07317_),
    .Y(_01776_),
    .B1(net613));
 sg13g2_nand2_1 _27519_ (.Y(_07318_),
    .A(_12890_),
    .B(net55));
 sg13g2_xnor2_1 _27520_ (.Y(_07319_),
    .A(_07180_),
    .B(_07190_));
 sg13g2_nor3_1 _27521_ (.A(_11257_),
    .B(net70),
    .C(_07319_),
    .Y(_07320_));
 sg13g2_a21o_1 _27522_ (.A2(_07319_),
    .A1(_11257_),
    .B1(_07320_),
    .X(_07321_));
 sg13g2_a22oi_1 _27523_ (.Y(_07322_),
    .B1(_07321_),
    .B2(net637),
    .A2(net57),
    .A1(_11257_));
 sg13g2_a21oi_1 _27524_ (.A1(_07318_),
    .A2(_07322_),
    .Y(_01777_),
    .B1(net613));
 sg13g2_nand2b_1 _27525_ (.Y(_07323_),
    .B(net58),
    .A_N(_13013_));
 sg13g2_xnor2_1 _27526_ (.Y(_07324_),
    .A(_05898_),
    .B(_07193_));
 sg13g2_nor3_1 _27527_ (.A(_11279_),
    .B(net70),
    .C(_07324_),
    .Y(_07325_));
 sg13g2_a21o_1 _27528_ (.A2(_07324_),
    .A1(_11279_),
    .B1(_07325_),
    .X(_07326_));
 sg13g2_a22oi_1 _27529_ (.Y(_07327_),
    .B1(_07326_),
    .B2(net637),
    .A2(net57),
    .A1(_11279_));
 sg13g2_a21oi_1 _27530_ (.A1(_07323_),
    .A2(_07327_),
    .Y(_01778_),
    .B1(net613));
 sg13g2_nand2_1 _27531_ (.Y(_07328_),
    .A(_13142_),
    .B(net55));
 sg13g2_xnor2_1 _27532_ (.Y(_07329_),
    .A(_07179_),
    .B(_07196_));
 sg13g2_nor3_1 _27533_ (.A(_11254_),
    .B(_07166_),
    .C(_07329_),
    .Y(_07330_));
 sg13g2_a21o_1 _27534_ (.A2(_07329_),
    .A1(_11254_),
    .B1(_07330_),
    .X(_07331_));
 sg13g2_a22oi_1 _27535_ (.Y(_07332_),
    .B1(_07331_),
    .B2(net637),
    .A2(net57),
    .A1(_11254_));
 sg13g2_a21oi_1 _27536_ (.A1(_07328_),
    .A2(_07332_),
    .Y(_01779_),
    .B1(net613));
 sg13g2_nand2_1 _27537_ (.Y(_07333_),
    .A(_13282_),
    .B(net55));
 sg13g2_xnor2_1 _27538_ (.Y(_07334_),
    .A(_05904_),
    .B(_07199_));
 sg13g2_nor3_1 _27539_ (.A(_11248_),
    .B(net70),
    .C(_07334_),
    .Y(_07335_));
 sg13g2_a21o_1 _27540_ (.A2(_07334_),
    .A1(_11248_),
    .B1(_07335_),
    .X(_07336_));
 sg13g2_a22oi_1 _27541_ (.Y(_07337_),
    .B1(_07336_),
    .B2(net637),
    .A2(net66),
    .A1(_11248_));
 sg13g2_a21oi_1 _27542_ (.A1(_07333_),
    .A2(_07337_),
    .Y(_01780_),
    .B1(net613));
 sg13g2_nand2b_1 _27543_ (.Y(_07338_),
    .B(net58),
    .A_N(_13422_));
 sg13g2_xnor2_1 _27544_ (.Y(_07339_),
    .A(_05907_),
    .B(_07202_));
 sg13g2_nor3_1 _27545_ (.A(_11246_),
    .B(net70),
    .C(_07339_),
    .Y(_07340_));
 sg13g2_a21o_1 _27546_ (.A2(_07339_),
    .A1(_11246_),
    .B1(_07340_),
    .X(_07341_));
 sg13g2_a22oi_1 _27547_ (.Y(_07342_),
    .B1(_07341_),
    .B2(net637),
    .A2(net66),
    .A1(_11246_));
 sg13g2_a21oi_1 _27548_ (.A1(_07338_),
    .A2(_07342_),
    .Y(_01781_),
    .B1(net613));
 sg13g2_nand2_1 _27549_ (.Y(_07343_),
    .A(_13559_),
    .B(net58));
 sg13g2_xnor2_1 _27550_ (.Y(_07344_),
    .A(_05910_),
    .B(_07205_));
 sg13g2_nor3_1 _27551_ (.A(_11244_),
    .B(_07166_),
    .C(_07344_),
    .Y(_07345_));
 sg13g2_a21o_1 _27552_ (.A2(_07344_),
    .A1(_11244_),
    .B1(_07345_),
    .X(_07346_));
 sg13g2_a22oi_1 _27553_ (.Y(_07347_),
    .B1(_07346_),
    .B2(net637),
    .A2(net66),
    .A1(_11244_));
 sg13g2_a21oi_1 _27554_ (.A1(_07343_),
    .A2(_07347_),
    .Y(_01782_),
    .B1(_07312_));
 sg13g2_nor2_1 _27555_ (.A(_11323_),
    .B(_08631_),
    .Y(_07348_));
 sg13g2_buf_1 _27556_ (.A(_07348_),
    .X(_07349_));
 sg13g2_buf_1 _27557_ (.A(_07349_),
    .X(_07350_));
 sg13g2_nor2_1 _27558_ (.A(_11846_),
    .B(net322),
    .Y(_07351_));
 sg13g2_mux2_1 _27559_ (.A0(_11268_),
    .A1(_11267_),
    .S(_05722_),
    .X(_07352_));
 sg13g2_nor2_1 _27560_ (.A(net323),
    .B(_07352_),
    .Y(_07353_));
 sg13g2_nor3_1 _27561_ (.A(net629),
    .B(_07351_),
    .C(_07353_),
    .Y(_01783_));
 sg13g2_nor2_1 _27562_ (.A(_08533_),
    .B(net322),
    .Y(_07354_));
 sg13g2_mux2_1 _27563_ (.A0(_11242_),
    .A1(_11291_),
    .S(net73),
    .X(_07355_));
 sg13g2_nor2_1 _27564_ (.A(net323),
    .B(_07355_),
    .Y(_07356_));
 sg13g2_nor3_1 _27565_ (.A(net629),
    .B(_07354_),
    .C(_07356_),
    .Y(_01784_));
 sg13g2_nor2_1 _27566_ (.A(_08532_),
    .B(net322),
    .Y(_07357_));
 sg13g2_nand2_1 _27567_ (.Y(_07358_),
    .A(_11239_),
    .B(_05721_));
 sg13g2_o21ai_1 _27568_ (.B1(_07358_),
    .Y(_07359_),
    .A1(_11241_),
    .A2(net73));
 sg13g2_nor2_1 _27569_ (.A(net323),
    .B(_07359_),
    .Y(_07360_));
 sg13g2_nor3_1 _27570_ (.A(net629),
    .B(_07357_),
    .C(_07360_),
    .Y(_01785_));
 sg13g2_nor2_1 _27571_ (.A(_08538_),
    .B(net322),
    .Y(_07361_));
 sg13g2_buf_1 _27572_ (.A(_11322_),
    .X(_07362_));
 sg13g2_mux2_1 _27573_ (.A0(_11236_),
    .A1(_11237_),
    .S(net75),
    .X(_07363_));
 sg13g2_nor2_1 _27574_ (.A(net323),
    .B(_07363_),
    .Y(_07364_));
 sg13g2_nor3_1 _27575_ (.A(net629),
    .B(_07361_),
    .C(_07364_),
    .Y(_01786_));
 sg13g2_nor2_1 _27576_ (.A(_08537_),
    .B(_07350_),
    .Y(_07365_));
 sg13g2_mux2_1 _27577_ (.A0(_11234_),
    .A1(_11233_),
    .S(net75),
    .X(_07366_));
 sg13g2_nor2_1 _27578_ (.A(net323),
    .B(_07366_),
    .Y(_07367_));
 sg13g2_nor3_1 _27579_ (.A(net629),
    .B(_07365_),
    .C(_07367_),
    .Y(_01787_));
 sg13g2_nor2_1 _27580_ (.A(_08536_),
    .B(net322),
    .Y(_07368_));
 sg13g2_mux2_1 _27581_ (.A0(_11232_),
    .A1(_11231_),
    .S(_07362_),
    .X(_07369_));
 sg13g2_nor2_1 _27582_ (.A(net323),
    .B(_07369_),
    .Y(_07370_));
 sg13g2_nor3_1 _27583_ (.A(net629),
    .B(_07368_),
    .C(_07370_),
    .Y(_01788_));
 sg13g2_nor2_1 _27584_ (.A(_08535_),
    .B(net322),
    .Y(_07371_));
 sg13g2_mux2_1 _27585_ (.A0(_11229_),
    .A1(_11228_),
    .S(_07362_),
    .X(_07372_));
 sg13g2_nor2_1 _27586_ (.A(_05720_),
    .B(_07372_),
    .Y(_07373_));
 sg13g2_nor3_1 _27587_ (.A(_12780_),
    .B(_07371_),
    .C(_07373_),
    .Y(_01789_));
 sg13g2_nor2_1 _27588_ (.A(_08547_),
    .B(net322),
    .Y(_07374_));
 sg13g2_mux2_1 _27589_ (.A0(_11226_),
    .A1(_11227_),
    .S(net75),
    .X(_07375_));
 sg13g2_nor2_1 _27590_ (.A(net323),
    .B(_07375_),
    .Y(_07376_));
 sg13g2_nor3_1 _27591_ (.A(_12780_),
    .B(_07374_),
    .C(_07376_),
    .Y(_01790_));
 sg13g2_buf_1 _27592_ (.A(_08746_),
    .X(_07377_));
 sg13g2_nor2_1 _27593_ (.A(_08546_),
    .B(net322),
    .Y(_07378_));
 sg13g2_buf_1 _27594_ (.A(_11325_),
    .X(_07379_));
 sg13g2_nand2_1 _27595_ (.Y(_07380_),
    .A(_11224_),
    .B(net76));
 sg13g2_o21ai_1 _27596_ (.B1(_07380_),
    .Y(_07381_),
    .A1(_11223_),
    .A2(net73));
 sg13g2_nor2_1 _27597_ (.A(net321),
    .B(_07381_),
    .Y(_07382_));
 sg13g2_nor3_1 _27598_ (.A(net612),
    .B(_07378_),
    .C(_07382_),
    .Y(_01791_));
 sg13g2_nor2_1 _27599_ (.A(_08545_),
    .B(_07350_),
    .Y(_07383_));
 sg13g2_mux2_1 _27600_ (.A0(_11221_),
    .A1(_11311_),
    .S(net75),
    .X(_07384_));
 sg13g2_nor2_1 _27601_ (.A(net321),
    .B(_07384_),
    .Y(_07385_));
 sg13g2_nor3_1 _27602_ (.A(net612),
    .B(_07383_),
    .C(_07385_),
    .Y(_01792_));
 sg13g2_buf_1 _27603_ (.A(_07349_),
    .X(_07386_));
 sg13g2_nor2_1 _27604_ (.A(_08542_),
    .B(_07386_),
    .Y(_07387_));
 sg13g2_mux2_1 _27605_ (.A0(_11218_),
    .A1(_11219_),
    .S(net75),
    .X(_07388_));
 sg13g2_nor2_1 _27606_ (.A(_07379_),
    .B(_07388_),
    .Y(_07389_));
 sg13g2_nor3_1 _27607_ (.A(_07377_),
    .B(_07387_),
    .C(_07389_),
    .Y(_01793_));
 sg13g2_nor2_1 _27608_ (.A(_11796_),
    .B(net320),
    .Y(_07390_));
 sg13g2_nand2_1 _27609_ (.Y(_07391_),
    .A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(net76));
 sg13g2_o21ai_1 _27610_ (.B1(_07391_),
    .Y(_07392_),
    .A1(_07182_),
    .A2(_05722_));
 sg13g2_nor2_1 _27611_ (.A(net321),
    .B(_07392_),
    .Y(_07393_));
 sg13g2_nor3_1 _27612_ (.A(net612),
    .B(_07390_),
    .C(_07393_),
    .Y(_01794_));
 sg13g2_nor2_1 _27613_ (.A(_08543_),
    .B(_07386_),
    .Y(_07394_));
 sg13g2_mux2_1 _27614_ (.A0(_11317_),
    .A1(_11216_),
    .S(net75),
    .X(_07395_));
 sg13g2_nor2_1 _27615_ (.A(_07379_),
    .B(_07395_),
    .Y(_07396_));
 sg13g2_nor3_1 _27616_ (.A(_07377_),
    .B(_07394_),
    .C(_07396_),
    .Y(_01795_));
 sg13g2_nand2_1 _27617_ (.Y(_07397_),
    .A(_08481_),
    .B(net323));
 sg13g2_nand3_1 _27618_ (.B(_11214_),
    .C(_07349_),
    .A(_11212_),
    .Y(_07398_));
 sg13g2_a21oi_1 _27619_ (.A1(_07397_),
    .A2(_07398_),
    .Y(_01796_),
    .B1(_07312_));
 sg13g2_nor2_1 _27620_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(net320),
    .Y(_07399_));
 sg13g2_nand2_1 _27621_ (.Y(_07400_),
    .A(_11262_),
    .B(net76));
 sg13g2_o21ai_1 _27622_ (.B1(_07400_),
    .Y(_07401_),
    .A1(_11265_),
    .A2(net73));
 sg13g2_nor2_1 _27623_ (.A(net321),
    .B(_07401_),
    .Y(_07402_));
 sg13g2_nor3_1 _27624_ (.A(net612),
    .B(_07399_),
    .C(_07402_),
    .Y(_01797_));
 sg13g2_nor2_1 _27625_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(net320),
    .Y(_07403_));
 sg13g2_mux2_1 _27626_ (.A0(_11274_),
    .A1(_11261_),
    .S(net75),
    .X(_07404_));
 sg13g2_nor2_1 _27627_ (.A(net321),
    .B(_07404_),
    .Y(_07405_));
 sg13g2_nor3_1 _27628_ (.A(net612),
    .B(_07403_),
    .C(_07405_),
    .Y(_01798_));
 sg13g2_nor2_1 _27629_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(net320),
    .Y(_07406_));
 sg13g2_nand2_1 _27630_ (.Y(_07407_),
    .A(_11258_),
    .B(net76));
 sg13g2_o21ai_1 _27631_ (.B1(_07407_),
    .Y(_07408_),
    .A1(_11260_),
    .A2(net73));
 sg13g2_nor2_1 _27632_ (.A(net321),
    .B(_07408_),
    .Y(_07409_));
 sg13g2_nor3_1 _27633_ (.A(net612),
    .B(_07406_),
    .C(_07409_),
    .Y(_01799_));
 sg13g2_nor2_1 _27634_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(net320),
    .Y(_07410_));
 sg13g2_mux2_1 _27635_ (.A0(_11279_),
    .A1(_11256_),
    .S(net75),
    .X(_07411_));
 sg13g2_nor2_1 _27636_ (.A(net321),
    .B(_07411_),
    .Y(_07412_));
 sg13g2_nor3_1 _27637_ (.A(net612),
    .B(_07410_),
    .C(_07412_),
    .Y(_01800_));
 sg13g2_nor2_1 _27638_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(net320),
    .Y(_07413_));
 sg13g2_nand2_1 _27639_ (.Y(_07414_),
    .A(_11252_),
    .B(net76));
 sg13g2_o21ai_1 _27640_ (.B1(_07414_),
    .Y(_07415_),
    .A1(_11255_),
    .A2(net73));
 sg13g2_nor2_1 _27641_ (.A(net321),
    .B(_07415_),
    .Y(_07416_));
 sg13g2_nor3_1 _27642_ (.A(net612),
    .B(_07413_),
    .C(_07416_),
    .Y(_01801_));
 sg13g2_nor2_1 _27643_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(net320),
    .Y(_07417_));
 sg13g2_nand2_1 _27644_ (.Y(_07418_),
    .A(_11249_),
    .B(net76));
 sg13g2_o21ai_1 _27645_ (.B1(_07418_),
    .Y(_07419_),
    .A1(_11251_),
    .A2(net73));
 sg13g2_nor2_1 _27646_ (.A(_11325_),
    .B(_07419_),
    .Y(_07420_));
 sg13g2_nor3_1 _27647_ (.A(net680),
    .B(_07417_),
    .C(_07420_),
    .Y(_01802_));
 sg13g2_nor2_1 _27648_ (.A(_08541_),
    .B(net320),
    .Y(_07421_));
 sg13g2_mux2_1 _27649_ (.A0(_11246_),
    .A1(_11247_),
    .S(net76),
    .X(_07422_));
 sg13g2_nor2_1 _27650_ (.A(_11325_),
    .B(_07422_),
    .Y(_07423_));
 sg13g2_nor3_1 _27651_ (.A(_08747_),
    .B(_07421_),
    .C(_07423_),
    .Y(_01803_));
 sg13g2_nor2_1 _27652_ (.A(_08540_),
    .B(_07349_),
    .Y(_07424_));
 sg13g2_mux2_1 _27653_ (.A0(_11244_),
    .A1(_11243_),
    .S(net76),
    .X(_07425_));
 sg13g2_nor2_1 _27654_ (.A(_11325_),
    .B(_07425_),
    .Y(_07426_));
 sg13g2_nor3_1 _27655_ (.A(_08747_),
    .B(_07424_),
    .C(_07426_),
    .Y(_01804_));
 sg13g2_nor2_1 _27656_ (.A(_08414_),
    .B(net684),
    .Y(_07427_));
 sg13g2_nor2_1 _27657_ (.A(_05716_),
    .B(_05717_),
    .Y(_07428_));
 sg13g2_a21oi_1 _27658_ (.A1(_05716_),
    .A2(_07427_),
    .Y(_07429_),
    .B1(_07428_));
 sg13g2_nand3_1 _27659_ (.B(_05716_),
    .C(_07429_),
    .A(_11721_),
    .Y(_07430_));
 sg13g2_nand2_1 _27660_ (.Y(_07431_),
    .A(_11720_),
    .B(_07429_));
 sg13g2_nor2_1 _27661_ (.A(_08415_),
    .B(_07431_),
    .Y(_07432_));
 sg13g2_a21oi_1 _27662_ (.A1(_08415_),
    .A2(_07430_),
    .Y(_07433_),
    .B1(_07432_));
 sg13g2_nor2_1 _27663_ (.A(_08676_),
    .B(_07433_),
    .Y(_01805_));
 sg13g2_a21oi_1 _27664_ (.A1(_08415_),
    .A2(_05716_),
    .Y(_07434_),
    .B1(_07431_));
 sg13g2_nand2b_1 _27665_ (.Y(_07435_),
    .B(_07434_),
    .A_N(\rbzero.wall_tracer.w[1] ));
 sg13g2_o21ai_1 _27666_ (.B1(\rbzero.wall_tracer.w[1] ),
    .Y(_07436_),
    .A1(_08415_),
    .A2(_07430_));
 sg13g2_a21oi_1 _27667_ (.A1(_07435_),
    .A2(_07436_),
    .Y(_01806_),
    .B1(net613));
 sg13g2_xor2_1 _27668_ (.B(_08416_),
    .A(_00015_),
    .X(_07437_));
 sg13g2_a21oi_1 _27669_ (.A1(_05716_),
    .A2(_07437_),
    .Y(_07438_),
    .B1(_07431_));
 sg13g2_a21oi_1 _27670_ (.A1(\rbzero.wall_tracer.w[2] ),
    .A2(_07431_),
    .Y(_07439_),
    .B1(_07438_));
 sg13g2_nor2_1 _27671_ (.A(_08676_),
    .B(_07439_),
    .Y(_01807_));
 sg13g2_nor2_1 _27672_ (.A(_08572_),
    .B(_11327_),
    .Y(_07440_));
 sg13g2_nor2_1 _27673_ (.A(_08588_),
    .B(_08626_),
    .Y(_07441_));
 sg13g2_a221oi_1 _27674_ (.B2(\rbzero.mapdyw[0] ),
    .C1(_07441_),
    .B1(_07440_),
    .A1(\rbzero.mapdxw[0] ),
    .Y(_07442_),
    .A2(_11333_));
 sg13g2_or2_1 _27675_ (.X(_07443_),
    .B(_07442_),
    .A(_08632_));
 sg13g2_nand2_1 _27676_ (.Y(_07444_),
    .A(\rbzero.wall_tracer.wall[0] ),
    .B(_08632_));
 sg13g2_a21oi_1 _27677_ (.A1(_07443_),
    .A2(_07444_),
    .Y(_01808_),
    .B1(net635));
 sg13g2_nor2_1 _27678_ (.A(_08588_),
    .B(_08601_),
    .Y(_07445_));
 sg13g2_a221oi_1 _27679_ (.B2(\rbzero.mapdyw[1] ),
    .C1(_07445_),
    .B1(_07440_),
    .A1(\rbzero.mapdxw[1] ),
    .Y(_07446_),
    .A2(_11333_));
 sg13g2_or2_1 _27680_ (.X(_07447_),
    .B(_07446_),
    .A(_08632_));
 sg13g2_nand2_1 _27681_ (.Y(_07448_),
    .A(\rbzero.wall_tracer.wall[1] ),
    .B(_08632_));
 sg13g2_a21oi_1 _27682_ (.A1(_07447_),
    .A2(_07448_),
    .Y(_01809_),
    .B1(net635));
 sg13g2_inv_1 _27683_ (.Y(_07449_),
    .A(_00029_));
 sg13g2_mux4_1 _27684_ (.S0(net695),
    .A0(\rbzero.spi_registers.texadd3[22] ),
    .A1(\rbzero.spi_registers.texadd1[22] ),
    .A2(_07449_),
    .A3(\rbzero.spi_registers.texadd2[22] ),
    .S1(net628),
    .X(_07450_));
 sg13g2_inv_1 _27685_ (.Y(_07451_),
    .A(_00030_));
 sg13g2_mux4_1 _27686_ (.S0(_02002_),
    .A0(\rbzero.spi_registers.texadd3[21] ),
    .A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(_07451_),
    .A3(\rbzero.spi_registers.texadd2[21] ),
    .S1(_01996_),
    .X(_07452_));
 sg13g2_inv_1 _27687_ (.Y(_07453_),
    .A(_00031_));
 sg13g2_mux4_1 _27688_ (.S0(net695),
    .A0(\rbzero.spi_registers.texadd3[20] ),
    .A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(_07453_),
    .A3(\rbzero.spi_registers.texadd2[20] ),
    .S1(net696),
    .X(_07454_));
 sg13g2_inv_1 _27689_ (.Y(_07455_),
    .A(_00032_));
 sg13g2_mux4_1 _27690_ (.S0(net695),
    .A0(\rbzero.spi_registers.texadd3[19] ),
    .A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(_07455_),
    .A3(\rbzero.spi_registers.texadd2[19] ),
    .S1(net696),
    .X(_07456_));
 sg13g2_inv_1 _27691_ (.Y(_07457_),
    .A(_00034_));
 sg13g2_mux4_1 _27692_ (.S0(net695),
    .A0(\rbzero.spi_registers.texadd3[17] ),
    .A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(_07457_),
    .A3(\rbzero.spi_registers.texadd2[17] ),
    .S1(net696),
    .X(_07458_));
 sg13g2_inv_1 _27693_ (.Y(_07459_),
    .A(\rbzero.spi_registers.texadd3[16] ));
 sg13g2_inv_1 _27694_ (.Y(_07460_),
    .A(\rbzero.spi_registers.texadd1[16] ));
 sg13g2_inv_1 _27695_ (.Y(_07461_),
    .A(\rbzero.spi_registers.texadd2[16] ));
 sg13g2_mux4_1 _27696_ (.S0(net695),
    .A0(_07459_),
    .A1(_07460_),
    .A2(_00035_),
    .A3(_07461_),
    .S1(net696),
    .X(_07462_));
 sg13g2_inv_1 _27697_ (.Y(_07463_),
    .A(_00036_));
 sg13g2_mux4_1 _27698_ (.S0(net738),
    .A0(\rbzero.spi_registers.texadd3[15] ),
    .A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(_07463_),
    .A3(\rbzero.spi_registers.texadd2[15] ),
    .S1(net696),
    .X(_07464_));
 sg13g2_buf_1 _27699_ (.A(_07464_),
    .X(_07465_));
 sg13g2_and2_1 _27700_ (.A(net739),
    .B(net738),
    .X(_07466_));
 sg13g2_buf_1 _27701_ (.A(_07466_),
    .X(_07467_));
 sg13g2_nor2_1 _27702_ (.A(net696),
    .B(net738),
    .Y(_07468_));
 sg13g2_a22oi_1 _27703_ (.Y(_07469_),
    .B1(_07468_),
    .B2(\rbzero.spi_registers.texadd3[14] ),
    .A2(_07467_),
    .A1(\rbzero.spi_registers.texadd2[14] ));
 sg13g2_buf_1 _27704_ (.A(_07469_),
    .X(_07470_));
 sg13g2_inv_1 _27705_ (.Y(_07471_),
    .A(\rbzero.spi_registers.texadd2[13] ));
 sg13g2_mux2_1 _27706_ (.A0(_00038_),
    .A1(_07471_),
    .S(net738),
    .X(_07472_));
 sg13g2_mux2_1 _27707_ (.A0(\rbzero.spi_registers.texadd3[13] ),
    .A1(\rbzero.spi_registers.texadd1[13] ),
    .S(net738),
    .X(_07473_));
 sg13g2_nand2b_1 _27708_ (.Y(_07474_),
    .B(_07473_),
    .A_N(net739));
 sg13g2_inv_1 _27709_ (.Y(_07475_),
    .A(_00039_));
 sg13g2_mux4_1 _27710_ (.S0(net738),
    .A0(\rbzero.spi_registers.texadd3[12] ),
    .A1(\rbzero.spi_registers.texadd1[12] ),
    .A2(_07475_),
    .A3(\rbzero.spi_registers.texadd2[12] ),
    .S1(net739),
    .X(_07476_));
 sg13g2_inv_1 _27711_ (.Y(_07477_),
    .A(\rbzero.side_hot ));
 sg13g2_inv_1 _27712_ (.Y(_07478_),
    .A(_07476_));
 sg13g2_inv_1 _27713_ (.Y(_07479_),
    .A(_00040_));
 sg13g2_mux4_1 _27714_ (.S0(net738),
    .A0(\rbzero.spi_registers.texadd3[11] ),
    .A1(\rbzero.spi_registers.texadd1[11] ),
    .A2(_07479_),
    .A3(\rbzero.spi_registers.texadd2[11] ),
    .S1(net739),
    .X(_07480_));
 sg13g2_inv_1 _27715_ (.Y(_07481_),
    .A(_00042_));
 sg13g2_mux4_1 _27716_ (.S0(_02000_),
    .A0(\rbzero.spi_registers.texadd3[9] ),
    .A1(\rbzero.spi_registers.texadd1[9] ),
    .A2(_07481_),
    .A3(\rbzero.spi_registers.texadd2[9] ),
    .S1(_01995_),
    .X(_07482_));
 sg13g2_nor2_1 _27717_ (.A(_01979_),
    .B(_07482_),
    .Y(_07483_));
 sg13g2_inv_1 _27718_ (.Y(_07484_),
    .A(_00043_));
 sg13g2_mux4_1 _27719_ (.S0(_02000_),
    .A0(\rbzero.spi_registers.texadd3[8] ),
    .A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(_07484_),
    .A3(\rbzero.spi_registers.texadd2[8] ),
    .S1(_01995_),
    .X(_07485_));
 sg13g2_inv_1 _27720_ (.Y(_07486_),
    .A(_00044_));
 sg13g2_mux4_1 _27721_ (.S0(_02000_),
    .A0(\rbzero.spi_registers.texadd3[7] ),
    .A1(\rbzero.spi_registers.texadd1[7] ),
    .A2(_07486_),
    .A3(\rbzero.spi_registers.texadd2[7] ),
    .S1(_01994_),
    .X(_07487_));
 sg13g2_nand2_1 _27722_ (.Y(_07488_),
    .A(_01974_),
    .B(_07487_));
 sg13g2_inv_1 _27723_ (.Y(_07489_),
    .A(_00045_));
 sg13g2_mux4_1 _27724_ (.S0(_02000_),
    .A0(\rbzero.spi_registers.texadd3[6] ),
    .A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(_07489_),
    .A3(\rbzero.spi_registers.texadd2[6] ),
    .S1(_01994_),
    .X(_07490_));
 sg13g2_and2_1 _27725_ (.A(\rbzero.texu_hot[0] ),
    .B(_07490_),
    .X(_07491_));
 sg13g2_o21ai_1 _27726_ (.B1(_07491_),
    .Y(_07492_),
    .A1(_01974_),
    .A2(_07487_));
 sg13g2_nand2_1 _27727_ (.Y(_07493_),
    .A(_07488_),
    .B(_07492_));
 sg13g2_nand2_1 _27728_ (.Y(_07494_),
    .A(_07485_),
    .B(_07493_));
 sg13g2_o21ai_1 _27729_ (.B1(\rbzero.texu_hot[2] ),
    .Y(_07495_),
    .A1(_07485_),
    .A2(_07493_));
 sg13g2_nand2_1 _27730_ (.Y(_07496_),
    .A(_07494_),
    .B(_07495_));
 sg13g2_a21oi_1 _27731_ (.A1(_01979_),
    .A2(_07482_),
    .Y(_07497_),
    .B1(_07496_));
 sg13g2_nor2_1 _27732_ (.A(_07483_),
    .B(_07497_),
    .Y(_07498_));
 sg13g2_inv_1 _27733_ (.Y(_07499_),
    .A(_00041_));
 sg13g2_mux4_1 _27734_ (.S0(_02000_),
    .A0(\rbzero.spi_registers.texadd3[10] ),
    .A1(\rbzero.spi_registers.texadd1[10] ),
    .A2(_07499_),
    .A3(\rbzero.spi_registers.texadd2[10] ),
    .S1(net739),
    .X(_07500_));
 sg13g2_a21o_1 _27735_ (.A2(_07500_),
    .A1(_07498_),
    .B1(\rbzero.texu_hot[4] ),
    .X(_07501_));
 sg13g2_o21ai_1 _27736_ (.B1(_07501_),
    .Y(_07502_),
    .A1(_07498_),
    .A2(_07500_));
 sg13g2_nand2_1 _27737_ (.Y(_07503_),
    .A(_01984_),
    .B(_07480_));
 sg13g2_nand2_1 _27738_ (.Y(_07504_),
    .A(_07502_),
    .B(_07503_));
 sg13g2_o21ai_1 _27739_ (.B1(_07504_),
    .Y(_07505_),
    .A1(_01984_),
    .A2(_07480_));
 sg13g2_a21oi_1 _27740_ (.A1(_07477_),
    .A2(_07478_),
    .Y(_07506_),
    .B1(_07505_));
 sg13g2_a21oi_1 _27741_ (.A1(\rbzero.side_hot ),
    .A2(_07476_),
    .Y(_07507_),
    .B1(_07506_));
 sg13g2_a22oi_1 _27742_ (.Y(_07508_),
    .B1(_07474_),
    .B2(_07507_),
    .A2(_07472_),
    .A1(net696));
 sg13g2_nor2b_1 _27743_ (.A(_02001_),
    .B_N(net739),
    .Y(_07509_));
 sg13g2_nand2b_1 _27744_ (.Y(_07510_),
    .B(net738),
    .A_N(net739));
 sg13g2_nor2_1 _27745_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_07510_),
    .Y(_07511_));
 sg13g2_a21oi_2 _27746_ (.B1(_07511_),
    .Y(_07512_),
    .A2(_07509_),
    .A1(_00037_));
 sg13g2_nand2_1 _27747_ (.Y(_07513_),
    .A(_07508_),
    .B(_07512_));
 sg13g2_nand2_1 _27748_ (.Y(_07514_),
    .A(_07470_),
    .B(_07513_));
 sg13g2_nand2_1 _27749_ (.Y(_07515_),
    .A(_07465_),
    .B(_07514_));
 sg13g2_nor2_1 _27750_ (.A(_07462_),
    .B(_07515_),
    .Y(_07516_));
 sg13g2_and2_1 _27751_ (.A(_07458_),
    .B(_07516_),
    .X(_07517_));
 sg13g2_buf_1 _27752_ (.A(_07517_),
    .X(_07518_));
 sg13g2_inv_1 _27753_ (.Y(_07519_),
    .A(_00033_));
 sg13g2_mux4_1 _27754_ (.S0(net695),
    .A0(\rbzero.spi_registers.texadd3[18] ),
    .A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(_07519_),
    .A3(\rbzero.spi_registers.texadd2[18] ),
    .S1(net696),
    .X(_07520_));
 sg13g2_and3_1 _27755_ (.X(_07521_),
    .A(_07456_),
    .B(_07518_),
    .C(_07520_));
 sg13g2_buf_1 _27756_ (.A(_07521_),
    .X(_07522_));
 sg13g2_and3_1 _27757_ (.X(_07523_),
    .A(_07452_),
    .B(_07454_),
    .C(_07522_));
 sg13g2_xnor2_1 _27758_ (.Y(_07524_),
    .A(_07450_),
    .B(_07523_));
 sg13g2_mux4_1 _27759_ (.S0(_02002_),
    .A0(\rbzero.spi_registers.texadd3[23] ),
    .A1(\rbzero.spi_registers.texadd1[23] ),
    .A2(\rbzero.spi_registers.texadd0[23] ),
    .A3(\rbzero.spi_registers.texadd2[23] ),
    .S1(net628),
    .X(_07525_));
 sg13g2_and2_1 _27760_ (.A(_07450_),
    .B(_07523_),
    .X(_07526_));
 sg13g2_nor3_1 _27761_ (.A(net783),
    .B(_07525_),
    .C(_07526_),
    .Y(_07527_));
 sg13g2_a21o_1 _27762_ (.A2(_07526_),
    .A1(_07525_),
    .B1(_07527_),
    .X(_07528_));
 sg13g2_a21o_1 _27763_ (.A2(_07524_),
    .A1(net723),
    .B1(_07528_),
    .X(_07529_));
 sg13g2_nor2_1 _27764_ (.A(net783),
    .B(_07452_),
    .Y(_07530_));
 sg13g2_inv_1 _27765_ (.Y(_07531_),
    .A(_07454_));
 sg13g2_nand2_1 _27766_ (.Y(_07532_),
    .A(_07530_),
    .B(_07531_));
 sg13g2_nor2_1 _27767_ (.A(_07530_),
    .B(_07531_),
    .Y(_07533_));
 sg13g2_a21oi_1 _27768_ (.A1(net783),
    .A2(_07531_),
    .Y(_07534_),
    .B1(_07530_));
 sg13g2_nor2_1 _27769_ (.A(_07522_),
    .B(_07534_),
    .Y(_07535_));
 sg13g2_a21oi_1 _27770_ (.A1(_07522_),
    .A2(_07533_),
    .Y(_07536_),
    .B1(_07535_));
 sg13g2_nand3_1 _27771_ (.B(_07532_),
    .C(_07536_),
    .A(net754),
    .Y(_07537_));
 sg13g2_o21ai_1 _27772_ (.B1(_07537_),
    .Y(_07538_),
    .A1(net754),
    .A2(_07529_));
 sg13g2_buf_1 _27773_ (.A(net783),
    .X(_07539_));
 sg13g2_nor3_1 _27774_ (.A(net687),
    .B(_07458_),
    .C(_07516_),
    .Y(_07540_));
 sg13g2_xnor2_1 _27775_ (.Y(_07541_),
    .A(_07462_),
    .B(_07515_));
 sg13g2_and2_1 _27776_ (.A(net687),
    .B(_07541_),
    .X(_07542_));
 sg13g2_nor3_1 _27777_ (.A(_07518_),
    .B(_07540_),
    .C(_07542_),
    .Y(_07543_));
 sg13g2_nand2_1 _27778_ (.Y(_07544_),
    .A(_07518_),
    .B(_07520_));
 sg13g2_nor2_1 _27779_ (.A(net687),
    .B(_07456_),
    .Y(_07545_));
 sg13g2_xnor2_1 _27780_ (.Y(_07546_),
    .A(_07518_),
    .B(_07520_));
 sg13g2_a221oi_1 _27781_ (.B2(net723),
    .C1(_07522_),
    .B1(_07546_),
    .A1(_07544_),
    .Y(_07547_),
    .A2(_07545_));
 sg13g2_mux2_1 _27782_ (.A0(_07543_),
    .A1(_07547_),
    .S(_09696_),
    .X(_07548_));
 sg13g2_or2_1 _27783_ (.X(_07549_),
    .B(_07487_),
    .A(_01974_));
 sg13g2_a21o_1 _27784_ (.A2(_07549_),
    .A1(_07488_),
    .B1(_08709_),
    .X(_07550_));
 sg13g2_inv_1 _27785_ (.Y(_07551_),
    .A(\rbzero.texu_hot[0] ));
 sg13g2_nand2_1 _27786_ (.Y(_07552_),
    .A(_08709_),
    .B(_07551_));
 sg13g2_a21oi_1 _27787_ (.A1(_07550_),
    .A2(_07552_),
    .Y(_07553_),
    .B1(_07490_));
 sg13g2_mux2_1 _27788_ (.A0(_07551_),
    .A1(_07491_),
    .S(_07550_),
    .X(_07554_));
 sg13g2_or2_1 _27789_ (.X(_07555_),
    .B(_07554_),
    .A(_07553_));
 sg13g2_mux2_1 _27790_ (.A0(\rbzero.spi_registers.texadd0[5] ),
    .A1(\rbzero.spi_registers.texadd0[4] ),
    .S(net687),
    .X(_07556_));
 sg13g2_o21ai_1 _27791_ (.B1(_07509_),
    .Y(_07557_),
    .A1(_09696_),
    .A2(_07556_));
 sg13g2_nor2b_1 _27792_ (.A(net627),
    .B_N(\rbzero.spi_registers.texadd3[4] ),
    .Y(_07558_));
 sg13g2_a21oi_1 _27793_ (.A1(net627),
    .A2(\rbzero.spi_registers.texadd1[4] ),
    .Y(_07559_),
    .B1(_07558_));
 sg13g2_nand2_1 _27794_ (.Y(_07560_),
    .A(\rbzero.spi_registers.texadd2[4] ),
    .B(_07467_));
 sg13g2_o21ai_1 _27795_ (.B1(_07560_),
    .Y(_07561_),
    .A1(net628),
    .A2(_07559_));
 sg13g2_o21ai_1 _27796_ (.B1(net627),
    .Y(_07562_),
    .A1(\rbzero.spi_registers.texadd2[5] ),
    .A2(_09699_));
 sg13g2_or2_1 _27797_ (.X(_07563_),
    .B(\rbzero.spi_registers.texadd3[5] ),
    .A(net695));
 sg13g2_o21ai_1 _27798_ (.B1(_07563_),
    .Y(_07564_),
    .A1(\rbzero.spi_registers.texadd1[5] ),
    .A2(_07510_));
 sg13g2_nor2b_1 _27799_ (.A(_09699_),
    .B_N(_07564_),
    .Y(_07565_));
 sg13g2_a21oi_1 _27800_ (.A1(_01997_),
    .A2(_07562_),
    .Y(_07566_),
    .B1(_07565_));
 sg13g2_o21ai_1 _27801_ (.B1(_07566_),
    .Y(_07567_),
    .A1(_09703_),
    .A2(_07561_));
 sg13g2_a22oi_1 _27802_ (.Y(_07568_),
    .B1(_07557_),
    .B2(_07567_),
    .A2(_07555_),
    .A1(_09696_));
 sg13g2_nor2b_1 _27803_ (.A(net627),
    .B_N(\rbzero.spi_registers.texadd3[2] ),
    .Y(_07569_));
 sg13g2_a21oi_1 _27804_ (.A1(net627),
    .A2(\rbzero.spi_registers.texadd1[2] ),
    .Y(_07570_),
    .B1(_07569_));
 sg13g2_nand2_1 _27805_ (.Y(_07571_),
    .A(\rbzero.spi_registers.texadd2[2] ),
    .B(_07467_));
 sg13g2_o21ai_1 _27806_ (.B1(_07571_),
    .Y(_07572_),
    .A1(net628),
    .A2(_07570_));
 sg13g2_nor3_1 _27807_ (.A(net754),
    .B(net783),
    .C(\rbzero.spi_registers.texadd2[3] ),
    .Y(_07573_));
 sg13g2_nand2b_1 _27808_ (.Y(_07574_),
    .B(net627),
    .A_N(_07573_));
 sg13g2_or2_1 _27809_ (.X(_07575_),
    .B(\rbzero.spi_registers.texadd3[3] ),
    .A(net627));
 sg13g2_o21ai_1 _27810_ (.B1(_07575_),
    .Y(_07576_),
    .A1(\rbzero.spi_registers.texadd1[3] ),
    .A2(_07510_));
 sg13g2_nor2_1 _27811_ (.A(net754),
    .B(net687),
    .Y(_07577_));
 sg13g2_a22oi_1 _27812_ (.Y(_07578_),
    .B1(_07576_),
    .B2(_07577_),
    .A2(_07574_),
    .A1(net628));
 sg13g2_o21ai_1 _27813_ (.B1(_07578_),
    .Y(_07579_),
    .A1(_09697_),
    .A2(_07572_));
 sg13g2_mux2_1 _27814_ (.A0(\rbzero.spi_registers.texadd0[3] ),
    .A1(\rbzero.spi_registers.texadd0[2] ),
    .S(net687),
    .X(_07580_));
 sg13g2_o21ai_1 _27815_ (.B1(_07509_),
    .Y(_07581_),
    .A1(net754),
    .A2(_07580_));
 sg13g2_mux4_1 _27816_ (.S0(net627),
    .A0(\rbzero.spi_registers.texadd3[1] ),
    .A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(\rbzero.spi_registers.texadd0[1] ),
    .A3(\rbzero.spi_registers.texadd2[1] ),
    .S1(net628),
    .X(_07582_));
 sg13g2_mux4_1 _27817_ (.S0(_02003_),
    .A0(\rbzero.spi_registers.texadd3[0] ),
    .A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(\rbzero.spi_registers.texadd0[0] ),
    .A3(\rbzero.spi_registers.texadd2[0] ),
    .S1(net628),
    .X(_07583_));
 sg13g2_nand2b_1 _27818_ (.Y(_07584_),
    .B(net723),
    .A_N(_07583_));
 sg13g2_o21ai_1 _27819_ (.B1(_07584_),
    .Y(_07585_),
    .A1(net723),
    .A2(_07582_));
 sg13g2_a22oi_1 _27820_ (.Y(_07586_),
    .B1(_07585_),
    .B2(net754),
    .A2(_07581_),
    .A1(_07579_));
 sg13g2_mux4_1 _27821_ (.S0(net829),
    .A0(_07538_),
    .A1(_07548_),
    .A2(_07568_),
    .A3(_07586_),
    .S1(net796),
    .X(_07587_));
 sg13g2_xnor2_1 _27822_ (.Y(_07588_),
    .A(_07477_),
    .B(_07476_));
 sg13g2_xnor2_1 _27823_ (.Y(_07589_),
    .A(_07505_),
    .B(_07588_));
 sg13g2_mux2_1 _27824_ (.A0(_07473_),
    .A1(_07472_),
    .S(_01997_),
    .X(_07590_));
 sg13g2_xnor2_1 _27825_ (.Y(_07591_),
    .A(_07507_),
    .B(_07590_));
 sg13g2_nor2_1 _27826_ (.A(net687),
    .B(_07591_),
    .Y(_07592_));
 sg13g2_a21oi_1 _27827_ (.A1(net723),
    .A2(_07589_),
    .Y(_07593_),
    .B1(_07592_));
 sg13g2_mux2_1 _27828_ (.A0(_07512_),
    .A1(_07470_),
    .S(_07465_),
    .X(_07594_));
 sg13g2_nor2b_1 _27829_ (.A(_07465_),
    .B_N(_07470_),
    .Y(_07595_));
 sg13g2_nand3_1 _27830_ (.B(_07470_),
    .C(_07512_),
    .A(net828),
    .Y(_07596_));
 sg13g2_o21ai_1 _27831_ (.B1(_07596_),
    .Y(_07597_),
    .A1(net783),
    .A2(_07595_));
 sg13g2_mux2_1 _27832_ (.A0(_07465_),
    .A1(_07470_),
    .S(net828),
    .X(_07598_));
 sg13g2_nand2_1 _27833_ (.Y(_07599_),
    .A(_07512_),
    .B(_07598_));
 sg13g2_mux2_1 _27834_ (.A0(_07597_),
    .A1(_07599_),
    .S(_07508_),
    .X(_07600_));
 sg13g2_o21ai_1 _27835_ (.B1(_07600_),
    .Y(_07601_),
    .A1(net723),
    .A2(_07594_));
 sg13g2_xnor2_1 _27836_ (.Y(_07602_),
    .A(_01979_),
    .B(_07482_));
 sg13g2_xnor2_1 _27837_ (.Y(_07603_),
    .A(_07496_),
    .B(_07602_));
 sg13g2_xor2_1 _27838_ (.B(_07485_),
    .A(\rbzero.texu_hot[2] ),
    .X(_07604_));
 sg13g2_xnor2_1 _27839_ (.Y(_07605_),
    .A(_07493_),
    .B(_07604_));
 sg13g2_nand2_1 _27840_ (.Y(_07606_),
    .A(net687),
    .B(_07605_));
 sg13g2_o21ai_1 _27841_ (.B1(_07606_),
    .Y(_07607_),
    .A1(_07539_),
    .A2(_07603_));
 sg13g2_xor2_1 _27842_ (.B(_07480_),
    .A(_01984_),
    .X(_07608_));
 sg13g2_xnor2_1 _27843_ (.Y(_07609_),
    .A(_07502_),
    .B(_07608_));
 sg13g2_xor2_1 _27844_ (.B(_07500_),
    .A(\rbzero.texu_hot[4] ),
    .X(_07610_));
 sg13g2_xnor2_1 _27845_ (.Y(_07611_),
    .A(_07498_),
    .B(_07610_));
 sg13g2_nand2_1 _27846_ (.Y(_07612_),
    .A(_07539_),
    .B(_07611_));
 sg13g2_o21ai_1 _27847_ (.B1(_07612_),
    .Y(_07613_),
    .A1(_08710_),
    .A2(_07609_));
 sg13g2_mux4_1 _27848_ (.S0(_09696_),
    .A0(_07593_),
    .A1(_07601_),
    .A2(_07607_),
    .A3(_07613_),
    .S1(net829),
    .X(_07614_));
 sg13g2_or2_1 _27849_ (.X(_07615_),
    .B(_07614_),
    .A(net796));
 sg13g2_xnor2_1 _27850_ (.Y(_07616_),
    .A(net785),
    .B(_08664_));
 sg13g2_xnor2_1 _27851_ (.Y(_07617_),
    .A(net786),
    .B(_07616_));
 sg13g2_a21oi_1 _27852_ (.A1(net830),
    .A2(_07615_),
    .Y(_07618_),
    .B1(_07617_));
 sg13g2_o21ai_1 _27853_ (.B1(_07618_),
    .Y(_07619_),
    .A1(net830),
    .A2(_07587_));
 sg13g2_nor3_1 _27854_ (.A(net830),
    .B(net796),
    .C(_09718_),
    .Y(_07620_));
 sg13g2_nor2_1 _27855_ (.A(_08653_),
    .B(_07620_),
    .Y(_07621_));
 sg13g2_nor2_1 _27856_ (.A(_00014_),
    .B(_07621_),
    .Y(_07622_));
 sg13g2_o21ai_1 _27857_ (.B1(_09703_),
    .Y(_07623_),
    .A1(_09698_),
    .A2(_09693_));
 sg13g2_nand2_1 _27858_ (.Y(_07624_),
    .A(net829),
    .B(_09697_));
 sg13g2_o21ai_1 _27859_ (.B1(_07624_),
    .Y(_07625_),
    .A1(net829),
    .A2(_07623_));
 sg13g2_nand3_1 _27860_ (.B(_07622_),
    .C(_07625_),
    .A(_08653_),
    .Y(_07626_));
 sg13g2_o21ai_1 _27861_ (.B1(_07626_),
    .Y(_07627_),
    .A1(_07619_),
    .A2(_07622_));
 sg13g2_and2_1 _27862_ (.A(net13),
    .B(_07627_),
    .X(\rbzero.o_tex_out0 ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_or2_1 _27864_ (.X(_07628_),
    .B(_08461_),
    .A(_08456_));
 sg13g2_o21ai_1 _27865_ (.B1(_00051_),
    .Y(_07629_),
    .A1(_08453_),
    .A2(_07628_));
 sg13g2_o21ai_1 _27866_ (.B1(_08465_),
    .Y(_07630_),
    .A1(_08468_),
    .A2(_07629_));
 sg13g2_xor2_1 _27867_ (.B(_07630_),
    .A(_08466_),
    .X(_07631_));
 sg13g2_buf_1 _27868_ (.A(_07631_),
    .X(_07632_));
 sg13g2_and2_1 _27869_ (.A(_00014_),
    .B(_07632_),
    .X(_07633_));
 sg13g2_and3_1 _27870_ (.X(_07634_),
    .A(net796),
    .B(_09693_),
    .C(_09718_));
 sg13g2_xor2_1 _27871_ (.B(_07629_),
    .A(_08664_),
    .X(_07635_));
 sg13g2_buf_2 _27872_ (.A(_07635_),
    .X(_07636_));
 sg13g2_or3_1 _27873_ (.A(_08468_),
    .B(_08453_),
    .C(_08462_),
    .X(_07637_));
 sg13g2_xnor2_1 _27874_ (.Y(_07638_),
    .A(_09709_),
    .B(_07637_));
 sg13g2_buf_1 _27875_ (.A(_07638_),
    .X(_07639_));
 sg13g2_nor2_1 _27876_ (.A(_07636_),
    .B(net493),
    .Y(_07640_));
 sg13g2_and3_1 _27877_ (.X(_07641_),
    .A(_08465_),
    .B(_08466_),
    .C(_07637_));
 sg13g2_buf_1 _27878_ (.A(_07641_),
    .X(_07642_));
 sg13g2_buf_2 _27879_ (.A(_00052_),
    .X(_07643_));
 sg13g2_inv_1 _27880_ (.Y(_07644_),
    .A(_07643_));
 sg13g2_o21ai_1 _27881_ (.B1(_07644_),
    .Y(_07645_),
    .A1(net831),
    .A2(_07642_));
 sg13g2_nand4_1 _27882_ (.B(_07634_),
    .C(_07640_),
    .A(_07633_),
    .Y(_07646_),
    .D(_07645_));
 sg13g2_nand3_1 _27883_ (.B(net831),
    .C(_07642_),
    .A(_08470_),
    .Y(_07647_));
 sg13g2_nand3_1 _27884_ (.B(_09406_),
    .C(_11185_),
    .A(_09404_),
    .Y(_07648_));
 sg13g2_nand3b_1 _27885_ (.B(net4),
    .C(_11182_),
    .Y(_07649_),
    .A_N(_09399_));
 sg13g2_a221oi_1 _27886_ (.B2(_09412_),
    .C1(_07649_),
    .B1(_07648_),
    .A1(_07643_),
    .Y(_07650_),
    .A2(_07647_));
 sg13g2_nand2_1 _27887_ (.Y(_07651_),
    .A(_07646_),
    .B(_07650_));
 sg13g2_buf_2 _27888_ (.A(_07651_),
    .X(_07652_));
 sg13g2_inv_1 _27889_ (.Y(_07653_),
    .A(_11758_));
 sg13g2_inv_1 _27890_ (.Y(_07654_),
    .A(_11724_));
 sg13g2_nor4_1 _27891_ (.A(_11742_),
    .B(_11739_),
    .C(_11736_),
    .D(net811),
    .Y(_07655_));
 sg13g2_nand3b_1 _27892_ (.B(_07654_),
    .C(_07655_),
    .Y(_07656_),
    .A_N(_11746_));
 sg13g2_a21oi_2 _27893_ (.B1(_11754_),
    .Y(_07657_),
    .A2(_07656_),
    .A1(_11750_));
 sg13g2_nor2_1 _27894_ (.A(_07653_),
    .B(_11729_),
    .Y(_07658_));
 sg13g2_a22oi_1 _27895_ (.Y(_07659_),
    .B1(_07657_),
    .B2(_07658_),
    .A2(_00047_),
    .A1(net730));
 sg13g2_or2_1 _27896_ (.X(_07660_),
    .B(_07659_),
    .A(_11762_));
 sg13g2_nand2_1 _27897_ (.Y(_07661_),
    .A(_00050_),
    .B(_07655_));
 sg13g2_nor2_1 _27898_ (.A(_11746_),
    .B(_07661_),
    .Y(_07662_));
 sg13g2_a21oi_1 _27899_ (.A1(_11750_),
    .A2(_07662_),
    .Y(_07663_),
    .B1(_00049_));
 sg13g2_nor3_1 _27900_ (.A(net730),
    .B(_11754_),
    .C(_07663_),
    .Y(_07664_));
 sg13g2_nor2_1 _27901_ (.A(net730),
    .B(_07664_),
    .Y(_07665_));
 sg13g2_xnor2_1 _27902_ (.Y(_07666_),
    .A(_11762_),
    .B(_07665_));
 sg13g2_xnor2_1 _27903_ (.Y(_07667_),
    .A(_07643_),
    .B(_07666_));
 sg13g2_buf_1 _27904_ (.A(_00053_),
    .X(_07668_));
 sg13g2_inv_1 _27905_ (.Y(_07669_),
    .A(_11750_));
 sg13g2_nor2_1 _27906_ (.A(_07669_),
    .B(_07662_),
    .Y(_07670_));
 sg13g2_xnor2_1 _27907_ (.Y(_07671_),
    .A(_11754_),
    .B(_07670_));
 sg13g2_xor2_1 _27908_ (.B(_07656_),
    .A(_00049_),
    .X(_07672_));
 sg13g2_nand2_1 _27909_ (.Y(_07673_),
    .A(_09709_),
    .B(_07672_));
 sg13g2_xnor2_1 _27910_ (.Y(_07674_),
    .A(_11746_),
    .B(_07661_));
 sg13g2_xnor2_1 _27911_ (.Y(_07675_),
    .A(_08664_),
    .B(_07674_));
 sg13g2_nor4_1 _27912_ (.A(_11739_),
    .B(_11736_),
    .C(_11724_),
    .D(_11732_),
    .Y(_07676_));
 sg13g2_xnor2_1 _27913_ (.Y(_07677_),
    .A(_11742_),
    .B(_07676_));
 sg13g2_inv_1 _27914_ (.Y(_07678_),
    .A(_00050_));
 sg13g2_nor3_1 _27915_ (.A(_11736_),
    .B(_11732_),
    .C(_07678_),
    .Y(_07679_));
 sg13g2_xnor2_1 _27916_ (.Y(_07680_),
    .A(_11739_),
    .B(_07679_));
 sg13g2_inv_1 _27917_ (.Y(_07681_),
    .A(_07680_));
 sg13g2_buf_1 _27918_ (.A(_00028_),
    .X(_07682_));
 sg13g2_nor3_1 _27919_ (.A(_08458_),
    .B(net811),
    .C(_07682_),
    .Y(_07683_));
 sg13g2_a21oi_1 _27920_ (.A1(net811),
    .A2(_07682_),
    .Y(_07684_),
    .B1(_07683_));
 sg13g2_inv_1 _27921_ (.Y(_07685_),
    .A(\rbzero.row_render.size[1] ));
 sg13g2_o21ai_1 _27922_ (.B1(net828),
    .Y(_07686_),
    .A1(_07685_),
    .A2(_07682_));
 sg13g2_nand2b_1 _27923_ (.Y(_07687_),
    .B(net828),
    .A_N(_07682_));
 sg13g2_a221oi_1 _27924_ (.B2(_07685_),
    .C1(_07654_),
    .B1(_07687_),
    .A1(_09696_),
    .Y(_07688_),
    .A2(_07686_));
 sg13g2_a21oi_1 _27925_ (.A1(_07654_),
    .A2(_07684_),
    .Y(_07689_),
    .B1(_07688_));
 sg13g2_nor2b_1 _27926_ (.A(_07689_),
    .B_N(_00027_),
    .Y(_07690_));
 sg13g2_nor2_1 _27927_ (.A(_11724_),
    .B(net811),
    .Y(_07691_));
 sg13g2_xor2_1 _27928_ (.B(_07691_),
    .A(_11736_),
    .X(_07692_));
 sg13g2_o21ai_1 _27929_ (.B1(_07692_),
    .Y(_07693_),
    .A1(net829),
    .A2(_07690_));
 sg13g2_or3_1 _27930_ (.A(_00027_),
    .B(_07689_),
    .C(_07692_),
    .X(_07694_));
 sg13g2_a22oi_1 _27931_ (.Y(_07695_),
    .B1(_07680_),
    .B2(_08456_),
    .A2(_07694_),
    .A1(_07693_));
 sg13g2_a21oi_1 _27932_ (.A1(net830),
    .A2(_07681_),
    .Y(_07696_),
    .B1(_07695_));
 sg13g2_a21o_1 _27933_ (.A2(_07696_),
    .A1(_07677_),
    .B1(_00051_),
    .X(_07697_));
 sg13g2_o21ai_1 _27934_ (.B1(_07697_),
    .Y(_07698_),
    .A1(_07677_),
    .A2(_07696_));
 sg13g2_a22oi_1 _27935_ (.Y(_07699_),
    .B1(_07675_),
    .B2(_07698_),
    .A2(_07674_),
    .A1(_08468_));
 sg13g2_o21ai_1 _27936_ (.B1(_07699_),
    .Y(_07700_),
    .A1(_09709_),
    .A2(_07672_));
 sg13g2_a22oi_1 _27937_ (.Y(_07701_),
    .B1(_07673_),
    .B2(_07700_),
    .A2(_07671_),
    .A1(net787));
 sg13g2_inv_1 _27938_ (.Y(_07702_),
    .A(_07701_));
 sg13g2_o21ai_1 _27939_ (.B1(_07702_),
    .Y(_07703_),
    .A1(net787),
    .A2(_07671_));
 sg13g2_xnor2_1 _27940_ (.Y(_07704_),
    .A(net730),
    .B(_07657_));
 sg13g2_a21o_1 _27941_ (.A2(_07703_),
    .A1(_07668_),
    .B1(_07704_),
    .X(_07705_));
 sg13g2_o21ai_1 _27942_ (.B1(_07705_),
    .Y(_07706_),
    .A1(_07668_),
    .A2(_07703_));
 sg13g2_a22oi_1 _27943_ (.Y(_07707_),
    .B1(_07667_),
    .B2(_07706_),
    .A2(_07666_),
    .A1(_08469_));
 sg13g2_nor2_1 _27944_ (.A(_00048_),
    .B(_07664_),
    .Y(_07708_));
 sg13g2_nor2_1 _27945_ (.A(_11762_),
    .B(_11729_),
    .Y(_07709_));
 sg13g2_o21ai_1 _27946_ (.B1(_07709_),
    .Y(_07710_),
    .A1(net730),
    .A2(_07657_));
 sg13g2_nand2_2 _27947_ (.Y(_07711_),
    .A(_11754_),
    .B(_11750_));
 sg13g2_nand2_1 _27948_ (.Y(_07712_),
    .A(net730),
    .B(_07711_));
 sg13g2_nor2b_1 _27949_ (.A(_00048_),
    .B_N(_11729_),
    .Y(_07713_));
 sg13g2_a21o_1 _27950_ (.A2(_07712_),
    .A1(_00047_),
    .B1(_07713_),
    .X(_07714_));
 sg13g2_xnor2_1 _27951_ (.Y(_07715_),
    .A(net730),
    .B(_07711_));
 sg13g2_o21ai_1 _27952_ (.B1(_00048_),
    .Y(_07716_),
    .A1(_11758_),
    .A2(_07711_));
 sg13g2_xor2_1 _27953_ (.B(_07716_),
    .A(_11762_),
    .X(_07717_));
 sg13g2_xnor2_1 _27954_ (.Y(_07718_),
    .A(_07643_),
    .B(_07717_));
 sg13g2_a21oi_1 _27955_ (.A1(_07668_),
    .A2(_07715_),
    .Y(_07719_),
    .B1(_07718_));
 sg13g2_xnor2_1 _27956_ (.Y(_07720_),
    .A(_08457_),
    .B(_11736_));
 sg13g2_xnor2_1 _27957_ (.Y(_07721_),
    .A(net828),
    .B(_11724_));
 sg13g2_xnor2_1 _27958_ (.Y(_07722_),
    .A(net796),
    .B(_11742_));
 sg13g2_xor2_1 _27959_ (.B(_11739_),
    .A(net830),
    .X(_07723_));
 sg13g2_nor2b_1 _27960_ (.A(_08468_),
    .B_N(_11746_),
    .Y(_07724_));
 sg13g2_nand2b_1 _27961_ (.Y(_07725_),
    .B(_08468_),
    .A_N(_11746_));
 sg13g2_nand2b_1 _27962_ (.Y(_07726_),
    .B(_07725_),
    .A_N(_07724_));
 sg13g2_xnor2_1 _27963_ (.Y(_07727_),
    .A(_08465_),
    .B(_11750_));
 sg13g2_xor2_1 _27964_ (.B(net811),
    .A(_08458_),
    .X(_07728_));
 sg13g2_nor4_1 _27965_ (.A(_07723_),
    .B(_07726_),
    .C(_07727_),
    .D(_07728_),
    .Y(_07729_));
 sg13g2_nand4_1 _27966_ (.B(_07721_),
    .C(_07722_),
    .A(_07720_),
    .Y(_07730_),
    .D(_07729_));
 sg13g2_nor2_1 _27967_ (.A(_07668_),
    .B(_07715_),
    .Y(_07731_));
 sg13g2_xnor2_1 _27968_ (.Y(_07732_),
    .A(_11754_),
    .B(_11750_));
 sg13g2_xnor2_1 _27969_ (.Y(_07733_),
    .A(_08648_),
    .B(_07732_));
 sg13g2_nor3_1 _27970_ (.A(_07730_),
    .B(_07731_),
    .C(_07733_),
    .Y(_07734_));
 sg13g2_o21ai_1 _27971_ (.B1(net730),
    .Y(_07735_),
    .A1(_11729_),
    .A2(_07711_));
 sg13g2_a21oi_1 _27972_ (.A1(_11762_),
    .A2(_07735_),
    .Y(_07736_),
    .B1(_00047_));
 sg13g2_a221oi_1 _27973_ (.B2(_07734_),
    .C1(_07736_),
    .B1(_07719_),
    .A1(_11762_),
    .Y(_07737_),
    .A2(_07714_));
 sg13g2_inv_1 _27974_ (.Y(_07738_),
    .A(_11739_));
 sg13g2_nor2_1 _27975_ (.A(net828),
    .B(_07654_),
    .Y(_07739_));
 sg13g2_nor2_1 _27976_ (.A(net811),
    .B(_07739_),
    .Y(_07740_));
 sg13g2_a21oi_1 _27977_ (.A1(net811),
    .A2(_07739_),
    .Y(_07741_),
    .B1(_09696_));
 sg13g2_nor2_1 _27978_ (.A(_07740_),
    .B(_07741_),
    .Y(_07742_));
 sg13g2_nor2_1 _27979_ (.A(_11736_),
    .B(_07742_),
    .Y(_07743_));
 sg13g2_nor2_1 _27980_ (.A(_08457_),
    .B(_07743_),
    .Y(_07744_));
 sg13g2_a221oi_1 _27981_ (.B2(_07742_),
    .C1(_07744_),
    .B1(_11736_),
    .A1(_08456_),
    .Y(_07745_),
    .A2(_11739_));
 sg13g2_a21oi_1 _27982_ (.A1(net830),
    .A2(_07738_),
    .Y(_07746_),
    .B1(_07745_));
 sg13g2_nor2_1 _27983_ (.A(_11742_),
    .B(_07746_),
    .Y(_07747_));
 sg13g2_nand2_1 _27984_ (.Y(_07748_),
    .A(_11742_),
    .B(_07746_));
 sg13g2_o21ai_1 _27985_ (.B1(_07748_),
    .Y(_07749_),
    .A1(_08454_),
    .A2(_07747_));
 sg13g2_a21oi_2 _27986_ (.B1(_07724_),
    .Y(_07750_),
    .A2(_07749_),
    .A1(_07725_));
 sg13g2_o21ai_1 _27987_ (.B1(_08466_),
    .Y(_07751_),
    .A1(_07669_),
    .A2(_07750_));
 sg13g2_a21oi_1 _27988_ (.A1(_07669_),
    .A2(_07750_),
    .Y(_07752_),
    .B1(_08466_));
 sg13g2_a21oi_1 _27989_ (.A1(_09709_),
    .A2(_07751_),
    .Y(_07753_),
    .B1(_07752_));
 sg13g2_nand2_1 _27990_ (.Y(_07754_),
    .A(_11754_),
    .B(_07669_));
 sg13g2_o21ai_1 _27991_ (.B1(_07754_),
    .Y(_07755_),
    .A1(_08466_),
    .A2(_07750_));
 sg13g2_a21oi_1 _27992_ (.A1(_08648_),
    .A2(_07750_),
    .Y(_07756_),
    .B1(_07754_));
 sg13g2_a21oi_1 _27993_ (.A1(_09709_),
    .A2(_07755_),
    .Y(_07757_),
    .B1(_07756_));
 sg13g2_o21ai_1 _27994_ (.B1(_07757_),
    .Y(_07758_),
    .A1(_11754_),
    .A2(_07753_));
 sg13g2_nand2b_1 _27995_ (.Y(_07759_),
    .B(_07758_),
    .A_N(_07731_));
 sg13g2_nand2_1 _27996_ (.Y(_07760_),
    .A(_07719_),
    .B(_07759_));
 sg13g2_o21ai_1 _27997_ (.B1(_07760_),
    .Y(_07761_),
    .A1(_08470_),
    .A2(_07717_));
 sg13g2_and2_1 _27998_ (.A(_07737_),
    .B(_07761_),
    .X(_07762_));
 sg13g2_nor4_1 _27999_ (.A(_07707_),
    .B(_07708_),
    .C(_07710_),
    .D(_07762_),
    .Y(_07763_));
 sg13g2_xnor2_1 _28000_ (.Y(_07764_),
    .A(\rbzero.traced_texVinit[9] ),
    .B(_09668_));
 sg13g2_nor2_1 _28001_ (.A(_13882_),
    .B(_09646_),
    .Y(_07765_));
 sg13g2_a21oi_1 _28002_ (.A1(_13882_),
    .A2(_09646_),
    .Y(_07766_),
    .B1(_11179_));
 sg13g2_or2_1 _28003_ (.X(_07767_),
    .B(_07766_),
    .A(_07765_));
 sg13g2_nor2_1 _28004_ (.A(_07764_),
    .B(_07767_),
    .Y(_07768_));
 sg13g2_nor2_1 _28005_ (.A(_13726_),
    .B(_09642_),
    .Y(_07769_));
 sg13g2_a21oi_1 _28006_ (.A1(_13726_),
    .A2(_09642_),
    .Y(_07770_),
    .B1(\rbzero.spi_registers.vshift[4] ));
 sg13g2_nor2_1 _28007_ (.A(_07769_),
    .B(_07770_),
    .Y(_07771_));
 sg13g2_inv_1 _28008_ (.Y(_07772_),
    .A(_07771_));
 sg13g2_a21o_1 _28009_ (.A2(_09631_),
    .A1(_13561_),
    .B1(\rbzero.spi_registers.vshift[3] ),
    .X(_07773_));
 sg13g2_o21ai_1 _28010_ (.B1(_07773_),
    .Y(_07774_),
    .A1(_13561_),
    .A2(_09631_));
 sg13g2_buf_1 _28011_ (.A(_07774_),
    .X(_07775_));
 sg13g2_xor2_1 _28012_ (.B(_09631_),
    .A(_13561_),
    .X(_07776_));
 sg13g2_xnor2_1 _28013_ (.Y(_07777_),
    .A(\rbzero.spi_registers.vshift[3] ),
    .B(_07776_));
 sg13g2_inv_1 _28014_ (.Y(_07778_),
    .A(_07777_));
 sg13g2_xnor2_1 _28015_ (.Y(_07779_),
    .A(_13146_),
    .B(_09619_));
 sg13g2_xnor2_1 _28016_ (.Y(_07780_),
    .A(\rbzero.spi_registers.vshift[1] ),
    .B(_07779_));
 sg13g2_nor2_1 _28017_ (.A(\rbzero.traced_texVinit[2] ),
    .B(_09604_),
    .Y(_07781_));
 sg13g2_a21o_1 _28018_ (.A2(_09590_),
    .A1(\rbzero.traced_texVinit[0] ),
    .B1(_09594_),
    .X(_07782_));
 sg13g2_and3_1 _28019_ (.X(_07783_),
    .A(_09594_),
    .B(\rbzero.traced_texVinit[0] ),
    .C(_09590_));
 sg13g2_a221oi_1 _28020_ (.B2(_07782_),
    .C1(_07783_),
    .B1(\rbzero.traced_texVinit[1] ),
    .A1(\rbzero.traced_texVinit[2] ),
    .Y(_07784_),
    .A2(_09604_));
 sg13g2_nor2_1 _28021_ (.A(_07781_),
    .B(_07784_),
    .Y(_07785_));
 sg13g2_and2_1 _28022_ (.A(_09611_),
    .B(_07785_),
    .X(_07786_));
 sg13g2_buf_1 _28023_ (.A(_07786_),
    .X(_07787_));
 sg13g2_or2_1 _28024_ (.X(_07788_),
    .B(_07785_),
    .A(_09611_));
 sg13g2_buf_1 _28025_ (.A(_07788_),
    .X(_07789_));
 sg13g2_o21ai_1 _28026_ (.B1(_07789_),
    .Y(_07790_),
    .A1(_13144_),
    .A2(_07787_));
 sg13g2_inv_1 _28027_ (.Y(_07791_),
    .A(_07790_));
 sg13g2_o21ai_1 _28028_ (.B1(_13144_),
    .Y(_07792_),
    .A1(_07780_),
    .A2(_07787_));
 sg13g2_nand2_1 _28029_ (.Y(_07793_),
    .A(_07780_),
    .B(_07789_));
 sg13g2_nand2_1 _28030_ (.Y(_07794_),
    .A(_07792_),
    .B(_07793_));
 sg13g2_a22oi_1 _28031_ (.Y(_07795_),
    .B1(_07794_),
    .B2(_11167_),
    .A2(_07791_),
    .A1(_07780_));
 sg13g2_buf_1 _28032_ (.A(_07795_),
    .X(_07796_));
 sg13g2_nor2_1 _28033_ (.A(_13146_),
    .B(_09619_),
    .Y(_07797_));
 sg13g2_a21oi_1 _28034_ (.A1(_13146_),
    .A2(_09619_),
    .Y(_07798_),
    .B1(\rbzero.spi_registers.vshift[1] ));
 sg13g2_nor2_1 _28035_ (.A(_07797_),
    .B(_07798_),
    .Y(_07799_));
 sg13g2_nor2b_1 _28036_ (.A(_07796_),
    .B_N(_07799_),
    .Y(_07800_));
 sg13g2_buf_1 _28037_ (.A(_07800_),
    .X(_07801_));
 sg13g2_nand2_1 _28038_ (.Y(_07802_),
    .A(_13284_),
    .B(_09626_));
 sg13g2_or2_1 _28039_ (.X(_07803_),
    .B(_09626_),
    .A(_13284_));
 sg13g2_a21oi_1 _28040_ (.A1(_07803_),
    .A2(_07778_),
    .Y(_07804_),
    .B1(_11172_));
 sg13g2_a21oi_1 _28041_ (.A1(_07802_),
    .A2(_07777_),
    .Y(_07805_),
    .B1(_07804_));
 sg13g2_nand2b_1 _28042_ (.Y(_07806_),
    .B(_07796_),
    .A_N(_07799_));
 sg13g2_buf_1 _28043_ (.A(_07806_),
    .X(_07807_));
 sg13g2_nand2_1 _28044_ (.Y(_07808_),
    .A(_11172_),
    .B(_07803_));
 sg13g2_nor2_1 _28045_ (.A(_07778_),
    .B(_07801_),
    .Y(_07809_));
 sg13g2_a21oi_1 _28046_ (.A1(_07802_),
    .A2(_07808_),
    .Y(_07810_),
    .B1(_07809_));
 sg13g2_a221oi_1 _28047_ (.B2(_07807_),
    .C1(_07810_),
    .B1(_07805_),
    .A1(_07778_),
    .Y(_07811_),
    .A2(_07801_));
 sg13g2_buf_1 _28048_ (.A(_07811_),
    .X(_07812_));
 sg13g2_nor2_1 _28049_ (.A(_07775_),
    .B(_07812_),
    .Y(_07813_));
 sg13g2_xnor2_1 _28050_ (.Y(_07814_),
    .A(_13726_),
    .B(_09642_));
 sg13g2_xnor2_1 _28051_ (.Y(_07815_),
    .A(\rbzero.spi_registers.vshift[4] ),
    .B(_07814_));
 sg13g2_nand2_1 _28052_ (.Y(_07816_),
    .A(_07775_),
    .B(_07812_));
 sg13g2_o21ai_1 _28053_ (.B1(_07816_),
    .Y(_07817_),
    .A1(_07813_),
    .A2(_07815_));
 sg13g2_buf_1 _28054_ (.A(_07817_),
    .X(_07818_));
 sg13g2_a22oi_1 _28055_ (.Y(_07819_),
    .B1(_07764_),
    .B2(_07767_),
    .A2(_07818_),
    .A1(_07772_));
 sg13g2_nand2_1 _28056_ (.Y(_07820_),
    .A(_13882_),
    .B(_09646_));
 sg13g2_nand2_1 _28057_ (.Y(_07821_),
    .A(_07820_),
    .B(_07764_));
 sg13g2_nor2_1 _28058_ (.A(_07764_),
    .B(_07765_),
    .Y(_07822_));
 sg13g2_a21oi_1 _28059_ (.A1(_11179_),
    .A2(_07821_),
    .Y(_07823_),
    .B1(_07822_));
 sg13g2_o21ai_1 _28060_ (.B1(_07823_),
    .Y(_07824_),
    .A1(_07772_),
    .A2(_07818_));
 sg13g2_o21ai_1 _28061_ (.B1(_07824_),
    .Y(_07825_),
    .A1(_07768_),
    .A2(_07819_));
 sg13g2_xor2_1 _28062_ (.B(\rbzero.texV[10] ),
    .A(\rbzero.traced_texVinit[10] ),
    .X(_07826_));
 sg13g2_nand2_1 _28063_ (.Y(_07827_),
    .A(\rbzero.traced_texVinit[9] ),
    .B(_09668_));
 sg13g2_xnor2_1 _28064_ (.Y(_07828_),
    .A(_07826_),
    .B(_07827_));
 sg13g2_xnor2_1 _28065_ (.Y(_07829_),
    .A(_07825_),
    .B(_07828_));
 sg13g2_and2_1 _28066_ (.A(_00046_),
    .B(_07829_),
    .X(_07830_));
 sg13g2_buf_1 _28067_ (.A(_07830_),
    .X(_07831_));
 sg13g2_inv_1 _28068_ (.Y(_07832_),
    .A(_11167_));
 sg13g2_xnor2_1 _28069_ (.Y(_07833_),
    .A(_13144_),
    .B(_09611_));
 sg13g2_xnor2_1 _28070_ (.Y(_07834_),
    .A(_07832_),
    .B(_07833_));
 sg13g2_xnor2_1 _28071_ (.Y(_07835_),
    .A(_07785_),
    .B(_07834_));
 sg13g2_nand2b_1 _28072_ (.Y(_07836_),
    .B(_07835_),
    .A_N(_07831_));
 sg13g2_buf_1 _28073_ (.A(_07836_),
    .X(_07837_));
 sg13g2_buf_1 _28074_ (.A(_07837_),
    .X(_07838_));
 sg13g2_nand3_1 _28075_ (.B(_13144_),
    .C(_07787_),
    .A(_11167_),
    .Y(_07839_));
 sg13g2_o21ai_1 _28076_ (.B1(_07839_),
    .Y(_07840_),
    .A1(_13144_),
    .A2(_07789_));
 sg13g2_a21oi_1 _28077_ (.A1(_07832_),
    .A2(_07790_),
    .Y(_07841_),
    .B1(_07840_));
 sg13g2_xnor2_1 _28078_ (.Y(_07842_),
    .A(_07780_),
    .B(_07841_));
 sg13g2_or2_1 _28079_ (.X(_07843_),
    .B(_07842_),
    .A(_07831_));
 sg13g2_buf_1 _28080_ (.A(_07843_),
    .X(_07844_));
 sg13g2_xor2_1 _28081_ (.B(net755),
    .A(_13284_),
    .X(_07845_));
 sg13g2_xnor2_1 _28082_ (.Y(_07846_),
    .A(_11172_),
    .B(_07845_));
 sg13g2_xnor2_1 _28083_ (.Y(_07847_),
    .A(_07799_),
    .B(_07846_));
 sg13g2_xnor2_1 _28084_ (.Y(_07848_),
    .A(_07796_),
    .B(_07847_));
 sg13g2_nand2b_1 _28085_ (.Y(_07849_),
    .B(_07848_),
    .A_N(_07831_));
 sg13g2_buf_1 _28086_ (.A(_07849_),
    .X(_07850_));
 sg13g2_and2_1 _28087_ (.A(net177),
    .B(_07850_),
    .X(_07851_));
 sg13g2_buf_1 _28088_ (.A(_07851_),
    .X(_07852_));
 sg13g2_and2_1 _28089_ (.A(net159),
    .B(_07852_),
    .X(_07853_));
 sg13g2_buf_1 _28090_ (.A(_07853_),
    .X(_07854_));
 sg13g2_xnor2_1 _28091_ (.Y(_07855_),
    .A(_07775_),
    .B(_07815_));
 sg13g2_xnor2_1 _28092_ (.Y(_07856_),
    .A(_07812_),
    .B(_07855_));
 sg13g2_nand2b_1 _28093_ (.Y(_07857_),
    .B(_07856_),
    .A_N(_07831_));
 sg13g2_buf_1 _28094_ (.A(_07857_),
    .X(_07858_));
 sg13g2_xor2_1 _28095_ (.B(_09646_),
    .A(_13882_),
    .X(_07859_));
 sg13g2_xnor2_1 _28096_ (.Y(_07860_),
    .A(_11179_),
    .B(_07859_));
 sg13g2_xnor2_1 _28097_ (.Y(_07861_),
    .A(_07771_),
    .B(_07860_));
 sg13g2_xnor2_1 _28098_ (.Y(_07862_),
    .A(_07818_),
    .B(_07861_));
 sg13g2_nand2b_1 _28099_ (.Y(_07863_),
    .B(_07862_),
    .A_N(_07831_));
 sg13g2_buf_1 _28100_ (.A(_07863_),
    .X(_07864_));
 sg13g2_and2_1 _28101_ (.A(_07858_),
    .B(net176),
    .X(_07865_));
 sg13g2_buf_1 _28102_ (.A(_07865_),
    .X(_07866_));
 sg13g2_inv_1 _28103_ (.Y(_07867_),
    .A(_13284_));
 sg13g2_a21oi_1 _28104_ (.A1(net755),
    .A2(_07807_),
    .Y(_07868_),
    .B1(_07801_));
 sg13g2_nand2_1 _28105_ (.Y(_07869_),
    .A(net755),
    .B(_07801_));
 sg13g2_o21ai_1 _28106_ (.B1(_07869_),
    .Y(_07870_),
    .A1(_07867_),
    .A2(_07868_));
 sg13g2_nor2_1 _28107_ (.A(net755),
    .B(_07807_),
    .Y(_07871_));
 sg13g2_a21oi_1 _28108_ (.A1(_07867_),
    .A2(_07868_),
    .Y(_07872_),
    .B1(_07871_));
 sg13g2_nor3_1 _28109_ (.A(_13284_),
    .B(net755),
    .C(_07807_),
    .Y(_07873_));
 sg13g2_nand2b_1 _28110_ (.Y(_07874_),
    .B(_07801_),
    .A_N(_07802_));
 sg13g2_nor2b_1 _28111_ (.A(_07873_),
    .B_N(_07874_),
    .Y(_07875_));
 sg13g2_o21ai_1 _28112_ (.B1(_07875_),
    .Y(_07876_),
    .A1(_11172_),
    .A2(_07872_));
 sg13g2_a21oi_1 _28113_ (.A1(_11172_),
    .A2(_07870_),
    .Y(_07877_),
    .B1(_07876_));
 sg13g2_xnor2_1 _28114_ (.Y(_07878_),
    .A(_07778_),
    .B(_07877_));
 sg13g2_or2_1 _28115_ (.X(_07879_),
    .B(_07878_),
    .A(_07831_));
 sg13g2_buf_2 _28116_ (.A(_07879_),
    .X(_07880_));
 sg13g2_buf_1 _28117_ (.A(_07880_),
    .X(_07881_));
 sg13g2_o21ai_1 _28118_ (.B1(_08470_),
    .Y(_07882_),
    .A1(_08655_),
    .A2(_08467_));
 sg13g2_buf_2 _28119_ (.A(_07882_),
    .X(_07883_));
 sg13g2_nand4_1 _28120_ (.B(_07866_),
    .C(_07881_),
    .A(_07854_),
    .Y(_07884_),
    .D(_07883_));
 sg13g2_o21ai_1 _28121_ (.B1(_07884_),
    .Y(_07885_),
    .A1(_07660_),
    .A2(_07763_));
 sg13g2_buf_1 _28122_ (.A(_07858_),
    .X(_07886_));
 sg13g2_inv_1 _28123_ (.Y(_07887_),
    .A(\rbzero.floor_leak[3] ));
 sg13g2_nor2_1 _28124_ (.A(_07831_),
    .B(_07878_),
    .Y(_07888_));
 sg13g2_buf_1 _28125_ (.A(_07888_),
    .X(_07889_));
 sg13g2_buf_1 _28126_ (.A(_07850_),
    .X(_07890_));
 sg13g2_inv_1 _28127_ (.Y(_07891_),
    .A(\rbzero.floor_leak[2] ));
 sg13g2_inv_2 _28128_ (.Y(_07892_),
    .A(_07850_));
 sg13g2_nand2_1 _28129_ (.Y(_07893_),
    .A(\rbzero.floor_leak[0] ),
    .B(_07837_));
 sg13g2_inv_1 _28130_ (.Y(_07894_),
    .A(_07893_));
 sg13g2_nand2_1 _28131_ (.Y(_07895_),
    .A(net177),
    .B(_07894_));
 sg13g2_o21ai_1 _28132_ (.B1(\rbzero.floor_leak[1] ),
    .Y(_07896_),
    .A1(net177),
    .A2(_07894_));
 sg13g2_a22oi_1 _28133_ (.Y(_07897_),
    .B1(_07895_),
    .B2(_07896_),
    .A2(_07892_),
    .A1(_07891_));
 sg13g2_a221oi_1 _28134_ (.B2(\rbzero.floor_leak[3] ),
    .C1(_07897_),
    .B1(_07880_),
    .A1(\rbzero.floor_leak[2] ),
    .Y(_07898_),
    .A2(net156));
 sg13g2_a21oi_1 _28135_ (.A1(_07887_),
    .A2(net175),
    .Y(_07899_),
    .B1(_07898_));
 sg13g2_o21ai_1 _28136_ (.B1(_07899_),
    .Y(_07900_),
    .A1(\rbzero.floor_leak[4] ),
    .A2(net157));
 sg13g2_a22oi_1 _28137_ (.Y(_07901_),
    .B1(net176),
    .B2(\rbzero.floor_leak[5] ),
    .A2(net157),
    .A1(\rbzero.floor_leak[4] ));
 sg13g2_nor2_1 _28138_ (.A(\rbzero.floor_leak[5] ),
    .B(net176),
    .Y(_07902_));
 sg13g2_a21oi_1 _28139_ (.A1(_07900_),
    .A2(_07901_),
    .Y(_07903_),
    .B1(_07902_));
 sg13g2_a21oi_1 _28140_ (.A1(_00046_),
    .A2(_07885_),
    .Y(_07904_),
    .B1(_07903_));
 sg13g2_buf_2 _28141_ (.A(_07904_),
    .X(_07905_));
 sg13g2_buf_1 _28142_ (.A(ui_in[7]),
    .X(_07906_));
 sg13g2_buf_1 _28143_ (.A(_07906_),
    .X(_07907_));
 sg13g2_nor2_1 _28144_ (.A(\rbzero.row_render.texu[1] ),
    .B(_01965_),
    .Y(_07908_));
 sg13g2_buf_1 _28145_ (.A(net177),
    .X(_07909_));
 sg13g2_nor3_1 _28146_ (.A(net155),
    .B(net156),
    .C(_07878_),
    .Y(_07910_));
 sg13g2_a21oi_2 _28147_ (.B1(_07910_),
    .Y(_07911_),
    .A2(_07908_),
    .A1(_00056_));
 sg13g2_nand2_1 _28148_ (.Y(_07912_),
    .A(\rbzero.row_render.texu[1] ),
    .B(_01965_));
 sg13g2_buf_1 _28149_ (.A(_07852_),
    .X(_07913_));
 sg13g2_nand2_1 _28150_ (.Y(_07914_),
    .A(net116),
    .B(_07880_));
 sg13g2_o21ai_1 _28151_ (.B1(_07914_),
    .Y(_07915_),
    .A1(_00056_),
    .A2(_07912_));
 sg13g2_nand2_1 _28152_ (.Y(_07916_),
    .A(_07911_),
    .B(_07915_));
 sg13g2_xor2_1 _28153_ (.B(_07916_),
    .A(net812),
    .X(_07917_));
 sg13g2_and2_1 _28154_ (.A(net812),
    .B(_07854_),
    .X(_07918_));
 sg13g2_nand3_1 _28155_ (.B(\rbzero.row_render.texu[4] ),
    .C(_07908_),
    .A(\rbzero.row_render.texu[3] ),
    .Y(_07919_));
 sg13g2_inv_1 _28156_ (.Y(_07920_),
    .A(_00054_));
 sg13g2_or4_1 _28157_ (.A(_07920_),
    .B(\rbzero.row_render.texu[3] ),
    .C(_07888_),
    .D(_07912_),
    .X(_07921_));
 sg13g2_o21ai_1 _28158_ (.B1(_07921_),
    .Y(_07922_),
    .A1(_07880_),
    .A2(_07919_));
 sg13g2_or2_1 _28159_ (.X(_07923_),
    .B(_07922_),
    .A(_07854_));
 sg13g2_buf_1 _28160_ (.A(_07923_),
    .X(_07924_));
 sg13g2_nor2_1 _28161_ (.A(_01959_),
    .B(_11717_),
    .Y(_07925_));
 sg13g2_a221oi_1 _28162_ (.B2(_07925_),
    .C1(net810),
    .B1(_07924_),
    .A1(_01959_),
    .Y(_07926_),
    .A2(_07918_));
 sg13g2_a21oi_1 _28163_ (.A1(net810),
    .A2(_07917_),
    .Y(_07927_),
    .B1(_07926_));
 sg13g2_buf_1 _28164_ (.A(_00055_),
    .X(_07928_));
 sg13g2_nor2_1 _28165_ (.A(net809),
    .B(_07928_),
    .Y(_07929_));
 sg13g2_a21oi_1 _28166_ (.A1(_01991_),
    .A2(_07927_),
    .Y(_07930_),
    .B1(_07929_));
 sg13g2_buf_1 _28167_ (.A(net159),
    .X(_07931_));
 sg13g2_buf_2 _28168_ (.A(net134),
    .X(_07932_));
 sg13g2_buf_1 _28169_ (.A(_07909_),
    .X(_07933_));
 sg13g2_mux4_1 _28170_ (.S0(net115),
    .A0(_00228_),
    .A1(_00227_),
    .A2(_00226_),
    .A3(_00225_),
    .S1(net133),
    .X(_07934_));
 sg13g2_mux4_1 _28171_ (.S0(net115),
    .A0(_00224_),
    .A1(_00223_),
    .A2(_00222_),
    .A3(_00221_),
    .S1(net133),
    .X(_07935_));
 sg13g2_mux4_1 _28172_ (.S0(net115),
    .A0(_00212_),
    .A1(_00211_),
    .A2(_00210_),
    .A3(_00209_),
    .S1(net133),
    .X(_07936_));
 sg13g2_mux4_1 _28173_ (.S0(_07932_),
    .A0(_00208_),
    .A1(_00207_),
    .A2(_00206_),
    .A3(_00205_),
    .S1(net133),
    .X(_07937_));
 sg13g2_buf_1 _28174_ (.A(net156),
    .X(_07938_));
 sg13g2_buf_1 _28175_ (.A(net157),
    .X(_07939_));
 sg13g2_mux4_1 _28176_ (.S0(net132),
    .A0(_07934_),
    .A1(_07935_),
    .A2(_07936_),
    .A3(_07937_),
    .S1(net131),
    .X(_07940_));
 sg13g2_mux4_1 _28177_ (.S0(net115),
    .A0(_00220_),
    .A1(_00219_),
    .A2(_00218_),
    .A3(_00217_),
    .S1(net133),
    .X(_07941_));
 sg13g2_mux4_1 _28178_ (.S0(_07932_),
    .A0(_00216_),
    .A1(_00215_),
    .A2(_00214_),
    .A3(_00213_),
    .S1(net133),
    .X(_07942_));
 sg13g2_buf_1 _28179_ (.A(_07838_),
    .X(_07943_));
 sg13g2_buf_2 _28180_ (.A(net130),
    .X(_07944_));
 sg13g2_buf_1 _28181_ (.A(net155),
    .X(_07945_));
 sg13g2_mux4_1 _28182_ (.S0(net114),
    .A0(_00204_),
    .A1(_00203_),
    .A2(_00202_),
    .A3(_00201_),
    .S1(net129),
    .X(_07946_));
 sg13g2_mux4_1 _28183_ (.S0(net114),
    .A0(_00200_),
    .A1(_00199_),
    .A2(_00198_),
    .A3(_00197_),
    .S1(net129),
    .X(_07947_));
 sg13g2_mux4_1 _28184_ (.S0(net132),
    .A0(_07941_),
    .A1(_07942_),
    .A2(_07946_),
    .A3(_07947_),
    .S1(net131),
    .X(_07948_));
 sg13g2_mux2_1 _28185_ (.A0(_07940_),
    .A1(_07948_),
    .S(_07881_),
    .X(_07949_));
 sg13g2_buf_1 _28186_ (.A(net176),
    .X(_07950_));
 sg13g2_nor2b_1 _28187_ (.A(_07949_),
    .B_N(net154),
    .Y(_07951_));
 sg13g2_mux4_1 _28188_ (.S0(net115),
    .A0(_00256_),
    .A1(_00255_),
    .A2(_00254_),
    .A3(_00253_),
    .S1(net133),
    .X(_07952_));
 sg13g2_mux4_1 _28189_ (.S0(net115),
    .A0(_00248_),
    .A1(_00247_),
    .A2(_00246_),
    .A3(_00245_),
    .S1(_07933_),
    .X(_07953_));
 sg13g2_mux4_1 _28190_ (.S0(_07944_),
    .A0(_00260_),
    .A1(_00259_),
    .A2(_00258_),
    .A3(_00257_),
    .S1(_07945_),
    .X(_07954_));
 sg13g2_mux4_1 _28191_ (.S0(_07944_),
    .A0(_00252_),
    .A1(_00251_),
    .A2(_00250_),
    .A3(_00249_),
    .S1(_07945_),
    .X(_07955_));
 sg13g2_buf_2 _28192_ (.A(_07880_),
    .X(_07956_));
 sg13g2_buf_1 _28193_ (.A(_07892_),
    .X(_07957_));
 sg13g2_mux4_1 _28194_ (.S0(_07956_),
    .A0(_07952_),
    .A1(_07953_),
    .A2(_07954_),
    .A3(_07955_),
    .S1(_07957_),
    .X(_07958_));
 sg13g2_nor2b_1 _28195_ (.A(_07939_),
    .B_N(_07958_),
    .Y(_07959_));
 sg13g2_buf_1 _28196_ (.A(_07837_),
    .X(_07960_));
 sg13g2_buf_1 _28197_ (.A(net152),
    .X(_07961_));
 sg13g2_buf_2 _28198_ (.A(net127),
    .X(_07962_));
 sg13g2_buf_1 _28199_ (.A(net177),
    .X(_07963_));
 sg13g2_buf_1 _28200_ (.A(net151),
    .X(_07964_));
 sg13g2_mux4_1 _28201_ (.S0(net113),
    .A0(_00244_),
    .A1(_00243_),
    .A2(_00242_),
    .A3(_00241_),
    .S1(net126),
    .X(_07965_));
 sg13g2_mux2_1 _28202_ (.A0(_00238_),
    .A1(_00237_),
    .S(net134),
    .X(_07966_));
 sg13g2_nor2_1 _28203_ (.A(net177),
    .B(_07892_),
    .Y(_07967_));
 sg13g2_buf_1 _28204_ (.A(_07967_),
    .X(_07968_));
 sg13g2_buf_2 _28205_ (.A(net152),
    .X(_07969_));
 sg13g2_mux2_1 _28206_ (.A0(_00240_),
    .A1(_00239_),
    .S(net125),
    .X(_07970_));
 sg13g2_a221oi_1 _28207_ (.B2(_07970_),
    .C1(net153),
    .B1(net112),
    .A1(_07913_),
    .Y(_07971_),
    .A2(_07966_));
 sg13g2_nand2b_1 _28208_ (.Y(_07972_),
    .B(_07971_),
    .A_N(_07965_));
 sg13g2_mux4_1 _28209_ (.S0(net113),
    .A0(_00236_),
    .A1(_00235_),
    .A2(_00234_),
    .A3(_00233_),
    .S1(net126),
    .X(_07973_));
 sg13g2_mux2_1 _28210_ (.A0(_00232_),
    .A1(_00231_),
    .S(_07931_),
    .X(_07974_));
 sg13g2_mux2_1 _28211_ (.A0(_00230_),
    .A1(_00229_),
    .S(_07961_),
    .X(_07975_));
 sg13g2_a221oi_1 _28212_ (.B2(_07913_),
    .C1(_07889_),
    .B1(_07975_),
    .A1(net112),
    .Y(_07976_),
    .A2(_07974_));
 sg13g2_nand2b_1 _28213_ (.Y(_07977_),
    .B(_07976_),
    .A_N(_07973_));
 sg13g2_o21ai_1 _28214_ (.B1(_07938_),
    .Y(_07978_),
    .A1(_07971_),
    .A2(_07976_));
 sg13g2_and4_1 _28215_ (.A(_07939_),
    .B(_07972_),
    .C(_07977_),
    .D(_07978_),
    .X(_07979_));
 sg13g2_nor3_1 _28216_ (.A(_07950_),
    .B(_07959_),
    .C(_07979_),
    .Y(_07980_));
 sg13g2_nor3_1 _28217_ (.A(net801),
    .B(_07951_),
    .C(_07980_),
    .Y(_07981_));
 sg13g2_a21oi_1 _28218_ (.A1(net801),
    .A2(_07930_),
    .Y(_07982_),
    .B1(_07981_));
 sg13g2_mux2_1 _28219_ (.A0(_00195_),
    .A1(_00196_),
    .S(_07883_),
    .X(_07983_));
 sg13g2_nor2_1 _28220_ (.A(_07905_),
    .B(_07983_),
    .Y(_07984_));
 sg13g2_a21oi_1 _28221_ (.A1(_07905_),
    .A2(_07982_),
    .Y(_07985_),
    .B1(_07984_));
 sg13g2_nand2_1 _28222_ (.Y(_07986_),
    .A(_09404_),
    .B(_09398_));
 sg13g2_inv_1 _28223_ (.Y(_07987_),
    .A(_11200_));
 sg13g2_nor2_1 _28224_ (.A(_09402_),
    .B(_07987_),
    .Y(_07988_));
 sg13g2_a21oi_1 _28225_ (.A1(_09403_),
    .A2(_09726_),
    .Y(_07989_),
    .B1(_07988_));
 sg13g2_o21ai_1 _28226_ (.B1(_08461_),
    .Y(_07990_),
    .A1(_09405_),
    .A2(_11184_));
 sg13g2_a21oi_1 _28227_ (.A1(_07986_),
    .A2(_07989_),
    .Y(_07991_),
    .B1(_07990_));
 sg13g2_or4_1 _28228_ (.A(_09405_),
    .B(net753),
    .C(_11184_),
    .D(_07986_),
    .X(_07992_));
 sg13g2_a21oi_1 _28229_ (.A1(_11200_),
    .A2(_07992_),
    .Y(_07993_),
    .B1(_09414_));
 sg13g2_nand2_1 _28230_ (.Y(_07994_),
    .A(_08655_),
    .B(_08649_));
 sg13g2_a21oi_1 _28231_ (.A1(_08469_),
    .A2(_07994_),
    .Y(_07995_),
    .B1(_09399_));
 sg13g2_nand2b_1 _28232_ (.Y(_07996_),
    .B(_07995_),
    .A_N(_07993_));
 sg13g2_inv_1 _28233_ (.Y(_07997_),
    .A(_07996_));
 sg13g2_o21ai_1 _28234_ (.B1(_07997_),
    .Y(_07998_),
    .A1(_07652_),
    .A2(_07991_));
 sg13g2_a21oi_1 _28235_ (.A1(_07652_),
    .A2(_07985_),
    .Y(\rbzero.rgb[0] ),
    .B1(_07998_));
 sg13g2_mux2_1 _28236_ (.A0(\rbzero.color_floor[1] ),
    .A1(\rbzero.color_sky[1] ),
    .S(_07883_),
    .X(_07999_));
 sg13g2_xnor2_1 _28237_ (.Y(_08000_),
    .A(_07920_),
    .B(_07886_));
 sg13g2_nand4_1 _28238_ (.B(_07928_),
    .C(_07911_),
    .A(_01991_),
    .Y(_08001_),
    .D(_07915_));
 sg13g2_o21ai_1 _28239_ (.B1(_08001_),
    .Y(_08002_),
    .A1(net809),
    .A2(_08000_));
 sg13g2_nor2b_1 _28240_ (.A(_01959_),
    .B_N(net812),
    .Y(_08003_));
 sg13g2_nand2_1 _28241_ (.Y(_08004_),
    .A(_07924_),
    .B(_08003_));
 sg13g2_nor2b_1 _28242_ (.A(net810),
    .B_N(\rbzero.row_render.wall[1] ),
    .Y(_08005_));
 sg13g2_buf_1 _28243_ (.A(_08005_),
    .X(_08006_));
 sg13g2_a22oi_1 _28244_ (.Y(_08007_),
    .B1(_08004_),
    .B2(_08006_),
    .A2(_08002_),
    .A1(net810));
 sg13g2_inv_1 _28245_ (.Y(_08008_),
    .A(_08007_));
 sg13g2_mux2_1 _28246_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_07838_),
    .X(_08009_));
 sg13g2_mux2_1 _28247_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(net159),
    .X(_08010_));
 sg13g2_a221oi_1 _28248_ (.B2(net112),
    .C1(_07889_),
    .B1(_08010_),
    .A1(_07852_),
    .Y(_08011_),
    .A2(_08009_));
 sg13g2_mux2_1 _28249_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(net159),
    .X(_08012_));
 sg13g2_mux2_1 _28250_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(net159),
    .X(_08013_));
 sg13g2_a221oi_1 _28251_ (.B2(net116),
    .C1(_07880_),
    .B1(_08013_),
    .A1(_07968_),
    .Y(_08014_),
    .A2(_08012_));
 sg13g2_o21ai_1 _28252_ (.B1(_07938_),
    .Y(_08015_),
    .A1(_08011_),
    .A2(_08014_));
 sg13g2_mux4_1 _28253_ (.S0(_07969_),
    .A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[54] ),
    .A2(\rbzero.tex_r1[53] ),
    .A3(\rbzero.tex_r1[52] ),
    .S1(_07963_),
    .X(_08016_));
 sg13g2_nand2b_1 _28254_ (.Y(_08017_),
    .B(_08011_),
    .A_N(_08016_));
 sg13g2_mux4_1 _28255_ (.S0(net125),
    .A0(\rbzero.tex_r1[63] ),
    .A1(\rbzero.tex_r1[62] ),
    .A2(\rbzero.tex_r1[61] ),
    .A3(\rbzero.tex_r1[60] ),
    .S1(net151),
    .X(_08018_));
 sg13g2_nand2b_1 _28256_ (.Y(_08019_),
    .B(_08014_),
    .A_N(_08018_));
 sg13g2_nand3_1 _28257_ (.B(_08017_),
    .C(_08019_),
    .A(_08015_),
    .Y(_08020_));
 sg13g2_nor2_1 _28258_ (.A(_07950_),
    .B(_08020_),
    .Y(_08021_));
 sg13g2_mux4_1 _28259_ (.S0(_07931_),
    .A0(\rbzero.tex_r1[39] ),
    .A1(\rbzero.tex_r1[38] ),
    .A2(\rbzero.tex_r1[37] ),
    .A3(\rbzero.tex_r1[36] ),
    .S1(net155),
    .X(_08022_));
 sg13g2_mux2_1 _28260_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_07837_),
    .X(_08023_));
 sg13g2_mux2_1 _28261_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(net159),
    .X(_08024_));
 sg13g2_a221oi_1 _28262_ (.B2(_07852_),
    .C1(_07888_),
    .B1(_08024_),
    .A1(_07967_),
    .Y(_08025_),
    .A2(_08023_));
 sg13g2_nand2b_1 _28263_ (.Y(_08026_),
    .B(_08025_),
    .A_N(_08022_));
 sg13g2_mux4_1 _28264_ (.S0(_07943_),
    .A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[46] ),
    .A2(\rbzero.tex_r1[45] ),
    .A3(\rbzero.tex_r1[44] ),
    .S1(_07909_),
    .X(_08027_));
 sg13g2_mux2_1 _28265_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[40] ),
    .S(net159),
    .X(_08028_));
 sg13g2_mux2_1 _28266_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(net159),
    .X(_08029_));
 sg13g2_a221oi_1 _28267_ (.B2(_07968_),
    .C1(_07880_),
    .B1(_08029_),
    .A1(_07852_),
    .Y(_08030_),
    .A2(_08028_));
 sg13g2_nand2b_1 _28268_ (.Y(_08031_),
    .B(_08030_),
    .A_N(_08027_));
 sg13g2_o21ai_1 _28269_ (.B1(_07890_),
    .Y(_08032_),
    .A1(_08025_),
    .A2(_08030_));
 sg13g2_nand3_1 _28270_ (.B(_08031_),
    .C(_08032_),
    .A(_08026_),
    .Y(_08033_));
 sg13g2_mux4_1 _28271_ (.S0(net152),
    .A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[10] ),
    .A2(\rbzero.tex_r1[9] ),
    .A3(\rbzero.tex_r1[8] ),
    .S1(net177),
    .X(_08034_));
 sg13g2_mux4_1 _28272_ (.S0(net152),
    .A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[2] ),
    .A2(\rbzero.tex_r1[1] ),
    .A3(\rbzero.tex_r1[0] ),
    .S1(net155),
    .X(_08035_));
 sg13g2_mux4_1 _28273_ (.S0(net152),
    .A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[14] ),
    .A2(\rbzero.tex_r1[13] ),
    .A3(\rbzero.tex_r1[12] ),
    .S1(net177),
    .X(_08036_));
 sg13g2_mux4_1 _28274_ (.S0(_07960_),
    .A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[6] ),
    .A2(\rbzero.tex_r1[5] ),
    .A3(\rbzero.tex_r1[4] ),
    .S1(_07844_),
    .X(_08037_));
 sg13g2_mux4_1 _28275_ (.S0(_07880_),
    .A0(_08034_),
    .A1(_08035_),
    .A2(_08036_),
    .A3(_08037_),
    .S1(_07892_),
    .X(_08038_));
 sg13g2_nand2_1 _28276_ (.Y(_08039_),
    .A(net176),
    .B(_08038_));
 sg13g2_o21ai_1 _28277_ (.B1(_08039_),
    .Y(_08040_),
    .A1(_07864_),
    .A2(_08033_));
 sg13g2_mux2_1 _28278_ (.A0(_08021_),
    .A1(_08040_),
    .S(net131),
    .X(_08041_));
 sg13g2_buf_1 _28279_ (.A(net112),
    .X(_08042_));
 sg13g2_mux2_1 _28280_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(net125),
    .X(_08043_));
 sg13g2_mux2_1 _28281_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(net127),
    .X(_08044_));
 sg13g2_buf_1 _28282_ (.A(net116),
    .X(_08045_));
 sg13g2_a22oi_1 _28283_ (.Y(_08046_),
    .B1(_08044_),
    .B2(net98),
    .A2(_08043_),
    .A1(net99));
 sg13g2_nand2_1 _28284_ (.Y(_08047_),
    .A(_07956_),
    .B(_08046_));
 sg13g2_mux2_1 _28285_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(net125),
    .X(_08048_));
 sg13g2_mux2_1 _28286_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_07961_),
    .X(_08049_));
 sg13g2_a22oi_1 _28287_ (.Y(_08050_),
    .B1(_08049_),
    .B2(net99),
    .A2(_08048_),
    .A1(net116));
 sg13g2_nand2_1 _28288_ (.Y(_08051_),
    .A(net175),
    .B(_08050_));
 sg13g2_a21oi_1 _28289_ (.A1(_08047_),
    .A2(_08051_),
    .Y(_08052_),
    .B1(net128));
 sg13g2_nand2b_1 _28290_ (.Y(_08053_),
    .B(net176),
    .A_N(net131));
 sg13g2_buf_2 _28291_ (.A(net114),
    .X(_08054_));
 sg13g2_buf_1 _28292_ (.A(net129),
    .X(_08055_));
 sg13g2_mux4_1 _28293_ (.S0(net97),
    .A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[22] ),
    .A2(\rbzero.tex_r1[21] ),
    .A3(\rbzero.tex_r1[20] ),
    .S1(net111),
    .X(_08056_));
 sg13g2_nor2_1 _28294_ (.A(_08047_),
    .B(_08056_),
    .Y(_08057_));
 sg13g2_mux4_1 _28295_ (.S0(net97),
    .A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[30] ),
    .A2(\rbzero.tex_r1[29] ),
    .A3(\rbzero.tex_r1[28] ),
    .S1(net111),
    .X(_08058_));
 sg13g2_nor2_1 _28296_ (.A(_08051_),
    .B(_08058_),
    .Y(_08059_));
 sg13g2_nor4_1 _28297_ (.A(_08052_),
    .B(_08053_),
    .C(_08057_),
    .D(_08059_),
    .Y(_08060_));
 sg13g2_nor3_1 _28298_ (.A(_07906_),
    .B(_08041_),
    .C(_08060_),
    .Y(_08061_));
 sg13g2_a21oi_1 _28299_ (.A1(net801),
    .A2(_08008_),
    .Y(_08062_),
    .B1(_08061_));
 sg13g2_mux2_1 _28300_ (.A0(_07999_),
    .A1(_08062_),
    .S(_07905_),
    .X(_08063_));
 sg13g2_inv_1 _28301_ (.Y(_08064_),
    .A(_08063_));
 sg13g2_xnor2_1 _28302_ (.Y(_08065_),
    .A(net831),
    .B(_07642_));
 sg13g2_and2_1 _28303_ (.A(_07632_),
    .B(_08065_),
    .X(_08066_));
 sg13g2_buf_1 _28304_ (.A(_08066_),
    .X(_08067_));
 sg13g2_nor2b_1 _28305_ (.A(_07636_),
    .B_N(net493),
    .Y(_08068_));
 sg13g2_nand2_1 _28306_ (.Y(_08069_),
    .A(_08067_),
    .B(_08068_));
 sg13g2_inv_1 _28307_ (.Y(_08070_),
    .A(_07647_));
 sg13g2_nor3_1 _28308_ (.A(net831),
    .B(_07643_),
    .C(_07642_),
    .Y(_08071_));
 sg13g2_a21oi_1 _28309_ (.A1(_07643_),
    .A2(_08070_),
    .Y(_08072_),
    .B1(_08071_));
 sg13g2_a21oi_1 _28310_ (.A1(_09706_),
    .A2(_07636_),
    .Y(_08073_),
    .B1(net493));
 sg13g2_nor2_1 _28311_ (.A(_07632_),
    .B(_08073_),
    .Y(_08074_));
 sg13g2_nor2_2 _28312_ (.A(_08072_),
    .B(_08074_),
    .Y(_08075_));
 sg13g2_nand3_1 _28313_ (.B(net543),
    .C(_08075_),
    .A(_09705_),
    .Y(_08076_));
 sg13g2_buf_1 _28314_ (.A(_08076_),
    .X(_08077_));
 sg13g2_nor2_1 _28315_ (.A(_08069_),
    .B(_08077_),
    .Y(_08078_));
 sg13g2_buf_1 _28316_ (.A(_08078_),
    .X(_08079_));
 sg13g2_nand2_1 _28317_ (.Y(_08080_),
    .A(_08485_),
    .B(_08079_));
 sg13g2_nand2b_1 _28318_ (.Y(_08081_),
    .B(_08075_),
    .A_N(_09705_));
 sg13g2_or2_1 _28319_ (.X(_08082_),
    .B(_08081_),
    .A(net543));
 sg13g2_xor2_1 _28320_ (.B(net493),
    .A(net543),
    .X(_08083_));
 sg13g2_nand3_1 _28321_ (.B(_08067_),
    .C(_08083_),
    .A(_07636_),
    .Y(_08084_));
 sg13g2_buf_1 _28322_ (.A(_08084_),
    .X(_08085_));
 sg13g2_nor2_1 _28323_ (.A(_08082_),
    .B(_08085_),
    .Y(_08086_));
 sg13g2_buf_2 _28324_ (.A(_08086_),
    .X(_08087_));
 sg13g2_nand3b_1 _28325_ (.B(net543),
    .C(_08075_),
    .Y(_08088_),
    .A_N(_09705_));
 sg13g2_buf_1 _28326_ (.A(_08088_),
    .X(_08089_));
 sg13g2_or2_1 _28327_ (.X(_08090_),
    .B(net493),
    .A(_07632_));
 sg13g2_nand3_1 _28328_ (.B(_07632_),
    .C(net493),
    .A(net543),
    .Y(_08091_));
 sg13g2_o21ai_1 _28329_ (.B1(_08091_),
    .Y(_08092_),
    .A1(net543),
    .A2(_08090_));
 sg13g2_nand3_1 _28330_ (.B(_08065_),
    .C(_08092_),
    .A(_07636_),
    .Y(_08093_));
 sg13g2_nor2_1 _28331_ (.A(_08089_),
    .B(_08093_),
    .Y(_08094_));
 sg13g2_buf_1 _28332_ (.A(_08094_),
    .X(_08095_));
 sg13g2_a22oi_1 _28333_ (.Y(_08096_),
    .B1(_08095_),
    .B2(_09935_),
    .A2(_08087_),
    .A1(_09934_));
 sg13g2_nand2_1 _28334_ (.Y(_08097_),
    .A(_09705_),
    .B(_08075_));
 sg13g2_or2_1 _28335_ (.X(_08098_),
    .B(_08097_),
    .A(net543));
 sg13g2_buf_1 _28336_ (.A(_08098_),
    .X(_08099_));
 sg13g2_nand3b_1 _28337_ (.B(_07640_),
    .C(_08065_),
    .Y(_08100_),
    .A_N(_07632_));
 sg13g2_buf_1 _28338_ (.A(_08100_),
    .X(_08101_));
 sg13g2_nor2_1 _28339_ (.A(_08099_),
    .B(_08101_),
    .Y(_08102_));
 sg13g2_buf_2 _28340_ (.A(_08102_),
    .X(_08103_));
 sg13g2_or2_1 _28341_ (.X(_08104_),
    .B(_08101_),
    .A(_08089_));
 sg13g2_buf_2 _28342_ (.A(_08104_),
    .X(_08105_));
 sg13g2_nor2_1 _28343_ (.A(_09926_),
    .B(_08105_),
    .Y(_08106_));
 sg13g2_a21oi_1 _28344_ (.A1(_09936_),
    .A2(_08103_),
    .Y(_08107_),
    .B1(_08106_));
 sg13g2_nor2_1 _28345_ (.A(_08085_),
    .B(_08099_),
    .Y(_08108_));
 sg13g2_buf_2 _28346_ (.A(_08108_),
    .X(_08109_));
 sg13g2_nor2_1 _28347_ (.A(_08069_),
    .B(_08089_),
    .Y(_08110_));
 sg13g2_buf_1 _28348_ (.A(_08110_),
    .X(_08111_));
 sg13g2_a22oi_1 _28349_ (.Y(_08112_),
    .B1(_08111_),
    .B2(_09931_),
    .A2(_08109_),
    .A1(_09932_));
 sg13g2_nand4_1 _28350_ (.B(_08096_),
    .C(_08107_),
    .A(_08080_),
    .Y(_08113_),
    .D(_08112_));
 sg13g2_nor2_1 _28351_ (.A(_08082_),
    .B(_08101_),
    .Y(_08114_));
 sg13g2_buf_2 _28352_ (.A(_08114_),
    .X(_08115_));
 sg13g2_nor2_1 _28353_ (.A(_08077_),
    .B(_08093_),
    .Y(_08116_));
 sg13g2_buf_2 _28354_ (.A(_08116_),
    .X(_08117_));
 sg13g2_a22oi_1 _28355_ (.Y(_08118_),
    .B1(_08117_),
    .B2(_09933_),
    .A2(_08115_),
    .A1(_09938_));
 sg13g2_nor2_1 _28356_ (.A(_08077_),
    .B(_08101_),
    .Y(_08119_));
 sg13g2_buf_1 _28357_ (.A(_08119_),
    .X(_08120_));
 sg13g2_nor2_1 _28358_ (.A(_08077_),
    .B(_08085_),
    .Y(_08121_));
 sg13g2_a22oi_1 _28359_ (.Y(_08122_),
    .B1(_08121_),
    .B2(_08492_),
    .A2(_08120_),
    .A1(_09937_));
 sg13g2_nand2_1 _28360_ (.Y(_08123_),
    .A(_08118_),
    .B(_08122_));
 sg13g2_nor2_1 _28361_ (.A(net543),
    .B(_08081_),
    .Y(_08124_));
 sg13g2_inv_1 _28362_ (.Y(_08125_),
    .A(_08099_));
 sg13g2_a22oi_1 _28363_ (.Y(_08126_),
    .B1(_08125_),
    .B2(_08518_),
    .A2(_08124_),
    .A1(_08507_));
 sg13g2_nor2_1 _28364_ (.A(_08085_),
    .B(_08089_),
    .Y(_08127_));
 sg13g2_nor2b_1 _28365_ (.A(net493),
    .B_N(_08498_),
    .Y(_08128_));
 sg13g2_nand4_1 _28366_ (.B(_08067_),
    .C(_08124_),
    .A(_07636_),
    .Y(_08129_),
    .D(_08128_));
 sg13g2_nand3_1 _28367_ (.B(_07988_),
    .C(_08129_),
    .A(_09403_),
    .Y(_08130_));
 sg13g2_a21oi_1 _28368_ (.A1(_08489_),
    .A2(_08127_),
    .Y(_08131_),
    .B1(_08130_));
 sg13g2_o21ai_1 _28369_ (.B1(_08131_),
    .Y(_08132_),
    .A1(_08069_),
    .A2(_08126_));
 sg13g2_nor3_1 _28370_ (.A(_08113_),
    .B(_08123_),
    .C(_08132_),
    .Y(_08133_));
 sg13g2_inv_1 _28371_ (.Y(_08134_),
    .A(_09739_));
 sg13g2_a22oi_1 _28372_ (.Y(_08135_),
    .B1(_08115_),
    .B2(_09754_),
    .A2(_08103_),
    .A1(_09757_));
 sg13g2_o21ai_1 _28373_ (.B1(_08135_),
    .Y(_08136_),
    .A1(_08134_),
    .A2(_08105_));
 sg13g2_o21ai_1 _28374_ (.B1(net493),
    .Y(_08137_),
    .A1(_09707_),
    .A2(_07636_));
 sg13g2_and3_1 _28375_ (.X(_08138_),
    .A(_08067_),
    .B(_08075_),
    .C(_08137_));
 sg13g2_buf_1 _28376_ (.A(_08138_),
    .X(_08139_));
 sg13g2_nand3_1 _28377_ (.B(net753),
    .C(_11200_),
    .A(_09403_),
    .Y(_08140_));
 sg13g2_a221oi_1 _28378_ (.B2(_09747_),
    .C1(_08140_),
    .B1(_08139_),
    .A1(_09777_),
    .Y(_08141_),
    .A2(_08111_));
 sg13g2_a22oi_1 _28379_ (.Y(_08142_),
    .B1(_08120_),
    .B2(_09751_),
    .A2(_08117_),
    .A1(_09767_));
 sg13g2_a22oi_1 _28380_ (.Y(_08143_),
    .B1(_08087_),
    .B2(_09770_),
    .A2(_08079_),
    .A1(_09781_));
 sg13g2_a22oi_1 _28381_ (.Y(_08144_),
    .B1(_08109_),
    .B2(_09774_),
    .A2(_08095_),
    .A1(_09762_));
 sg13g2_nand4_1 _28382_ (.B(_08142_),
    .C(_08143_),
    .A(_08141_),
    .Y(_08145_),
    .D(_08144_));
 sg13g2_nor2_1 _28383_ (.A(_08136_),
    .B(_08145_),
    .Y(_08146_));
 sg13g2_nor2b_1 _28384_ (.A(_09403_),
    .B_N(net753),
    .Y(_08147_));
 sg13g2_nor4_1 _28385_ (.A(_07987_),
    .B(_08133_),
    .C(_08146_),
    .D(_08147_),
    .Y(_08148_));
 sg13g2_and2_1 _28386_ (.A(net770),
    .B(_08095_),
    .X(_08149_));
 sg13g2_a221oi_1 _28387_ (.B2(net767),
    .C1(_08149_),
    .B1(_08117_),
    .A1(net763),
    .Y(_08150_),
    .A2(_08087_));
 sg13g2_nand2_1 _28388_ (.Y(_08151_),
    .A(net768),
    .B(_08120_));
 sg13g2_o21ai_1 _28389_ (.B1(_08151_),
    .Y(_08152_),
    .A1(_09146_),
    .A2(_08105_));
 sg13g2_a221oi_1 _28390_ (.B2(net820),
    .C1(_08152_),
    .B1(_08139_),
    .A1(net765),
    .Y(_08153_),
    .A2(_08103_));
 sg13g2_a22oi_1 _28391_ (.Y(_08154_),
    .B1(_08109_),
    .B2(net822),
    .A2(_08079_),
    .A1(net821));
 sg13g2_a22oi_1 _28392_ (.Y(_08155_),
    .B1(_08115_),
    .B2(net766),
    .A2(_08111_),
    .A1(net762));
 sg13g2_nand4_1 _28393_ (.B(_08153_),
    .C(_08154_),
    .A(_08150_),
    .Y(_08156_),
    .D(_08155_));
 sg13g2_nand4_1 _28394_ (.B(net753),
    .C(_07987_),
    .A(_09403_),
    .Y(_08157_),
    .D(_08156_));
 sg13g2_and2_1 _28395_ (.A(_09790_),
    .B(_08120_),
    .X(_08158_));
 sg13g2_a221oi_1 _28396_ (.B2(_09792_),
    .C1(_08158_),
    .B1(_08115_),
    .A1(_09805_),
    .Y(_08159_),
    .A2(_08087_));
 sg13g2_a22oi_1 _28397_ (.Y(_08160_),
    .B1(_08117_),
    .B2(_09802_),
    .A2(_08111_),
    .A1(_09811_));
 sg13g2_a22oi_1 _28398_ (.Y(_08161_),
    .B1(_08109_),
    .B2(_09807_),
    .A2(_08103_),
    .A1(_09795_));
 sg13g2_inv_1 _28399_ (.Y(_08162_),
    .A(_09783_));
 sg13g2_nor2_1 _28400_ (.A(net753),
    .B(_07986_),
    .Y(_08163_));
 sg13g2_o21ai_1 _28401_ (.B1(_08163_),
    .Y(_08164_),
    .A1(_08162_),
    .A2(_08105_));
 sg13g2_a221oi_1 _28402_ (.B2(_09798_),
    .C1(_08164_),
    .B1(_08095_),
    .A1(_09813_),
    .Y(_08165_),
    .A2(_08079_));
 sg13g2_nand4_1 _28403_ (.B(_08160_),
    .C(_08161_),
    .A(_08159_),
    .Y(_08166_),
    .D(_08165_));
 sg13g2_a22oi_1 _28404_ (.Y(_08167_),
    .B1(_08117_),
    .B2(net779),
    .A2(_08079_),
    .A1(net771));
 sg13g2_nand2_1 _28405_ (.Y(_08168_),
    .A(net775),
    .B(_08087_));
 sg13g2_nand2_1 _28406_ (.Y(_08169_),
    .A(_08768_),
    .B(_08103_));
 sg13g2_nand4_1 _28407_ (.B(_09398_),
    .C(_09726_),
    .A(_09404_),
    .Y(_08170_),
    .D(_08169_));
 sg13g2_a221oi_1 _28408_ (.B2(net781),
    .C1(_08170_),
    .B1(_08120_),
    .A1(net773),
    .Y(_08171_),
    .A2(_08109_));
 sg13g2_nand2_1 _28409_ (.Y(_08172_),
    .A(net780),
    .B(_08115_));
 sg13g2_o21ai_1 _28410_ (.B1(_08172_),
    .Y(_08173_),
    .A1(_08817_),
    .A2(_08105_));
 sg13g2_a221oi_1 _28411_ (.B2(net772),
    .C1(_08173_),
    .B1(_08111_),
    .A1(net722),
    .Y(_08174_),
    .A2(_08095_));
 sg13g2_nand4_1 _28412_ (.B(_08168_),
    .C(_08171_),
    .A(_08167_),
    .Y(_08175_),
    .D(_08174_));
 sg13g2_nand2_1 _28413_ (.Y(_08176_),
    .A(_08166_),
    .B(_08175_));
 sg13g2_o21ai_1 _28414_ (.B1(_08139_),
    .Y(_08177_),
    .A1(net825),
    .A2(_08175_));
 sg13g2_nor2_1 _28415_ (.A(_08133_),
    .B(_08146_),
    .Y(_08178_));
 sg13g2_o21ai_1 _28416_ (.B1(_08178_),
    .Y(_08179_),
    .A1(_09786_),
    .A2(_08166_));
 sg13g2_a221oi_1 _28417_ (.B2(_08177_),
    .C1(_08179_),
    .B1(_08176_),
    .A1(_07986_),
    .Y(_08180_),
    .A2(_08157_));
 sg13g2_a22oi_1 _28418_ (.Y(_08181_),
    .B1(_08103_),
    .B2(_09839_),
    .A2(_08079_),
    .A1(_08494_));
 sg13g2_nor2_1 _28419_ (.A(_08069_),
    .B(_08099_),
    .Y(_08182_));
 sg13g2_nor2b_1 _28420_ (.A(_07639_),
    .B_N(_08522_),
    .Y(_08183_));
 sg13g2_a22oi_1 _28421_ (.Y(_08184_),
    .B1(_08183_),
    .B2(_07636_),
    .A2(_08068_),
    .A1(_08511_));
 sg13g2_nor2b_1 _28422_ (.A(_08184_),
    .B_N(_08067_),
    .Y(_08185_));
 sg13g2_a22oi_1 _28423_ (.Y(_08186_),
    .B1(_08185_),
    .B2(_08124_),
    .A2(_08182_),
    .A1(_08501_));
 sg13g2_nand4_1 _28424_ (.B(_07988_),
    .C(_08181_),
    .A(_09404_),
    .Y(_08187_),
    .D(_08186_));
 sg13g2_a221oi_1 _28425_ (.B2(_09836_),
    .C1(_08187_),
    .B1(_08117_),
    .A1(_09841_),
    .Y(_08188_),
    .A2(_08115_));
 sg13g2_a22oi_1 _28426_ (.Y(_08189_),
    .B1(_08109_),
    .B2(_09835_),
    .A2(_08095_),
    .A1(_09838_));
 sg13g2_a22oi_1 _28427_ (.Y(_08190_),
    .B1(_08127_),
    .B2(_08483_),
    .A2(_08120_),
    .A1(_09840_));
 sg13g2_nor2_1 _28428_ (.A(_09820_),
    .B(_08105_),
    .Y(_08191_));
 sg13g2_a21oi_1 _28429_ (.A1(_09834_),
    .A2(_08111_),
    .Y(_08192_),
    .B1(_08191_));
 sg13g2_a22oi_1 _28430_ (.Y(_08193_),
    .B1(_08121_),
    .B2(_08514_),
    .A2(_08087_),
    .A1(_09837_));
 sg13g2_and4_1 _28431_ (.A(_08189_),
    .B(_08190_),
    .C(_08192_),
    .D(_08193_),
    .X(_08194_));
 sg13g2_a21oi_1 _28432_ (.A1(_08188_),
    .A2(_08194_),
    .Y(_08195_),
    .B1(_07990_));
 sg13g2_o21ai_1 _28433_ (.B1(_08195_),
    .Y(_08196_),
    .A1(_08148_),
    .A2(_08180_));
 sg13g2_inv_1 _28434_ (.Y(_08197_),
    .A(_08068_));
 sg13g2_xor2_1 _28435_ (.B(_08454_),
    .A(_08455_),
    .X(_08198_));
 sg13g2_nor4_1 _28436_ (.A(_08461_),
    .B(_08197_),
    .C(_08072_),
    .D(_08198_),
    .Y(_08199_));
 sg13g2_a21oi_1 _28437_ (.A1(_07633_),
    .A2(_08199_),
    .Y(_08200_),
    .B1(_07652_));
 sg13g2_a21oi_1 _28438_ (.A1(_08196_),
    .A2(_08200_),
    .Y(_08201_),
    .B1(_07996_));
 sg13g2_inv_1 _28439_ (.Y(_08202_),
    .A(_08201_));
 sg13g2_a21oi_1 _28440_ (.A1(_07652_),
    .A2(_08064_),
    .Y(\rbzero.rgb[1] ),
    .B1(_08202_));
 sg13g2_mux2_1 _28441_ (.A0(_00261_),
    .A1(_00262_),
    .S(_07883_),
    .X(_08203_));
 sg13g2_nand2b_1 _28442_ (.Y(_08204_),
    .B(net131),
    .A_N(net176));
 sg13g2_mux4_1 _28443_ (.S0(net113),
    .A0(_00306_),
    .A1(_00305_),
    .A2(_00304_),
    .A3(_00303_),
    .S1(net126),
    .X(_08205_));
 sg13g2_mux4_1 _28444_ (.S0(net113),
    .A0(_00298_),
    .A1(_00297_),
    .A2(_00296_),
    .A3(_00295_),
    .S1(net126),
    .X(_08206_));
 sg13g2_mux4_1 _28445_ (.S0(net113),
    .A0(_00310_),
    .A1(_00309_),
    .A2(_00308_),
    .A3(_00307_),
    .S1(net126),
    .X(_08207_));
 sg13g2_mux4_1 _28446_ (.S0(net113),
    .A0(_00302_),
    .A1(_00301_),
    .A2(_00300_),
    .A3(_00299_),
    .S1(net126),
    .X(_08208_));
 sg13g2_mux4_1 _28447_ (.S0(net158),
    .A0(_08205_),
    .A1(_08206_),
    .A2(_08207_),
    .A3(_08208_),
    .S1(net128),
    .X(_08209_));
 sg13g2_nor2b_1 _28448_ (.A(_08204_),
    .B_N(_08209_),
    .Y(_08210_));
 sg13g2_buf_1 _28449_ (.A(net152),
    .X(_08211_));
 sg13g2_mux2_1 _28450_ (.A0(_00280_),
    .A1(_00279_),
    .S(_08211_),
    .X(_08212_));
 sg13g2_buf_1 _28451_ (.A(net130),
    .X(_08213_));
 sg13g2_mux2_1 _28452_ (.A0(_00282_),
    .A1(_00281_),
    .S(net110),
    .X(_08214_));
 sg13g2_a22oi_1 _28453_ (.Y(_08215_),
    .B1(_08214_),
    .B2(net99),
    .A2(_08212_),
    .A1(net98));
 sg13g2_nand2_1 _28454_ (.Y(_08216_),
    .A(net158),
    .B(_08215_));
 sg13g2_mux4_1 _28455_ (.S0(net97),
    .A0(_00286_),
    .A1(_00285_),
    .A2(_00284_),
    .A3(_00283_),
    .S1(net111),
    .X(_08217_));
 sg13g2_nor2_1 _28456_ (.A(_08216_),
    .B(_08217_),
    .Y(_08218_));
 sg13g2_mux2_1 _28457_ (.A0(_00290_),
    .A1(_00289_),
    .S(_08211_),
    .X(_08219_));
 sg13g2_mux2_1 _28458_ (.A0(_00288_),
    .A1(_00287_),
    .S(_08213_),
    .X(_08220_));
 sg13g2_a22oi_1 _28459_ (.Y(_08221_),
    .B1(_08220_),
    .B2(net98),
    .A2(_08219_),
    .A1(net99));
 sg13g2_nand2_1 _28460_ (.Y(_08222_),
    .A(net175),
    .B(_08221_));
 sg13g2_mux4_1 _28461_ (.S0(net97),
    .A0(_00294_),
    .A1(_00293_),
    .A2(_00292_),
    .A3(_00291_),
    .S1(net111),
    .X(_08223_));
 sg13g2_nor2_1 _28462_ (.A(_08222_),
    .B(_08223_),
    .Y(_08224_));
 sg13g2_a21oi_1 _28463_ (.A1(_08216_),
    .A2(_08222_),
    .Y(_08225_),
    .B1(net128));
 sg13g2_nor4_1 _28464_ (.A(_08053_),
    .B(_08218_),
    .C(_08224_),
    .D(_08225_),
    .Y(_08226_));
 sg13g2_mux2_1 _28465_ (.A0(_00322_),
    .A1(_00321_),
    .S(net130),
    .X(_08227_));
 sg13g2_mux2_1 _28466_ (.A0(_00320_),
    .A1(_00319_),
    .S(net130),
    .X(_08228_));
 sg13g2_a22oi_1 _28467_ (.Y(_08229_),
    .B1(_08228_),
    .B2(net116),
    .A2(_08227_),
    .A1(net112));
 sg13g2_nand2_1 _28468_ (.Y(_08230_),
    .A(net175),
    .B(_08229_));
 sg13g2_mux4_1 _28469_ (.S0(net113),
    .A0(_00326_),
    .A1(_00325_),
    .A2(_00324_),
    .A3(_00323_),
    .S1(net126),
    .X(_08231_));
 sg13g2_nor2_1 _28470_ (.A(_08230_),
    .B(_08231_),
    .Y(_08232_));
 sg13g2_mux2_1 _28471_ (.A0(_00314_),
    .A1(_00313_),
    .S(net152),
    .X(_08233_));
 sg13g2_mux2_1 _28472_ (.A0(_00312_),
    .A1(_00311_),
    .S(_07943_),
    .X(_08234_));
 sg13g2_a22oi_1 _28473_ (.Y(_08235_),
    .B1(_08234_),
    .B2(net116),
    .A2(_08233_),
    .A1(net112));
 sg13g2_nand2_1 _28474_ (.Y(_08236_),
    .A(net153),
    .B(_08235_));
 sg13g2_mux4_1 _28475_ (.S0(net115),
    .A0(_00318_),
    .A1(_00317_),
    .A2(_00316_),
    .A3(_00315_),
    .S1(net133),
    .X(_08237_));
 sg13g2_nor2_1 _28476_ (.A(_07858_),
    .B(net176),
    .Y(_08238_));
 sg13g2_o21ai_1 _28477_ (.B1(_08238_),
    .Y(_08239_),
    .A1(_08236_),
    .A2(_08237_));
 sg13g2_or2_1 _28478_ (.X(_08240_),
    .B(_08239_),
    .A(_08232_));
 sg13g2_a21oi_1 _28479_ (.A1(_08230_),
    .A2(_08236_),
    .Y(_08241_),
    .B1(_07957_));
 sg13g2_mux4_1 _28480_ (.S0(_07962_),
    .A0(_00278_),
    .A1(_00277_),
    .A2(_00276_),
    .A3(_00275_),
    .S1(_07964_),
    .X(_08242_));
 sg13g2_mux2_1 _28481_ (.A0(_00272_),
    .A1(_00271_),
    .S(_07969_),
    .X(_08243_));
 sg13g2_mux2_1 _28482_ (.A0(_00274_),
    .A1(_00273_),
    .S(net127),
    .X(_08244_));
 sg13g2_a221oi_1 _28483_ (.B2(net112),
    .C1(net153),
    .B1(_08244_),
    .A1(net116),
    .Y(_08245_),
    .A2(_08243_));
 sg13g2_nand2b_1 _28484_ (.Y(_08246_),
    .B(_08245_),
    .A_N(_08242_));
 sg13g2_mux4_1 _28485_ (.S0(_07962_),
    .A0(_00270_),
    .A1(_00269_),
    .A2(_00268_),
    .A3(_00267_),
    .S1(_07964_),
    .X(_08247_));
 sg13g2_mux2_1 _28486_ (.A0(_00266_),
    .A1(_00265_),
    .S(net125),
    .X(_08248_));
 sg13g2_mux2_1 _28487_ (.A0(_00264_),
    .A1(_00263_),
    .S(net127),
    .X(_08249_));
 sg13g2_a221oi_1 _28488_ (.B2(net116),
    .C1(net175),
    .B1(_08249_),
    .A1(_08042_),
    .Y(_08250_),
    .A2(_08248_));
 sg13g2_nand2b_1 _28489_ (.Y(_08251_),
    .B(_08250_),
    .A_N(_08247_));
 sg13g2_o21ai_1 _28490_ (.B1(net132),
    .Y(_08252_),
    .A1(_08245_),
    .A2(_08250_));
 sg13g2_nand4_1 _28491_ (.B(_08246_),
    .C(_08251_),
    .A(_07866_),
    .Y(_08253_),
    .D(_08252_));
 sg13g2_o21ai_1 _28492_ (.B1(_08253_),
    .Y(_08254_),
    .A1(_08240_),
    .A2(_08241_));
 sg13g2_nor3_1 _28493_ (.A(_08210_),
    .B(_08226_),
    .C(_08254_),
    .Y(_08255_));
 sg13g2_nor3_1 _28494_ (.A(net115),
    .B(_07963_),
    .C(_07890_),
    .Y(_08256_));
 sg13g2_nand2b_1 _28495_ (.Y(_08257_),
    .B(_08256_),
    .A_N(_07922_));
 sg13g2_o21ai_1 _28496_ (.B1(net812),
    .Y(_08258_),
    .A1(_07854_),
    .A2(_08256_));
 sg13g2_o21ai_1 _28497_ (.B1(_08006_),
    .Y(_08259_),
    .A1(net812),
    .A2(_07924_));
 sg13g2_a221oi_1 _28498_ (.B2(_01959_),
    .C1(_08259_),
    .B1(_08258_),
    .A1(_08003_),
    .Y(_08260_),
    .A2(_08257_));
 sg13g2_nand2_1 _28499_ (.Y(_08261_),
    .A(net809),
    .B(_07911_));
 sg13g2_nand3b_1 _28500_ (.B(_08261_),
    .C(net810),
    .Y(_08262_),
    .A_N(_07928_));
 sg13g2_nand3b_1 _28501_ (.B(_08262_),
    .C(_07907_),
    .Y(_08263_),
    .A_N(_08260_));
 sg13g2_o21ai_1 _28502_ (.B1(_08263_),
    .Y(_08264_),
    .A1(net801),
    .A2(_08255_));
 sg13g2_mux2_1 _28503_ (.A0(_08203_),
    .A1(_08264_),
    .S(_07905_),
    .X(_08265_));
 sg13g2_a21oi_1 _28504_ (.A1(_07652_),
    .A2(_08265_),
    .Y(\rbzero.rgb[2] ),
    .B1(_07998_));
 sg13g2_mux2_1 _28505_ (.A0(_00062_),
    .A1(_00063_),
    .S(_07883_),
    .X(_08266_));
 sg13g2_xor2_1 _28506_ (.B(net132),
    .A(_01965_),
    .X(_08267_));
 sg13g2_nand2b_1 _28507_ (.Y(_08268_),
    .B(net810),
    .A_N(net809));
 sg13g2_nand3_1 _28508_ (.B(_08003_),
    .C(_08006_),
    .A(_07924_),
    .Y(_08269_));
 sg13g2_o21ai_1 _28509_ (.B1(_08269_),
    .Y(_08270_),
    .A1(_08267_),
    .A2(_08268_));
 sg13g2_mux2_1 _28510_ (.A0(_00107_),
    .A1(_00106_),
    .S(net124),
    .X(_08271_));
 sg13g2_mux2_1 _28511_ (.A0(_00105_),
    .A1(_00104_),
    .S(net110),
    .X(_08272_));
 sg13g2_a22oi_1 _28512_ (.Y(_08273_),
    .B1(_08272_),
    .B2(net98),
    .A2(_08271_),
    .A1(net99));
 sg13g2_nand2_1 _28513_ (.Y(_08274_),
    .A(net175),
    .B(_08273_));
 sg13g2_mux4_1 _28514_ (.S0(net97),
    .A0(_00111_),
    .A1(_00110_),
    .A2(_00109_),
    .A3(_00108_),
    .S1(net111),
    .X(_08275_));
 sg13g2_nor2_1 _28515_ (.A(_08274_),
    .B(_08275_),
    .Y(_08276_));
 sg13g2_mux2_1 _28516_ (.A0(_00099_),
    .A1(_00098_),
    .S(net124),
    .X(_08277_));
 sg13g2_mux2_1 _28517_ (.A0(_00097_),
    .A1(_00096_),
    .S(net110),
    .X(_08278_));
 sg13g2_a22oi_1 _28518_ (.Y(_08279_),
    .B1(_08278_),
    .B2(net98),
    .A2(_08277_),
    .A1(net99));
 sg13g2_nand2_1 _28519_ (.Y(_08280_),
    .A(net158),
    .B(_08279_));
 sg13g2_mux4_1 _28520_ (.S0(net97),
    .A0(_00103_),
    .A1(_00102_),
    .A2(_00101_),
    .A3(_00100_),
    .S1(net111),
    .X(_08281_));
 sg13g2_nor2_1 _28521_ (.A(_08280_),
    .B(_08281_),
    .Y(_08282_));
 sg13g2_a21oi_1 _28522_ (.A1(_08274_),
    .A2(_08280_),
    .Y(_08283_),
    .B1(net128));
 sg13g2_nor4_1 _28523_ (.A(_08204_),
    .B(_08276_),
    .C(_08282_),
    .D(_08283_),
    .Y(_08284_));
 sg13g2_mux4_1 _28524_ (.S0(net114),
    .A0(_00123_),
    .A1(_00122_),
    .A2(_00121_),
    .A3(_00120_),
    .S1(net129),
    .X(_08285_));
 sg13g2_mux4_1 _28525_ (.S0(net114),
    .A0(_00115_),
    .A1(_00114_),
    .A2(_00113_),
    .A3(_00112_),
    .S1(net129),
    .X(_08286_));
 sg13g2_buf_1 _28526_ (.A(net155),
    .X(_08287_));
 sg13g2_mux4_1 _28527_ (.S0(_08213_),
    .A0(_00127_),
    .A1(_00126_),
    .A2(_00125_),
    .A3(_00124_),
    .S1(_08287_),
    .X(_08288_));
 sg13g2_mux4_1 _28528_ (.S0(net114),
    .A0(_00119_),
    .A1(_00118_),
    .A2(_00117_),
    .A3(_00116_),
    .S1(net129),
    .X(_08289_));
 sg13g2_mux4_1 _28529_ (.S0(net153),
    .A0(_08285_),
    .A1(_08286_),
    .A2(_08288_),
    .A3(_08289_),
    .S1(net128),
    .X(_08290_));
 sg13g2_nand2b_1 _28530_ (.Y(_08291_),
    .B(_08290_),
    .A_N(net154));
 sg13g2_mux4_1 _28531_ (.S0(net114),
    .A0(_00091_),
    .A1(_00090_),
    .A2(_00089_),
    .A3(_00088_),
    .S1(net129),
    .X(_08292_));
 sg13g2_mux4_1 _28532_ (.S0(net114),
    .A0(_00083_),
    .A1(_00082_),
    .A2(_00081_),
    .A3(_00080_),
    .S1(net129),
    .X(_08293_));
 sg13g2_mux4_1 _28533_ (.S0(net110),
    .A0(_00095_),
    .A1(_00094_),
    .A2(_00093_),
    .A3(_00092_),
    .S1(net123),
    .X(_08294_));
 sg13g2_mux4_1 _28534_ (.S0(net110),
    .A0(_00087_),
    .A1(_00086_),
    .A2(_00085_),
    .A3(_00084_),
    .S1(net123),
    .X(_08295_));
 sg13g2_mux4_1 _28535_ (.S0(net153),
    .A0(_08292_),
    .A1(_08293_),
    .A2(_08294_),
    .A3(_08295_),
    .S1(net128),
    .X(_08296_));
 sg13g2_nand2_1 _28536_ (.Y(_08297_),
    .A(net154),
    .B(_08296_));
 sg13g2_a21oi_1 _28537_ (.A1(_08291_),
    .A2(_08297_),
    .Y(_08298_),
    .B1(net131));
 sg13g2_buf_2 _28538_ (.A(net124),
    .X(_08299_));
 sg13g2_buf_1 _28539_ (.A(_08287_),
    .X(_08300_));
 sg13g2_mux4_1 _28540_ (.S0(net109),
    .A0(_00075_),
    .A1(_00074_),
    .A2(_00073_),
    .A3(_00072_),
    .S1(net108),
    .X(_08301_));
 sg13g2_mux4_1 _28541_ (.S0(net109),
    .A0(_00067_),
    .A1(_00066_),
    .A2(_00065_),
    .A3(_00064_),
    .S1(net108),
    .X(_08302_));
 sg13g2_mux4_1 _28542_ (.S0(net113),
    .A0(_00079_),
    .A1(_00078_),
    .A2(_00077_),
    .A3(_00076_),
    .S1(net126),
    .X(_08303_));
 sg13g2_mux4_1 _28543_ (.S0(net109),
    .A0(_00071_),
    .A1(_00070_),
    .A2(_00069_),
    .A3(_00068_),
    .S1(net108),
    .X(_08304_));
 sg13g2_mux4_1 _28544_ (.S0(net158),
    .A0(_08301_),
    .A1(_08302_),
    .A2(_08303_),
    .A3(_08304_),
    .S1(net128),
    .X(_08305_));
 sg13g2_and2_1 _28545_ (.A(_07866_),
    .B(_08305_),
    .X(_08306_));
 sg13g2_nor4_1 _28546_ (.A(_07906_),
    .B(_08284_),
    .C(_08298_),
    .D(_08306_),
    .Y(_08307_));
 sg13g2_a21oi_1 _28547_ (.A1(net801),
    .A2(_08270_),
    .Y(_08308_),
    .B1(_08307_));
 sg13g2_mux2_1 _28548_ (.A0(_08266_),
    .A1(_08308_),
    .S(_07905_),
    .X(_08309_));
 sg13g2_a21oi_1 _28549_ (.A1(_07652_),
    .A2(_08309_),
    .Y(\rbzero.rgb[3] ),
    .B1(_08202_));
 sg13g2_mux2_1 _28550_ (.A0(_00327_),
    .A1(_00328_),
    .S(_07883_),
    .X(_08310_));
 sg13g2_mux4_1 _28551_ (.S0(net97),
    .A0(_00368_),
    .A1(_00367_),
    .A2(_00366_),
    .A3(_00365_),
    .S1(_08055_),
    .X(_08311_));
 sg13g2_mux2_1 _28552_ (.A0(_00364_),
    .A1(_00363_),
    .S(net134),
    .X(_08312_));
 sg13g2_mux2_1 _28553_ (.A0(_00362_),
    .A1(_00361_),
    .S(net125),
    .X(_08313_));
 sg13g2_a22oi_1 _28554_ (.Y(_08314_),
    .B1(_08313_),
    .B2(net98),
    .A2(_08312_),
    .A1(net112));
 sg13g2_and2_1 _28555_ (.A(net157),
    .B(_08314_),
    .X(_08315_));
 sg13g2_nor2b_1 _28556_ (.A(_08311_),
    .B_N(_08315_),
    .Y(_08316_));
 sg13g2_mux4_1 _28557_ (.S0(_08054_),
    .A0(_00384_),
    .A1(_00383_),
    .A2(_00382_),
    .A3(_00381_),
    .S1(_08055_),
    .X(_08317_));
 sg13g2_mux2_1 _28558_ (.A0(_00380_),
    .A1(_00379_),
    .S(net124),
    .X(_08318_));
 sg13g2_mux2_1 _28559_ (.A0(_00378_),
    .A1(_00377_),
    .S(net124),
    .X(_08319_));
 sg13g2_a221oi_1 _28560_ (.B2(_08045_),
    .C1(net157),
    .B1(_08319_),
    .A1(_08042_),
    .Y(_08320_),
    .A2(_08318_));
 sg13g2_nor2b_1 _28561_ (.A(_08317_),
    .B_N(_08320_),
    .Y(_08321_));
 sg13g2_nor4_1 _28562_ (.A(net154),
    .B(net175),
    .C(_08316_),
    .D(_08321_),
    .Y(_08322_));
 sg13g2_o21ai_1 _28563_ (.B1(net132),
    .Y(_08323_),
    .A1(_08315_),
    .A2(_08320_));
 sg13g2_mux4_1 _28564_ (.S0(_08299_),
    .A0(_00336_),
    .A1(_00335_),
    .A2(_00334_),
    .A3(_00333_),
    .S1(_08300_),
    .X(_08324_));
 sg13g2_mux2_1 _28565_ (.A0(_00330_),
    .A1(_00329_),
    .S(net127),
    .X(_08325_));
 sg13g2_mux2_1 _28566_ (.A0(_00332_),
    .A1(_00331_),
    .S(net127),
    .X(_08326_));
 sg13g2_a22oi_1 _28567_ (.Y(_08327_),
    .B1(_08326_),
    .B2(net99),
    .A2(_08325_),
    .A1(net98));
 sg13g2_and2_1 _28568_ (.A(net157),
    .B(_08327_),
    .X(_08328_));
 sg13g2_nand2b_1 _28569_ (.Y(_08329_),
    .B(_08328_),
    .A_N(_08324_));
 sg13g2_mux4_1 _28570_ (.S0(_08299_),
    .A0(_00352_),
    .A1(_00351_),
    .A2(_00350_),
    .A3(_00349_),
    .S1(_08300_),
    .X(_08330_));
 sg13g2_mux2_1 _28571_ (.A0(_00346_),
    .A1(_00345_),
    .S(net127),
    .X(_08331_));
 sg13g2_mux2_1 _28572_ (.A0(_00348_),
    .A1(_00347_),
    .S(net124),
    .X(_08332_));
 sg13g2_a221oi_1 _28573_ (.B2(net99),
    .C1(net157),
    .B1(_08332_),
    .A1(net98),
    .Y(_08333_),
    .A2(_08331_));
 sg13g2_nand2b_1 _28574_ (.Y(_08334_),
    .B(_08333_),
    .A_N(_08330_));
 sg13g2_and4_1 _28575_ (.A(net154),
    .B(net158),
    .C(_08329_),
    .D(_08334_),
    .X(_08335_));
 sg13g2_o21ai_1 _28576_ (.B1(net132),
    .Y(_08336_),
    .A1(_08328_),
    .A2(_08333_));
 sg13g2_mux4_1 _28577_ (.S0(net124),
    .A0(_00340_),
    .A1(_00339_),
    .A2(_00338_),
    .A3(_00337_),
    .S1(net123),
    .X(_08337_));
 sg13g2_mux4_1 _28578_ (.S0(net130),
    .A0(_00344_),
    .A1(_00343_),
    .A2(_00342_),
    .A3(_00341_),
    .S1(net155),
    .X(_08338_));
 sg13g2_and2_1 _28579_ (.A(_07892_),
    .B(_08338_),
    .X(_08339_));
 sg13g2_a21oi_1 _28580_ (.A1(net132),
    .A2(_08337_),
    .Y(_08340_),
    .B1(_08339_));
 sg13g2_mux4_1 _28581_ (.S0(net134),
    .A0(_00360_),
    .A1(_00359_),
    .A2(_00356_),
    .A3(_00355_),
    .S1(net156),
    .X(_08341_));
 sg13g2_mux4_1 _28582_ (.S0(net130),
    .A0(_00358_),
    .A1(_00357_),
    .A2(_00354_),
    .A3(_00353_),
    .S1(net156),
    .X(_08342_));
 sg13g2_mux2_1 _28583_ (.A0(_08341_),
    .A1(_08342_),
    .S(net123),
    .X(_08343_));
 sg13g2_nor2_1 _28584_ (.A(net157),
    .B(_08343_),
    .Y(_08344_));
 sg13g2_a21oi_1 _28585_ (.A1(net131),
    .A2(_08340_),
    .Y(_08345_),
    .B1(_08344_));
 sg13g2_mux4_1 _28586_ (.S0(net125),
    .A0(_00392_),
    .A1(_00391_),
    .A2(_00390_),
    .A3(_00389_),
    .S1(net151),
    .X(_08346_));
 sg13g2_mux4_1 _28587_ (.S0(net125),
    .A0(_00388_),
    .A1(_00387_),
    .A2(_00386_),
    .A3(_00385_),
    .S1(net151),
    .X(_08347_));
 sg13g2_mux4_1 _28588_ (.S0(net134),
    .A0(_00376_),
    .A1(_00375_),
    .A2(_00374_),
    .A3(_00373_),
    .S1(net151),
    .X(_08348_));
 sg13g2_mux4_1 _28589_ (.S0(net134),
    .A0(_00372_),
    .A1(_00371_),
    .A2(_00370_),
    .A3(_00369_),
    .S1(net151),
    .X(_08349_));
 sg13g2_mux4_1 _28590_ (.S0(net156),
    .A0(_08346_),
    .A1(_08347_),
    .A2(_08348_),
    .A3(_08349_),
    .S1(_07886_),
    .X(_08350_));
 sg13g2_nor2b_1 _28591_ (.A(net154),
    .B_N(_08350_),
    .Y(_08351_));
 sg13g2_a21oi_1 _28592_ (.A1(net154),
    .A2(_08345_),
    .Y(_08352_),
    .B1(_08351_));
 sg13g2_nor2_1 _28593_ (.A(net158),
    .B(_08352_),
    .Y(_08353_));
 sg13g2_a221oi_1 _28594_ (.B2(_08336_),
    .C1(_08353_),
    .B1(_08335_),
    .A1(_08322_),
    .Y(_08354_),
    .A2(_08323_));
 sg13g2_and2_1 _28595_ (.A(_00194_),
    .B(_07854_),
    .X(_08355_));
 sg13g2_nor2b_1 _28596_ (.A(_01959_),
    .B_N(_07922_),
    .Y(_08356_));
 sg13g2_or3_1 _28597_ (.A(net812),
    .B(_08256_),
    .C(_08356_),
    .X(_08357_));
 sg13g2_o21ai_1 _28598_ (.B1(_08004_),
    .Y(_08358_),
    .A1(_08355_),
    .A2(_08357_));
 sg13g2_nand3_1 _28599_ (.B(_07928_),
    .C(_07911_),
    .A(_01987_),
    .Y(_08359_));
 sg13g2_o21ai_1 _28600_ (.B1(_08359_),
    .Y(_08360_),
    .A1(_01987_),
    .A2(_08358_));
 sg13g2_nand2_1 _28601_ (.Y(_08361_),
    .A(net809),
    .B(_08360_));
 sg13g2_nand3_1 _28602_ (.B(_08262_),
    .C(_08361_),
    .A(_07907_),
    .Y(_08362_));
 sg13g2_o21ai_1 _28603_ (.B1(_08362_),
    .Y(_08363_),
    .A1(net801),
    .A2(_08354_));
 sg13g2_mux2_1 _28604_ (.A0(_08310_),
    .A1(_08363_),
    .S(_07905_),
    .X(_08364_));
 sg13g2_a21oi_1 _28605_ (.A1(_07652_),
    .A2(_08364_),
    .Y(\rbzero.rgb[4] ),
    .B1(_07998_));
 sg13g2_xnor2_1 _28606_ (.Y(_08365_),
    .A(_00194_),
    .B(_08054_));
 sg13g2_inv_1 _28607_ (.Y(_08366_),
    .A(_07911_));
 sg13g2_o21ai_1 _28608_ (.B1(net809),
    .Y(_08367_),
    .A1(net812),
    .A2(_08366_));
 sg13g2_o21ai_1 _28609_ (.B1(_08367_),
    .Y(_08368_),
    .A1(net809),
    .A2(_08365_));
 sg13g2_o21ai_1 _28610_ (.B1(_08004_),
    .Y(_08369_),
    .A1(_08045_),
    .A2(_08356_));
 sg13g2_a22oi_1 _28611_ (.Y(_08370_),
    .B1(_08369_),
    .B2(_08006_),
    .A2(_08368_),
    .A1(net810));
 sg13g2_mux4_1 _28612_ (.S0(net110),
    .A0(_00173_),
    .A1(_00172_),
    .A2(_00171_),
    .A3(_00170_),
    .S1(net123),
    .X(_08371_));
 sg13g2_mux4_1 _28613_ (.S0(net110),
    .A0(_00165_),
    .A1(_00164_),
    .A2(_00163_),
    .A3(_00162_),
    .S1(net123),
    .X(_08372_));
 sg13g2_mux4_1 _28614_ (.S0(net124),
    .A0(_00177_),
    .A1(_00176_),
    .A2(_00175_),
    .A3(_00174_),
    .S1(net123),
    .X(_08373_));
 sg13g2_mux4_1 _28615_ (.S0(net110),
    .A0(_00169_),
    .A1(_00168_),
    .A2(_00167_),
    .A3(_00166_),
    .S1(net123),
    .X(_08374_));
 sg13g2_mux4_1 _28616_ (.S0(net153),
    .A0(_08371_),
    .A1(_08372_),
    .A2(_08373_),
    .A3(_08374_),
    .S1(_07892_),
    .X(_08375_));
 sg13g2_mux4_1 _28617_ (.S0(net127),
    .A0(_00135_),
    .A1(_00134_),
    .A2(_00131_),
    .A3(_00130_),
    .S1(net156),
    .X(_08376_));
 sg13g2_mux4_1 _28618_ (.S0(net152),
    .A0(_00137_),
    .A1(_00136_),
    .A2(_00133_),
    .A3(_00132_),
    .S1(_07850_),
    .X(_08377_));
 sg13g2_nor2b_1 _28619_ (.A(_07933_),
    .B_N(_08377_),
    .Y(_08378_));
 sg13g2_a21oi_1 _28620_ (.A1(net108),
    .A2(_08376_),
    .Y(_08379_),
    .B1(_08378_));
 sg13g2_mux4_1 _28621_ (.S0(net130),
    .A0(_00145_),
    .A1(_00144_),
    .A2(_00143_),
    .A3(_00142_),
    .S1(net155),
    .X(_08380_));
 sg13g2_mux4_1 _28622_ (.S0(net130),
    .A0(_00141_),
    .A1(_00140_),
    .A2(_00139_),
    .A3(_00138_),
    .S1(net155),
    .X(_08381_));
 sg13g2_mux2_1 _28623_ (.A0(_08380_),
    .A1(_08381_),
    .S(net156),
    .X(_08382_));
 sg13g2_nor2_1 _28624_ (.A(net153),
    .B(_08382_),
    .Y(_08383_));
 sg13g2_a21oi_1 _28625_ (.A1(net158),
    .A2(_08379_),
    .Y(_08384_),
    .B1(_08383_));
 sg13g2_mux2_1 _28626_ (.A0(_08375_),
    .A1(_08384_),
    .S(net154),
    .X(_08385_));
 sg13g2_mux4_1 _28627_ (.S0(net109),
    .A0(_00189_),
    .A1(_00188_),
    .A2(_00187_),
    .A3(_00186_),
    .S1(net111),
    .X(_08386_));
 sg13g2_mux4_1 _28628_ (.S0(net97),
    .A0(_00181_),
    .A1(_00180_),
    .A2(_00179_),
    .A3(_00178_),
    .S1(net111),
    .X(_08387_));
 sg13g2_mux4_1 _28629_ (.S0(net109),
    .A0(_00193_),
    .A1(_00192_),
    .A2(_00191_),
    .A3(_00190_),
    .S1(net108),
    .X(_08388_));
 sg13g2_mux4_1 _28630_ (.S0(net109),
    .A0(_00185_),
    .A1(_00184_),
    .A2(_00183_),
    .A3(_00182_),
    .S1(net108),
    .X(_08389_));
 sg13g2_mux4_1 _28631_ (.S0(net158),
    .A0(_08386_),
    .A1(_08387_),
    .A2(_08388_),
    .A3(_08389_),
    .S1(net128),
    .X(_08390_));
 sg13g2_mux4_1 _28632_ (.S0(net109),
    .A0(_00149_),
    .A1(_00148_),
    .A2(_00147_),
    .A3(_00146_),
    .S1(net108),
    .X(_08391_));
 sg13g2_mux4_1 _28633_ (.S0(net134),
    .A0(_00153_),
    .A1(_00152_),
    .A2(_00151_),
    .A3(_00150_),
    .S1(net151),
    .X(_08392_));
 sg13g2_a21oi_1 _28634_ (.A1(_07892_),
    .A2(_08392_),
    .Y(_08393_),
    .B1(net175));
 sg13g2_nor2b_1 _28635_ (.A(_08391_),
    .B_N(_08393_),
    .Y(_08394_));
 sg13g2_mux4_1 _28636_ (.S0(net109),
    .A0(_00157_),
    .A1(_00156_),
    .A2(_00155_),
    .A3(_00154_),
    .S1(net108),
    .X(_08395_));
 sg13g2_mux4_1 _28637_ (.S0(net134),
    .A0(_00161_),
    .A1(_00160_),
    .A2(_00159_),
    .A3(_00158_),
    .S1(net151),
    .X(_08396_));
 sg13g2_a21oi_1 _28638_ (.A1(_07892_),
    .A2(_08396_),
    .Y(_08397_),
    .B1(net153));
 sg13g2_nor2b_1 _28639_ (.A(_08395_),
    .B_N(_08397_),
    .Y(_08398_));
 sg13g2_nor2_1 _28640_ (.A(_08393_),
    .B(_08397_),
    .Y(_08399_));
 sg13g2_nor2_1 _28641_ (.A(net132),
    .B(_08399_),
    .Y(_08400_));
 sg13g2_nor4_1 _28642_ (.A(_08053_),
    .B(_08394_),
    .C(_08398_),
    .D(_08400_),
    .Y(_08401_));
 sg13g2_a221oi_1 _28643_ (.B2(_08238_),
    .C1(_08401_),
    .B1(_08390_),
    .A1(net131),
    .Y(_08402_),
    .A2(_08385_));
 sg13g2_nor2_1 _28644_ (.A(net801),
    .B(_08402_),
    .Y(_08403_));
 sg13g2_a21oi_1 _28645_ (.A1(net801),
    .A2(_08370_),
    .Y(_08404_),
    .B1(_08403_));
 sg13g2_mux2_1 _28646_ (.A0(_00128_),
    .A1(_00129_),
    .S(_07883_),
    .X(_08405_));
 sg13g2_nor2_1 _28647_ (.A(_07905_),
    .B(_08405_),
    .Y(_08406_));
 sg13g2_a21oi_1 _28648_ (.A1(_07905_),
    .A2(_08404_),
    .Y(_08407_),
    .B1(_08406_));
 sg13g2_a21oi_1 _28649_ (.A1(_07652_),
    .A2(_08407_),
    .Y(\rbzero.rgb[5] ),
    .B1(_08202_));
 sg13g2_buf_4 _28650_ (.X(_08408_),
    .A(ui_in[6]));
 sg13g2_mux2_1 _28651_ (.A0(\rbzero.rgb[1] ),
    .A1(\registered_vga_output[0] ),
    .S(_08408_),
    .X(net17));
 sg13g2_mux2_1 _28652_ (.A0(\rbzero.rgb[3] ),
    .A1(\registered_vga_output[1] ),
    .S(_08408_),
    .X(net18));
 sg13g2_mux2_1 _28653_ (.A0(\rbzero.rgb[5] ),
    .A1(\registered_vga_output[2] ),
    .S(_08408_),
    .X(net19));
 sg13g2_mux2_1 _28654_ (.A0(\rbzero.vsync_n ),
    .A1(\registered_vga_output[3] ),
    .S(_08408_),
    .X(net20));
 sg13g2_mux2_1 _28655_ (.A0(\rbzero.rgb[0] ),
    .A1(\registered_vga_output[4] ),
    .S(_08408_),
    .X(net21));
 sg13g2_mux2_1 _28656_ (.A0(\rbzero.rgb[2] ),
    .A1(\registered_vga_output[5] ),
    .S(_08408_),
    .X(net22));
 sg13g2_mux2_1 _28657_ (.A0(\rbzero.rgb[4] ),
    .A1(\registered_vga_output[6] ),
    .S(_08408_),
    .X(net23));
 sg13g2_mux2_1 _28658_ (.A0(hsync_n),
    .A1(\registered_vga_output[7] ),
    .S(_08408_),
    .X(net24));
 sg13g2_inv_1 _27863__1 (.Y(net2202),
    .A(clknet_leaf_76_clk));
 sg13g2_tiehi _28661__844 (.L_HI(net844));
 sg13g2_buf_1 _28661_ (.A(net844),
    .X(uio_oe[0]));
 sg13g2_buf_1 _28662_ (.A(net845),
    .X(uio_oe[1]));
 sg13g2_buf_1 _28663_ (.A(net834),
    .X(uio_oe[2]));
 sg13g2_buf_1 _28664_ (.A(net835),
    .X(uio_oe[3]));
 sg13g2_buf_1 _28665_ (.A(net836),
    .X(uio_oe[4]));
 sg13g2_buf_1 _28666_ (.A(net837),
    .X(uio_oe[6]));
 sg13g2_buf_1 _28667_ (.A(net838),
    .X(uio_oe[7]));
 sg13g2_buf_1 _28668_ (.A(\rbzero.o_tex_csb ),
    .X(net14));
 sg13g2_buf_1 _28669_ (.A(net2586),
    .X(net15));
 sg13g2_buf_1 _28670_ (.A(net839),
    .X(uio_out[2]));
 sg13g2_buf_1 _28671_ (.A(net840),
    .X(uio_out[3]));
 sg13g2_buf_1 _28672_ (.A(net841),
    .X(uio_out[4]));
 sg13g2_buf_1 _28673_ (.A(\rbzero.o_tex_out0 ),
    .X(net16));
 sg13g2_buf_1 _28674_ (.A(net842),
    .X(uio_out[6]));
 sg13g2_buf_1 _28675_ (.A(net843),
    .X(uio_out[7]));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net846),
    .D(_00476_),
    .Q_N(_14975_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net847),
    .D(_00477_),
    .Q_N(_14974_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net848),
    .D(_00478_),
    .Q_N(_14973_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net849),
    .D(_00479_),
    .Q_N(_14972_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net850),
    .D(_00480_),
    .Q_N(_14971_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net851),
    .D(_00481_),
    .Q_N(_14970_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net852),
    .D(_00482_),
    .Q_N(_14969_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[6]$_SDFFE_PN1P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net853),
    .D(_00483_),
    .Q_N(_14968_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net854),
    .D(_00484_),
    .Q_N(_14967_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net855),
    .D(_00485_),
    .Q_N(_14966_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRX[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net856),
    .D(_00486_),
    .Q_N(_14965_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net857),
    .D(_00487_),
    .Q_N(_14964_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[10]$_SDFFE_PN1P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net858),
    .D(_00488_),
    .Q_N(_14963_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net859),
    .D(_00489_),
    .Q_N(_14962_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net860),
    .D(_00490_),
    .Q_N(_14961_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net861),
    .D(_00491_),
    .Q_N(_14960_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net862),
    .D(_00492_),
    .Q_N(_14959_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net863),
    .D(_00493_),
    .Q_N(_14958_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net864),
    .D(_00494_),
    .Q_N(_14957_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net865),
    .D(_00495_),
    .Q_N(_14956_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net866),
    .D(_00496_),
    .Q_N(_14955_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.facingRY[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net867),
    .D(_00497_),
    .Q_N(_14954_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.mosi_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net868),
    .D(_00498_),
    .Q_N(_14953_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.mosi_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net869),
    .D(_00499_),
    .Q_N(_14952_),
    .Q(\rbzero.pov.mosi ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net870),
    .D(_00500_),
    .Q_N(_00057_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[10]$_SDFFE_PN1P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net871),
    .D(_00501_),
    .Q_N(_14951_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net872),
    .D(_00502_),
    .Q_N(_14950_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[12]$_SDFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net873),
    .D(_00503_),
    .Q_N(_14949_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net874),
    .D(_00504_),
    .Q_N(_14948_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net875),
    .D(_00505_),
    .Q_N(_14947_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net876),
    .D(_00506_),
    .Q_N(_00443_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net877),
    .D(_00507_),
    .Q_N(_00437_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net878),
    .D(_00508_),
    .Q_N(_00431_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net879),
    .D(_00509_),
    .Q_N(_00425_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net880),
    .D(_00510_),
    .Q_N(_00419_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net881),
    .D(_00511_),
    .Q_N(_00413_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net882),
    .D(_00512_),
    .Q_N(_00408_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net883),
    .D(_00513_),
    .Q_N(_00402_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRX[9]$_SDFFE_PN1P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net884),
    .D(_00514_),
    .Q_N(_14946_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net885),
    .D(_00515_),
    .Q_N(_00059_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[10]$_SDFFE_PN1P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net886),
    .D(_00516_),
    .Q_N(_14945_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net887),
    .D(_00517_),
    .Q_N(_14944_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[12]$_SDFFE_PN1P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net888),
    .D(_00518_),
    .Q_N(_14943_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net889),
    .D(_00519_),
    .Q_N(_14942_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net890),
    .D(_00520_),
    .Q_N(_14941_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net891),
    .D(_00521_),
    .Q_N(_00442_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net892),
    .D(_00522_),
    .Q_N(_00436_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net893),
    .D(_00523_),
    .Q_N(_00430_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net894),
    .D(_00524_),
    .Q_N(_00424_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net895),
    .D(_00525_),
    .Q_N(_00418_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net896),
    .D(_00526_),
    .Q_N(_00412_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net897),
    .D(_00527_),
    .Q_N(_00407_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[8]$_SDFFE_PN1P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net898),
    .D(_00528_),
    .Q_N(_00401_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.playerRY[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net899),
    .D(_00529_),
    .Q_N(_14940_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready$_SDFFE_PP0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net900),
    .D(_00530_),
    .Q_N(_14939_),
    .Q(\rbzero.pov.ready ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net901),
    .D(_00531_),
    .Q_N(_14938_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net902),
    .D(_00532_),
    .Q_N(_14937_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net903),
    .D(_00533_),
    .Q_N(_14936_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net904),
    .D(_00534_),
    .Q_N(_14935_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net905),
    .D(_00535_),
    .Q_N(_14934_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net906),
    .D(_00536_),
    .Q_N(_14933_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net907),
    .D(_00537_),
    .Q_N(_14932_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net908),
    .D(_00538_),
    .Q_N(_14931_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net909),
    .D(_00539_),
    .Q_N(_14930_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net910),
    .D(_00540_),
    .Q_N(_14929_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net911),
    .D(_00541_),
    .Q_N(_14928_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net912),
    .D(_00542_),
    .Q_N(_14927_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net913),
    .D(_00543_),
    .Q_N(_14926_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net914),
    .D(_00544_),
    .Q_N(_14925_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net915),
    .D(_00545_),
    .Q_N(_14924_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net916),
    .D(_00546_),
    .Q_N(_14923_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net917),
    .D(_00547_),
    .Q_N(_14922_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net918),
    .D(_00548_),
    .Q_N(_14921_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net919),
    .D(_00549_),
    .Q_N(_14920_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net920),
    .D(_00550_),
    .Q_N(_14919_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net921),
    .D(_00551_),
    .Q_N(_14918_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net922),
    .D(_00552_),
    .Q_N(_14917_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net923),
    .D(_00553_),
    .Q_N(_14916_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net924),
    .D(_00554_),
    .Q_N(_14915_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net925),
    .D(_00555_),
    .Q_N(_14914_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net926),
    .D(_00556_),
    .Q_N(_14913_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net927),
    .D(_00557_),
    .Q_N(_14912_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net928),
    .D(_00558_),
    .Q_N(_14911_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net929),
    .D(_00559_),
    .Q_N(_14910_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net930),
    .D(_00560_),
    .Q_N(_14909_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net931),
    .D(_00561_),
    .Q_N(_14908_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net932),
    .D(_00562_),
    .Q_N(_14907_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net933),
    .D(_00563_),
    .Q_N(_14906_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net934),
    .D(_00564_),
    .Q_N(_14905_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net935),
    .D(_00565_),
    .Q_N(_14904_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net936),
    .D(_00566_),
    .Q_N(_14903_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net937),
    .D(_00567_),
    .Q_N(_14902_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net938),
    .D(_00568_),
    .Q_N(_14901_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net939),
    .D(_00569_),
    .Q_N(_14900_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net940),
    .D(_00570_),
    .Q_N(_14899_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net941),
    .D(_00571_),
    .Q_N(_14898_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net942),
    .D(_00572_),
    .Q_N(_14897_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net943),
    .D(_00573_),
    .Q_N(_14896_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net944),
    .D(_00574_),
    .Q_N(_14895_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net945),
    .D(_00575_),
    .Q_N(_14894_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net946),
    .D(_00576_),
    .Q_N(_14893_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net947),
    .D(_00577_),
    .Q_N(_14892_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net948),
    .D(_00578_),
    .Q_N(_14891_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net949),
    .D(_00579_),
    .Q_N(_14890_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net950),
    .D(_00580_),
    .Q_N(_14889_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net951),
    .D(_00581_),
    .Q_N(_14888_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net952),
    .D(_00582_),
    .Q_N(_14887_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net953),
    .D(_00583_),
    .Q_N(_14886_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net954),
    .D(_00584_),
    .Q_N(_14885_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net955),
    .D(_00585_),
    .Q_N(_14884_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net956),
    .D(_00586_),
    .Q_N(_14883_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net957),
    .D(_00587_),
    .Q_N(_14882_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net958),
    .D(_00588_),
    .Q_N(_14881_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net959),
    .D(_00589_),
    .Q_N(_14880_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net960),
    .D(_00590_),
    .Q_N(_14879_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[64]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net961),
    .D(_00591_),
    .Q_N(_14878_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[65]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net962),
    .D(_00592_),
    .Q_N(_14877_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[66]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net963),
    .D(_00593_),
    .Q_N(_14876_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[67]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net964),
    .D(_00594_),
    .Q_N(_14875_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[68]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net965),
    .D(_00595_),
    .Q_N(_14874_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[69]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net966),
    .D(_00596_),
    .Q_N(_14873_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net967),
    .D(_00597_),
    .Q_N(_14872_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[70]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net968),
    .D(_00598_),
    .Q_N(_14871_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[71]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net969),
    .D(_00599_),
    .Q_N(_14870_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[72]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net970),
    .D(_00600_),
    .Q_N(_14869_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[73]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net971),
    .D(_00601_),
    .Q_N(_14868_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net972),
    .D(_00602_),
    .Q_N(_14867_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net973),
    .D(_00603_),
    .Q_N(_14866_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sg13g2_dfrbp_1 \rbzero.pov.ready_buffer[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net974),
    .D(_00604_),
    .Q_N(_14865_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sg13g2_dfrbp_1 \rbzero.pov.sclk_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net975),
    .D(_00605_),
    .Q_N(_14864_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.sclk_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net976),
    .D(_00606_),
    .Q_N(_14863_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.sclk_buffer[2]$_SDFF_PN0_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net977),
    .D(_00607_),
    .Q_N(_14862_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net978),
    .D(_00608_),
    .Q_N(_14861_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net979),
    .D(_00609_),
    .Q_N(_14860_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net980),
    .D(_00610_),
    .Q_N(_14859_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net981),
    .D(_00611_),
    .Q_N(_14858_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net982),
    .D(_00612_),
    .Q_N(_14857_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net983),
    .D(_00613_),
    .Q_N(_14856_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net984),
    .D(_00614_),
    .Q_N(_14855_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net985),
    .D(_00615_),
    .Q_N(_14854_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net986),
    .D(_00616_),
    .Q_N(_14853_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net987),
    .D(_00617_),
    .Q_N(_14852_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net988),
    .D(_00618_),
    .Q_N(_14851_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net989),
    .D(_00619_),
    .Q_N(_14850_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net990),
    .D(_00620_),
    .Q_N(_14849_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net991),
    .D(_00621_),
    .Q_N(_14848_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net992),
    .D(_00622_),
    .Q_N(_14847_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net993),
    .D(_00623_),
    .Q_N(_14846_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net994),
    .D(_00624_),
    .Q_N(_14845_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net995),
    .D(_00625_),
    .Q_N(_14844_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net996),
    .D(_00626_),
    .Q_N(_14843_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net997),
    .D(_00627_),
    .Q_N(_14842_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net998),
    .D(_00628_),
    .Q_N(_14841_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net999),
    .D(_00629_),
    .Q_N(_14840_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1000),
    .D(_00630_),
    .Q_N(_14839_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1001),
    .D(_00631_),
    .Q_N(_14838_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1002),
    .D(_00632_),
    .Q_N(_14837_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1003),
    .D(_00633_),
    .Q_N(_14836_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1004),
    .D(_00634_),
    .Q_N(_14835_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1005),
    .D(_00635_),
    .Q_N(_14834_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1006),
    .D(_00636_),
    .Q_N(_14833_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1007),
    .D(_00637_),
    .Q_N(_14832_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1008),
    .D(_00638_),
    .Q_N(_14831_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1009),
    .D(_00639_),
    .Q_N(_14830_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1010),
    .D(_00640_),
    .Q_N(_14829_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1011),
    .D(_00641_),
    .Q_N(_14828_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[40]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1012),
    .D(_00642_),
    .Q_N(_14827_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1013),
    .D(_00643_),
    .Q_N(_14826_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1014),
    .D(_00644_),
    .Q_N(_14825_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1015),
    .D(_00645_),
    .Q_N(_14824_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1016),
    .D(_00646_),
    .Q_N(_14823_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1017),
    .D(_00647_),
    .Q_N(_14822_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1018),
    .D(_00648_),
    .Q_N(_14821_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1019),
    .D(_00649_),
    .Q_N(_14820_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1020),
    .D(_00650_),
    .Q_N(_14819_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1021),
    .D(_00651_),
    .Q_N(_14818_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1022),
    .D(_00652_),
    .Q_N(_14817_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1023),
    .D(_00653_),
    .Q_N(_14816_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1024),
    .D(_00654_),
    .Q_N(_14815_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1025),
    .D(_00655_),
    .Q_N(_14814_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1026),
    .D(_00656_),
    .Q_N(_14813_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1027),
    .D(_00657_),
    .Q_N(_14812_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1028),
    .D(_00658_),
    .Q_N(_14811_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1029),
    .D(_00659_),
    .Q_N(_14810_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1030),
    .D(_00660_),
    .Q_N(_14809_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1031),
    .D(_00661_),
    .Q_N(_14808_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1032),
    .D(_00662_),
    .Q_N(_14807_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1033),
    .D(_00663_),
    .Q_N(_14806_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1034),
    .D(_00664_),
    .Q_N(_14805_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1035),
    .D(_00665_),
    .Q_N(_14804_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1036),
    .D(_00666_),
    .Q_N(_14803_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1037),
    .D(_00667_),
    .Q_N(_14802_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[64]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1038),
    .D(_00668_),
    .Q_N(_14801_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[65]$_SDFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1039),
    .D(_00669_),
    .Q_N(_14800_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[66]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1040),
    .D(_00670_),
    .Q_N(_14799_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[67]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1041),
    .D(_00671_),
    .Q_N(_14798_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[68]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1042),
    .D(_00672_),
    .Q_N(_14797_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[69]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1043),
    .D(_00673_),
    .Q_N(_14796_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1044),
    .D(_00674_),
    .Q_N(_14795_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[70]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1045),
    .D(_00675_),
    .Q_N(_14794_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[71]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1046),
    .D(_00676_),
    .Q_N(_14793_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[72]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1047),
    .D(_00677_),
    .Q_N(_14792_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[73]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1048),
    .D(_00678_),
    .Q_N(_14791_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1049),
    .D(_00679_),
    .Q_N(_14790_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1050),
    .D(_00680_),
    .Q_N(_14789_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_buffer[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1051),
    .D(_00681_),
    .Q_N(_14788_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1052),
    .D(_00682_),
    .Q_N(_14787_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[1]$_SDFFE_PP0N_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1053),
    .D(_00683_),
    .Q_N(_14786_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[2]$_SDFFE_PP0N_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1054),
    .D(_00684_),
    .Q_N(_14785_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[3]$_SDFFE_PP0N_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1055),
    .D(_00685_),
    .Q_N(_14784_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[4]$_SDFFE_PP0N_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1056),
    .D(_00686_),
    .Q_N(_14783_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[5]$_SDFFE_PP0N_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1057),
    .D(_00687_),
    .Q_N(_14782_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_counter[6]$_SDFFE_PP0N_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1058),
    .D(_00688_),
    .Q_N(_00026_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sg13g2_dfrbp_1 \rbzero.pov.spi_done$_SDFF_PP0_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1059),
    .D(_00689_),
    .Q_N(_14781_),
    .Q(\rbzero.pov.spi_done ));
 sg13g2_dfrbp_1 \rbzero.pov.ss_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1060),
    .D(_00690_),
    .Q_N(_14780_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.ss_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1061),
    .D(_00691_),
    .Q_N(_14779_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1062),
    .D(_00692_),
    .Q_N(_00060_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1063),
    .D(_00693_),
    .Q_N(_14778_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1064),
    .D(_00694_),
    .Q_N(_14777_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1065),
    .D(_00695_),
    .Q_N(_14776_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1066),
    .D(_00696_),
    .Q_N(_14775_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1067),
    .D(_00697_),
    .Q_N(_14774_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1068),
    .D(_00698_),
    .Q_N(_14773_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1069),
    .D(_00699_),
    .Q_N(_14772_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1070),
    .D(_00700_),
    .Q_N(_14771_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1071),
    .D(_00701_),
    .Q_N(_14770_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRX[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1072),
    .D(_00702_),
    .Q_N(_14769_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1073),
    .D(_00703_),
    .Q_N(_00061_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1074),
    .D(_00704_),
    .Q_N(_14768_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1075),
    .D(_00705_),
    .Q_N(_14767_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1076),
    .D(_00706_),
    .Q_N(_14766_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1077),
    .D(_00707_),
    .Q_N(_14765_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1078),
    .D(_00708_),
    .Q_N(_14764_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1079),
    .D(_00709_),
    .Q_N(_14763_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1080),
    .D(_00710_),
    .Q_N(_14762_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[7]$_SDFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1081),
    .D(_00711_),
    .Q_N(_14761_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1082),
    .D(_00712_),
    .Q_N(_14760_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sg13g2_dfrbp_1 \rbzero.pov.vplaneRY[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1083),
    .D(_00713_),
    .Q_N(_14759_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1084),
    .D(_00714_),
    .Q_N(_14758_),
    .Q(\rbzero.spi_registers.buf_floor[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1085),
    .D(_00715_),
    .Q_N(_14757_),
    .Q(\rbzero.spi_registers.buf_floor[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1086),
    .D(_00716_),
    .Q_N(_14756_),
    .Q(\rbzero.spi_registers.buf_floor[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1087),
    .D(_00717_),
    .Q_N(_14755_),
    .Q(\rbzero.spi_registers.buf_floor[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1088),
    .D(_00718_),
    .Q_N(_14754_),
    .Q(\rbzero.spi_registers.buf_floor[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_floor[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1089),
    .D(_00719_),
    .Q_N(_14753_),
    .Q(\rbzero.spi_registers.buf_floor[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1090),
    .D(_00720_),
    .Q_N(_14752_),
    .Q(\rbzero.spi_registers.buf_leak[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1091),
    .D(_00721_),
    .Q_N(_14751_),
    .Q(\rbzero.spi_registers.buf_leak[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1092),
    .D(_00722_),
    .Q_N(_14750_),
    .Q(\rbzero.spi_registers.buf_leak[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1093),
    .D(_00723_),
    .Q_N(_14749_),
    .Q(\rbzero.spi_registers.buf_leak[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1094),
    .D(_00724_),
    .Q_N(_14748_),
    .Q(\rbzero.spi_registers.buf_leak[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_leak[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1095),
    .D(_00725_),
    .Q_N(_14747_),
    .Q(\rbzero.spi_registers.buf_leak[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1096),
    .D(_00726_),
    .Q_N(_14746_),
    .Q(\rbzero.spi_registers.buf_mapdx[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1097),
    .D(_00727_),
    .Q_N(_14745_),
    .Q(\rbzero.spi_registers.buf_mapdx[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1098),
    .D(_00728_),
    .Q_N(_14744_),
    .Q(\rbzero.spi_registers.buf_mapdx[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdx[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1099),
    .D(_00729_),
    .Q_N(_14743_),
    .Q(\rbzero.spi_registers.buf_mapdx[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdx[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1100),
    .D(_00730_),
    .Q_N(_14742_),
    .Q(\rbzero.spi_registers.buf_mapdx[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdxw[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1101),
    .D(_00731_),
    .Q_N(_14741_),
    .Q(\rbzero.spi_registers.buf_mapdxw[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdxw[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1102),
    .D(_00732_),
    .Q_N(_14740_),
    .Q(\rbzero.spi_registers.buf_mapdxw[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdy[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1103),
    .D(_00733_),
    .Q_N(_14739_),
    .Q(\rbzero.spi_registers.buf_mapdy[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdy[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1104),
    .D(_00734_),
    .Q_N(_14738_),
    .Q(\rbzero.spi_registers.buf_mapdy[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdy[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1105),
    .D(_00735_),
    .Q_N(_14737_),
    .Q(\rbzero.spi_registers.buf_mapdy[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdy[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1106),
    .D(_00736_),
    .Q_N(_14736_),
    .Q(\rbzero.spi_registers.buf_mapdy[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdy[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1107),
    .D(_00737_),
    .Q_N(_14735_),
    .Q(\rbzero.spi_registers.buf_mapdy[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdyw[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1108),
    .D(_00738_),
    .Q_N(_14734_),
    .Q(\rbzero.spi_registers.buf_mapdyw[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_mapdyw[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1109),
    .D(_00739_),
    .Q_N(_14733_),
    .Q(\rbzero.spi_registers.buf_mapdyw[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_otherx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1110),
    .D(_00740_),
    .Q_N(_14732_),
    .Q(\rbzero.spi_registers.buf_otherx[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_otherx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1111),
    .D(_00741_),
    .Q_N(_14731_),
    .Q(\rbzero.spi_registers.buf_otherx[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_otherx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1112),
    .D(_00742_),
    .Q_N(_14730_),
    .Q(\rbzero.spi_registers.buf_otherx[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_otherx[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1113),
    .D(_00743_),
    .Q_N(_14729_),
    .Q(\rbzero.spi_registers.buf_otherx[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_otherx[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1114),
    .D(_00744_),
    .Q_N(_14728_),
    .Q(\rbzero.spi_registers.buf_otherx[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_othery[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1115),
    .D(_00745_),
    .Q_N(_14727_),
    .Q(\rbzero.spi_registers.buf_othery[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_othery[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1116),
    .D(_00746_),
    .Q_N(_14726_),
    .Q(\rbzero.spi_registers.buf_othery[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_othery[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1117),
    .D(_00747_),
    .Q_N(_14725_),
    .Q(\rbzero.spi_registers.buf_othery[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_othery[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1118),
    .D(_00748_),
    .Q_N(_14724_),
    .Q(\rbzero.spi_registers.buf_othery[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_othery[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1119),
    .D(_00749_),
    .Q_N(_14723_),
    .Q(\rbzero.spi_registers.buf_othery[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1120),
    .D(_00750_),
    .Q_N(_14722_),
    .Q(\rbzero.spi_registers.buf_sky[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1121),
    .D(_00751_),
    .Q_N(_14721_),
    .Q(\rbzero.spi_registers.buf_sky[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1122),
    .D(_00752_),
    .Q_N(_14720_),
    .Q(\rbzero.spi_registers.buf_sky[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1123),
    .D(_00753_),
    .Q_N(_14719_),
    .Q(\rbzero.spi_registers.buf_sky[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1124),
    .D(_00754_),
    .Q_N(_14718_),
    .Q(\rbzero.spi_registers.buf_sky[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_sky[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1125),
    .D(_00755_),
    .Q_N(_14717_),
    .Q(\rbzero.spi_registers.buf_sky[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1126),
    .D(_00756_),
    .Q_N(_14716_),
    .Q(\rbzero.spi_registers.buf_texadd0[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1127),
    .D(_00757_),
    .Q_N(_14715_),
    .Q(\rbzero.spi_registers.buf_texadd0[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1128),
    .D(_00758_),
    .Q_N(_14714_),
    .Q(\rbzero.spi_registers.buf_texadd0[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1129),
    .D(_00759_),
    .Q_N(_14713_),
    .Q(\rbzero.spi_registers.buf_texadd0[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1130),
    .D(_00760_),
    .Q_N(_14712_),
    .Q(\rbzero.spi_registers.buf_texadd0[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1131),
    .D(_00761_),
    .Q_N(_14711_),
    .Q(\rbzero.spi_registers.buf_texadd0[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1132),
    .D(_00762_),
    .Q_N(_14710_),
    .Q(\rbzero.spi_registers.buf_texadd0[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1133),
    .D(_00763_),
    .Q_N(_14709_),
    .Q(\rbzero.spi_registers.buf_texadd0[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1134),
    .D(_00764_),
    .Q_N(_14708_),
    .Q(\rbzero.spi_registers.buf_texadd0[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1135),
    .D(_00765_),
    .Q_N(_14707_),
    .Q(\rbzero.spi_registers.buf_texadd0[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1136),
    .D(_00766_),
    .Q_N(_14706_),
    .Q(\rbzero.spi_registers.buf_texadd0[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1137),
    .D(_00767_),
    .Q_N(_14705_),
    .Q(\rbzero.spi_registers.buf_texadd0[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1138),
    .D(_00768_),
    .Q_N(_14704_),
    .Q(\rbzero.spi_registers.buf_texadd0[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1139),
    .D(_00769_),
    .Q_N(_14703_),
    .Q(\rbzero.spi_registers.buf_texadd0[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1140),
    .D(_00770_),
    .Q_N(_14702_),
    .Q(\rbzero.spi_registers.buf_texadd0[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1141),
    .D(_00771_),
    .Q_N(_14701_),
    .Q(\rbzero.spi_registers.buf_texadd0[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1142),
    .D(_00772_),
    .Q_N(_14700_),
    .Q(\rbzero.spi_registers.buf_texadd0[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1143),
    .D(_00773_),
    .Q_N(_14699_),
    .Q(\rbzero.spi_registers.buf_texadd0[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1144),
    .D(_00774_),
    .Q_N(_14698_),
    .Q(\rbzero.spi_registers.buf_texadd0[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1145),
    .D(_00775_),
    .Q_N(_14697_),
    .Q(\rbzero.spi_registers.buf_texadd0[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1146),
    .D(_00776_),
    .Q_N(_14696_),
    .Q(\rbzero.spi_registers.buf_texadd0[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1147),
    .D(_00777_),
    .Q_N(_14695_),
    .Q(\rbzero.spi_registers.buf_texadd0[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1148),
    .D(_00778_),
    .Q_N(_14694_),
    .Q(\rbzero.spi_registers.buf_texadd0[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd0[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1149),
    .D(_00779_),
    .Q_N(_14693_),
    .Q(\rbzero.spi_registers.buf_texadd0[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1150),
    .D(_00780_),
    .Q_N(_14692_),
    .Q(\rbzero.spi_registers.buf_texadd1[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1151),
    .D(_00781_),
    .Q_N(_14691_),
    .Q(\rbzero.spi_registers.buf_texadd1[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1152),
    .D(_00782_),
    .Q_N(_14690_),
    .Q(\rbzero.spi_registers.buf_texadd1[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1153),
    .D(_00783_),
    .Q_N(_14689_),
    .Q(\rbzero.spi_registers.buf_texadd1[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1154),
    .D(_00784_),
    .Q_N(_14688_),
    .Q(\rbzero.spi_registers.buf_texadd1[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1155),
    .D(_00785_),
    .Q_N(_14687_),
    .Q(\rbzero.spi_registers.buf_texadd1[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1156),
    .D(_00786_),
    .Q_N(_14686_),
    .Q(\rbzero.spi_registers.buf_texadd1[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1157),
    .D(_00787_),
    .Q_N(_14685_),
    .Q(\rbzero.spi_registers.buf_texadd1[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1158),
    .D(_00788_),
    .Q_N(_14684_),
    .Q(\rbzero.spi_registers.buf_texadd1[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1159),
    .D(_00789_),
    .Q_N(_14683_),
    .Q(\rbzero.spi_registers.buf_texadd1[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1160),
    .D(_00790_),
    .Q_N(_14682_),
    .Q(\rbzero.spi_registers.buf_texadd1[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1161),
    .D(_00791_),
    .Q_N(_14681_),
    .Q(\rbzero.spi_registers.buf_texadd1[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1162),
    .D(_00792_),
    .Q_N(_14680_),
    .Q(\rbzero.spi_registers.buf_texadd1[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1163),
    .D(_00793_),
    .Q_N(_14679_),
    .Q(\rbzero.spi_registers.buf_texadd1[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1164),
    .D(_00794_),
    .Q_N(_14678_),
    .Q(\rbzero.spi_registers.buf_texadd1[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1165),
    .D(_00795_),
    .Q_N(_14677_),
    .Q(\rbzero.spi_registers.buf_texadd1[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1166),
    .D(_00796_),
    .Q_N(_14676_),
    .Q(\rbzero.spi_registers.buf_texadd1[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1167),
    .D(_00797_),
    .Q_N(_14675_),
    .Q(\rbzero.spi_registers.buf_texadd1[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1168),
    .D(_00798_),
    .Q_N(_14674_),
    .Q(\rbzero.spi_registers.buf_texadd1[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1169),
    .D(_00799_),
    .Q_N(_14673_),
    .Q(\rbzero.spi_registers.buf_texadd1[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1170),
    .D(_00800_),
    .Q_N(_14672_),
    .Q(\rbzero.spi_registers.buf_texadd1[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1171),
    .D(_00801_),
    .Q_N(_14671_),
    .Q(\rbzero.spi_registers.buf_texadd1[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1172),
    .D(_00802_),
    .Q_N(_14670_),
    .Q(\rbzero.spi_registers.buf_texadd1[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1173),
    .D(_00803_),
    .Q_N(_14669_),
    .Q(\rbzero.spi_registers.buf_texadd1[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1174),
    .D(_00804_),
    .Q_N(_14668_),
    .Q(\rbzero.spi_registers.buf_texadd2[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1175),
    .D(_00805_),
    .Q_N(_14667_),
    .Q(\rbzero.spi_registers.buf_texadd2[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1176),
    .D(_00806_),
    .Q_N(_14666_),
    .Q(\rbzero.spi_registers.buf_texadd2[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1177),
    .D(_00807_),
    .Q_N(_14665_),
    .Q(\rbzero.spi_registers.buf_texadd2[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1178),
    .D(_00808_),
    .Q_N(_14664_),
    .Q(\rbzero.spi_registers.buf_texadd2[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1179),
    .D(_00809_),
    .Q_N(_14663_),
    .Q(\rbzero.spi_registers.buf_texadd2[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1180),
    .D(_00810_),
    .Q_N(_14662_),
    .Q(\rbzero.spi_registers.buf_texadd2[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1181),
    .D(_00811_),
    .Q_N(_14661_),
    .Q(\rbzero.spi_registers.buf_texadd2[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1182),
    .D(_00812_),
    .Q_N(_14660_),
    .Q(\rbzero.spi_registers.buf_texadd2[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1183),
    .D(_00813_),
    .Q_N(_14659_),
    .Q(\rbzero.spi_registers.buf_texadd2[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1184),
    .D(_00814_),
    .Q_N(_14658_),
    .Q(\rbzero.spi_registers.buf_texadd2[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1185),
    .D(_00815_),
    .Q_N(_14657_),
    .Q(\rbzero.spi_registers.buf_texadd2[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1186),
    .D(_00816_),
    .Q_N(_14656_),
    .Q(\rbzero.spi_registers.buf_texadd2[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1187),
    .D(_00817_),
    .Q_N(_14655_),
    .Q(\rbzero.spi_registers.buf_texadd2[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1188),
    .D(_00818_),
    .Q_N(_14654_),
    .Q(\rbzero.spi_registers.buf_texadd2[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1189),
    .D(_00819_),
    .Q_N(_14653_),
    .Q(\rbzero.spi_registers.buf_texadd2[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1190),
    .D(_00820_),
    .Q_N(_14652_),
    .Q(\rbzero.spi_registers.buf_texadd2[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1191),
    .D(_00821_),
    .Q_N(_14651_),
    .Q(\rbzero.spi_registers.buf_texadd2[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1192),
    .D(_00822_),
    .Q_N(_14650_),
    .Q(\rbzero.spi_registers.buf_texadd2[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1193),
    .D(_00823_),
    .Q_N(_14649_),
    .Q(\rbzero.spi_registers.buf_texadd2[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1194),
    .D(_00824_),
    .Q_N(_14648_),
    .Q(\rbzero.spi_registers.buf_texadd2[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1195),
    .D(_00825_),
    .Q_N(_14647_),
    .Q(\rbzero.spi_registers.buf_texadd2[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1196),
    .D(_00826_),
    .Q_N(_14646_),
    .Q(\rbzero.spi_registers.buf_texadd2[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1197),
    .D(_00827_),
    .Q_N(_14645_),
    .Q(\rbzero.spi_registers.buf_texadd2[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1198),
    .D(_00828_),
    .Q_N(_14644_),
    .Q(\rbzero.spi_registers.buf_texadd3[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1199),
    .D(_00829_),
    .Q_N(_14643_),
    .Q(\rbzero.spi_registers.buf_texadd3[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1200),
    .D(_00830_),
    .Q_N(_14642_),
    .Q(\rbzero.spi_registers.buf_texadd3[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1201),
    .D(_00831_),
    .Q_N(_14641_),
    .Q(\rbzero.spi_registers.buf_texadd3[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1202),
    .D(_00832_),
    .Q_N(_14640_),
    .Q(\rbzero.spi_registers.buf_texadd3[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1203),
    .D(_00833_),
    .Q_N(_14639_),
    .Q(\rbzero.spi_registers.buf_texadd3[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1204),
    .D(_00834_),
    .Q_N(_14638_),
    .Q(\rbzero.spi_registers.buf_texadd3[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1205),
    .D(_00835_),
    .Q_N(_14637_),
    .Q(\rbzero.spi_registers.buf_texadd3[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1206),
    .D(_00836_),
    .Q_N(_14636_),
    .Q(\rbzero.spi_registers.buf_texadd3[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1207),
    .D(_00837_),
    .Q_N(_14635_),
    .Q(\rbzero.spi_registers.buf_texadd3[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1208),
    .D(_00838_),
    .Q_N(_14634_),
    .Q(\rbzero.spi_registers.buf_texadd3[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1209),
    .D(_00839_),
    .Q_N(_14633_),
    .Q(\rbzero.spi_registers.buf_texadd3[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1210),
    .D(_00840_),
    .Q_N(_14632_),
    .Q(\rbzero.spi_registers.buf_texadd3[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1211),
    .D(_00841_),
    .Q_N(_14631_),
    .Q(\rbzero.spi_registers.buf_texadd3[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1212),
    .D(_00842_),
    .Q_N(_14630_),
    .Q(\rbzero.spi_registers.buf_texadd3[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1213),
    .D(_00843_),
    .Q_N(_14629_),
    .Q(\rbzero.spi_registers.buf_texadd3[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1214),
    .D(_00844_),
    .Q_N(_14628_),
    .Q(\rbzero.spi_registers.buf_texadd3[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1215),
    .D(_00845_),
    .Q_N(_14627_),
    .Q(\rbzero.spi_registers.buf_texadd3[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1216),
    .D(_00846_),
    .Q_N(_14626_),
    .Q(\rbzero.spi_registers.buf_texadd3[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1217),
    .D(_00847_),
    .Q_N(_14625_),
    .Q(\rbzero.spi_registers.buf_texadd3[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1218),
    .D(_00848_),
    .Q_N(_14624_),
    .Q(\rbzero.spi_registers.buf_texadd3[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1219),
    .D(_00849_),
    .Q_N(_14623_),
    .Q(\rbzero.spi_registers.buf_texadd3[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1220),
    .D(_00850_),
    .Q_N(_14622_),
    .Q(\rbzero.spi_registers.buf_texadd3[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_texadd3[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1221),
    .D(_00851_),
    .Q_N(_14621_),
    .Q(\rbzero.spi_registers.buf_texadd3[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vinf$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1222),
    .D(_00852_),
    .Q_N(_14620_),
    .Q(\rbzero.spi_registers.buf_vinf ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1223),
    .D(_00853_),
    .Q_N(_14619_),
    .Q(\rbzero.spi_registers.buf_vshift[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1224),
    .D(_00854_),
    .Q_N(_14618_),
    .Q(\rbzero.spi_registers.buf_vshift[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1225),
    .D(_00855_),
    .Q_N(_14617_),
    .Q(\rbzero.spi_registers.buf_vshift[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1226),
    .D(_00856_),
    .Q_N(_14616_),
    .Q(\rbzero.spi_registers.buf_vshift[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1227),
    .D(_00857_),
    .Q_N(_14615_),
    .Q(\rbzero.spi_registers.buf_vshift[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.buf_vshift[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1228),
    .D(_00858_),
    .Q_N(_14614_),
    .Q(\rbzero.spi_registers.buf_vshift[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1229),
    .D(_00859_),
    .Q_N(_00195_),
    .Q(\rbzero.color_floor[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1230),
    .D(_00860_),
    .Q_N(_14613_),
    .Q(\rbzero.color_floor[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1231),
    .D(_00861_),
    .Q_N(_00261_),
    .Q(\rbzero.color_floor[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1232),
    .D(_00862_),
    .Q_N(_00062_),
    .Q(\rbzero.color_floor[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1233),
    .D(_00863_),
    .Q_N(_00327_),
    .Q(\rbzero.color_floor[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.floor[5]$_SDFFE_PN1P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1234),
    .D(_00864_),
    .Q_N(_00128_),
    .Q(\rbzero.color_floor[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1235),
    .D(_00865_),
    .Q_N(_14612_),
    .Q(\rbzero.floor_leak[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1236),
    .D(_00866_),
    .Q_N(_14611_),
    .Q(\rbzero.floor_leak[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1237),
    .D(_00867_),
    .Q_N(_14610_),
    .Q(\rbzero.floor_leak[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1238),
    .D(_00868_),
    .Q_N(_14609_),
    .Q(\rbzero.floor_leak[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1239),
    .D(_00869_),
    .Q_N(_14608_),
    .Q(\rbzero.floor_leak[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.leak[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1240),
    .D(_00870_),
    .Q_N(_14607_),
    .Q(\rbzero.floor_leak[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1241),
    .D(_00871_),
    .Q_N(_14606_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1242),
    .D(_00872_),
    .Q_N(_14605_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1243),
    .D(_00873_),
    .Q_N(_14604_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdx[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1244),
    .D(_00874_),
    .Q_N(_14603_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdx[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1245),
    .D(_00875_),
    .Q_N(_14602_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdxw[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1246),
    .D(_00876_),
    .Q_N(_14601_),
    .Q(\rbzero.mapdxw[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdxw[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1247),
    .D(_00877_),
    .Q_N(_14600_),
    .Q(\rbzero.mapdxw[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdy[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1248),
    .D(_00878_),
    .Q_N(_14599_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdy[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1249),
    .D(_00879_),
    .Q_N(_14598_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdy[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1250),
    .D(_00880_),
    .Q_N(_14597_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdy[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1251),
    .D(_00881_),
    .Q_N(_14596_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdy[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1252),
    .D(_00882_),
    .Q_N(_14595_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdyw[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1253),
    .D(_00883_),
    .Q_N(_14594_),
    .Q(\rbzero.mapdyw[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mapdyw[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1254),
    .D(_00884_),
    .Q_N(_14593_),
    .Q(\rbzero.mapdyw[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mosi_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1255),
    .D(_00885_),
    .Q_N(_14592_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.mosi_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1256),
    .D(_00886_),
    .Q_N(_14591_),
    .Q(\rbzero.spi_registers.mosi ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.otherx[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1257),
    .D(_00887_),
    .Q_N(_14590_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.otherx[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1258),
    .D(_00888_),
    .Q_N(_14589_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.otherx[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1259),
    .D(_00889_),
    .Q_N(_14588_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.otherx[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1260),
    .D(_00890_),
    .Q_N(_14587_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.otherx[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1261),
    .D(_00891_),
    .Q_N(_14586_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.othery[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1262),
    .D(_00892_),
    .Q_N(_14585_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.othery[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1263),
    .D(_00893_),
    .Q_N(_14584_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.othery[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1264),
    .D(_00894_),
    .Q_N(_14583_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.othery[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1265),
    .D(_00895_),
    .Q_N(_14582_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.othery[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1266),
    .D(_00896_),
    .Q_N(_14581_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sclk_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1267),
    .D(_00897_),
    .Q_N(_14580_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sclk_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1268),
    .D(_00898_),
    .Q_N(_14579_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sclk_buffer[2]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1269),
    .D(_00899_),
    .Q_N(_14578_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1270),
    .D(_00900_),
    .Q_N(_00196_),
    .Q(\rbzero.color_sky[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1271),
    .D(_00901_),
    .Q_N(_14577_),
    .Q(\rbzero.color_sky[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1272),
    .D(_00902_),
    .Q_N(_00262_),
    .Q(\rbzero.color_sky[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1273),
    .D(_00903_),
    .Q_N(_00063_),
    .Q(\rbzero.color_sky[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[4]$_SDFFE_PN1P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1274),
    .D(_00904_),
    .Q_N(_00328_),
    .Q(\rbzero.color_sky[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.sky[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1275),
    .D(_00905_),
    .Q_N(_00129_),
    .Q(\rbzero.color_sky[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1276),
    .D(_00906_),
    .Q_N(_14576_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1277),
    .D(_00907_),
    .Q_N(_14575_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1278),
    .D(_00908_),
    .Q_N(_14574_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1279),
    .D(_00909_),
    .Q_N(_14573_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1280),
    .D(_00910_),
    .Q_N(_14572_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1281),
    .D(_00911_),
    .Q_N(_14571_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1282),
    .D(_00912_),
    .Q_N(_14570_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1283),
    .D(_00913_),
    .Q_N(_14569_),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1284),
    .D(_00914_),
    .Q_N(_14568_),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1285),
    .D(_00915_),
    .Q_N(_14567_),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1286),
    .D(_00916_),
    .Q_N(_14566_),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1287),
    .D(_00917_),
    .Q_N(_14565_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1288),
    .D(_00918_),
    .Q_N(_14564_),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1289),
    .D(_00919_),
    .Q_N(_14563_),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1290),
    .D(_00920_),
    .Q_N(_14562_),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1291),
    .D(_00921_),
    .Q_N(_14561_),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1292),
    .D(_00922_),
    .Q_N(_14560_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1293),
    .D(_00923_),
    .Q_N(_14559_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1294),
    .D(_00924_),
    .Q_N(_14558_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1295),
    .D(_00925_),
    .Q_N(_14557_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1296),
    .D(_00926_),
    .Q_N(_14556_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1297),
    .D(_00927_),
    .Q_N(_14555_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1298),
    .D(_00928_),
    .Q_N(_14554_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_buffer[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1299),
    .D(_00929_),
    .Q_N(_14553_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_cmd[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1300),
    .D(_00930_),
    .Q_N(_14552_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_cmd[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1301),
    .D(_00931_),
    .Q_N(_14551_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_cmd[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1302),
    .D(_00932_),
    .Q_N(_14550_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_cmd[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1303),
    .D(_00933_),
    .Q_N(_14549_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1304),
    .D(_00934_),
    .Q_N(_00475_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1305),
    .D(_00935_),
    .Q_N(_14548_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1306),
    .D(_00936_),
    .Q_N(_14547_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1307),
    .D(_00937_),
    .Q_N(_14546_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1308),
    .D(_00938_),
    .Q_N(_14545_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1309),
    .D(_00939_),
    .Q_N(_14544_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_counter[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1310),
    .D(_00940_),
    .Q_N(_14543_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.spi_done$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1311),
    .D(_00941_),
    .Q_N(_14542_),
    .Q(\rbzero.spi_registers.spi_done ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.ss_buffer[0]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1312),
    .D(_00942_),
    .Q_N(_14541_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.ss_buffer[1]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1313),
    .D(_00943_),
    .Q_N(_14540_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1314),
    .D(_00944_),
    .Q_N(_14539_),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1315),
    .D(_00945_),
    .Q_N(_00041_),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1316),
    .D(_00946_),
    .Q_N(_00040_),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1317),
    .D(_00947_),
    .Q_N(_00039_),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1318),
    .D(_00948_),
    .Q_N(_00038_),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1319),
    .D(_00949_),
    .Q_N(_00037_),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1320),
    .D(_00950_),
    .Q_N(_00036_),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1321),
    .D(_00951_),
    .Q_N(_00035_),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1322),
    .D(_00952_),
    .Q_N(_00034_),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1323),
    .D(_00953_),
    .Q_N(_00033_),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1324),
    .D(_00954_),
    .Q_N(_00032_),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1325),
    .D(_00955_),
    .Q_N(_14538_),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1326),
    .D(_00956_),
    .Q_N(_00031_),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1327),
    .D(_00957_),
    .Q_N(_00030_),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1328),
    .D(_00958_),
    .Q_N(_00029_),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1329),
    .D(_00959_),
    .Q_N(_14537_),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1330),
    .D(_00960_),
    .Q_N(_14536_),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1331),
    .D(_00961_),
    .Q_N(_14535_),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1332),
    .D(_00962_),
    .Q_N(_14534_),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1333),
    .D(_00963_),
    .Q_N(_14533_),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1334),
    .D(_00964_),
    .Q_N(_00045_),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1335),
    .D(_00965_),
    .Q_N(_00044_),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1336),
    .D(_00966_),
    .Q_N(_00043_),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd0[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1337),
    .D(_00967_),
    .Q_N(_00042_),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1338),
    .D(_00968_),
    .Q_N(_14532_),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1339),
    .D(_00969_),
    .Q_N(_14531_),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1340),
    .D(_00970_),
    .Q_N(_14530_),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1341),
    .D(_00971_),
    .Q_N(_14529_),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1342),
    .D(_00972_),
    .Q_N(_14528_),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1343),
    .D(_00973_),
    .Q_N(_14527_),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1344),
    .D(_00974_),
    .Q_N(_14526_),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1345),
    .D(_00975_),
    .Q_N(_14525_),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1346),
    .D(_00976_),
    .Q_N(_14524_),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1347),
    .D(_00977_),
    .Q_N(_14523_),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1348),
    .D(_00978_),
    .Q_N(_14522_),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1349),
    .D(_00979_),
    .Q_N(_14521_),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1350),
    .D(_00980_),
    .Q_N(_14520_),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1351),
    .D(_00981_),
    .Q_N(_14519_),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1352),
    .D(_00982_),
    .Q_N(_14518_),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1353),
    .D(_00983_),
    .Q_N(_14517_),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1354),
    .D(_00984_),
    .Q_N(_14516_),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1355),
    .D(_00985_),
    .Q_N(_14515_),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1356),
    .D(_00986_),
    .Q_N(_14514_),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1357),
    .D(_00987_),
    .Q_N(_14513_),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1358),
    .D(_00988_),
    .Q_N(_14512_),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1359),
    .D(_00989_),
    .Q_N(_14511_),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1360),
    .D(_00990_),
    .Q_N(_14510_),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1361),
    .D(_00991_),
    .Q_N(_14509_),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1362),
    .D(_00992_),
    .Q_N(_14508_),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1363),
    .D(_00993_),
    .Q_N(_14507_),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1364),
    .D(_00994_),
    .Q_N(_14506_),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1365),
    .D(_00995_),
    .Q_N(_14505_),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1366),
    .D(_00996_),
    .Q_N(_14504_),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1367),
    .D(_00997_),
    .Q_N(_14503_),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1368),
    .D(_00998_),
    .Q_N(_14502_),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1369),
    .D(_00999_),
    .Q_N(_14501_),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1370),
    .D(_01000_),
    .Q_N(_14500_),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1371),
    .D(_01001_),
    .Q_N(_14499_),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1372),
    .D(_01002_),
    .Q_N(_14498_),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1373),
    .D(_01003_),
    .Q_N(_14497_),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1374),
    .D(_01004_),
    .Q_N(_14496_),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1375),
    .D(_01005_),
    .Q_N(_14495_),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1376),
    .D(_01006_),
    .Q_N(_14494_),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1377),
    .D(_01007_),
    .Q_N(_14493_),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1378),
    .D(_01008_),
    .Q_N(_14492_),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1379),
    .D(_01009_),
    .Q_N(_14491_),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1380),
    .D(_01010_),
    .Q_N(_14490_),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1381),
    .D(_01011_),
    .Q_N(_14489_),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1382),
    .D(_01012_),
    .Q_N(_14488_),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1383),
    .D(_01013_),
    .Q_N(_14487_),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1384),
    .D(_01014_),
    .Q_N(_14486_),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1385),
    .D(_01015_),
    .Q_N(_14485_),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1386),
    .D(_01016_),
    .Q_N(_14484_),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1387),
    .D(_01017_),
    .Q_N(_14483_),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1388),
    .D(_01018_),
    .Q_N(_14482_),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1389),
    .D(_01019_),
    .Q_N(_14481_),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1390),
    .D(_01020_),
    .Q_N(_14480_),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1391),
    .D(_01021_),
    .Q_N(_14479_),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1392),
    .D(_01022_),
    .Q_N(_14478_),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1393),
    .D(_01023_),
    .Q_N(_14477_),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1394),
    .D(_01024_),
    .Q_N(_14476_),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1395),
    .D(_01025_),
    .Q_N(_14475_),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1396),
    .D(_01026_),
    .Q_N(_14474_),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1397),
    .D(_01027_),
    .Q_N(_14473_),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1398),
    .D(_01028_),
    .Q_N(_14472_),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1399),
    .D(_01029_),
    .Q_N(_14471_),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1400),
    .D(_01030_),
    .Q_N(_14470_),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1401),
    .D(_01031_),
    .Q_N(_14469_),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1402),
    .D(_01032_),
    .Q_N(_14468_),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1403),
    .D(_01033_),
    .Q_N(_14467_),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1404),
    .D(_01034_),
    .Q_N(_14466_),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1405),
    .D(_01035_),
    .Q_N(_14465_),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1406),
    .D(_01036_),
    .Q_N(_14464_),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1407),
    .D(_01037_),
    .Q_N(_14463_),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1408),
    .D(_01038_),
    .Q_N(_14462_),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.texadd3[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1409),
    .D(_01039_),
    .Q_N(_14461_),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vinf$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1410),
    .D(_01040_),
    .Q_N(_00046_),
    .Q(\rbzero.o_vinf ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1411),
    .D(_01041_),
    .Q_N(_14460_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1412),
    .D(_01042_),
    .Q_N(_14459_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1413),
    .D(_01043_),
    .Q_N(_14458_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1414),
    .D(_01044_),
    .Q_N(_14457_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1415),
    .D(_01045_),
    .Q_N(_14456_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sg13g2_dfrbp_1 \rbzero.spi_registers.vshift[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1416),
    .D(_01046_),
    .Q_N(_14455_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sg13g2_dfrbp_1 \rbzero.texV[0]$_SDFF_PP0_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1417),
    .D(_01047_),
    .Q_N(_14454_),
    .Q(\rbzero.texV[-11] ));
 sg13g2_dfrbp_1 \rbzero.texV[10]$_SDFF_PP0_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1418),
    .D(_01048_),
    .Q_N(_14453_),
    .Q(\rbzero.texV[-1] ));
 sg13g2_dfrbp_1 \rbzero.texV[11]$_SDFF_PP0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1419),
    .D(_01049_),
    .Q_N(_14452_),
    .Q(\rbzero.texV[0] ));
 sg13g2_dfrbp_1 \rbzero.texV[12]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1420),
    .D(_01050_),
    .Q_N(_14451_),
    .Q(\rbzero.texV[1] ));
 sg13g2_dfrbp_1 \rbzero.texV[13]$_SDFF_PP0_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1421),
    .D(_01051_),
    .Q_N(_14450_),
    .Q(\rbzero.texV[2] ));
 sg13g2_dfrbp_1 \rbzero.texV[14]$_SDFF_PP0_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1422),
    .D(_01052_),
    .Q_N(_14449_),
    .Q(\rbzero.texV[3] ));
 sg13g2_dfrbp_1 \rbzero.texV[15]$_SDFF_PP0_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1423),
    .D(_01053_),
    .Q_N(_14448_),
    .Q(\rbzero.texV[4] ));
 sg13g2_dfrbp_1 \rbzero.texV[16]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1424),
    .D(_01054_),
    .Q_N(_14447_),
    .Q(\rbzero.texV[5] ));
 sg13g2_dfrbp_1 \rbzero.texV[17]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1425),
    .D(_01055_),
    .Q_N(_14446_),
    .Q(\rbzero.texV[6] ));
 sg13g2_dfrbp_1 \rbzero.texV[18]$_SDFF_PP0_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1426),
    .D(_01056_),
    .Q_N(_14445_),
    .Q(\rbzero.texV[7] ));
 sg13g2_dfrbp_1 \rbzero.texV[19]$_SDFF_PP0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1427),
    .D(_01057_),
    .Q_N(_14444_),
    .Q(\rbzero.texV[8] ));
 sg13g2_dfrbp_1 \rbzero.texV[1]$_SDFF_PP0_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1428),
    .D(_01058_),
    .Q_N(_14443_),
    .Q(\rbzero.texV[-10] ));
 sg13g2_dfrbp_1 \rbzero.texV[20]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1429),
    .D(_01059_),
    .Q_N(_14442_),
    .Q(\rbzero.texV[9] ));
 sg13g2_dfrbp_1 \rbzero.texV[21]$_SDFF_PP0_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1430),
    .D(_01060_),
    .Q_N(_14441_),
    .Q(\rbzero.texV[10] ));
 sg13g2_dfrbp_1 \rbzero.texV[2]$_SDFF_PP0_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1431),
    .D(_01061_),
    .Q_N(_14440_),
    .Q(\rbzero.texV[-9] ));
 sg13g2_dfrbp_1 \rbzero.texV[3]$_SDFF_PP0_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1432),
    .D(_01062_),
    .Q_N(_14439_),
    .Q(\rbzero.texV[-8] ));
 sg13g2_dfrbp_1 \rbzero.texV[4]$_SDFF_PP0_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1433),
    .D(_01063_),
    .Q_N(_14438_),
    .Q(\rbzero.texV[-7] ));
 sg13g2_dfrbp_1 \rbzero.texV[5]$_SDFF_PP0_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1434),
    .D(_01064_),
    .Q_N(_14437_),
    .Q(\rbzero.texV[-6] ));
 sg13g2_dfrbp_1 \rbzero.texV[6]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1435),
    .D(_01065_),
    .Q_N(_14436_),
    .Q(\rbzero.texV[-5] ));
 sg13g2_dfrbp_1 \rbzero.texV[7]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1436),
    .D(_01066_),
    .Q_N(_14435_),
    .Q(\rbzero.texV[-4] ));
 sg13g2_dfrbp_1 \rbzero.texV[8]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1437),
    .D(_01067_),
    .Q_N(_14434_),
    .Q(\rbzero.texV[-3] ));
 sg13g2_dfrbp_1 \rbzero.texV[9]$_SDFF_PP0_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1438),
    .D(_01068_),
    .Q_N(_14433_),
    .Q(\rbzero.texV[-2] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[0]$_DFFE_NP_  (.CLK(net2585),
    .RESET_B(net1439),
    .D(_01069_),
    .Q_N(_00329_),
    .Q(\rbzero.tex_b0[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[10]$_DFFE_NP_  (.CLK(net2584),
    .RESET_B(net1440),
    .D(_01070_),
    .Q_N(_00339_),
    .Q(\rbzero.tex_b0[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[11]$_DFFE_NP_  (.CLK(net2583),
    .RESET_B(net1441),
    .D(_01071_),
    .Q_N(_00340_),
    .Q(\rbzero.tex_b0[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[12]$_DFFE_NP_  (.CLK(net2582),
    .RESET_B(net1442),
    .D(_01072_),
    .Q_N(_00341_),
    .Q(\rbzero.tex_b0[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[13]$_DFFE_NP_  (.CLK(net2581),
    .RESET_B(net1443),
    .D(_01073_),
    .Q_N(_00342_),
    .Q(\rbzero.tex_b0[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[14]$_DFFE_NP_  (.CLK(net2580),
    .RESET_B(net1444),
    .D(_01074_),
    .Q_N(_00343_),
    .Q(\rbzero.tex_b0[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[15]$_DFFE_NP_  (.CLK(net2579),
    .RESET_B(net1445),
    .D(_01075_),
    .Q_N(_00344_),
    .Q(\rbzero.tex_b0[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[16]$_DFFE_NP_  (.CLK(net2578),
    .RESET_B(net1446),
    .D(_01076_),
    .Q_N(_00345_),
    .Q(\rbzero.tex_b0[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[17]$_DFFE_NP_  (.CLK(net2577),
    .RESET_B(net1447),
    .D(_01077_),
    .Q_N(_00346_),
    .Q(\rbzero.tex_b0[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[18]$_DFFE_NP_  (.CLK(net2576),
    .RESET_B(net1448),
    .D(_01078_),
    .Q_N(_00347_),
    .Q(\rbzero.tex_b0[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[19]$_DFFE_NP_  (.CLK(net2575),
    .RESET_B(net1449),
    .D(_01079_),
    .Q_N(_00348_),
    .Q(\rbzero.tex_b0[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[1]$_DFFE_NP_  (.CLK(net2574),
    .RESET_B(net1450),
    .D(_01080_),
    .Q_N(_00330_),
    .Q(\rbzero.tex_b0[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[20]$_DFFE_NP_  (.CLK(net2573),
    .RESET_B(net1451),
    .D(_01081_),
    .Q_N(_00349_),
    .Q(\rbzero.tex_b0[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[21]$_DFFE_NP_  (.CLK(net2572),
    .RESET_B(net1452),
    .D(_01082_),
    .Q_N(_00350_),
    .Q(\rbzero.tex_b0[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[22]$_DFFE_NP_  (.CLK(net2571),
    .RESET_B(net1453),
    .D(_01083_),
    .Q_N(_00351_),
    .Q(\rbzero.tex_b0[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[23]$_DFFE_NP_  (.CLK(net2570),
    .RESET_B(net1454),
    .D(_01084_),
    .Q_N(_00352_),
    .Q(\rbzero.tex_b0[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[24]$_DFFE_NP_  (.CLK(net2569),
    .RESET_B(net1455),
    .D(_01085_),
    .Q_N(_00353_),
    .Q(\rbzero.tex_b0[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[25]$_DFFE_NP_  (.CLK(net2568),
    .RESET_B(net1456),
    .D(_01086_),
    .Q_N(_00354_),
    .Q(\rbzero.tex_b0[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[26]$_DFFE_NP_  (.CLK(net2567),
    .RESET_B(net1457),
    .D(_01087_),
    .Q_N(_00355_),
    .Q(\rbzero.tex_b0[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[27]$_DFFE_NP_  (.CLK(net2566),
    .RESET_B(net1458),
    .D(_01088_),
    .Q_N(_00356_),
    .Q(\rbzero.tex_b0[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[28]$_DFFE_NP_  (.CLK(net2565),
    .RESET_B(net1459),
    .D(_01089_),
    .Q_N(_00357_),
    .Q(\rbzero.tex_b0[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[29]$_DFFE_NP_  (.CLK(net2564),
    .RESET_B(net1460),
    .D(_01090_),
    .Q_N(_00358_),
    .Q(\rbzero.tex_b0[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[2]$_DFFE_NP_  (.CLK(net2563),
    .RESET_B(net1461),
    .D(_01091_),
    .Q_N(_00331_),
    .Q(\rbzero.tex_b0[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[30]$_DFFE_NP_  (.CLK(net2562),
    .RESET_B(net1462),
    .D(_01092_),
    .Q_N(_00359_),
    .Q(\rbzero.tex_b0[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[31]$_DFFE_NP_  (.CLK(net2561),
    .RESET_B(net1463),
    .D(_01093_),
    .Q_N(_00360_),
    .Q(\rbzero.tex_b0[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[32]$_DFFE_NP_  (.CLK(net2560),
    .RESET_B(net1464),
    .D(_01094_),
    .Q_N(_00361_),
    .Q(\rbzero.tex_b0[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[33]$_DFFE_NP_  (.CLK(net2559),
    .RESET_B(net1465),
    .D(_01095_),
    .Q_N(_00362_),
    .Q(\rbzero.tex_b0[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[34]$_DFFE_NP_  (.CLK(net2558),
    .RESET_B(net1466),
    .D(_01096_),
    .Q_N(_00363_),
    .Q(\rbzero.tex_b0[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[35]$_DFFE_NP_  (.CLK(net2557),
    .RESET_B(net1467),
    .D(_01097_),
    .Q_N(_00364_),
    .Q(\rbzero.tex_b0[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[36]$_DFFE_NP_  (.CLK(net2556),
    .RESET_B(net1468),
    .D(_01098_),
    .Q_N(_00365_),
    .Q(\rbzero.tex_b0[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[37]$_DFFE_NP_  (.CLK(net2555),
    .RESET_B(net1469),
    .D(_01099_),
    .Q_N(_00366_),
    .Q(\rbzero.tex_b0[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[38]$_DFFE_NP_  (.CLK(net2554),
    .RESET_B(net1470),
    .D(_01100_),
    .Q_N(_00367_),
    .Q(\rbzero.tex_b0[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[39]$_DFFE_NP_  (.CLK(net2553),
    .RESET_B(net1471),
    .D(_01101_),
    .Q_N(_00368_),
    .Q(\rbzero.tex_b0[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[3]$_DFFE_NP_  (.CLK(net2552),
    .RESET_B(net1472),
    .D(_01102_),
    .Q_N(_00332_),
    .Q(\rbzero.tex_b0[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[40]$_DFFE_NP_  (.CLK(net2551),
    .RESET_B(net1473),
    .D(_01103_),
    .Q_N(_00369_),
    .Q(\rbzero.tex_b0[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[41]$_DFFE_NP_  (.CLK(net2550),
    .RESET_B(net1474),
    .D(_01104_),
    .Q_N(_00370_),
    .Q(\rbzero.tex_b0[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[42]$_DFFE_NP_  (.CLK(net2549),
    .RESET_B(net1475),
    .D(_01105_),
    .Q_N(_00371_),
    .Q(\rbzero.tex_b0[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[43]$_DFFE_NP_  (.CLK(net2548),
    .RESET_B(net1476),
    .D(_01106_),
    .Q_N(_00372_),
    .Q(\rbzero.tex_b0[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[44]$_DFFE_NP_  (.CLK(net2547),
    .RESET_B(net1477),
    .D(_01107_),
    .Q_N(_00373_),
    .Q(\rbzero.tex_b0[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[45]$_DFFE_NP_  (.CLK(net2546),
    .RESET_B(net1478),
    .D(_01108_),
    .Q_N(_00374_),
    .Q(\rbzero.tex_b0[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[46]$_DFFE_NP_  (.CLK(net2545),
    .RESET_B(net1479),
    .D(_01109_),
    .Q_N(_00375_),
    .Q(\rbzero.tex_b0[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[47]$_DFFE_NP_  (.CLK(net2544),
    .RESET_B(net1480),
    .D(_01110_),
    .Q_N(_00376_),
    .Q(\rbzero.tex_b0[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[48]$_DFFE_NP_  (.CLK(net2543),
    .RESET_B(net1481),
    .D(_01111_),
    .Q_N(_00377_),
    .Q(\rbzero.tex_b0[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[49]$_DFFE_NP_  (.CLK(net2542),
    .RESET_B(net1482),
    .D(_01112_),
    .Q_N(_00378_),
    .Q(\rbzero.tex_b0[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[4]$_DFFE_NP_  (.CLK(net2541),
    .RESET_B(net1483),
    .D(_01113_),
    .Q_N(_00333_),
    .Q(\rbzero.tex_b0[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[50]$_DFFE_NP_  (.CLK(net2540),
    .RESET_B(net1484),
    .D(_01114_),
    .Q_N(_00379_),
    .Q(\rbzero.tex_b0[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[51]$_DFFE_NP_  (.CLK(net2539),
    .RESET_B(net1485),
    .D(_01115_),
    .Q_N(_00380_),
    .Q(\rbzero.tex_b0[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[52]$_DFFE_NP_  (.CLK(net2538),
    .RESET_B(net1486),
    .D(_01116_),
    .Q_N(_00381_),
    .Q(\rbzero.tex_b0[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[53]$_DFFE_NP_  (.CLK(net2537),
    .RESET_B(net1487),
    .D(_01117_),
    .Q_N(_00382_),
    .Q(\rbzero.tex_b0[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[54]$_DFFE_NP_  (.CLK(net2536),
    .RESET_B(net1488),
    .D(_01118_),
    .Q_N(_00383_),
    .Q(\rbzero.tex_b0[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[55]$_DFFE_NP_  (.CLK(net2535),
    .RESET_B(net1489),
    .D(_01119_),
    .Q_N(_00384_),
    .Q(\rbzero.tex_b0[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[56]$_DFFE_NP_  (.CLK(net2534),
    .RESET_B(net1490),
    .D(_01120_),
    .Q_N(_00385_),
    .Q(\rbzero.tex_b0[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[57]$_DFFE_NP_  (.CLK(net2533),
    .RESET_B(net1491),
    .D(_01121_),
    .Q_N(_00386_),
    .Q(\rbzero.tex_b0[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[58]$_DFFE_NP_  (.CLK(net2532),
    .RESET_B(net1492),
    .D(_01122_),
    .Q_N(_00387_),
    .Q(\rbzero.tex_b0[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[59]$_DFFE_NP_  (.CLK(net2531),
    .RESET_B(net1493),
    .D(_01123_),
    .Q_N(_00388_),
    .Q(\rbzero.tex_b0[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[5]$_DFFE_NP_  (.CLK(net2530),
    .RESET_B(net1494),
    .D(_01124_),
    .Q_N(_00334_),
    .Q(\rbzero.tex_b0[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[60]$_DFFE_NP_  (.CLK(net2529),
    .RESET_B(net1495),
    .D(_01125_),
    .Q_N(_00389_),
    .Q(\rbzero.tex_b0[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[61]$_DFFE_NP_  (.CLK(net2528),
    .RESET_B(net1496),
    .D(_01126_),
    .Q_N(_00390_),
    .Q(\rbzero.tex_b0[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[62]$_DFFE_NP_  (.CLK(net2527),
    .RESET_B(net1497),
    .D(_01127_),
    .Q_N(_00391_),
    .Q(\rbzero.tex_b0[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[63]$_DFFE_NP_  (.CLK(net2526),
    .RESET_B(net1498),
    .D(_01128_),
    .Q_N(_00392_),
    .Q(\rbzero.tex_b0[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[6]$_DFFE_NP_  (.CLK(net2525),
    .RESET_B(net1499),
    .D(_01129_),
    .Q_N(_00335_),
    .Q(\rbzero.tex_b0[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[7]$_DFFE_NP_  (.CLK(net2524),
    .RESET_B(net1500),
    .D(_01130_),
    .Q_N(_00336_),
    .Q(\rbzero.tex_b0[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[8]$_DFFE_NP_  (.CLK(net2523),
    .RESET_B(net1501),
    .D(_01131_),
    .Q_N(_00337_),
    .Q(\rbzero.tex_b0[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_b0[9]$_DFFE_NP_  (.CLK(net2522),
    .RESET_B(net1502),
    .D(_01132_),
    .Q_N(_00338_),
    .Q(\rbzero.tex_b0[9] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[0]$_DFFE_NP_  (.CLK(net2521),
    .RESET_B(net1503),
    .D(_01133_),
    .Q_N(_00130_),
    .Q(\rbzero.tex_b1[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[10]$_DFFE_NP_  (.CLK(net2520),
    .RESET_B(net1504),
    .D(_01134_),
    .Q_N(_00140_),
    .Q(\rbzero.tex_b1[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[11]$_DFFE_NP_  (.CLK(net2519),
    .RESET_B(net1505),
    .D(_01135_),
    .Q_N(_00141_),
    .Q(\rbzero.tex_b1[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[12]$_DFFE_NP_  (.CLK(net2518),
    .RESET_B(net1506),
    .D(_01136_),
    .Q_N(_00142_),
    .Q(\rbzero.tex_b1[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[13]$_DFFE_NP_  (.CLK(net2517),
    .RESET_B(net1507),
    .D(_01137_),
    .Q_N(_00143_),
    .Q(\rbzero.tex_b1[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[14]$_DFFE_NP_  (.CLK(net2516),
    .RESET_B(net1508),
    .D(_01138_),
    .Q_N(_00144_),
    .Q(\rbzero.tex_b1[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[15]$_DFFE_NP_  (.CLK(net2515),
    .RESET_B(net1509),
    .D(_01139_),
    .Q_N(_00145_),
    .Q(\rbzero.tex_b1[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[16]$_DFFE_NP_  (.CLK(net2514),
    .RESET_B(net1510),
    .D(_01140_),
    .Q_N(_00146_),
    .Q(\rbzero.tex_b1[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[17]$_DFFE_NP_  (.CLK(net2513),
    .RESET_B(net1511),
    .D(_01141_),
    .Q_N(_00147_),
    .Q(\rbzero.tex_b1[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[18]$_DFFE_NP_  (.CLK(net2512),
    .RESET_B(net1512),
    .D(_01142_),
    .Q_N(_00148_),
    .Q(\rbzero.tex_b1[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[19]$_DFFE_NP_  (.CLK(net2511),
    .RESET_B(net1513),
    .D(_01143_),
    .Q_N(_00149_),
    .Q(\rbzero.tex_b1[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[1]$_DFFE_NP_  (.CLK(net2510),
    .RESET_B(net1514),
    .D(_01144_),
    .Q_N(_00131_),
    .Q(\rbzero.tex_b1[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[20]$_DFFE_NP_  (.CLK(net2509),
    .RESET_B(net1515),
    .D(_01145_),
    .Q_N(_00150_),
    .Q(\rbzero.tex_b1[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[21]$_DFFE_NP_  (.CLK(net2508),
    .RESET_B(net1516),
    .D(_01146_),
    .Q_N(_00151_),
    .Q(\rbzero.tex_b1[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[22]$_DFFE_NP_  (.CLK(net2507),
    .RESET_B(net1517),
    .D(_01147_),
    .Q_N(_00152_),
    .Q(\rbzero.tex_b1[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[23]$_DFFE_NP_  (.CLK(net2506),
    .RESET_B(net1518),
    .D(_01148_),
    .Q_N(_00153_),
    .Q(\rbzero.tex_b1[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[24]$_DFFE_NP_  (.CLK(net2505),
    .RESET_B(net1519),
    .D(_01149_),
    .Q_N(_00154_),
    .Q(\rbzero.tex_b1[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[25]$_DFFE_NP_  (.CLK(net2504),
    .RESET_B(net1520),
    .D(_01150_),
    .Q_N(_00155_),
    .Q(\rbzero.tex_b1[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[26]$_DFFE_NP_  (.CLK(net2503),
    .RESET_B(net1521),
    .D(_01151_),
    .Q_N(_00156_),
    .Q(\rbzero.tex_b1[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[27]$_DFFE_NP_  (.CLK(net2502),
    .RESET_B(net1522),
    .D(_01152_),
    .Q_N(_00157_),
    .Q(\rbzero.tex_b1[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[28]$_DFFE_NP_  (.CLK(net2501),
    .RESET_B(net1523),
    .D(_01153_),
    .Q_N(_00158_),
    .Q(\rbzero.tex_b1[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[29]$_DFFE_NP_  (.CLK(net2500),
    .RESET_B(net1524),
    .D(_01154_),
    .Q_N(_00159_),
    .Q(\rbzero.tex_b1[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[2]$_DFFE_NP_  (.CLK(net2499),
    .RESET_B(net1525),
    .D(_01155_),
    .Q_N(_00132_),
    .Q(\rbzero.tex_b1[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[30]$_DFFE_NP_  (.CLK(net2498),
    .RESET_B(net1526),
    .D(_01156_),
    .Q_N(_00160_),
    .Q(\rbzero.tex_b1[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[31]$_DFFE_NP_  (.CLK(net2497),
    .RESET_B(net1527),
    .D(_01157_),
    .Q_N(_00161_),
    .Q(\rbzero.tex_b1[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[32]$_DFFE_NP_  (.CLK(net2496),
    .RESET_B(net1528),
    .D(_01158_),
    .Q_N(_00162_),
    .Q(\rbzero.tex_b1[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[33]$_DFFE_NP_  (.CLK(net2495),
    .RESET_B(net1529),
    .D(_01159_),
    .Q_N(_00163_),
    .Q(\rbzero.tex_b1[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[34]$_DFFE_NP_  (.CLK(net2494),
    .RESET_B(net1530),
    .D(_01160_),
    .Q_N(_00164_),
    .Q(\rbzero.tex_b1[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[35]$_DFFE_NP_  (.CLK(net2493),
    .RESET_B(net1531),
    .D(_01161_),
    .Q_N(_00165_),
    .Q(\rbzero.tex_b1[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[36]$_DFFE_NP_  (.CLK(net2492),
    .RESET_B(net1532),
    .D(_01162_),
    .Q_N(_00166_),
    .Q(\rbzero.tex_b1[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[37]$_DFFE_NP_  (.CLK(net2491),
    .RESET_B(net1533),
    .D(_01163_),
    .Q_N(_00167_),
    .Q(\rbzero.tex_b1[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[38]$_DFFE_NP_  (.CLK(net2490),
    .RESET_B(net1534),
    .D(_01164_),
    .Q_N(_00168_),
    .Q(\rbzero.tex_b1[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[39]$_DFFE_NP_  (.CLK(net2489),
    .RESET_B(net1535),
    .D(_01165_),
    .Q_N(_00169_),
    .Q(\rbzero.tex_b1[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[3]$_DFFE_NP_  (.CLK(net2488),
    .RESET_B(net1536),
    .D(_01166_),
    .Q_N(_00133_),
    .Q(\rbzero.tex_b1[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[40]$_DFFE_NP_  (.CLK(net2487),
    .RESET_B(net1537),
    .D(_01167_),
    .Q_N(_00170_),
    .Q(\rbzero.tex_b1[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[41]$_DFFE_NP_  (.CLK(net2486),
    .RESET_B(net1538),
    .D(_01168_),
    .Q_N(_00171_),
    .Q(\rbzero.tex_b1[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[42]$_DFFE_NP_  (.CLK(net2485),
    .RESET_B(net1539),
    .D(_01169_),
    .Q_N(_00172_),
    .Q(\rbzero.tex_b1[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[43]$_DFFE_NP_  (.CLK(net2484),
    .RESET_B(net1540),
    .D(_01170_),
    .Q_N(_00173_),
    .Q(\rbzero.tex_b1[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[44]$_DFFE_NP_  (.CLK(net2483),
    .RESET_B(net1541),
    .D(_01171_),
    .Q_N(_00174_),
    .Q(\rbzero.tex_b1[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[45]$_DFFE_NP_  (.CLK(net2482),
    .RESET_B(net1542),
    .D(_01172_),
    .Q_N(_00175_),
    .Q(\rbzero.tex_b1[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[46]$_DFFE_NP_  (.CLK(net2481),
    .RESET_B(net1543),
    .D(_01173_),
    .Q_N(_00176_),
    .Q(\rbzero.tex_b1[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[47]$_DFFE_NP_  (.CLK(net2480),
    .RESET_B(net1544),
    .D(_01174_),
    .Q_N(_00177_),
    .Q(\rbzero.tex_b1[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[48]$_DFFE_NP_  (.CLK(net2479),
    .RESET_B(net1545),
    .D(_01175_),
    .Q_N(_00178_),
    .Q(\rbzero.tex_b1[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[49]$_DFFE_NP_  (.CLK(net2478),
    .RESET_B(net1546),
    .D(_01176_),
    .Q_N(_00179_),
    .Q(\rbzero.tex_b1[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[4]$_DFFE_NP_  (.CLK(net2477),
    .RESET_B(net1547),
    .D(_01177_),
    .Q_N(_00134_),
    .Q(\rbzero.tex_b1[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[50]$_DFFE_NP_  (.CLK(net2476),
    .RESET_B(net1548),
    .D(_01178_),
    .Q_N(_00180_),
    .Q(\rbzero.tex_b1[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[51]$_DFFE_NP_  (.CLK(net2475),
    .RESET_B(net1549),
    .D(_01179_),
    .Q_N(_00181_),
    .Q(\rbzero.tex_b1[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[52]$_DFFE_NP_  (.CLK(net2474),
    .RESET_B(net1550),
    .D(_01180_),
    .Q_N(_00182_),
    .Q(\rbzero.tex_b1[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[53]$_DFFE_NP_  (.CLK(net2473),
    .RESET_B(net1551),
    .D(_01181_),
    .Q_N(_00183_),
    .Q(\rbzero.tex_b1[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[54]$_DFFE_NP_  (.CLK(net2472),
    .RESET_B(net1552),
    .D(_01182_),
    .Q_N(_00184_),
    .Q(\rbzero.tex_b1[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[55]$_DFFE_NP_  (.CLK(net2471),
    .RESET_B(net1553),
    .D(_01183_),
    .Q_N(_00185_),
    .Q(\rbzero.tex_b1[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[56]$_DFFE_NP_  (.CLK(net2470),
    .RESET_B(net1554),
    .D(_01184_),
    .Q_N(_00186_),
    .Q(\rbzero.tex_b1[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[57]$_DFFE_NP_  (.CLK(net2469),
    .RESET_B(net1555),
    .D(_01185_),
    .Q_N(_00187_),
    .Q(\rbzero.tex_b1[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[58]$_DFFE_NP_  (.CLK(net2468),
    .RESET_B(net1556),
    .D(_01186_),
    .Q_N(_00188_),
    .Q(\rbzero.tex_b1[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[59]$_DFFE_NP_  (.CLK(net2467),
    .RESET_B(net1557),
    .D(_01187_),
    .Q_N(_00189_),
    .Q(\rbzero.tex_b1[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[5]$_DFFE_NP_  (.CLK(net2466),
    .RESET_B(net1558),
    .D(_01188_),
    .Q_N(_00135_),
    .Q(\rbzero.tex_b1[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[60]$_DFFE_NP_  (.CLK(net2465),
    .RESET_B(net1559),
    .D(_01189_),
    .Q_N(_00190_),
    .Q(\rbzero.tex_b1[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[61]$_DFFE_NP_  (.CLK(net2464),
    .RESET_B(net1560),
    .D(_01190_),
    .Q_N(_00191_),
    .Q(\rbzero.tex_b1[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[62]$_DFFE_NP_  (.CLK(net2463),
    .RESET_B(net1561),
    .D(_01191_),
    .Q_N(_00192_),
    .Q(\rbzero.tex_b1[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[63]$_DFFE_NP_  (.CLK(net2462),
    .RESET_B(net1562),
    .D(_01192_),
    .Q_N(_00193_),
    .Q(\rbzero.tex_b1[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[6]$_DFFE_NP_  (.CLK(net2461),
    .RESET_B(net1563),
    .D(_01193_),
    .Q_N(_00136_),
    .Q(\rbzero.tex_b1[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[7]$_DFFE_NP_  (.CLK(net2460),
    .RESET_B(net1564),
    .D(_01194_),
    .Q_N(_00137_),
    .Q(\rbzero.tex_b1[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[8]$_DFFE_NP_  (.CLK(net2459),
    .RESET_B(net1565),
    .D(_01195_),
    .Q_N(_00138_),
    .Q(\rbzero.tex_b1[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_b1[9]$_DFFE_NP_  (.CLK(net2458),
    .RESET_B(net1566),
    .D(_01196_),
    .Q_N(_00139_),
    .Q(\rbzero.tex_b1[9] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[0]$_DFFE_NP_  (.CLK(net2457),
    .RESET_B(net1567),
    .D(_01197_),
    .Q_N(_00263_),
    .Q(\rbzero.tex_g0[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[10]$_DFFE_NP_  (.CLK(net2456),
    .RESET_B(net1568),
    .D(_01198_),
    .Q_N(_00273_),
    .Q(\rbzero.tex_g0[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[11]$_DFFE_NP_  (.CLK(net2455),
    .RESET_B(net1569),
    .D(_01199_),
    .Q_N(_00274_),
    .Q(\rbzero.tex_g0[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[12]$_DFFE_NP_  (.CLK(net2454),
    .RESET_B(net1570),
    .D(_01200_),
    .Q_N(_00275_),
    .Q(\rbzero.tex_g0[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[13]$_DFFE_NP_  (.CLK(net2453),
    .RESET_B(net1571),
    .D(_01201_),
    .Q_N(_00276_),
    .Q(\rbzero.tex_g0[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[14]$_DFFE_NP_  (.CLK(net2452),
    .RESET_B(net1572),
    .D(_01202_),
    .Q_N(_00277_),
    .Q(\rbzero.tex_g0[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[15]$_DFFE_NP_  (.CLK(net2451),
    .RESET_B(net1573),
    .D(_01203_),
    .Q_N(_00278_),
    .Q(\rbzero.tex_g0[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[16]$_DFFE_NP_  (.CLK(net2450),
    .RESET_B(net1574),
    .D(_01204_),
    .Q_N(_00279_),
    .Q(\rbzero.tex_g0[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[17]$_DFFE_NP_  (.CLK(net2449),
    .RESET_B(net1575),
    .D(_01205_),
    .Q_N(_00280_),
    .Q(\rbzero.tex_g0[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[18]$_DFFE_NP_  (.CLK(net2448),
    .RESET_B(net1576),
    .D(_01206_),
    .Q_N(_00281_),
    .Q(\rbzero.tex_g0[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[19]$_DFFE_NP_  (.CLK(net2447),
    .RESET_B(net1577),
    .D(_01207_),
    .Q_N(_00282_),
    .Q(\rbzero.tex_g0[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[1]$_DFFE_NP_  (.CLK(net2446),
    .RESET_B(net1578),
    .D(_01208_),
    .Q_N(_00264_),
    .Q(\rbzero.tex_g0[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[20]$_DFFE_NP_  (.CLK(net2445),
    .RESET_B(net1579),
    .D(_01209_),
    .Q_N(_00283_),
    .Q(\rbzero.tex_g0[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[21]$_DFFE_NP_  (.CLK(net2444),
    .RESET_B(net1580),
    .D(_01210_),
    .Q_N(_00284_),
    .Q(\rbzero.tex_g0[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[22]$_DFFE_NP_  (.CLK(net2443),
    .RESET_B(net1581),
    .D(_01211_),
    .Q_N(_00285_),
    .Q(\rbzero.tex_g0[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[23]$_DFFE_NP_  (.CLK(net2442),
    .RESET_B(net1582),
    .D(_01212_),
    .Q_N(_00286_),
    .Q(\rbzero.tex_g0[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[24]$_DFFE_NP_  (.CLK(net2441),
    .RESET_B(net1583),
    .D(_01213_),
    .Q_N(_00287_),
    .Q(\rbzero.tex_g0[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[25]$_DFFE_NP_  (.CLK(net2440),
    .RESET_B(net1584),
    .D(_01214_),
    .Q_N(_00288_),
    .Q(\rbzero.tex_g0[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[26]$_DFFE_NP_  (.CLK(net2439),
    .RESET_B(net1585),
    .D(_01215_),
    .Q_N(_00289_),
    .Q(\rbzero.tex_g0[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[27]$_DFFE_NP_  (.CLK(net2438),
    .RESET_B(net1586),
    .D(_01216_),
    .Q_N(_00290_),
    .Q(\rbzero.tex_g0[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[28]$_DFFE_NP_  (.CLK(net2437),
    .RESET_B(net1587),
    .D(_01217_),
    .Q_N(_00291_),
    .Q(\rbzero.tex_g0[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[29]$_DFFE_NP_  (.CLK(net2436),
    .RESET_B(net1588),
    .D(_01218_),
    .Q_N(_00292_),
    .Q(\rbzero.tex_g0[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[2]$_DFFE_NP_  (.CLK(net2435),
    .RESET_B(net1589),
    .D(_01219_),
    .Q_N(_00265_),
    .Q(\rbzero.tex_g0[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[30]$_DFFE_NP_  (.CLK(net2434),
    .RESET_B(net1590),
    .D(_01220_),
    .Q_N(_00293_),
    .Q(\rbzero.tex_g0[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[31]$_DFFE_NP_  (.CLK(net2433),
    .RESET_B(net1591),
    .D(_01221_),
    .Q_N(_00294_),
    .Q(\rbzero.tex_g0[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[32]$_DFFE_NP_  (.CLK(net2432),
    .RESET_B(net1592),
    .D(_01222_),
    .Q_N(_00295_),
    .Q(\rbzero.tex_g0[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[33]$_DFFE_NP_  (.CLK(net2431),
    .RESET_B(net1593),
    .D(_01223_),
    .Q_N(_00296_),
    .Q(\rbzero.tex_g0[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[34]$_DFFE_NP_  (.CLK(net2430),
    .RESET_B(net1594),
    .D(_01224_),
    .Q_N(_00297_),
    .Q(\rbzero.tex_g0[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[35]$_DFFE_NP_  (.CLK(net2429),
    .RESET_B(net1595),
    .D(_01225_),
    .Q_N(_00298_),
    .Q(\rbzero.tex_g0[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[36]$_DFFE_NP_  (.CLK(net2428),
    .RESET_B(net1596),
    .D(_01226_),
    .Q_N(_00299_),
    .Q(\rbzero.tex_g0[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[37]$_DFFE_NP_  (.CLK(net2427),
    .RESET_B(net1597),
    .D(_01227_),
    .Q_N(_00300_),
    .Q(\rbzero.tex_g0[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[38]$_DFFE_NP_  (.CLK(net2426),
    .RESET_B(net1598),
    .D(_01228_),
    .Q_N(_00301_),
    .Q(\rbzero.tex_g0[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[39]$_DFFE_NP_  (.CLK(net2425),
    .RESET_B(net1599),
    .D(_01229_),
    .Q_N(_00302_),
    .Q(\rbzero.tex_g0[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[3]$_DFFE_NP_  (.CLK(net2424),
    .RESET_B(net1600),
    .D(_01230_),
    .Q_N(_00266_),
    .Q(\rbzero.tex_g0[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[40]$_DFFE_NP_  (.CLK(net2423),
    .RESET_B(net1601),
    .D(_01231_),
    .Q_N(_00303_),
    .Q(\rbzero.tex_g0[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[41]$_DFFE_NP_  (.CLK(net2422),
    .RESET_B(net1602),
    .D(_01232_),
    .Q_N(_00304_),
    .Q(\rbzero.tex_g0[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[42]$_DFFE_NP_  (.CLK(net2421),
    .RESET_B(net1603),
    .D(_01233_),
    .Q_N(_00305_),
    .Q(\rbzero.tex_g0[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[43]$_DFFE_NP_  (.CLK(net2420),
    .RESET_B(net1604),
    .D(_01234_),
    .Q_N(_00306_),
    .Q(\rbzero.tex_g0[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[44]$_DFFE_NP_  (.CLK(net2419),
    .RESET_B(net1605),
    .D(_01235_),
    .Q_N(_00307_),
    .Q(\rbzero.tex_g0[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[45]$_DFFE_NP_  (.CLK(net2418),
    .RESET_B(net1606),
    .D(_01236_),
    .Q_N(_00308_),
    .Q(\rbzero.tex_g0[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[46]$_DFFE_NP_  (.CLK(net2417),
    .RESET_B(net1607),
    .D(_01237_),
    .Q_N(_00309_),
    .Q(\rbzero.tex_g0[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[47]$_DFFE_NP_  (.CLK(net2416),
    .RESET_B(net1608),
    .D(_01238_),
    .Q_N(_00310_),
    .Q(\rbzero.tex_g0[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[48]$_DFFE_NP_  (.CLK(net2415),
    .RESET_B(net1609),
    .D(_01239_),
    .Q_N(_00311_),
    .Q(\rbzero.tex_g0[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[49]$_DFFE_NP_  (.CLK(net2414),
    .RESET_B(net1610),
    .D(_01240_),
    .Q_N(_00312_),
    .Q(\rbzero.tex_g0[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[4]$_DFFE_NP_  (.CLK(net2413),
    .RESET_B(net1611),
    .D(_01241_),
    .Q_N(_00267_),
    .Q(\rbzero.tex_g0[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[50]$_DFFE_NP_  (.CLK(net2412),
    .RESET_B(net1612),
    .D(_01242_),
    .Q_N(_00313_),
    .Q(\rbzero.tex_g0[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[51]$_DFFE_NP_  (.CLK(net2411),
    .RESET_B(net1613),
    .D(_01243_),
    .Q_N(_00314_),
    .Q(\rbzero.tex_g0[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[52]$_DFFE_NP_  (.CLK(net2410),
    .RESET_B(net1614),
    .D(_01244_),
    .Q_N(_00315_),
    .Q(\rbzero.tex_g0[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[53]$_DFFE_NP_  (.CLK(net2409),
    .RESET_B(net1615),
    .D(_01245_),
    .Q_N(_00316_),
    .Q(\rbzero.tex_g0[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[54]$_DFFE_NP_  (.CLK(net2408),
    .RESET_B(net1616),
    .D(_01246_),
    .Q_N(_00317_),
    .Q(\rbzero.tex_g0[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[55]$_DFFE_NP_  (.CLK(net2407),
    .RESET_B(net1617),
    .D(_01247_),
    .Q_N(_00318_),
    .Q(\rbzero.tex_g0[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[56]$_DFFE_NP_  (.CLK(net2406),
    .RESET_B(net1618),
    .D(_01248_),
    .Q_N(_00319_),
    .Q(\rbzero.tex_g0[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[57]$_DFFE_NP_  (.CLK(net2405),
    .RESET_B(net1619),
    .D(_01249_),
    .Q_N(_00320_),
    .Q(\rbzero.tex_g0[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[58]$_DFFE_NP_  (.CLK(net2404),
    .RESET_B(net1620),
    .D(_01250_),
    .Q_N(_00321_),
    .Q(\rbzero.tex_g0[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[59]$_DFFE_NP_  (.CLK(net2403),
    .RESET_B(net1621),
    .D(_01251_),
    .Q_N(_00322_),
    .Q(\rbzero.tex_g0[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[5]$_DFFE_NP_  (.CLK(net2402),
    .RESET_B(net1622),
    .D(_01252_),
    .Q_N(_00268_),
    .Q(\rbzero.tex_g0[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[60]$_DFFE_NP_  (.CLK(net2401),
    .RESET_B(net1623),
    .D(_01253_),
    .Q_N(_00323_),
    .Q(\rbzero.tex_g0[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[61]$_DFFE_NP_  (.CLK(net2400),
    .RESET_B(net1624),
    .D(_01254_),
    .Q_N(_00324_),
    .Q(\rbzero.tex_g0[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[62]$_DFFE_NP_  (.CLK(net2399),
    .RESET_B(net1625),
    .D(_01255_),
    .Q_N(_00325_),
    .Q(\rbzero.tex_g0[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[63]$_DFFE_NP_  (.CLK(net2398),
    .RESET_B(net1626),
    .D(_01256_),
    .Q_N(_00326_),
    .Q(\rbzero.tex_g0[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[6]$_DFFE_NP_  (.CLK(net2397),
    .RESET_B(net1627),
    .D(_01257_),
    .Q_N(_00269_),
    .Q(\rbzero.tex_g0[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[7]$_DFFE_NP_  (.CLK(net2396),
    .RESET_B(net1628),
    .D(_01258_),
    .Q_N(_00270_),
    .Q(\rbzero.tex_g0[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[8]$_DFFE_NP_  (.CLK(net2395),
    .RESET_B(net1629),
    .D(_01259_),
    .Q_N(_00271_),
    .Q(\rbzero.tex_g0[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_g0[9]$_DFFE_NP_  (.CLK(net2394),
    .RESET_B(net1630),
    .D(_01260_),
    .Q_N(_00272_),
    .Q(\rbzero.tex_g0[9] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[0]$_DFFE_NP_  (.CLK(net2393),
    .RESET_B(net1631),
    .D(_01261_),
    .Q_N(_00064_),
    .Q(\rbzero.tex_g1[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[10]$_DFFE_NP_  (.CLK(net2392),
    .RESET_B(net1632),
    .D(_01262_),
    .Q_N(_00074_),
    .Q(\rbzero.tex_g1[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[11]$_DFFE_NP_  (.CLK(net2391),
    .RESET_B(net1633),
    .D(_01263_),
    .Q_N(_00075_),
    .Q(\rbzero.tex_g1[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[12]$_DFFE_NP_  (.CLK(net2390),
    .RESET_B(net1634),
    .D(_01264_),
    .Q_N(_00076_),
    .Q(\rbzero.tex_g1[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[13]$_DFFE_NP_  (.CLK(net2389),
    .RESET_B(net1635),
    .D(_01265_),
    .Q_N(_00077_),
    .Q(\rbzero.tex_g1[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[14]$_DFFE_NP_  (.CLK(net2388),
    .RESET_B(net1636),
    .D(_01266_),
    .Q_N(_00078_),
    .Q(\rbzero.tex_g1[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[15]$_DFFE_NP_  (.CLK(net2387),
    .RESET_B(net1637),
    .D(_01267_),
    .Q_N(_00079_),
    .Q(\rbzero.tex_g1[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[16]$_DFFE_NP_  (.CLK(net2386),
    .RESET_B(net1638),
    .D(_01268_),
    .Q_N(_00080_),
    .Q(\rbzero.tex_g1[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[17]$_DFFE_NP_  (.CLK(net2385),
    .RESET_B(net1639),
    .D(_01269_),
    .Q_N(_00081_),
    .Q(\rbzero.tex_g1[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[18]$_DFFE_NP_  (.CLK(net2384),
    .RESET_B(net1640),
    .D(_01270_),
    .Q_N(_00082_),
    .Q(\rbzero.tex_g1[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[19]$_DFFE_NP_  (.CLK(net2383),
    .RESET_B(net1641),
    .D(_01271_),
    .Q_N(_00083_),
    .Q(\rbzero.tex_g1[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[1]$_DFFE_NP_  (.CLK(net2382),
    .RESET_B(net1642),
    .D(_01272_),
    .Q_N(_00065_),
    .Q(\rbzero.tex_g1[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[20]$_DFFE_NP_  (.CLK(net2381),
    .RESET_B(net1643),
    .D(_01273_),
    .Q_N(_00084_),
    .Q(\rbzero.tex_g1[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[21]$_DFFE_NP_  (.CLK(net2380),
    .RESET_B(net1644),
    .D(_01274_),
    .Q_N(_00085_),
    .Q(\rbzero.tex_g1[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[22]$_DFFE_NP_  (.CLK(net2379),
    .RESET_B(net1645),
    .D(_01275_),
    .Q_N(_00086_),
    .Q(\rbzero.tex_g1[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[23]$_DFFE_NP_  (.CLK(net2378),
    .RESET_B(net1646),
    .D(_01276_),
    .Q_N(_00087_),
    .Q(\rbzero.tex_g1[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[24]$_DFFE_NP_  (.CLK(net2377),
    .RESET_B(net1647),
    .D(_01277_),
    .Q_N(_00088_),
    .Q(\rbzero.tex_g1[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[25]$_DFFE_NP_  (.CLK(net2376),
    .RESET_B(net1648),
    .D(_01278_),
    .Q_N(_00089_),
    .Q(\rbzero.tex_g1[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[26]$_DFFE_NP_  (.CLK(net2375),
    .RESET_B(net1649),
    .D(_01279_),
    .Q_N(_00090_),
    .Q(\rbzero.tex_g1[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[27]$_DFFE_NP_  (.CLK(net2374),
    .RESET_B(net1650),
    .D(_01280_),
    .Q_N(_00091_),
    .Q(\rbzero.tex_g1[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[28]$_DFFE_NP_  (.CLK(net2373),
    .RESET_B(net1651),
    .D(_01281_),
    .Q_N(_00092_),
    .Q(\rbzero.tex_g1[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[29]$_DFFE_NP_  (.CLK(net2372),
    .RESET_B(net1652),
    .D(_01282_),
    .Q_N(_00093_),
    .Q(\rbzero.tex_g1[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[2]$_DFFE_NP_  (.CLK(net2371),
    .RESET_B(net1653),
    .D(_01283_),
    .Q_N(_00066_),
    .Q(\rbzero.tex_g1[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[30]$_DFFE_NP_  (.CLK(net2370),
    .RESET_B(net1654),
    .D(_01284_),
    .Q_N(_00094_),
    .Q(\rbzero.tex_g1[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[31]$_DFFE_NP_  (.CLK(net2369),
    .RESET_B(net1655),
    .D(_01285_),
    .Q_N(_00095_),
    .Q(\rbzero.tex_g1[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[32]$_DFFE_NP_  (.CLK(net2368),
    .RESET_B(net1656),
    .D(_01286_),
    .Q_N(_00096_),
    .Q(\rbzero.tex_g1[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[33]$_DFFE_NP_  (.CLK(net2367),
    .RESET_B(net1657),
    .D(_01287_),
    .Q_N(_00097_),
    .Q(\rbzero.tex_g1[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[34]$_DFFE_NP_  (.CLK(net2366),
    .RESET_B(net1658),
    .D(_01288_),
    .Q_N(_00098_),
    .Q(\rbzero.tex_g1[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[35]$_DFFE_NP_  (.CLK(net2365),
    .RESET_B(net1659),
    .D(_01289_),
    .Q_N(_00099_),
    .Q(\rbzero.tex_g1[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[36]$_DFFE_NP_  (.CLK(net2364),
    .RESET_B(net1660),
    .D(_01290_),
    .Q_N(_00100_),
    .Q(\rbzero.tex_g1[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[37]$_DFFE_NP_  (.CLK(net2363),
    .RESET_B(net1661),
    .D(_01291_),
    .Q_N(_00101_),
    .Q(\rbzero.tex_g1[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[38]$_DFFE_NP_  (.CLK(net2362),
    .RESET_B(net1662),
    .D(_01292_),
    .Q_N(_00102_),
    .Q(\rbzero.tex_g1[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[39]$_DFFE_NP_  (.CLK(net2361),
    .RESET_B(net1663),
    .D(_01293_),
    .Q_N(_00103_),
    .Q(\rbzero.tex_g1[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[3]$_DFFE_NP_  (.CLK(net2360),
    .RESET_B(net1664),
    .D(_01294_),
    .Q_N(_00067_),
    .Q(\rbzero.tex_g1[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[40]$_DFFE_NP_  (.CLK(net2359),
    .RESET_B(net1665),
    .D(_01295_),
    .Q_N(_00104_),
    .Q(\rbzero.tex_g1[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[41]$_DFFE_NP_  (.CLK(net2358),
    .RESET_B(net1666),
    .D(_01296_),
    .Q_N(_00105_),
    .Q(\rbzero.tex_g1[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[42]$_DFFE_NP_  (.CLK(net2357),
    .RESET_B(net1667),
    .D(_01297_),
    .Q_N(_00106_),
    .Q(\rbzero.tex_g1[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[43]$_DFFE_NP_  (.CLK(net2356),
    .RESET_B(net1668),
    .D(_01298_),
    .Q_N(_00107_),
    .Q(\rbzero.tex_g1[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[44]$_DFFE_NP_  (.CLK(net2355),
    .RESET_B(net1669),
    .D(_01299_),
    .Q_N(_00108_),
    .Q(\rbzero.tex_g1[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[45]$_DFFE_NP_  (.CLK(net2354),
    .RESET_B(net1670),
    .D(_01300_),
    .Q_N(_00109_),
    .Q(\rbzero.tex_g1[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[46]$_DFFE_NP_  (.CLK(net2353),
    .RESET_B(net1671),
    .D(_01301_),
    .Q_N(_00110_),
    .Q(\rbzero.tex_g1[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[47]$_DFFE_NP_  (.CLK(net2352),
    .RESET_B(net1672),
    .D(_01302_),
    .Q_N(_00111_),
    .Q(\rbzero.tex_g1[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[48]$_DFFE_NP_  (.CLK(net2351),
    .RESET_B(net1673),
    .D(_01303_),
    .Q_N(_00112_),
    .Q(\rbzero.tex_g1[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[49]$_DFFE_NP_  (.CLK(net2350),
    .RESET_B(net1674),
    .D(_01304_),
    .Q_N(_00113_),
    .Q(\rbzero.tex_g1[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[4]$_DFFE_NP_  (.CLK(net2349),
    .RESET_B(net1675),
    .D(_01305_),
    .Q_N(_00068_),
    .Q(\rbzero.tex_g1[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[50]$_DFFE_NP_  (.CLK(net2348),
    .RESET_B(net1676),
    .D(_01306_),
    .Q_N(_00114_),
    .Q(\rbzero.tex_g1[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[51]$_DFFE_NP_  (.CLK(net2347),
    .RESET_B(net1677),
    .D(_01307_),
    .Q_N(_00115_),
    .Q(\rbzero.tex_g1[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[52]$_DFFE_NP_  (.CLK(net2346),
    .RESET_B(net1678),
    .D(_01308_),
    .Q_N(_00116_),
    .Q(\rbzero.tex_g1[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[53]$_DFFE_NP_  (.CLK(net2345),
    .RESET_B(net1679),
    .D(_01309_),
    .Q_N(_00117_),
    .Q(\rbzero.tex_g1[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[54]$_DFFE_NP_  (.CLK(net2344),
    .RESET_B(net1680),
    .D(_01310_),
    .Q_N(_00118_),
    .Q(\rbzero.tex_g1[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[55]$_DFFE_NP_  (.CLK(net2343),
    .RESET_B(net1681),
    .D(_01311_),
    .Q_N(_00119_),
    .Q(\rbzero.tex_g1[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[56]$_DFFE_NP_  (.CLK(net2342),
    .RESET_B(net1682),
    .D(_01312_),
    .Q_N(_00120_),
    .Q(\rbzero.tex_g1[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[57]$_DFFE_NP_  (.CLK(net2341),
    .RESET_B(net1683),
    .D(_01313_),
    .Q_N(_00121_),
    .Q(\rbzero.tex_g1[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[58]$_DFFE_NP_  (.CLK(net2340),
    .RESET_B(net1684),
    .D(_01314_),
    .Q_N(_00122_),
    .Q(\rbzero.tex_g1[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[59]$_DFFE_NP_  (.CLK(net2339),
    .RESET_B(net1685),
    .D(_01315_),
    .Q_N(_00123_),
    .Q(\rbzero.tex_g1[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[5]$_DFFE_NP_  (.CLK(net2338),
    .RESET_B(net1686),
    .D(_01316_),
    .Q_N(_00069_),
    .Q(\rbzero.tex_g1[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[60]$_DFFE_NP_  (.CLK(net2337),
    .RESET_B(net1687),
    .D(_01317_),
    .Q_N(_00124_),
    .Q(\rbzero.tex_g1[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[61]$_DFFE_NP_  (.CLK(net2336),
    .RESET_B(net1688),
    .D(_01318_),
    .Q_N(_00125_),
    .Q(\rbzero.tex_g1[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[62]$_DFFE_NP_  (.CLK(net2335),
    .RESET_B(net1689),
    .D(_01319_),
    .Q_N(_00126_),
    .Q(\rbzero.tex_g1[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[63]$_DFFE_NP_  (.CLK(net2334),
    .RESET_B(net1690),
    .D(_01320_),
    .Q_N(_00127_),
    .Q(\rbzero.tex_g1[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[6]$_DFFE_NP_  (.CLK(net2333),
    .RESET_B(net1691),
    .D(_01321_),
    .Q_N(_00070_),
    .Q(\rbzero.tex_g1[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[7]$_DFFE_NP_  (.CLK(net2332),
    .RESET_B(net1692),
    .D(_01322_),
    .Q_N(_00071_),
    .Q(\rbzero.tex_g1[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[8]$_DFFE_NP_  (.CLK(net2331),
    .RESET_B(net1693),
    .D(_01323_),
    .Q_N(_00072_),
    .Q(\rbzero.tex_g1[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_g1[9]$_DFFE_NP_  (.CLK(net2330),
    .RESET_B(net1694),
    .D(_01324_),
    .Q_N(_00073_),
    .Q(\rbzero.tex_g1[9] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[0]$_DFFE_NP_  (.CLK(net2329),
    .RESET_B(net1695),
    .D(_01325_),
    .Q_N(_00197_),
    .Q(\rbzero.tex_r0[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[10]$_DFFE_NP_  (.CLK(net2328),
    .RESET_B(net1696),
    .D(_01326_),
    .Q_N(_00207_),
    .Q(\rbzero.tex_r0[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[11]$_DFFE_NP_  (.CLK(net2327),
    .RESET_B(net1697),
    .D(_01327_),
    .Q_N(_00208_),
    .Q(\rbzero.tex_r0[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[12]$_DFFE_NP_  (.CLK(net2326),
    .RESET_B(net1698),
    .D(_01328_),
    .Q_N(_00209_),
    .Q(\rbzero.tex_r0[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[13]$_DFFE_NP_  (.CLK(net2325),
    .RESET_B(net1699),
    .D(_01329_),
    .Q_N(_00210_),
    .Q(\rbzero.tex_r0[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[14]$_DFFE_NP_  (.CLK(net2324),
    .RESET_B(net1700),
    .D(_01330_),
    .Q_N(_00211_),
    .Q(\rbzero.tex_r0[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[15]$_DFFE_NP_  (.CLK(net2323),
    .RESET_B(net1701),
    .D(_01331_),
    .Q_N(_00212_),
    .Q(\rbzero.tex_r0[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[16]$_DFFE_NP_  (.CLK(net2322),
    .RESET_B(net1702),
    .D(_01332_),
    .Q_N(_00213_),
    .Q(\rbzero.tex_r0[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[17]$_DFFE_NP_  (.CLK(net2321),
    .RESET_B(net1703),
    .D(_01333_),
    .Q_N(_00214_),
    .Q(\rbzero.tex_r0[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[18]$_DFFE_NP_  (.CLK(net2320),
    .RESET_B(net1704),
    .D(_01334_),
    .Q_N(_00215_),
    .Q(\rbzero.tex_r0[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[19]$_DFFE_NP_  (.CLK(net2319),
    .RESET_B(net1705),
    .D(_01335_),
    .Q_N(_00216_),
    .Q(\rbzero.tex_r0[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[1]$_DFFE_NP_  (.CLK(net2318),
    .RESET_B(net1706),
    .D(_01336_),
    .Q_N(_00198_),
    .Q(\rbzero.tex_r0[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[20]$_DFFE_NP_  (.CLK(net2317),
    .RESET_B(net1707),
    .D(_01337_),
    .Q_N(_00217_),
    .Q(\rbzero.tex_r0[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[21]$_DFFE_NP_  (.CLK(net2316),
    .RESET_B(net1708),
    .D(_01338_),
    .Q_N(_00218_),
    .Q(\rbzero.tex_r0[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[22]$_DFFE_NP_  (.CLK(net2315),
    .RESET_B(net1709),
    .D(_01339_),
    .Q_N(_00219_),
    .Q(\rbzero.tex_r0[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[23]$_DFFE_NP_  (.CLK(net2314),
    .RESET_B(net1710),
    .D(_01340_),
    .Q_N(_00220_),
    .Q(\rbzero.tex_r0[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[24]$_DFFE_NP_  (.CLK(net2313),
    .RESET_B(net1711),
    .D(_01341_),
    .Q_N(_00221_),
    .Q(\rbzero.tex_r0[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[25]$_DFFE_NP_  (.CLK(net2312),
    .RESET_B(net1712),
    .D(_01342_),
    .Q_N(_00222_),
    .Q(\rbzero.tex_r0[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[26]$_DFFE_NP_  (.CLK(net2311),
    .RESET_B(net1713),
    .D(_01343_),
    .Q_N(_00223_),
    .Q(\rbzero.tex_r0[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[27]$_DFFE_NP_  (.CLK(net2310),
    .RESET_B(net1714),
    .D(_01344_),
    .Q_N(_00224_),
    .Q(\rbzero.tex_r0[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[28]$_DFFE_NP_  (.CLK(net2309),
    .RESET_B(net1715),
    .D(_01345_),
    .Q_N(_00225_),
    .Q(\rbzero.tex_r0[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[29]$_DFFE_NP_  (.CLK(net2308),
    .RESET_B(net1716),
    .D(_01346_),
    .Q_N(_00226_),
    .Q(\rbzero.tex_r0[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[2]$_DFFE_NP_  (.CLK(net2307),
    .RESET_B(net1717),
    .D(_01347_),
    .Q_N(_00199_),
    .Q(\rbzero.tex_r0[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[30]$_DFFE_NP_  (.CLK(net2306),
    .RESET_B(net1718),
    .D(_01348_),
    .Q_N(_00227_),
    .Q(\rbzero.tex_r0[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[31]$_DFFE_NP_  (.CLK(net2305),
    .RESET_B(net1719),
    .D(_01349_),
    .Q_N(_00228_),
    .Q(\rbzero.tex_r0[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[32]$_DFFE_NP_  (.CLK(net2304),
    .RESET_B(net1720),
    .D(_01350_),
    .Q_N(_00229_),
    .Q(\rbzero.tex_r0[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[33]$_DFFE_NP_  (.CLK(net2303),
    .RESET_B(net1721),
    .D(_01351_),
    .Q_N(_00230_),
    .Q(\rbzero.tex_r0[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[34]$_DFFE_NP_  (.CLK(net2302),
    .RESET_B(net1722),
    .D(_01352_),
    .Q_N(_00231_),
    .Q(\rbzero.tex_r0[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[35]$_DFFE_NP_  (.CLK(net2301),
    .RESET_B(net1723),
    .D(_01353_),
    .Q_N(_00232_),
    .Q(\rbzero.tex_r0[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[36]$_DFFE_NP_  (.CLK(net2300),
    .RESET_B(net1724),
    .D(_01354_),
    .Q_N(_00233_),
    .Q(\rbzero.tex_r0[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[37]$_DFFE_NP_  (.CLK(net2299),
    .RESET_B(net1725),
    .D(_01355_),
    .Q_N(_00234_),
    .Q(\rbzero.tex_r0[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[38]$_DFFE_NP_  (.CLK(net2298),
    .RESET_B(net1726),
    .D(_01356_),
    .Q_N(_00235_),
    .Q(\rbzero.tex_r0[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[39]$_DFFE_NP_  (.CLK(net2297),
    .RESET_B(net1727),
    .D(_01357_),
    .Q_N(_00236_),
    .Q(\rbzero.tex_r0[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[3]$_DFFE_NP_  (.CLK(net2296),
    .RESET_B(net1728),
    .D(_01358_),
    .Q_N(_00200_),
    .Q(\rbzero.tex_r0[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[40]$_DFFE_NP_  (.CLK(net2295),
    .RESET_B(net1729),
    .D(_01359_),
    .Q_N(_00237_),
    .Q(\rbzero.tex_r0[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[41]$_DFFE_NP_  (.CLK(net2294),
    .RESET_B(net1730),
    .D(_01360_),
    .Q_N(_00238_),
    .Q(\rbzero.tex_r0[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[42]$_DFFE_NP_  (.CLK(net2293),
    .RESET_B(net1731),
    .D(_01361_),
    .Q_N(_00239_),
    .Q(\rbzero.tex_r0[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[43]$_DFFE_NP_  (.CLK(net2292),
    .RESET_B(net1732),
    .D(_01362_),
    .Q_N(_00240_),
    .Q(\rbzero.tex_r0[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[44]$_DFFE_NP_  (.CLK(net2291),
    .RESET_B(net1733),
    .D(_01363_),
    .Q_N(_00241_),
    .Q(\rbzero.tex_r0[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[45]$_DFFE_NP_  (.CLK(net2290),
    .RESET_B(net1734),
    .D(_01364_),
    .Q_N(_00242_),
    .Q(\rbzero.tex_r0[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[46]$_DFFE_NP_  (.CLK(net2289),
    .RESET_B(net1735),
    .D(_01365_),
    .Q_N(_00243_),
    .Q(\rbzero.tex_r0[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[47]$_DFFE_NP_  (.CLK(net2288),
    .RESET_B(net1736),
    .D(_01366_),
    .Q_N(_00244_),
    .Q(\rbzero.tex_r0[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[48]$_DFFE_NP_  (.CLK(net2287),
    .RESET_B(net1737),
    .D(_01367_),
    .Q_N(_00245_),
    .Q(\rbzero.tex_r0[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[49]$_DFFE_NP_  (.CLK(net2286),
    .RESET_B(net1738),
    .D(_01368_),
    .Q_N(_00246_),
    .Q(\rbzero.tex_r0[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[4]$_DFFE_NP_  (.CLK(net2285),
    .RESET_B(net1739),
    .D(_01369_),
    .Q_N(_00201_),
    .Q(\rbzero.tex_r0[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[50]$_DFFE_NP_  (.CLK(net2284),
    .RESET_B(net1740),
    .D(_01370_),
    .Q_N(_00247_),
    .Q(\rbzero.tex_r0[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[51]$_DFFE_NP_  (.CLK(net2283),
    .RESET_B(net1741),
    .D(_01371_),
    .Q_N(_00248_),
    .Q(\rbzero.tex_r0[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[52]$_DFFE_NP_  (.CLK(net2282),
    .RESET_B(net1742),
    .D(_01372_),
    .Q_N(_00249_),
    .Q(\rbzero.tex_r0[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[53]$_DFFE_NP_  (.CLK(net2281),
    .RESET_B(net1743),
    .D(_01373_),
    .Q_N(_00250_),
    .Q(\rbzero.tex_r0[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[54]$_DFFE_NP_  (.CLK(net2280),
    .RESET_B(net1744),
    .D(_01374_),
    .Q_N(_00251_),
    .Q(\rbzero.tex_r0[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[55]$_DFFE_NP_  (.CLK(net2279),
    .RESET_B(net1745),
    .D(_01375_),
    .Q_N(_00252_),
    .Q(\rbzero.tex_r0[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[56]$_DFFE_NP_  (.CLK(net2278),
    .RESET_B(net1746),
    .D(_01376_),
    .Q_N(_00253_),
    .Q(\rbzero.tex_r0[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[57]$_DFFE_NP_  (.CLK(net2277),
    .RESET_B(net1747),
    .D(_01377_),
    .Q_N(_00254_),
    .Q(\rbzero.tex_r0[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[58]$_DFFE_NP_  (.CLK(net2276),
    .RESET_B(net1748),
    .D(_01378_),
    .Q_N(_00255_),
    .Q(\rbzero.tex_r0[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[59]$_DFFE_NP_  (.CLK(net2275),
    .RESET_B(net1749),
    .D(_01379_),
    .Q_N(_00256_),
    .Q(\rbzero.tex_r0[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[5]$_DFFE_NP_  (.CLK(net2274),
    .RESET_B(net1750),
    .D(_01380_),
    .Q_N(_00202_),
    .Q(\rbzero.tex_r0[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[60]$_DFFE_NP_  (.CLK(net2273),
    .RESET_B(net1751),
    .D(_01381_),
    .Q_N(_00257_),
    .Q(\rbzero.tex_r0[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[61]$_DFFE_NP_  (.CLK(net2272),
    .RESET_B(net1752),
    .D(_01382_),
    .Q_N(_00258_),
    .Q(\rbzero.tex_r0[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[62]$_DFFE_NP_  (.CLK(net2271),
    .RESET_B(net1753),
    .D(_01383_),
    .Q_N(_00259_),
    .Q(\rbzero.tex_r0[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[63]$_DFFE_NP_  (.CLK(net2270),
    .RESET_B(net1754),
    .D(_01384_),
    .Q_N(_00260_),
    .Q(\rbzero.tex_r0[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[6]$_DFFE_NP_  (.CLK(net2269),
    .RESET_B(net1755),
    .D(_01385_),
    .Q_N(_00203_),
    .Q(\rbzero.tex_r0[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[7]$_DFFE_NP_  (.CLK(net2268),
    .RESET_B(net1756),
    .D(_01386_),
    .Q_N(_00204_),
    .Q(\rbzero.tex_r0[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[8]$_DFFE_NP_  (.CLK(net2267),
    .RESET_B(net1757),
    .D(_01387_),
    .Q_N(_00205_),
    .Q(\rbzero.tex_r0[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_r0[9]$_DFFE_NP_  (.CLK(net2266),
    .RESET_B(net1758),
    .D(_01388_),
    .Q_N(_00206_),
    .Q(\rbzero.tex_r0[9] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[0]$_DFFE_NP_  (.CLK(net2265),
    .RESET_B(net1759),
    .D(_01389_),
    .Q_N(_14432_),
    .Q(\rbzero.tex_r1[0] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[10]$_DFFE_NP_  (.CLK(net2264),
    .RESET_B(net1760),
    .D(_01390_),
    .Q_N(_14431_),
    .Q(\rbzero.tex_r1[10] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[11]$_DFFE_NP_  (.CLK(net2263),
    .RESET_B(net1761),
    .D(_01391_),
    .Q_N(_14430_),
    .Q(\rbzero.tex_r1[11] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[12]$_DFFE_NP_  (.CLK(net2262),
    .RESET_B(net1762),
    .D(_01392_),
    .Q_N(_14429_),
    .Q(\rbzero.tex_r1[12] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[13]$_DFFE_NP_  (.CLK(net2261),
    .RESET_B(net1763),
    .D(_01393_),
    .Q_N(_14428_),
    .Q(\rbzero.tex_r1[13] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[14]$_DFFE_NP_  (.CLK(net2260),
    .RESET_B(net1764),
    .D(_01394_),
    .Q_N(_14427_),
    .Q(\rbzero.tex_r1[14] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[15]$_DFFE_NP_  (.CLK(net2259),
    .RESET_B(net1765),
    .D(_01395_),
    .Q_N(_14426_),
    .Q(\rbzero.tex_r1[15] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[16]$_DFFE_NP_  (.CLK(net2258),
    .RESET_B(net1766),
    .D(_01396_),
    .Q_N(_14425_),
    .Q(\rbzero.tex_r1[16] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[17]$_DFFE_NP_  (.CLK(net2257),
    .RESET_B(net1767),
    .D(_01397_),
    .Q_N(_14424_),
    .Q(\rbzero.tex_r1[17] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[18]$_DFFE_NP_  (.CLK(net2256),
    .RESET_B(net1768),
    .D(_01398_),
    .Q_N(_14423_),
    .Q(\rbzero.tex_r1[18] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[19]$_DFFE_NP_  (.CLK(net2255),
    .RESET_B(net1769),
    .D(_01399_),
    .Q_N(_14422_),
    .Q(\rbzero.tex_r1[19] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[1]$_DFFE_NP_  (.CLK(net2254),
    .RESET_B(net1770),
    .D(_01400_),
    .Q_N(_14421_),
    .Q(\rbzero.tex_r1[1] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[20]$_DFFE_NP_  (.CLK(net2253),
    .RESET_B(net1771),
    .D(_01401_),
    .Q_N(_14420_),
    .Q(\rbzero.tex_r1[20] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[21]$_DFFE_NP_  (.CLK(net2252),
    .RESET_B(net1772),
    .D(_01402_),
    .Q_N(_14419_),
    .Q(\rbzero.tex_r1[21] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[22]$_DFFE_NP_  (.CLK(net2251),
    .RESET_B(net1773),
    .D(_01403_),
    .Q_N(_14418_),
    .Q(\rbzero.tex_r1[22] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[23]$_DFFE_NP_  (.CLK(net2250),
    .RESET_B(net1774),
    .D(_01404_),
    .Q_N(_14417_),
    .Q(\rbzero.tex_r1[23] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[24]$_DFFE_NP_  (.CLK(net2249),
    .RESET_B(net1775),
    .D(_01405_),
    .Q_N(_14416_),
    .Q(\rbzero.tex_r1[24] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[25]$_DFFE_NP_  (.CLK(net2248),
    .RESET_B(net1776),
    .D(_01406_),
    .Q_N(_14415_),
    .Q(\rbzero.tex_r1[25] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[26]$_DFFE_NP_  (.CLK(net2247),
    .RESET_B(net1777),
    .D(_01407_),
    .Q_N(_14414_),
    .Q(\rbzero.tex_r1[26] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[27]$_DFFE_NP_  (.CLK(net2246),
    .RESET_B(net1778),
    .D(_01408_),
    .Q_N(_14413_),
    .Q(\rbzero.tex_r1[27] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[28]$_DFFE_NP_  (.CLK(net2245),
    .RESET_B(net1779),
    .D(_01409_),
    .Q_N(_14412_),
    .Q(\rbzero.tex_r1[28] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[29]$_DFFE_NP_  (.CLK(net2244),
    .RESET_B(net1780),
    .D(_01410_),
    .Q_N(_14411_),
    .Q(\rbzero.tex_r1[29] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[2]$_DFFE_NP_  (.CLK(net2243),
    .RESET_B(net1781),
    .D(_01411_),
    .Q_N(_14410_),
    .Q(\rbzero.tex_r1[2] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[30]$_DFFE_NP_  (.CLK(net2242),
    .RESET_B(net1782),
    .D(_01412_),
    .Q_N(_14409_),
    .Q(\rbzero.tex_r1[30] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[31]$_DFFE_NP_  (.CLK(net2241),
    .RESET_B(net1783),
    .D(_01413_),
    .Q_N(_14408_),
    .Q(\rbzero.tex_r1[31] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[32]$_DFFE_NP_  (.CLK(net2240),
    .RESET_B(net1784),
    .D(_01414_),
    .Q_N(_14407_),
    .Q(\rbzero.tex_r1[32] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[33]$_DFFE_NP_  (.CLK(net2239),
    .RESET_B(net1785),
    .D(_01415_),
    .Q_N(_14406_),
    .Q(\rbzero.tex_r1[33] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[34]$_DFFE_NP_  (.CLK(net2238),
    .RESET_B(net1786),
    .D(_01416_),
    .Q_N(_14405_),
    .Q(\rbzero.tex_r1[34] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[35]$_DFFE_NP_  (.CLK(net2237),
    .RESET_B(net1787),
    .D(_01417_),
    .Q_N(_14404_),
    .Q(\rbzero.tex_r1[35] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[36]$_DFFE_NP_  (.CLK(net2236),
    .RESET_B(net1788),
    .D(_01418_),
    .Q_N(_14403_),
    .Q(\rbzero.tex_r1[36] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[37]$_DFFE_NP_  (.CLK(net2235),
    .RESET_B(net1789),
    .D(_01419_),
    .Q_N(_14402_),
    .Q(\rbzero.tex_r1[37] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[38]$_DFFE_NP_  (.CLK(net2234),
    .RESET_B(net1790),
    .D(_01420_),
    .Q_N(_14401_),
    .Q(\rbzero.tex_r1[38] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[39]$_DFFE_NP_  (.CLK(net2233),
    .RESET_B(net1791),
    .D(_01421_),
    .Q_N(_14400_),
    .Q(\rbzero.tex_r1[39] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[3]$_DFFE_NP_  (.CLK(net2232),
    .RESET_B(net1792),
    .D(_01422_),
    .Q_N(_14399_),
    .Q(\rbzero.tex_r1[3] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[40]$_DFFE_NP_  (.CLK(net2231),
    .RESET_B(net1793),
    .D(_01423_),
    .Q_N(_14398_),
    .Q(\rbzero.tex_r1[40] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[41]$_DFFE_NP_  (.CLK(net2230),
    .RESET_B(net1794),
    .D(_01424_),
    .Q_N(_14397_),
    .Q(\rbzero.tex_r1[41] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[42]$_DFFE_NP_  (.CLK(net2229),
    .RESET_B(net1795),
    .D(_01425_),
    .Q_N(_14396_),
    .Q(\rbzero.tex_r1[42] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[43]$_DFFE_NP_  (.CLK(net2228),
    .RESET_B(net1796),
    .D(_01426_),
    .Q_N(_14395_),
    .Q(\rbzero.tex_r1[43] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[44]$_DFFE_NP_  (.CLK(net2227),
    .RESET_B(net1797),
    .D(_01427_),
    .Q_N(_14394_),
    .Q(\rbzero.tex_r1[44] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[45]$_DFFE_NP_  (.CLK(net2226),
    .RESET_B(net1798),
    .D(_01428_),
    .Q_N(_14393_),
    .Q(\rbzero.tex_r1[45] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[46]$_DFFE_NP_  (.CLK(net2225),
    .RESET_B(net1799),
    .D(_01429_),
    .Q_N(_14392_),
    .Q(\rbzero.tex_r1[46] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[47]$_DFFE_NP_  (.CLK(net2224),
    .RESET_B(net1800),
    .D(_01430_),
    .Q_N(_14391_),
    .Q(\rbzero.tex_r1[47] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[48]$_DFFE_NP_  (.CLK(net2223),
    .RESET_B(net1801),
    .D(_01431_),
    .Q_N(_14390_),
    .Q(\rbzero.tex_r1[48] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[49]$_DFFE_NP_  (.CLK(net2222),
    .RESET_B(net1802),
    .D(_01432_),
    .Q_N(_14389_),
    .Q(\rbzero.tex_r1[49] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[4]$_DFFE_NP_  (.CLK(net2221),
    .RESET_B(net1803),
    .D(_01433_),
    .Q_N(_14388_),
    .Q(\rbzero.tex_r1[4] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[50]$_DFFE_NP_  (.CLK(net2220),
    .RESET_B(net1804),
    .D(_01434_),
    .Q_N(_14387_),
    .Q(\rbzero.tex_r1[50] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[51]$_DFFE_NP_  (.CLK(net2219),
    .RESET_B(net1805),
    .D(_01435_),
    .Q_N(_14386_),
    .Q(\rbzero.tex_r1[51] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[52]$_DFFE_NP_  (.CLK(net2218),
    .RESET_B(net1806),
    .D(_01436_),
    .Q_N(_14385_),
    .Q(\rbzero.tex_r1[52] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[53]$_DFFE_NP_  (.CLK(net2217),
    .RESET_B(net1807),
    .D(_01437_),
    .Q_N(_14384_),
    .Q(\rbzero.tex_r1[53] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[54]$_DFFE_NP_  (.CLK(net2216),
    .RESET_B(net1808),
    .D(_01438_),
    .Q_N(_14383_),
    .Q(\rbzero.tex_r1[54] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[55]$_DFFE_NP_  (.CLK(net2215),
    .RESET_B(net1809),
    .D(_01439_),
    .Q_N(_14382_),
    .Q(\rbzero.tex_r1[55] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[56]$_DFFE_NP_  (.CLK(net2214),
    .RESET_B(net1810),
    .D(_01440_),
    .Q_N(_14381_),
    .Q(\rbzero.tex_r1[56] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[57]$_DFFE_NP_  (.CLK(net2213),
    .RESET_B(net1811),
    .D(_01441_),
    .Q_N(_14380_),
    .Q(\rbzero.tex_r1[57] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[58]$_DFFE_NP_  (.CLK(net2212),
    .RESET_B(net1812),
    .D(_01442_),
    .Q_N(_14379_),
    .Q(\rbzero.tex_r1[58] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[59]$_DFFE_NP_  (.CLK(net2211),
    .RESET_B(net1813),
    .D(_01443_),
    .Q_N(_14378_),
    .Q(\rbzero.tex_r1[59] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[5]$_DFFE_NP_  (.CLK(net2210),
    .RESET_B(net1814),
    .D(_01444_),
    .Q_N(_14377_),
    .Q(\rbzero.tex_r1[5] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[60]$_DFFE_NP_  (.CLK(net2209),
    .RESET_B(net1815),
    .D(_01445_),
    .Q_N(_14376_),
    .Q(\rbzero.tex_r1[60] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[61]$_DFFE_NP_  (.CLK(net2208),
    .RESET_B(net1816),
    .D(_01446_),
    .Q_N(_14375_),
    .Q(\rbzero.tex_r1[61] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[62]$_DFFE_NP_  (.CLK(net2207),
    .RESET_B(net1817),
    .D(_01447_),
    .Q_N(_14374_),
    .Q(\rbzero.tex_r1[62] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[63]$_DFFE_NP_  (.CLK(net2206),
    .RESET_B(net1818),
    .D(_01448_),
    .Q_N(_14373_),
    .Q(\rbzero.tex_r1[63] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[6]$_DFFE_NP_  (.CLK(net2205),
    .RESET_B(net1819),
    .D(_01449_),
    .Q_N(_14372_),
    .Q(\rbzero.tex_r1[6] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[7]$_DFFE_NP_  (.CLK(net2204),
    .RESET_B(net1820),
    .D(_01450_),
    .Q_N(_14371_),
    .Q(\rbzero.tex_r1[7] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[8]$_DFFE_NP_  (.CLK(net2203),
    .RESET_B(net1821),
    .D(_01451_),
    .Q_N(_14370_),
    .Q(\rbzero.tex_r1[8] ));
 sg13g2_dfrbp_1 \rbzero.tex_r1[9]$_DFFE_NP_  (.CLK(net2202),
    .RESET_B(net1822),
    .D(_01452_),
    .Q_N(_14369_),
    .Q(\rbzero.tex_r1[9] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[0]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1823),
    .D(_01453_),
    .Q_N(\rbzero.debug_overlay.h[0] ),
    .Q(\hpos[0] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[1]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1824),
    .D(_01454_),
    .Q_N(_00028_),
    .Q(\hpos[1] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[2]$_SDFF_PP0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1825),
    .D(_01455_),
    .Q_N(_00027_),
    .Q(\hpos[2] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[3]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1826),
    .D(_01456_),
    .Q_N(_00014_),
    .Q(\hpos[3] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[4]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1827),
    .D(_01457_),
    .Q_N(_00051_),
    .Q(\hpos[4] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[5]$_SDFF_PP0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1828),
    .D(_01458_),
    .Q_N(_00025_),
    .Q(\hpos[5] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[6]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1829),
    .D(_01459_),
    .Q_N(_14368_),
    .Q(\hpos[6] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[7]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1830),
    .D(_01460_),
    .Q_N(_00024_),
    .Q(\hpos[7] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[8]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1831),
    .D(_01461_),
    .Q_N(_00053_),
    .Q(\hpos[8] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hpos[9]$_SDFF_PP0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1832),
    .D(_01462_),
    .Q_N(_00052_),
    .Q(\hpos[9] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.hsync$_SDFFE_PP0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1833),
    .D(_01463_),
    .Q_N(hsync_n),
    .Q(\rbzero.hsync ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1834),
    .D(_01464_),
    .Q_N(_14367_),
    .Q(\rbzero.debug_overlay.vpos[0] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1835),
    .D(_01465_),
    .Q_N(_14366_),
    .Q(\rbzero.debug_overlay.vpos[1] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1836),
    .D(_01466_),
    .Q_N(_14365_),
    .Q(\rbzero.debug_overlay.vpos[2] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1837),
    .D(_01467_),
    .Q_N(_14364_),
    .Q(\rbzero.debug_overlay.vpos[3] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1838),
    .D(_01468_),
    .Q_N(_14363_),
    .Q(\rbzero.debug_overlay.vpos[4] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1839),
    .D(_01469_),
    .Q_N(_00058_),
    .Q(\rbzero.debug_overlay.vpos[5] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1840),
    .D(_01470_),
    .Q_N(_14362_),
    .Q(\rbzero.debug_overlay.vpos[6] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1841),
    .D(_01471_),
    .Q_N(_14361_),
    .Q(\rbzero.debug_overlay.vpos[7] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1842),
    .D(_01472_),
    .Q_N(_14360_),
    .Q(\rbzero.debug_overlay.vpos[8] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vpos[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1843),
    .D(_01473_),
    .Q_N(_14359_),
    .Q(\rbzero.debug_overlay.vpos[9] ));
 sg13g2_dfrbp_1 \rbzero.vga_sync.vsync$_SDFFE_PP0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1844),
    .D(_01474_),
    .Q_N(\rbzero.vsync_n ),
    .Q(\rbzero.vga_sync.vsync ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1845),
    .D(_01475_),
    .Q_N(_00394_),
    .Q(\rbzero.map_rom.i_col[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1846),
    .D(_01476_),
    .Q_N(_14358_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1847),
    .D(_01477_),
    .Q_N(_14357_),
    .Q(\rbzero.map_rom.i_col[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1848),
    .D(_01478_),
    .Q_N(_14356_),
    .Q(\rbzero.map_rom.i_col[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1849),
    .D(_01479_),
    .Q_N(_00021_),
    .Q(\rbzero.map_rom.i_col[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1850),
    .D(_01480_),
    .Q_N(_00019_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1851),
    .D(_01481_),
    .Q_N(_14355_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1852),
    .D(_01482_),
    .Q_N(_00395_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1853),
    .D(_01483_),
    .Q_N(_00396_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1854),
    .D(_01484_),
    .Q_N(_00397_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapX[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1855),
    .D(_01485_),
    .Q_N(_00398_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1856),
    .D(_01486_),
    .Q_N(_00393_),
    .Q(\rbzero.map_rom.i_row[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1857),
    .D(_01487_),
    .Q_N(_14354_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1858),
    .D(_01488_),
    .Q_N(_14353_),
    .Q(\rbzero.map_rom.i_row[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1859),
    .D(_01489_),
    .Q_N(_00022_),
    .Q(\rbzero.map_rom.i_row[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1860),
    .D(_01490_),
    .Q_N(_14352_),
    .Q(\rbzero.map_rom.i_row[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1861),
    .D(_01491_),
    .Q_N(_00020_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1862),
    .D(_01492_),
    .Q_N(_14351_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1863),
    .D(_01493_),
    .Q_N(_14350_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1864),
    .D(_01494_),
    .Q_N(_14349_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1865),
    .D(_01495_),
    .Q_N(_14348_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.mapY[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1866),
    .D(_01496_),
    .Q_N(_14347_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_side$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1867),
    .D(_01497_),
    .Q_N(_00055_),
    .Q(\rbzero.row_render.side ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_side_hot$_SDFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1868),
    .D(_01498_),
    .Q_N(_14346_),
    .Q(\rbzero.side_hot ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1869),
    .D(_01499_),
    .Q_N(_00050_),
    .Q(\rbzero.row_render.size[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1870),
    .D(_01500_),
    .Q_N(_00047_),
    .Q(\rbzero.row_render.size[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1871),
    .D(_01501_),
    .Q_N(_14345_),
    .Q(\rbzero.row_render.size[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1872),
    .D(_01502_),
    .Q_N(_14344_),
    .Q(\rbzero.row_render.size[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1873),
    .D(_01503_),
    .Q_N(_14343_),
    .Q(\rbzero.row_render.size[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1874),
    .D(_01504_),
    .Q_N(_14342_),
    .Q(\rbzero.row_render.size[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1875),
    .D(_01505_),
    .Q_N(_14341_),
    .Q(\rbzero.row_render.size[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1876),
    .D(_01506_),
    .Q_N(_00049_),
    .Q(\rbzero.row_render.size[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1877),
    .D(_01507_),
    .Q_N(_14340_),
    .Q(\rbzero.row_render.size[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1878),
    .D(_01508_),
    .Q_N(_00048_),
    .Q(\rbzero.row_render.size[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_size[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1879),
    .D(_01509_),
    .Q_N(_14339_),
    .Q(\rbzero.row_render.size[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1880),
    .D(_01510_),
    .Q_N(_14338_),
    .Q(\rbzero.traced_texVinit[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1881),
    .D(_01511_),
    .Q_N(_14337_),
    .Q(\rbzero.traced_texVinit[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1882),
    .D(_01512_),
    .Q_N(_14336_),
    .Q(\rbzero.traced_texVinit[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1883),
    .D(_01513_),
    .Q_N(_14335_),
    .Q(\rbzero.traced_texVinit[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1884),
    .D(_01514_),
    .Q_N(_14334_),
    .Q(\rbzero.traced_texVinit[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1885),
    .D(_01515_),
    .Q_N(_14333_),
    .Q(\rbzero.traced_texVinit[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1886),
    .D(_01516_),
    .Q_N(_14332_),
    .Q(\rbzero.traced_texVinit[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1887),
    .D(_01517_),
    .Q_N(_14331_),
    .Q(\rbzero.traced_texVinit[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1888),
    .D(_01518_),
    .Q_N(_14330_),
    .Q(\rbzero.traced_texVinit[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1889),
    .D(_01519_),
    .Q_N(_14329_),
    .Q(\rbzero.traced_texVinit[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texVinit[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1890),
    .D(_01520_),
    .Q_N(_14328_),
    .Q(\rbzero.traced_texVinit[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1891),
    .D(_01521_),
    .Q_N(_14327_),
    .Q(\rbzero.traced_texa[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1892),
    .D(_01522_),
    .Q_N(_14326_),
    .Q(\rbzero.traced_texa[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1893),
    .D(_01523_),
    .Q_N(_14325_),
    .Q(\rbzero.traced_texa[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1894),
    .D(_01524_),
    .Q_N(_14324_),
    .Q(\rbzero.traced_texa[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1895),
    .D(_01525_),
    .Q_N(_14323_),
    .Q(\rbzero.traced_texa[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1896),
    .D(_01526_),
    .Q_N(_14322_),
    .Q(\rbzero.traced_texa[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1897),
    .D(_01527_),
    .Q_N(_14321_),
    .Q(\rbzero.traced_texa[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1898),
    .D(_01528_),
    .Q_N(_14320_),
    .Q(\rbzero.traced_texa[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1899),
    .D(_01529_),
    .Q_N(_14319_),
    .Q(\rbzero.traced_texa[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1900),
    .D(_01530_),
    .Q_N(_14318_),
    .Q(\rbzero.traced_texa[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1901),
    .D(_01531_),
    .Q_N(_14317_),
    .Q(\rbzero.traced_texa[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1902),
    .D(_01532_),
    .Q_N(_14316_),
    .Q(\rbzero.traced_texa[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1903),
    .D(_01533_),
    .Q_N(_14315_),
    .Q(\rbzero.traced_texa[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1904),
    .D(_01534_),
    .Q_N(_14314_),
    .Q(\rbzero.traced_texa[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1905),
    .D(_01535_),
    .Q_N(_14313_),
    .Q(\rbzero.traced_texa[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1906),
    .D(_01536_),
    .Q_N(_14312_),
    .Q(\rbzero.traced_texa[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1907),
    .D(_01537_),
    .Q_N(_14311_),
    .Q(\rbzero.traced_texa[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1908),
    .D(_01538_),
    .Q_N(_14310_),
    .Q(\rbzero.traced_texa[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1909),
    .D(_01539_),
    .Q_N(_14309_),
    .Q(\rbzero.traced_texa[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1910),
    .D(_01540_),
    .Q_N(_14308_),
    .Q(\rbzero.traced_texa[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1911),
    .D(_01541_),
    .Q_N(_14307_),
    .Q(\rbzero.traced_texa[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texa[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1912),
    .D(_01542_),
    .Q_N(_14306_),
    .Q(\rbzero.traced_texa[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1913),
    .D(_01543_),
    .Q_N(_00194_),
    .Q(\rbzero.row_render.texu[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1914),
    .D(_01544_),
    .Q_N(_14305_),
    .Q(\rbzero.row_render.texu[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1915),
    .D(_01545_),
    .Q_N(_14304_),
    .Q(\rbzero.row_render.texu[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1916),
    .D(_01546_),
    .Q_N(_00056_),
    .Q(\rbzero.row_render.texu[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1917),
    .D(_01547_),
    .Q_N(_00054_),
    .Q(\rbzero.row_render.texu[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1918),
    .D(_01548_),
    .Q_N(_14303_),
    .Q(\rbzero.texu_hot[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1919),
    .D(_01549_),
    .Q_N(_14302_),
    .Q(\rbzero.texu_hot[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1920),
    .D(_01550_),
    .Q_N(_14301_),
    .Q(\rbzero.texu_hot[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1921),
    .D(_01551_),
    .Q_N(_14300_),
    .Q(\rbzero.texu_hot[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1922),
    .D(_01552_),
    .Q_N(_14299_),
    .Q(\rbzero.texu_hot[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_texu_hot[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1923),
    .D(_01553_),
    .Q_N(_14298_),
    .Q(\rbzero.texu_hot[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_wall[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1924),
    .D(_01554_),
    .Q_N(_14297_),
    .Q(\rbzero.row_render.wall[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_wall[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1925),
    .D(_01555_),
    .Q_N(_14296_),
    .Q(\rbzero.row_render.wall[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_wall_hot[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1926),
    .D(_01556_),
    .Q_N(_14295_),
    .Q(\rbzero.wall_hot[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.o_wall_hot[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1927),
    .D(_01557_),
    .Q_N(_14294_),
    .Q(\rbzero.wall_hot[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[10]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1928),
    .D(_01558_),
    .Q_N(_14293_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[11]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1929),
    .D(_01559_),
    .Q_N(_14292_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1930),
    .D(_01560_),
    .Q_N(_14291_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[13]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1931),
    .D(_01561_),
    .Q_N(_14290_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[14]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1932),
    .D(_01562_),
    .Q_N(_14289_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[15]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1933),
    .D(_01563_),
    .Q_N(_14288_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[16]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1934),
    .D(_01564_),
    .Q_N(_14287_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[17]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1935),
    .D(_01565_),
    .Q_N(_14286_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[18]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1936),
    .D(_01566_),
    .Q_N(_14285_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[19]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1937),
    .D(_01567_),
    .Q_N(_14284_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[20]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1938),
    .D(_01568_),
    .Q_N(_14283_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[21]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1939),
    .D(_01569_),
    .Q_N(_14282_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1940),
    .D(_01570_),
    .Q_N(_14281_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1941),
    .D(_01571_),
    .Q_N(_14280_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1942),
    .D(_01572_),
    .Q_N(_14279_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1943),
    .D(_01573_),
    .Q_N(_14278_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[6]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1944),
    .D(_01574_),
    .Q_N(_14277_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[7]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1945),
    .D(_01575_),
    .Q_N(_14276_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[8]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1946),
    .D(_01576_),
    .Q_N(_14275_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendX[9]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1947),
    .D(_01577_),
    .Q_N(_14274_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1948),
    .D(_01578_),
    .Q_N(_14273_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[11]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1949),
    .D(_01579_),
    .Q_N(_14272_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[12]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1950),
    .D(_01580_),
    .Q_N(_14271_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1951),
    .D(_01581_),
    .Q_N(_14270_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[14]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1952),
    .D(_01582_),
    .Q_N(_14269_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[15]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1953),
    .D(_01583_),
    .Q_N(_14268_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1954),
    .D(_01584_),
    .Q_N(_14267_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[17]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1955),
    .D(_01585_),
    .Q_N(_14266_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[18]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1956),
    .D(_01586_),
    .Q_N(_14265_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[19]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1957),
    .D(_01587_),
    .Q_N(_14264_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[20]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1958),
    .D(_01588_),
    .Q_N(_14263_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[21]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1959),
    .D(_01589_),
    .Q_N(_14262_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1960),
    .D(_01590_),
    .Q_N(_14261_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1961),
    .D(_01591_),
    .Q_N(_14260_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1962),
    .D(_01592_),
    .Q_N(_14259_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1963),
    .D(_01593_),
    .Q_N(_14258_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[6]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1964),
    .D(_01594_),
    .Q_N(_14257_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[7]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1965),
    .D(_01595_),
    .Q_N(_14256_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1966),
    .D(_01596_),
    .Q_N(_14255_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rayAddendY[9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1967),
    .D(_01597_),
    .Q_N(_14254_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1968),
    .D(_01598_),
    .Q_N(_14253_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1969),
    .D(_01599_),
    .Q_N(_14252_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1970),
    .D(_01600_),
    .Q_N(_14251_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1971),
    .D(_01601_),
    .Q_N(_14250_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1972),
    .D(_01602_),
    .Q_N(_14249_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1973),
    .D(_01603_),
    .Q_N(_14248_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1974),
    .D(_01604_),
    .Q_N(_14247_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1975),
    .D(_01605_),
    .Q_N(_14246_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1976),
    .D(_01606_),
    .Q_N(_14245_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1977),
    .D(_01607_),
    .Q_N(_14244_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1978),
    .D(_01608_),
    .Q_N(_14243_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1979),
    .D(_01609_),
    .Q_N(_14242_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1980),
    .D(_01610_),
    .Q_N(_14241_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1981),
    .D(_01611_),
    .Q_N(_14240_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1982),
    .D(_01612_),
    .Q_N(_14239_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1983),
    .D(_01613_),
    .Q_N(_14238_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1984),
    .D(_01614_),
    .Q_N(_14237_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1985),
    .D(_01615_),
    .Q_N(_14236_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1986),
    .D(_01616_),
    .Q_N(_14235_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1987),
    .D(_01617_),
    .Q_N(_14234_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1988),
    .D(_01618_),
    .Q_N(_14233_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_data[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1989),
    .D(_01619_),
    .Q_N(_14232_),
    .Q(\rbzero.wall_tracer.rcp_fsm.o_data[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.o_done$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1990),
    .D(_01620_),
    .Q_N(_14231_),
    .Q(\rbzero.wall_tracer.rcp_done ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1991),
    .D(_01621_),
    .Q_N(_00474_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1992),
    .D(_01622_),
    .Q_N(_14230_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1993),
    .D(_01623_),
    .Q_N(_14229_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1994),
    .D(_01624_),
    .Q_N(_14228_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1995),
    .D(_01625_),
    .Q_N(_14227_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1996),
    .D(_01626_),
    .Q_N(_14226_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1997),
    .D(_01627_),
    .Q_N(_14225_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1998),
    .D(_01628_),
    .Q_N(_14224_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1999),
    .D(_01629_),
    .Q_N(_14223_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2000),
    .D(_01630_),
    .Q_N(_14222_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2001),
    .D(_01631_),
    .Q_N(_14221_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2002),
    .D(_01632_),
    .Q_N(_00472_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2003),
    .D(_01633_),
    .Q_N(_14220_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2004),
    .D(_01634_),
    .Q_N(_00473_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2005),
    .D(_01635_),
    .Q_N(_14219_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2006),
    .D(_01636_),
    .Q_N(_14218_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2007),
    .D(_01637_),
    .Q_N(_14217_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2008),
    .D(_01638_),
    .Q_N(_14216_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2009),
    .D(_01639_),
    .Q_N(_14215_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2010),
    .D(_01640_),
    .Q_N(_14214_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2011),
    .D(_01641_),
    .Q_N(_14213_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.operand[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2012),
    .D(_01642_),
    .Q_N(_14976_),
    .Q(\rbzero.wall_tracer.rcp_fsm.operand[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.state[0]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2013),
    .D(_00004_),
    .Q_N(_14977_),
    .Q(\rbzero.wall_tracer.rcp_fsm.state[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.state[1]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2014),
    .D(_00000_),
    .Q_N(_14978_),
    .Q(\rbzero.wall_tracer.rcp_fsm.state[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.state[2]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2015),
    .D(_00001_),
    .Q_N(_14979_),
    .Q(\rbzero.wall_tracer.rcp_fsm.state[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.state[3]$_DFF_P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2016),
    .D(_00002_),
    .Q_N(_14980_),
    .Q(\rbzero.wall_tracer.rcp_fsm.state[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_fsm.state[4]$_DFF_P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2017),
    .D(_00003_),
    .Q_N(_14212_),
    .Q(\rbzero.wall_tracer.rcp_fsm.state[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2018),
    .D(_01643_),
    .Q_N(_14211_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2019),
    .D(_01644_),
    .Q_N(_14210_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2020),
    .D(_01645_),
    .Q_N(_14209_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2021),
    .D(_01646_),
    .Q_N(_14208_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2022),
    .D(_01647_),
    .Q_N(_14207_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2023),
    .D(_01648_),
    .Q_N(_14206_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2024),
    .D(_01649_),
    .Q_N(_14205_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2025),
    .D(_01650_),
    .Q_N(_14204_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net2026),
    .D(_01651_),
    .Q_N(_14203_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2027),
    .D(_01652_),
    .Q_N(_14202_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2028),
    .D(_01653_),
    .Q_N(_14201_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2029),
    .D(_01654_),
    .Q_N(_14200_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2030),
    .D(_01655_),
    .Q_N(_14199_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2031),
    .D(_01656_),
    .Q_N(_14198_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2032),
    .D(_01657_),
    .Q_N(_14197_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2033),
    .D(_01658_),
    .Q_N(_14196_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2034),
    .D(_01659_),
    .Q_N(_14195_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2035),
    .D(_01660_),
    .Q_N(_14194_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2036),
    .D(_01661_),
    .Q_N(_14193_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2037),
    .D(_01662_),
    .Q_N(_14192_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2038),
    .D(_01663_),
    .Q_N(_14191_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_in[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2039),
    .D(_01664_),
    .Q_N(_14190_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_data[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.rcp_start$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2040),
    .D(_01665_),
    .Q_N(_00016_),
    .Q(\rbzero.wall_tracer.rcp_fsm.i_start ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.side$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2041),
    .D(_01666_),
    .Q_N(_14189_),
    .Q(\rbzero.wall_tracer.side ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2042),
    .D(_01667_),
    .Q_N(_14188_),
    .Q(\rbzero.wall_tracer.size_full[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net2043),
    .D(_01668_),
    .Q_N(_14187_),
    .Q(\rbzero.wall_tracer.size[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2044),
    .D(_01669_),
    .Q_N(_14186_),
    .Q(\rbzero.wall_tracer.size[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2045),
    .D(_01670_),
    .Q_N(_00453_),
    .Q(\rbzero.wall_tracer.size[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net2046),
    .D(_01671_),
    .Q_N(_14185_),
    .Q(\rbzero.wall_tracer.size[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2047),
    .D(_01672_),
    .Q_N(_14184_),
    .Q(\rbzero.wall_tracer.size_full[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2048),
    .D(_01673_),
    .Q_N(_14183_),
    .Q(\rbzero.wall_tracer.size_full[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2049),
    .D(_01674_),
    .Q_N(_14182_),
    .Q(\rbzero.wall_tracer.size_full[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2050),
    .D(_01675_),
    .Q_N(_14181_),
    .Q(\rbzero.wall_tracer.size_full[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2051),
    .D(_01676_),
    .Q_N(_14180_),
    .Q(\rbzero.wall_tracer.size_full[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2052),
    .D(_01677_),
    .Q_N(_14179_),
    .Q(\rbzero.wall_tracer.size_full[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2053),
    .D(_01678_),
    .Q_N(_14178_),
    .Q(\rbzero.wall_tracer.size_full[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2054),
    .D(_01679_),
    .Q_N(_14177_),
    .Q(\rbzero.wall_tracer.size_full[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2055),
    .D(_01680_),
    .Q_N(_14176_),
    .Q(\rbzero.wall_tracer.size_full[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2056),
    .D(_01681_),
    .Q_N(_00405_),
    .Q(\rbzero.wall_tracer.size_full[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2057),
    .D(_01682_),
    .Q_N(_00411_),
    .Q(\rbzero.wall_tracer.size[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2058),
    .D(_01683_),
    .Q_N(_00416_),
    .Q(\rbzero.wall_tracer.size[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2059),
    .D(_01684_),
    .Q_N(_00422_),
    .Q(\rbzero.wall_tracer.size[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2060),
    .D(_01685_),
    .Q_N(_00428_),
    .Q(\rbzero.wall_tracer.size[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2061),
    .D(_01686_),
    .Q_N(_00434_),
    .Q(\rbzero.wall_tracer.size[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2062),
    .D(_01687_),
    .Q_N(_00440_),
    .Q(\rbzero.wall_tracer.size[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.size_full[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2063),
    .D(_01688_),
    .Q_N(_14981_),
    .Q(\rbzero.wall_tracer.size[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[0]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2064),
    .D(_00005_),
    .Q_N(_14982_),
    .Q(\rbzero.wall_tracer.state[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[1]$_DFF_P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2065),
    .D(_00006_),
    .Q_N(_00017_),
    .Q(\rbzero.wall_tracer.state[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[2]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2066),
    .D(_00007_),
    .Q_N(_14983_),
    .Q(\rbzero.wall_tracer.state[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[3]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2067),
    .D(_00008_),
    .Q_N(_00023_),
    .Q(\rbzero.wall_tracer.state[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[4]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2068),
    .D(_00009_),
    .Q_N(_14984_),
    .Q(\rbzero.wall_tracer.state[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[5]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2069),
    .D(_00010_),
    .Q_N(_14985_),
    .Q(\rbzero.wall_tracer.state[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[6]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2070),
    .D(_00011_),
    .Q_N(_14986_),
    .Q(\rbzero.wall_tracer.state[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[7]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net2071),
    .D(_00012_),
    .Q_N(_14987_),
    .Q(\rbzero.wall_tracer.state[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.state[8]$_DFF_P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2072),
    .D(_00013_),
    .Q_N(_14175_),
    .Q(\rbzero.wall_tracer.state[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2073),
    .D(_01689_),
    .Q_N(_14174_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2074),
    .D(_01690_),
    .Q_N(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2075),
    .D(_01691_),
    .Q_N(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2076),
    .D(_01692_),
    .Q_N(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2077),
    .D(_01693_),
    .Q_N(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2078),
    .D(_01694_),
    .Q_N(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2079),
    .D(_01695_),
    .Q_N(_00458_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2080),
    .D(_01696_),
    .Q_N(_00460_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2081),
    .D(_01697_),
    .Q_N(_00462_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2082),
    .D(_01698_),
    .Q_N(_00464_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2083),
    .D(_01699_),
    .Q_N(_00466_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2084),
    .D(_01700_),
    .Q_N(_14173_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2085),
    .D(_01701_),
    .Q_N(_00468_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2086),
    .D(_01702_),
    .Q_N(_00470_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2087),
    .D(_01703_),
    .Q_N(_00403_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2088),
    .D(_01704_),
    .Q_N(_00409_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2089),
    .D(_01705_),
    .Q_N(_00414_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2090),
    .D(_01706_),
    .Q_N(_00420_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2091),
    .D(_01707_),
    .Q_N(_00426_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2092),
    .D(_01708_),
    .Q_N(_00432_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2093),
    .D(_01709_),
    .Q_N(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistX[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2094),
    .D(_01710_),
    .Q_N(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2095),
    .D(_01711_),
    .Q_N(_14172_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2096),
    .D(_01712_),
    .Q_N(_00448_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2097),
    .D(_01713_),
    .Q_N(_00450_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2098),
    .D(_01714_),
    .Q_N(_00452_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2099),
    .D(_01715_),
    .Q_N(_00455_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2100),
    .D(_01716_),
    .Q_N(_00457_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2101),
    .D(_01717_),
    .Q_N(_00459_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2102),
    .D(_01718_),
    .Q_N(_00461_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2103),
    .D(_01719_),
    .Q_N(_00463_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2104),
    .D(_01720_),
    .Q_N(_00465_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2105),
    .D(_01721_),
    .Q_N(_00467_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2106),
    .D(_01722_),
    .Q_N(_14171_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2107),
    .D(_01723_),
    .Q_N(_00469_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2108),
    .D(_01724_),
    .Q_N(_00471_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net2109),
    .D(_01725_),
    .Q_N(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2110),
    .D(_01726_),
    .Q_N(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2111),
    .D(_01727_),
    .Q_N(_00415_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2112),
    .D(_01728_),
    .Q_N(_00421_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2113),
    .D(_01729_),
    .Q_N(_00427_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2114),
    .D(_01730_),
    .Q_N(_00433_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2115),
    .D(_01731_),
    .Q_N(_00439_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.stepDistY[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net2116),
    .D(_01732_),
    .Q_N(_00445_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net2117),
    .D(_01733_),
    .Q_N(_14170_),
    .Q(\rbzero.wall_tracer.texu[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2118),
    .D(_01734_),
    .Q_N(_14169_),
    .Q(\rbzero.wall_tracer.texu[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2119),
    .D(_01735_),
    .Q_N(_14168_),
    .Q(\rbzero.wall_tracer.texu[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2120),
    .D(_01736_),
    .Q_N(_14167_),
    .Q(\rbzero.wall_tracer.texu[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net2121),
    .D(_01737_),
    .Q_N(_14166_),
    .Q(\rbzero.wall_tracer.texu[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.texu[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2122),
    .D(_01738_),
    .Q_N(_14165_),
    .Q(\rbzero.wall_tracer.texu[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2123),
    .D(_01739_),
    .Q_N(_14164_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2124),
    .D(_01740_),
    .Q_N(_14163_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2125),
    .D(_01741_),
    .Q_N(_14162_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2126),
    .D(_01742_),
    .Q_N(_14161_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2127),
    .D(_01743_),
    .Q_N(_14160_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2128),
    .D(_01744_),
    .Q_N(_14159_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2129),
    .D(_01745_),
    .Q_N(_14158_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2130),
    .D(_01746_),
    .Q_N(_14157_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2131),
    .D(_01747_),
    .Q_N(_14156_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2132),
    .D(_01748_),
    .Q_N(_14155_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2133),
    .D(_01749_),
    .Q_N(_14154_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2134),
    .D(_01750_),
    .Q_N(_14153_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2135),
    .D(_01751_),
    .Q_N(_14152_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2136),
    .D(_01752_),
    .Q_N(_14151_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2137),
    .D(_01753_),
    .Q_N(_14150_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net2138),
    .D(_01754_),
    .Q_N(_14149_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2139),
    .D(_01755_),
    .Q_N(_14148_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2140),
    .D(_01756_),
    .Q_N(_14147_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2141),
    .D(_01757_),
    .Q_N(_14146_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2142),
    .D(_01758_),
    .Q_N(_14145_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2143),
    .D(_01759_),
    .Q_N(_14144_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistX[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2144),
    .D(_01760_),
    .Q_N(_14143_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2145),
    .D(_01761_),
    .Q_N(_14142_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2146),
    .D(_01762_),
    .Q_N(_14141_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2147),
    .D(_01763_),
    .Q_N(_14140_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2148),
    .D(_01764_),
    .Q_N(_14139_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2149),
    .D(_01765_),
    .Q_N(_14138_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2150),
    .D(_01766_),
    .Q_N(_14137_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2151),
    .D(_01767_),
    .Q_N(_14136_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2152),
    .D(_01768_),
    .Q_N(_14135_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2153),
    .D(_01769_),
    .Q_N(_14134_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2154),
    .D(_01770_),
    .Q_N(_14133_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2155),
    .D(_01771_),
    .Q_N(_14132_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2156),
    .D(_01772_),
    .Q_N(_14131_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2157),
    .D(_01773_),
    .Q_N(_14130_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2158),
    .D(_01774_),
    .Q_N(_14129_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2159),
    .D(_01775_),
    .Q_N(_14128_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2160),
    .D(_01776_),
    .Q_N(_14127_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2161),
    .D(_01777_),
    .Q_N(_14126_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2162),
    .D(_01778_),
    .Q_N(_14125_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2163),
    .D(_01779_),
    .Q_N(_14124_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2164),
    .D(_01780_),
    .Q_N(_14123_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2165),
    .D(_01781_),
    .Q_N(_14122_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.trackDistY[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2166),
    .D(_01782_),
    .Q_N(_14121_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2167),
    .D(_01783_),
    .Q_N(_14120_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2168),
    .D(_01784_),
    .Q_N(_00400_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2169),
    .D(_01785_),
    .Q_N(_00399_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2170),
    .D(_01786_),
    .Q_N(_14119_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2171),
    .D(_01787_),
    .Q_N(_14118_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2172),
    .D(_01788_),
    .Q_N(_14117_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2173),
    .D(_01789_),
    .Q_N(_14116_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2174),
    .D(_01790_),
    .Q_N(_14115_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2175),
    .D(_01791_),
    .Q_N(_14114_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2176),
    .D(_01792_),
    .Q_N(_14113_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2177),
    .D(_01793_),
    .Q_N(_14112_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2178),
    .D(_01794_),
    .Q_N(_14111_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2179),
    .D(_01795_),
    .Q_N(_14110_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2180),
    .D(_01796_),
    .Q_N(_14109_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2181),
    .D(_01797_),
    .Q_N(_00446_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2182),
    .D(_01798_),
    .Q_N(_00441_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2183),
    .D(_01799_),
    .Q_N(_00435_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2184),
    .D(_01800_),
    .Q_N(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2185),
    .D(_01801_),
    .Q_N(_00423_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2186),
    .D(_01802_),
    .Q_N(_00417_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2187),
    .D(_01803_),
    .Q_N(_00018_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.visualWallDist[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net2188),
    .D(_01804_),
    .Q_N(_00406_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.w[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2189),
    .D(_01805_),
    .Q_N(_14108_),
    .Q(\rbzero.wall_tracer.w[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.w[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net2190),
    .D(_01806_),
    .Q_N(_14107_),
    .Q(\rbzero.wall_tracer.w[1] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.w[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net2191),
    .D(_01807_),
    .Q_N(_00015_),
    .Q(\rbzero.wall_tracer.w[2] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.wall[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2192),
    .D(_01808_),
    .Q_N(_14106_),
    .Q(\rbzero.wall_tracer.wall[0] ));
 sg13g2_dfrbp_1 \rbzero.wall_tracer.wall[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2193),
    .D(_01809_),
    .Q_N(_14988_),
    .Q(\rbzero.wall_tracer.wall[1] ));
 sg13g2_dfrbp_1 \registered_vga_output[0]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2194),
    .D(\rbzero.rgb[1] ),
    .Q_N(_14989_),
    .Q(\registered_vga_output[0] ));
 sg13g2_dfrbp_1 \registered_vga_output[1]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2195),
    .D(\rbzero.rgb[3] ),
    .Q_N(_14990_),
    .Q(\registered_vga_output[1] ));
 sg13g2_dfrbp_1 \registered_vga_output[2]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2196),
    .D(\rbzero.rgb[5] ),
    .Q_N(_14991_),
    .Q(\registered_vga_output[2] ));
 sg13g2_dfrbp_1 \registered_vga_output[3]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2197),
    .D(\rbzero.vsync_n ),
    .Q_N(_14992_),
    .Q(\registered_vga_output[3] ));
 sg13g2_dfrbp_1 \registered_vga_output[4]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2198),
    .D(\rbzero.rgb[0] ),
    .Q_N(_14993_),
    .Q(\registered_vga_output[4] ));
 sg13g2_dfrbp_1 \registered_vga_output[5]$_DFF_P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2199),
    .D(\rbzero.rgb[2] ),
    .Q_N(_14994_),
    .Q(\registered_vga_output[5] ));
 sg13g2_dfrbp_1 \registered_vga_output[6]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net2200),
    .D(\rbzero.rgb[4] ),
    .Q_N(_14995_),
    .Q(\registered_vga_output[6] ));
 sg13g2_dfrbp_1 \registered_vga_output[7]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2201),
    .D(hsync_n),
    .Q_N(_14105_),
    .Q(\registered_vga_output[7] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[3]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[7]),
    .X(net12));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[0]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[1]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout25 (.A(_05486_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_05465_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_05278_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_04259_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_04553_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04459_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_04590_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_03987_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_04039_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04153_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_04081_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_04047_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_04004_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_04003_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_04209_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_04123_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_04054_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_04036_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_04726_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_04203_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_04128_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04018_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_04280_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_03880_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_04527_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_04197_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_04048_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_04033_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_04547_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_04281_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_07176_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_04741_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_07249_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_07175_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_07169_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_05997_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_05988_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_04337_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_11478_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_11344_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_07218_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_07167_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_11531_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_11346_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_11343_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_07166_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_11345_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_11342_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_05722_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_02974_),
    .X(net74));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_07362_));
 sg13g2_buf_2 fanout76 (.A(_05721_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_03211_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_03206_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_03502_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_03996_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_06772_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_06593_));
 sg13g2_buf_2 fanout83 (.A(_02695_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_06644_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_04139_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_04138_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_04093_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03394_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_06232_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_04695_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_04145_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_04092_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_04043_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_03409_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03128_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_03070_),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(_08054_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_08045_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_08042_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04380_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04045_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04017_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04001_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03458_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_03397_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_02926_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_02619_),
    .X(net107));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_08300_));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(_08299_));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_08213_));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_08055_));
 sg13g2_buf_2 fanout112 (.A(_07968_),
    .X(net112));
 sg13g2_buf_8 fanout113 (.A(_07962_),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_07944_));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_07932_));
 sg13g2_buf_2 fanout116 (.A(_07913_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_06371_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_04500_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03258_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03083_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_02861_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02680_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_08287_));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_08211_));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_07969_));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_07964_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_07961_));
 sg13g2_buf_2 fanout128 (.A(_07957_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_07945_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_07943_));
 sg13g2_buf_2 fanout131 (.A(_07939_),
    .X(net131));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_07938_));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_07933_));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_07931_));
 sg13g2_buf_2 fanout135 (.A(_06520_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_06317_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04355_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04321_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04231_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04223_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_03067_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_02860_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_02853_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_02851_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_02790_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_02774_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_02761_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_02706_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_01890_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_13913_),
    .X(net150));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_07963_));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_07960_));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_07956_));
 sg13g2_buf_2 fanout154 (.A(_07950_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_07909_),
    .X(net155));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_07890_));
 sg13g2_buf_2 fanout157 (.A(_07886_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_07881_));
 sg13g2_buf_2 fanout159 (.A(_07838_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04419_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04362_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03073_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_02857_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_02760_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_02749_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_02734_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_02722_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_02705_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_02686_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_02616_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_02457_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_13954_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_13948_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_13903_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_07889_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_07864_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_07844_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03744_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_03573_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_03526_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03081_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03074_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03040_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02981_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_02933_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_02856_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_02792_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_02783_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_02772_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_02770_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_02759_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_02740_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_02733_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_02730_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_02728_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_02721_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_02712_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_02704_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_02685_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_02669_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_02615_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_02548_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_02456_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_14071_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_13920_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_13904_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_13758_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_13191_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_13174_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_13049_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_12905_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_06090_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_03645_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03171_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03080_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_03069_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_03049_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03010_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_02914_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_02913_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_02889_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_02745_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_02727_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_02711_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_02703_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_02684_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02641_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_02590_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_02455_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_02407_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_01891_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_13950_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_13947_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_13791_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_13748_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_13351_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_13160_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_12391_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_12383_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_12335_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_04100_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_03129_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_03079_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_03068_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_03048_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_03038_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_03009_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_02683_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_02681_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_02675_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_02673_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_02672_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_02640_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_02406_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_01812_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_01810_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_13910_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_13179_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_12959_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_12456_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_12452_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_12388_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_12337_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_12135_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_12066_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_11999_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_11938_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_11781_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_03041_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_02892_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_02767_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_02756_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_02755_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_02688_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_02682_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_12925_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_12762_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_12709_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_12226_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_12172_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_12012_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_11977_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_11780_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_06125_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_02687_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_02452_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_02421_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_01839_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_05234_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_05189_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_02577_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_12928_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_12813_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_11447_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_05307_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_05140_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_02558_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_02373_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_02367_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_13788_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_13221_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_11440_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_02518_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_02384_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_02377_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_12209_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_11794_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_11439_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_05306_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_05231_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_02432_));
 sg13g2_buf_2 fanout312 (.A(_02422_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_02376_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_11629_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_05230_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_02660_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_02565_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_02479_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_13216_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_07386_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_07379_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_07350_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_05720_),
    .X(net323));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_02569_));
 sg13g2_buf_2 fanout325 (.A(_02557_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_02494_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_02492_),
    .X(net327));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_02411_));
 sg13g2_buf_2 fanout329 (.A(_02368_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_02359_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_02254_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_12739_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_11837_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_09959_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_09956_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_09867_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_09861_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_09859_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_09831_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_09421_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_02495_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_02487_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_02395_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_02390_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_02361_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_02307_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_10369_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_10367_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_09860_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_09832_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_09825_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_09821_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_09765_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_09763_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_09748_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_09745_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_09743_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_09737_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_09420_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_02469_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_02355_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_13367_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_12362_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_11102_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_11100_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_11079_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_11077_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_11056_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_11054_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_11033_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_11031_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_11010_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_11008_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_10987_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_10985_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_10964_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_10961_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_10907_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_10905_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_10879_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_10877_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_10856_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_10854_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_10833_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_10831_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_10816_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_10813_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_09736_),
    .X(net388));
 sg13g2_buf_4 fanout389 (.X(net389),
    .A(_08733_));
 sg13g2_buf_4 fanout390 (.X(net390),
    .A(_08732_));
 sg13g2_buf_4 fanout391 (.X(net391),
    .A(_08731_));
 sg13g2_buf_4 fanout392 (.X(net392),
    .A(_08730_));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(_08729_));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(_08728_));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_08727_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_08726_));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_08725_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_08724_));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(_08723_));
 sg13g2_buf_4 fanout400 (.X(net400),
    .A(_08722_));
 sg13g2_buf_4 fanout401 (.X(net401),
    .A(_08721_));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_08708_));
 sg13g2_buf_2 fanout403 (.A(_02282_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_12974_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_12410_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_12217_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_11940_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_11148_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_11146_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_11125_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_11123_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_10815_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_10812_),
    .X(net413));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(_08745_));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(_08744_));
 sg13g2_buf_4 fanout416 (.X(net416),
    .A(_08743_));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(_08742_));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_08741_));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(_08740_));
 sg13g2_buf_4 fanout420 (.X(net420),
    .A(_08739_));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_08738_));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_08737_));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(_08736_));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(_08735_));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(_08734_));
 sg13g2_buf_4 fanout426 (.X(net426),
    .A(_08718_));
 sg13g2_buf_4 fanout427 (.X(net427),
    .A(_08717_));
 sg13g2_buf_4 fanout428 (.X(net428),
    .A(_08716_));
 sg13g2_buf_4 fanout429 (.X(net429),
    .A(_08715_));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_08714_));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(_08713_));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(_08705_));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_08704_));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(_08703_));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(_08702_));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(_08701_));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(_08700_));
 sg13g2_buf_2 fanout438 (.A(_01950_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_01935_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_01927_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_01912_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_13883_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_12423_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_12398_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_12244_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_12166_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_12124_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_11743_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_11734_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_11715_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_09740_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_08682_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_02249_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_12239_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_12138_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_12120_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_11988_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_11958_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_11714_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_09063_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_08981_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_08808_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_08749_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_08681_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_02218_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_12177_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_12144_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_12034_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_06133_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_10645_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_10621_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_09653_),
    .X(net472));
 sg13g2_buf_2 fanout473 (.A(_09538_),
    .X(net473));
 sg13g2_buf_2 fanout474 (.A(_05880_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_05874_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_05848_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_01863_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_01846_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_13391_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_13384_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_13023_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_12987_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_10763_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_10739_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_10703_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_10678_),
    .X(net486));
 sg13g2_buf_1 fanout487 (.A(_10637_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_10623_),
    .X(net488));
 sg13g2_buf_1 fanout489 (.A(_10620_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_08678_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_08450_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_08429_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_07639_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_05749_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_05739_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_05728_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_02187_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_01841_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_13807_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_13789_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_13368_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_13246_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_12732_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_12403_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_12363_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_11841_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_10705_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_10681_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_10580_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_10551_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_10468_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_08428_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_05812_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_05806_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_05780_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_05727_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_13712_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_12841_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_12837_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_12424_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_12415_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_12262_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_12169_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_11848_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_11721_),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_10928_));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(_10916_));
 sg13g2_buf_2 fanout528 (.A(_10799_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_10755_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_10729_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_10680_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_10536_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_10510_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_10335_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_10312_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_10288_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_10265_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_10242_),
    .X(net538));
 sg13g2_buf_1 fanout539 (.A(_10233_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_10219_),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(_10210_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_10194_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_09707_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_08693_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_08642_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_08635_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_08477_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_05902_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_05873_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_05841_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_05814_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_05782_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_05758_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_05735_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_05679_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_05664_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_05652_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_05639_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_05622_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_05599_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_02069_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_01989_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_01963_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_01940_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_01917_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_13630_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_12727_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_12199_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_11928_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_11866_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_11839_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_11765_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_11713_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_10765_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_10741_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_10714_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_10690_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_10600_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_10568_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_10499_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_10484_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_10470_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_10451_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_10450_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_10423_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_10422_),
    .X(net586));
 sg13g2_buf_1 fanout587 (.A(_10326_),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(_10302_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_10287_),
    .X(net589));
 sg13g2_buf_1 fanout590 (.A(_10279_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_10264_),
    .X(net591));
 sg13g2_buf_1 fanout592 (.A(_10256_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_10241_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_10218_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_10196_),
    .X(net595));
 sg13g2_buf_1 fanout596 (.A(_10193_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_10189_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_10167_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_10144_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_10120_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_10097_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_10074_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_10051_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_10027_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_09901_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_09760_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_09702_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_09078_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_09043_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_08641_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_08447_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_07377_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_07312_),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(_07223_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_07221_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_07126_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_07124_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_05994_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_05992_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_05648_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_05608_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_05606_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_05584_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_02046_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_02029_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_02008_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_02003_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_01997_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_12780_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_11798_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_11768_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_11726_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_11712_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_11690_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_11527_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_11507_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_11471_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_11353_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_11143_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_11120_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_11097_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_11074_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_11051_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_11028_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_11005_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_10982_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_10957_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_10898_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_10874_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_10851_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_10826_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_10794_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_10773_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_10749_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_10723_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_10698_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_10671_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10650_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10627_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_10598_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_10582_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10565_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_10553_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_10532_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_10512_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_10506_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_10478_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_10446_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_10433_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_10388_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_10356_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_10334_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_10311_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_09724_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_09701_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_09071_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_09058_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_09051_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_08791_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_08747_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_08692_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_08676_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_08446_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_08442_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_08421_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_08413_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_07539_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_05472_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_05452_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_02056_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_02028_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_02023_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_02018_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_02007_),
    .X(net694));
 sg13g2_buf_4 fanout695 (.X(net695),
    .A(_02002_));
 sg13g2_buf_2 fanout696 (.A(_01996_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_12129_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_11767_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_11711_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_11486_),
    .X(net700));
 sg13g2_buf_2 fanout701 (.A(_11470_),
    .X(net701));
 sg13g2_buf_2 fanout702 (.A(_11352_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_11347_),
    .X(net703));
 sg13g2_buf_1 fanout704 (.A(_10169_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_10156_),
    .X(net705));
 sg13g2_buf_1 fanout706 (.A(_10146_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_10132_),
    .X(net707));
 sg13g2_buf_1 fanout708 (.A(_10122_),
    .X(net708));
 sg13g2_buf_2 fanout709 (.A(_10109_),
    .X(net709));
 sg13g2_buf_1 fanout710 (.A(_10099_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_10086_),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(_10076_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_10063_),
    .X(net713));
 sg13g2_buf_1 fanout714 (.A(_10053_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_10040_),
    .X(net715));
 sg13g2_buf_1 fanout716 (.A(_10030_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_09776_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_09513_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_09460_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_09457_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_09177_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_08793_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_08710_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_08646_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_08445_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_08441_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_08433_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_08420_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_08412_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_07653_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_05646_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_02198_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_02171_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_02064_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_02035_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_02027_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_02013_),
    .X(net737));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(_02001_));
 sg13g2_buf_2 fanout739 (.A(_01995_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_11771_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_11710_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_10927_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_10913_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_10439_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_10436_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_10430_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_10427_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_10414_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_10379_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_10190_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_09816_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_09761_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_09726_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_09698_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_09627_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_09480_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_09476_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_09425_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_09423_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_09292_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_09248_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_09242_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_09164_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_09158_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_09144_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_09142_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_09141_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_09127_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_09126_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_09125_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_08928_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_08911_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_08890_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_08874_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_08865_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_08831_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_08815_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_08814_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_08812_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_08795_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_08794_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_08792_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_08709_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_08670_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_08663_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_08651_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_08648_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_08645_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_08591_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_08590_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_08558_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_08517_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_08510_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_08506_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_08480_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_08454_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_08444_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_08440_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_08432_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_08419_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_07907_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_02199_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_02140_),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(_02139_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_02138_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_02088_),
    .X(net806));
 sg13g2_buf_2 fanout807 (.A(_02031_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_02021_),
    .X(net808));
 sg13g2_buf_2 fanout809 (.A(_01991_),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(_01987_),
    .X(net810));
 sg13g2_buf_2 fanout811 (.A(_11732_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_11717_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_11709_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_10443_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_09461_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_09401_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_09207_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_09190_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_09174_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_09157_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_09133_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_09086_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_08997_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_08898_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_08830_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_08759_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_08495_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_08459_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_08457_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_08455_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_08452_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_08435_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_08418_),
    .X(net833));
 sg13g2_tielo _28663__834 (.L_LO(net834));
 sg13g2_tielo _28664__835 (.L_LO(net835));
 sg13g2_tielo _28665__836 (.L_LO(net836));
 sg13g2_tielo _28666__837 (.L_LO(net837));
 sg13g2_tielo _28667__838 (.L_LO(net838));
 sg13g2_tielo _28670__839 (.L_LO(net839));
 sg13g2_tielo _28671__840 (.L_LO(net840));
 sg13g2_tielo _28672__841 (.L_LO(net841));
 sg13g2_tielo _28674__842 (.L_LO(net842));
 sg13g2_tielo _28675__843 (.L_LO(net843));
 sg13g2_tiehi _28662__845 (.L_HI(net845));
 sg13g2_tiehi \rbzero.pov.facingRX[0]$_SDFFE_PN0P__846  (.L_HI(net846));
 sg13g2_tiehi \rbzero.pov.facingRX[10]$_SDFFE_PN0P__847  (.L_HI(net847));
 sg13g2_tiehi \rbzero.pov.facingRX[1]$_SDFFE_PN0P__848  (.L_HI(net848));
 sg13g2_tiehi \rbzero.pov.facingRX[2]$_SDFFE_PN0P__849  (.L_HI(net849));
 sg13g2_tiehi \rbzero.pov.facingRX[3]$_SDFFE_PN0P__850  (.L_HI(net850));
 sg13g2_tiehi \rbzero.pov.facingRX[4]$_SDFFE_PN1P__851  (.L_HI(net851));
 sg13g2_tiehi \rbzero.pov.facingRX[5]$_SDFFE_PN1P__852  (.L_HI(net852));
 sg13g2_tiehi \rbzero.pov.facingRX[6]$_SDFFE_PN1P__853  (.L_HI(net853));
 sg13g2_tiehi \rbzero.pov.facingRX[7]$_SDFFE_PN0P__854  (.L_HI(net854));
 sg13g2_tiehi \rbzero.pov.facingRX[8]$_SDFFE_PN1P__855  (.L_HI(net855));
 sg13g2_tiehi \rbzero.pov.facingRX[9]$_SDFFE_PN0P__856  (.L_HI(net856));
 sg13g2_tiehi \rbzero.pov.facingRY[0]$_SDFFE_PN1P__857  (.L_HI(net857));
 sg13g2_tiehi \rbzero.pov.facingRY[10]$_SDFFE_PN1P__858  (.L_HI(net858));
 sg13g2_tiehi \rbzero.pov.facingRY[1]$_SDFFE_PN0P__859  (.L_HI(net859));
 sg13g2_tiehi \rbzero.pov.facingRY[2]$_SDFFE_PN1P__860  (.L_HI(net860));
 sg13g2_tiehi \rbzero.pov.facingRY[3]$_SDFFE_PN1P__861  (.L_HI(net861));
 sg13g2_tiehi \rbzero.pov.facingRY[4]$_SDFFE_PN1P__862  (.L_HI(net862));
 sg13g2_tiehi \rbzero.pov.facingRY[5]$_SDFFE_PN0P__863  (.L_HI(net863));
 sg13g2_tiehi \rbzero.pov.facingRY[6]$_SDFFE_PN0P__864  (.L_HI(net864));
 sg13g2_tiehi \rbzero.pov.facingRY[7]$_SDFFE_PN1P__865  (.L_HI(net865));
 sg13g2_tiehi \rbzero.pov.facingRY[8]$_SDFFE_PN0P__866  (.L_HI(net866));
 sg13g2_tiehi \rbzero.pov.facingRY[9]$_SDFFE_PN1P__867  (.L_HI(net867));
 sg13g2_tiehi \rbzero.pov.mosi_buffer[0]$_SDFF_PN0__868  (.L_HI(net868));
 sg13g2_tiehi \rbzero.pov.mosi_buffer[1]$_SDFF_PN0__869  (.L_HI(net869));
 sg13g2_tiehi \rbzero.pov.playerRX[0]$_SDFFE_PN0P__870  (.L_HI(net870));
 sg13g2_tiehi \rbzero.pov.playerRX[10]$_SDFFE_PN1P__871  (.L_HI(net871));
 sg13g2_tiehi \rbzero.pov.playerRX[11]$_SDFFE_PN0P__872  (.L_HI(net872));
 sg13g2_tiehi \rbzero.pov.playerRX[12]$_SDFFE_PN1P__873  (.L_HI(net873));
 sg13g2_tiehi \rbzero.pov.playerRX[13]$_SDFFE_PN0P__874  (.L_HI(net874));
 sg13g2_tiehi \rbzero.pov.playerRX[14]$_SDFFE_PN0P__875  (.L_HI(net875));
 sg13g2_tiehi \rbzero.pov.playerRX[1]$_SDFFE_PN0P__876  (.L_HI(net876));
 sg13g2_tiehi \rbzero.pov.playerRX[2]$_SDFFE_PN0P__877  (.L_HI(net877));
 sg13g2_tiehi \rbzero.pov.playerRX[3]$_SDFFE_PN0P__878  (.L_HI(net878));
 sg13g2_tiehi \rbzero.pov.playerRX[4]$_SDFFE_PN0P__879  (.L_HI(net879));
 sg13g2_tiehi \rbzero.pov.playerRX[5]$_SDFFE_PN0P__880  (.L_HI(net880));
 sg13g2_tiehi \rbzero.pov.playerRX[6]$_SDFFE_PN0P__881  (.L_HI(net881));
 sg13g2_tiehi \rbzero.pov.playerRX[7]$_SDFFE_PN0P__882  (.L_HI(net882));
 sg13g2_tiehi \rbzero.pov.playerRX[8]$_SDFFE_PN1P__883  (.L_HI(net883));
 sg13g2_tiehi \rbzero.pov.playerRX[9]$_SDFFE_PN1P__884  (.L_HI(net884));
 sg13g2_tiehi \rbzero.pov.playerRY[0]$_SDFFE_PN0P__885  (.L_HI(net885));
 sg13g2_tiehi \rbzero.pov.playerRY[10]$_SDFFE_PN1P__886  (.L_HI(net886));
 sg13g2_tiehi \rbzero.pov.playerRY[11]$_SDFFE_PN0P__887  (.L_HI(net887));
 sg13g2_tiehi \rbzero.pov.playerRY[12]$_SDFFE_PN1P__888  (.L_HI(net888));
 sg13g2_tiehi \rbzero.pov.playerRY[13]$_SDFFE_PN0P__889  (.L_HI(net889));
 sg13g2_tiehi \rbzero.pov.playerRY[14]$_SDFFE_PN0P__890  (.L_HI(net890));
 sg13g2_tiehi \rbzero.pov.playerRY[1]$_SDFFE_PN0P__891  (.L_HI(net891));
 sg13g2_tiehi \rbzero.pov.playerRY[2]$_SDFFE_PN0P__892  (.L_HI(net892));
 sg13g2_tiehi \rbzero.pov.playerRY[3]$_SDFFE_PN0P__893  (.L_HI(net893));
 sg13g2_tiehi \rbzero.pov.playerRY[4]$_SDFFE_PN0P__894  (.L_HI(net894));
 sg13g2_tiehi \rbzero.pov.playerRY[5]$_SDFFE_PN0P__895  (.L_HI(net895));
 sg13g2_tiehi \rbzero.pov.playerRY[6]$_SDFFE_PN0P__896  (.L_HI(net896));
 sg13g2_tiehi \rbzero.pov.playerRY[7]$_SDFFE_PN0P__897  (.L_HI(net897));
 sg13g2_tiehi \rbzero.pov.playerRY[8]$_SDFFE_PN1P__898  (.L_HI(net898));
 sg13g2_tiehi \rbzero.pov.playerRY[9]$_SDFFE_PN0P__899  (.L_HI(net899));
 sg13g2_tiehi \rbzero.pov.ready$_SDFFE_PP0P__900  (.L_HI(net900));
 sg13g2_tiehi \rbzero.pov.ready_buffer[0]$_SDFFE_PN0P__901  (.L_HI(net901));
 sg13g2_tiehi \rbzero.pov.ready_buffer[10]$_SDFFE_PN0P__902  (.L_HI(net902));
 sg13g2_tiehi \rbzero.pov.ready_buffer[11]$_SDFFE_PN0P__903  (.L_HI(net903));
 sg13g2_tiehi \rbzero.pov.ready_buffer[12]$_SDFFE_PN0P__904  (.L_HI(net904));
 sg13g2_tiehi \rbzero.pov.ready_buffer[13]$_SDFFE_PN0P__905  (.L_HI(net905));
 sg13g2_tiehi \rbzero.pov.ready_buffer[14]$_SDFFE_PN0P__906  (.L_HI(net906));
 sg13g2_tiehi \rbzero.pov.ready_buffer[15]$_SDFFE_PN0P__907  (.L_HI(net907));
 sg13g2_tiehi \rbzero.pov.ready_buffer[16]$_SDFFE_PN0P__908  (.L_HI(net908));
 sg13g2_tiehi \rbzero.pov.ready_buffer[17]$_SDFFE_PN0P__909  (.L_HI(net909));
 sg13g2_tiehi \rbzero.pov.ready_buffer[18]$_SDFFE_PN0P__910  (.L_HI(net910));
 sg13g2_tiehi \rbzero.pov.ready_buffer[19]$_SDFFE_PN0P__911  (.L_HI(net911));
 sg13g2_tiehi \rbzero.pov.ready_buffer[1]$_SDFFE_PN0P__912  (.L_HI(net912));
 sg13g2_tiehi \rbzero.pov.ready_buffer[20]$_SDFFE_PN0P__913  (.L_HI(net913));
 sg13g2_tiehi \rbzero.pov.ready_buffer[21]$_SDFFE_PN0P__914  (.L_HI(net914));
 sg13g2_tiehi \rbzero.pov.ready_buffer[22]$_SDFFE_PN0P__915  (.L_HI(net915));
 sg13g2_tiehi \rbzero.pov.ready_buffer[23]$_SDFFE_PN0P__916  (.L_HI(net916));
 sg13g2_tiehi \rbzero.pov.ready_buffer[24]$_SDFFE_PN0P__917  (.L_HI(net917));
 sg13g2_tiehi \rbzero.pov.ready_buffer[25]$_SDFFE_PN0P__918  (.L_HI(net918));
 sg13g2_tiehi \rbzero.pov.ready_buffer[26]$_SDFFE_PN0P__919  (.L_HI(net919));
 sg13g2_tiehi \rbzero.pov.ready_buffer[27]$_SDFFE_PN0P__920  (.L_HI(net920));
 sg13g2_tiehi \rbzero.pov.ready_buffer[28]$_SDFFE_PN0P__921  (.L_HI(net921));
 sg13g2_tiehi \rbzero.pov.ready_buffer[29]$_SDFFE_PN0P__922  (.L_HI(net922));
 sg13g2_tiehi \rbzero.pov.ready_buffer[2]$_SDFFE_PN0P__923  (.L_HI(net923));
 sg13g2_tiehi \rbzero.pov.ready_buffer[30]$_SDFFE_PN0P__924  (.L_HI(net924));
 sg13g2_tiehi \rbzero.pov.ready_buffer[31]$_SDFFE_PN0P__925  (.L_HI(net925));
 sg13g2_tiehi \rbzero.pov.ready_buffer[32]$_SDFFE_PN0P__926  (.L_HI(net926));
 sg13g2_tiehi \rbzero.pov.ready_buffer[33]$_SDFFE_PN0P__927  (.L_HI(net927));
 sg13g2_tiehi \rbzero.pov.ready_buffer[34]$_SDFFE_PN0P__928  (.L_HI(net928));
 sg13g2_tiehi \rbzero.pov.ready_buffer[35]$_SDFFE_PN0P__929  (.L_HI(net929));
 sg13g2_tiehi \rbzero.pov.ready_buffer[36]$_SDFFE_PN0P__930  (.L_HI(net930));
 sg13g2_tiehi \rbzero.pov.ready_buffer[37]$_SDFFE_PN0P__931  (.L_HI(net931));
 sg13g2_tiehi \rbzero.pov.ready_buffer[38]$_SDFFE_PN0P__932  (.L_HI(net932));
 sg13g2_tiehi \rbzero.pov.ready_buffer[39]$_SDFFE_PN0P__933  (.L_HI(net933));
 sg13g2_tiehi \rbzero.pov.ready_buffer[3]$_SDFFE_PN0P__934  (.L_HI(net934));
 sg13g2_tiehi \rbzero.pov.ready_buffer[40]$_SDFFE_PN0P__935  (.L_HI(net935));
 sg13g2_tiehi \rbzero.pov.ready_buffer[41]$_SDFFE_PN0P__936  (.L_HI(net936));
 sg13g2_tiehi \rbzero.pov.ready_buffer[42]$_SDFFE_PN0P__937  (.L_HI(net937));
 sg13g2_tiehi \rbzero.pov.ready_buffer[43]$_SDFFE_PN0P__938  (.L_HI(net938));
 sg13g2_tiehi \rbzero.pov.ready_buffer[44]$_SDFFE_PN0P__939  (.L_HI(net939));
 sg13g2_tiehi \rbzero.pov.ready_buffer[45]$_SDFFE_PN0P__940  (.L_HI(net940));
 sg13g2_tiehi \rbzero.pov.ready_buffer[46]$_SDFFE_PN0P__941  (.L_HI(net941));
 sg13g2_tiehi \rbzero.pov.ready_buffer[47]$_SDFFE_PN0P__942  (.L_HI(net942));
 sg13g2_tiehi \rbzero.pov.ready_buffer[48]$_SDFFE_PN0P__943  (.L_HI(net943));
 sg13g2_tiehi \rbzero.pov.ready_buffer[49]$_SDFFE_PN0P__944  (.L_HI(net944));
 sg13g2_tiehi \rbzero.pov.ready_buffer[4]$_SDFFE_PN0P__945  (.L_HI(net945));
 sg13g2_tiehi \rbzero.pov.ready_buffer[50]$_SDFFE_PN0P__946  (.L_HI(net946));
 sg13g2_tiehi \rbzero.pov.ready_buffer[51]$_SDFFE_PN0P__947  (.L_HI(net947));
 sg13g2_tiehi \rbzero.pov.ready_buffer[52]$_SDFFE_PN0P__948  (.L_HI(net948));
 sg13g2_tiehi \rbzero.pov.ready_buffer[53]$_SDFFE_PN0P__949  (.L_HI(net949));
 sg13g2_tiehi \rbzero.pov.ready_buffer[54]$_SDFFE_PN0P__950  (.L_HI(net950));
 sg13g2_tiehi \rbzero.pov.ready_buffer[55]$_SDFFE_PN0P__951  (.L_HI(net951));
 sg13g2_tiehi \rbzero.pov.ready_buffer[56]$_SDFFE_PN0P__952  (.L_HI(net952));
 sg13g2_tiehi \rbzero.pov.ready_buffer[57]$_SDFFE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \rbzero.pov.ready_buffer[58]$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \rbzero.pov.ready_buffer[59]$_SDFFE_PN0P__955  (.L_HI(net955));
 sg13g2_tiehi \rbzero.pov.ready_buffer[5]$_SDFFE_PN0P__956  (.L_HI(net956));
 sg13g2_tiehi \rbzero.pov.ready_buffer[60]$_SDFFE_PN0P__957  (.L_HI(net957));
 sg13g2_tiehi \rbzero.pov.ready_buffer[61]$_SDFFE_PN0P__958  (.L_HI(net958));
 sg13g2_tiehi \rbzero.pov.ready_buffer[62]$_SDFFE_PN0P__959  (.L_HI(net959));
 sg13g2_tiehi \rbzero.pov.ready_buffer[63]$_SDFFE_PN0P__960  (.L_HI(net960));
 sg13g2_tiehi \rbzero.pov.ready_buffer[64]$_SDFFE_PN0P__961  (.L_HI(net961));
 sg13g2_tiehi \rbzero.pov.ready_buffer[65]$_SDFFE_PN0P__962  (.L_HI(net962));
 sg13g2_tiehi \rbzero.pov.ready_buffer[66]$_SDFFE_PN0P__963  (.L_HI(net963));
 sg13g2_tiehi \rbzero.pov.ready_buffer[67]$_SDFFE_PN0P__964  (.L_HI(net964));
 sg13g2_tiehi \rbzero.pov.ready_buffer[68]$_SDFFE_PN0P__965  (.L_HI(net965));
 sg13g2_tiehi \rbzero.pov.ready_buffer[69]$_SDFFE_PN0P__966  (.L_HI(net966));
 sg13g2_tiehi \rbzero.pov.ready_buffer[6]$_SDFFE_PN0P__967  (.L_HI(net967));
 sg13g2_tiehi \rbzero.pov.ready_buffer[70]$_SDFFE_PN0P__968  (.L_HI(net968));
 sg13g2_tiehi \rbzero.pov.ready_buffer[71]$_SDFFE_PN0P__969  (.L_HI(net969));
 sg13g2_tiehi \rbzero.pov.ready_buffer[72]$_SDFFE_PN0P__970  (.L_HI(net970));
 sg13g2_tiehi \rbzero.pov.ready_buffer[73]$_SDFFE_PN0P__971  (.L_HI(net971));
 sg13g2_tiehi \rbzero.pov.ready_buffer[7]$_SDFFE_PN0P__972  (.L_HI(net972));
 sg13g2_tiehi \rbzero.pov.ready_buffer[8]$_SDFFE_PN0P__973  (.L_HI(net973));
 sg13g2_tiehi \rbzero.pov.ready_buffer[9]$_SDFFE_PN0P__974  (.L_HI(net974));
 sg13g2_tiehi \rbzero.pov.sclk_buffer[0]$_SDFF_PN0__975  (.L_HI(net975));
 sg13g2_tiehi \rbzero.pov.sclk_buffer[1]$_SDFF_PN0__976  (.L_HI(net976));
 sg13g2_tiehi \rbzero.pov.sclk_buffer[2]$_SDFF_PN0__977  (.L_HI(net977));
 sg13g2_tiehi \rbzero.pov.spi_buffer[0]$_SDFFE_PN0P__978  (.L_HI(net978));
 sg13g2_tiehi \rbzero.pov.spi_buffer[10]$_SDFFE_PN0P__979  (.L_HI(net979));
 sg13g2_tiehi \rbzero.pov.spi_buffer[11]$_SDFFE_PN0P__980  (.L_HI(net980));
 sg13g2_tiehi \rbzero.pov.spi_buffer[12]$_SDFFE_PN0P__981  (.L_HI(net981));
 sg13g2_tiehi \rbzero.pov.spi_buffer[13]$_SDFFE_PN0P__982  (.L_HI(net982));
 sg13g2_tiehi \rbzero.pov.spi_buffer[14]$_SDFFE_PN0P__983  (.L_HI(net983));
 sg13g2_tiehi \rbzero.pov.spi_buffer[15]$_SDFFE_PN0P__984  (.L_HI(net984));
 sg13g2_tiehi \rbzero.pov.spi_buffer[16]$_SDFFE_PN0P__985  (.L_HI(net985));
 sg13g2_tiehi \rbzero.pov.spi_buffer[17]$_SDFFE_PN0P__986  (.L_HI(net986));
 sg13g2_tiehi \rbzero.pov.spi_buffer[18]$_SDFFE_PN0P__987  (.L_HI(net987));
 sg13g2_tiehi \rbzero.pov.spi_buffer[19]$_SDFFE_PN0P__988  (.L_HI(net988));
 sg13g2_tiehi \rbzero.pov.spi_buffer[1]$_SDFFE_PN0P__989  (.L_HI(net989));
 sg13g2_tiehi \rbzero.pov.spi_buffer[20]$_SDFFE_PN0P__990  (.L_HI(net990));
 sg13g2_tiehi \rbzero.pov.spi_buffer[21]$_SDFFE_PN0P__991  (.L_HI(net991));
 sg13g2_tiehi \rbzero.pov.spi_buffer[22]$_SDFFE_PN0P__992  (.L_HI(net992));
 sg13g2_tiehi \rbzero.pov.spi_buffer[23]$_SDFFE_PN0P__993  (.L_HI(net993));
 sg13g2_tiehi \rbzero.pov.spi_buffer[24]$_SDFFE_PN0P__994  (.L_HI(net994));
 sg13g2_tiehi \rbzero.pov.spi_buffer[25]$_SDFFE_PN0P__995  (.L_HI(net995));
 sg13g2_tiehi \rbzero.pov.spi_buffer[26]$_SDFFE_PN0P__996  (.L_HI(net996));
 sg13g2_tiehi \rbzero.pov.spi_buffer[27]$_SDFFE_PN0P__997  (.L_HI(net997));
 sg13g2_tiehi \rbzero.pov.spi_buffer[28]$_SDFFE_PN0P__998  (.L_HI(net998));
 sg13g2_tiehi \rbzero.pov.spi_buffer[29]$_SDFFE_PN0P__999  (.L_HI(net999));
 sg13g2_tiehi \rbzero.pov.spi_buffer[2]$_SDFFE_PN0P__1000  (.L_HI(net1000));
 sg13g2_tiehi \rbzero.pov.spi_buffer[30]$_SDFFE_PN0P__1001  (.L_HI(net1001));
 sg13g2_tiehi \rbzero.pov.spi_buffer[31]$_SDFFE_PN0P__1002  (.L_HI(net1002));
 sg13g2_tiehi \rbzero.pov.spi_buffer[32]$_SDFFE_PN0P__1003  (.L_HI(net1003));
 sg13g2_tiehi \rbzero.pov.spi_buffer[33]$_SDFFE_PN0P__1004  (.L_HI(net1004));
 sg13g2_tiehi \rbzero.pov.spi_buffer[34]$_SDFFE_PN0P__1005  (.L_HI(net1005));
 sg13g2_tiehi \rbzero.pov.spi_buffer[35]$_SDFFE_PN0P__1006  (.L_HI(net1006));
 sg13g2_tiehi \rbzero.pov.spi_buffer[36]$_SDFFE_PN0P__1007  (.L_HI(net1007));
 sg13g2_tiehi \rbzero.pov.spi_buffer[37]$_SDFFE_PN0P__1008  (.L_HI(net1008));
 sg13g2_tiehi \rbzero.pov.spi_buffer[38]$_SDFFE_PN0P__1009  (.L_HI(net1009));
 sg13g2_tiehi \rbzero.pov.spi_buffer[39]$_SDFFE_PN0P__1010  (.L_HI(net1010));
 sg13g2_tiehi \rbzero.pov.spi_buffer[3]$_SDFFE_PN0P__1011  (.L_HI(net1011));
 sg13g2_tiehi \rbzero.pov.spi_buffer[40]$_SDFFE_PN0P__1012  (.L_HI(net1012));
 sg13g2_tiehi \rbzero.pov.spi_buffer[41]$_SDFFE_PN0P__1013  (.L_HI(net1013));
 sg13g2_tiehi \rbzero.pov.spi_buffer[42]$_SDFFE_PN0P__1014  (.L_HI(net1014));
 sg13g2_tiehi \rbzero.pov.spi_buffer[43]$_SDFFE_PN0P__1015  (.L_HI(net1015));
 sg13g2_tiehi \rbzero.pov.spi_buffer[44]$_SDFFE_PN0P__1016  (.L_HI(net1016));
 sg13g2_tiehi \rbzero.pov.spi_buffer[45]$_SDFFE_PN0P__1017  (.L_HI(net1017));
 sg13g2_tiehi \rbzero.pov.spi_buffer[46]$_SDFFE_PN0P__1018  (.L_HI(net1018));
 sg13g2_tiehi \rbzero.pov.spi_buffer[47]$_SDFFE_PN0P__1019  (.L_HI(net1019));
 sg13g2_tiehi \rbzero.pov.spi_buffer[48]$_SDFFE_PN0P__1020  (.L_HI(net1020));
 sg13g2_tiehi \rbzero.pov.spi_buffer[49]$_SDFFE_PN0P__1021  (.L_HI(net1021));
 sg13g2_tiehi \rbzero.pov.spi_buffer[4]$_SDFFE_PN0P__1022  (.L_HI(net1022));
 sg13g2_tiehi \rbzero.pov.spi_buffer[50]$_SDFFE_PN0P__1023  (.L_HI(net1023));
 sg13g2_tiehi \rbzero.pov.spi_buffer[51]$_SDFFE_PN0P__1024  (.L_HI(net1024));
 sg13g2_tiehi \rbzero.pov.spi_buffer[52]$_SDFFE_PN0P__1025  (.L_HI(net1025));
 sg13g2_tiehi \rbzero.pov.spi_buffer[53]$_SDFFE_PN0P__1026  (.L_HI(net1026));
 sg13g2_tiehi \rbzero.pov.spi_buffer[54]$_SDFFE_PN0P__1027  (.L_HI(net1027));
 sg13g2_tiehi \rbzero.pov.spi_buffer[55]$_SDFFE_PN0P__1028  (.L_HI(net1028));
 sg13g2_tiehi \rbzero.pov.spi_buffer[56]$_SDFFE_PN0P__1029  (.L_HI(net1029));
 sg13g2_tiehi \rbzero.pov.spi_buffer[57]$_SDFFE_PN0P__1030  (.L_HI(net1030));
 sg13g2_tiehi \rbzero.pov.spi_buffer[58]$_SDFFE_PN0P__1031  (.L_HI(net1031));
 sg13g2_tiehi \rbzero.pov.spi_buffer[59]$_SDFFE_PN0P__1032  (.L_HI(net1032));
 sg13g2_tiehi \rbzero.pov.spi_buffer[5]$_SDFFE_PN0P__1033  (.L_HI(net1033));
 sg13g2_tiehi \rbzero.pov.spi_buffer[60]$_SDFFE_PN0P__1034  (.L_HI(net1034));
 sg13g2_tiehi \rbzero.pov.spi_buffer[61]$_SDFFE_PN0P__1035  (.L_HI(net1035));
 sg13g2_tiehi \rbzero.pov.spi_buffer[62]$_SDFFE_PN0P__1036  (.L_HI(net1036));
 sg13g2_tiehi \rbzero.pov.spi_buffer[63]$_SDFFE_PN0P__1037  (.L_HI(net1037));
 sg13g2_tiehi \rbzero.pov.spi_buffer[64]$_SDFFE_PN0P__1038  (.L_HI(net1038));
 sg13g2_tiehi \rbzero.pov.spi_buffer[65]$_SDFFE_PN0P__1039  (.L_HI(net1039));
 sg13g2_tiehi \rbzero.pov.spi_buffer[66]$_SDFFE_PN0P__1040  (.L_HI(net1040));
 sg13g2_tiehi \rbzero.pov.spi_buffer[67]$_SDFFE_PN0P__1041  (.L_HI(net1041));
 sg13g2_tiehi \rbzero.pov.spi_buffer[68]$_SDFFE_PN0P__1042  (.L_HI(net1042));
 sg13g2_tiehi \rbzero.pov.spi_buffer[69]$_SDFFE_PN0P__1043  (.L_HI(net1043));
 sg13g2_tiehi \rbzero.pov.spi_buffer[6]$_SDFFE_PN0P__1044  (.L_HI(net1044));
 sg13g2_tiehi \rbzero.pov.spi_buffer[70]$_SDFFE_PN0P__1045  (.L_HI(net1045));
 sg13g2_tiehi \rbzero.pov.spi_buffer[71]$_SDFFE_PN0P__1046  (.L_HI(net1046));
 sg13g2_tiehi \rbzero.pov.spi_buffer[72]$_SDFFE_PN0P__1047  (.L_HI(net1047));
 sg13g2_tiehi \rbzero.pov.spi_buffer[73]$_SDFFE_PN0P__1048  (.L_HI(net1048));
 sg13g2_tiehi \rbzero.pov.spi_buffer[7]$_SDFFE_PN0P__1049  (.L_HI(net1049));
 sg13g2_tiehi \rbzero.pov.spi_buffer[8]$_SDFFE_PN0P__1050  (.L_HI(net1050));
 sg13g2_tiehi \rbzero.pov.spi_buffer[9]$_SDFFE_PN0P__1051  (.L_HI(net1051));
 sg13g2_tiehi \rbzero.pov.spi_counter[0]$_SDFFE_PP0N__1052  (.L_HI(net1052));
 sg13g2_tiehi \rbzero.pov.spi_counter[1]$_SDFFE_PP0N__1053  (.L_HI(net1053));
 sg13g2_tiehi \rbzero.pov.spi_counter[2]$_SDFFE_PP0N__1054  (.L_HI(net1054));
 sg13g2_tiehi \rbzero.pov.spi_counter[3]$_SDFFE_PP0N__1055  (.L_HI(net1055));
 sg13g2_tiehi \rbzero.pov.spi_counter[4]$_SDFFE_PP0N__1056  (.L_HI(net1056));
 sg13g2_tiehi \rbzero.pov.spi_counter[5]$_SDFFE_PP0N__1057  (.L_HI(net1057));
 sg13g2_tiehi \rbzero.pov.spi_counter[6]$_SDFFE_PP0N__1058  (.L_HI(net1058));
 sg13g2_tiehi \rbzero.pov.spi_done$_SDFF_PP0__1059  (.L_HI(net1059));
 sg13g2_tiehi \rbzero.pov.ss_buffer[0]$_SDFF_PN0__1060  (.L_HI(net1060));
 sg13g2_tiehi \rbzero.pov.ss_buffer[1]$_SDFF_PN0__1061  (.L_HI(net1061));
 sg13g2_tiehi \rbzero.pov.vplaneRX[0]$_SDFFE_PN1P__1062  (.L_HI(net1062));
 sg13g2_tiehi \rbzero.pov.vplaneRX[10]$_SDFFE_PN0P__1063  (.L_HI(net1063));
 sg13g2_tiehi \rbzero.pov.vplaneRX[1]$_SDFFE_PN0P__1064  (.L_HI(net1064));
 sg13g2_tiehi \rbzero.pov.vplaneRX[2]$_SDFFE_PN0P__1065  (.L_HI(net1065));
 sg13g2_tiehi \rbzero.pov.vplaneRX[3]$_SDFFE_PN0P__1066  (.L_HI(net1066));
 sg13g2_tiehi \rbzero.pov.vplaneRX[4]$_SDFFE_PN1P__1067  (.L_HI(net1067));
 sg13g2_tiehi \rbzero.pov.vplaneRX[5]$_SDFFE_PN1P__1068  (.L_HI(net1068));
 sg13g2_tiehi \rbzero.pov.vplaneRX[6]$_SDFFE_PN0P__1069  (.L_HI(net1069));
 sg13g2_tiehi \rbzero.pov.vplaneRX[7]$_SDFFE_PN1P__1070  (.L_HI(net1070));
 sg13g2_tiehi \rbzero.pov.vplaneRX[8]$_SDFFE_PN0P__1071  (.L_HI(net1071));
 sg13g2_tiehi \rbzero.pov.vplaneRX[9]$_SDFFE_PN0P__1072  (.L_HI(net1072));
 sg13g2_tiehi \rbzero.pov.vplaneRY[0]$_SDFFE_PN0P__1073  (.L_HI(net1073));
 sg13g2_tiehi \rbzero.pov.vplaneRY[10]$_SDFFE_PN0P__1074  (.L_HI(net1074));
 sg13g2_tiehi \rbzero.pov.vplaneRY[1]$_SDFFE_PN0P__1075  (.L_HI(net1075));
 sg13g2_tiehi \rbzero.pov.vplaneRY[2]$_SDFFE_PN0P__1076  (.L_HI(net1076));
 sg13g2_tiehi \rbzero.pov.vplaneRY[3]$_SDFFE_PN1P__1077  (.L_HI(net1077));
 sg13g2_tiehi \rbzero.pov.vplaneRY[4]$_SDFFE_PN1P__1078  (.L_HI(net1078));
 sg13g2_tiehi \rbzero.pov.vplaneRY[5]$_SDFFE_PN1P__1079  (.L_HI(net1079));
 sg13g2_tiehi \rbzero.pov.vplaneRY[6]$_SDFFE_PN0P__1080  (.L_HI(net1080));
 sg13g2_tiehi \rbzero.pov.vplaneRY[7]$_SDFFE_PN1P__1081  (.L_HI(net1081));
 sg13g2_tiehi \rbzero.pov.vplaneRY[8]$_SDFFE_PN0P__1082  (.L_HI(net1082));
 sg13g2_tiehi \rbzero.pov.vplaneRY[9]$_SDFFE_PN0P__1083  (.L_HI(net1083));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[0]$_SDFFE_PN0P__1084  (.L_HI(net1084));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[1]$_SDFFE_PN1P__1085  (.L_HI(net1085));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[2]$_SDFFE_PN0P__1086  (.L_HI(net1086));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[3]$_SDFFE_PN1P__1087  (.L_HI(net1087));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[4]$_SDFFE_PN0P__1088  (.L_HI(net1088));
 sg13g2_tiehi \rbzero.spi_registers.buf_floor[5]$_SDFFE_PN1P__1089  (.L_HI(net1089));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[0]$_SDFFE_PN0P__1090  (.L_HI(net1090));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[1]$_SDFFE_PN0P__1091  (.L_HI(net1091));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[2]$_SDFFE_PN0P__1092  (.L_HI(net1092));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[3]$_SDFFE_PN0P__1093  (.L_HI(net1093));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[4]$_SDFFE_PN0P__1094  (.L_HI(net1094));
 sg13g2_tiehi \rbzero.spi_registers.buf_leak[5]$_SDFFE_PN0P__1095  (.L_HI(net1095));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdx[0]$_SDFFE_PN0P__1096  (.L_HI(net1096));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdx[1]$_SDFFE_PN0P__1097  (.L_HI(net1097));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdx[2]$_SDFFE_PN0P__1098  (.L_HI(net1098));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdx[3]$_SDFFE_PN0P__1099  (.L_HI(net1099));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdx[4]$_SDFFE_PN0P__1100  (.L_HI(net1100));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdxw[0]$_SDFFE_PN0P__1101  (.L_HI(net1101));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdxw[1]$_SDFFE_PN0P__1102  (.L_HI(net1102));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdy[0]$_SDFFE_PN0P__1103  (.L_HI(net1103));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdy[1]$_SDFFE_PN0P__1104  (.L_HI(net1104));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdy[2]$_SDFFE_PN0P__1105  (.L_HI(net1105));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdy[3]$_SDFFE_PN0P__1106  (.L_HI(net1106));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdy[4]$_SDFFE_PN0P__1107  (.L_HI(net1107));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdyw[0]$_SDFFE_PN0P__1108  (.L_HI(net1108));
 sg13g2_tiehi \rbzero.spi_registers.buf_mapdyw[1]$_SDFFE_PN0P__1109  (.L_HI(net1109));
 sg13g2_tiehi \rbzero.spi_registers.buf_otherx[0]$_SDFFE_PN0P__1110  (.L_HI(net1110));
 sg13g2_tiehi \rbzero.spi_registers.buf_otherx[1]$_SDFFE_PN0P__1111  (.L_HI(net1111));
 sg13g2_tiehi \rbzero.spi_registers.buf_otherx[2]$_SDFFE_PN0P__1112  (.L_HI(net1112));
 sg13g2_tiehi \rbzero.spi_registers.buf_otherx[3]$_SDFFE_PN0P__1113  (.L_HI(net1113));
 sg13g2_tiehi \rbzero.spi_registers.buf_otherx[4]$_SDFFE_PN0P__1114  (.L_HI(net1114));
 sg13g2_tiehi \rbzero.spi_registers.buf_othery[0]$_SDFFE_PN0P__1115  (.L_HI(net1115));
 sg13g2_tiehi \rbzero.spi_registers.buf_othery[1]$_SDFFE_PN0P__1116  (.L_HI(net1116));
 sg13g2_tiehi \rbzero.spi_registers.buf_othery[2]$_SDFFE_PN0P__1117  (.L_HI(net1117));
 sg13g2_tiehi \rbzero.spi_registers.buf_othery[3]$_SDFFE_PN0P__1118  (.L_HI(net1118));
 sg13g2_tiehi \rbzero.spi_registers.buf_othery[4]$_SDFFE_PN0P__1119  (.L_HI(net1119));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[0]$_SDFFE_PN1P__1120  (.L_HI(net1120));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[1]$_SDFFE_PN0P__1121  (.L_HI(net1121));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[2]$_SDFFE_PN1P__1122  (.L_HI(net1122));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[3]$_SDFFE_PN0P__1123  (.L_HI(net1123));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[4]$_SDFFE_PN1P__1124  (.L_HI(net1124));
 sg13g2_tiehi \rbzero.spi_registers.buf_sky[5]$_SDFFE_PN0P__1125  (.L_HI(net1125));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[0]$_SDFFE_PN0P__1126  (.L_HI(net1126));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[10]$_SDFFE_PN0P__1127  (.L_HI(net1127));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[11]$_SDFFE_PN0P__1128  (.L_HI(net1128));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[12]$_SDFFE_PN0P__1129  (.L_HI(net1129));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[13]$_SDFFE_PN0P__1130  (.L_HI(net1130));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[14]$_SDFFE_PN0P__1131  (.L_HI(net1131));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[15]$_SDFFE_PN0P__1132  (.L_HI(net1132));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[16]$_SDFFE_PN0P__1133  (.L_HI(net1133));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[17]$_SDFFE_PN0P__1134  (.L_HI(net1134));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[18]$_SDFFE_PN0P__1135  (.L_HI(net1135));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[19]$_SDFFE_PN0P__1136  (.L_HI(net1136));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[1]$_SDFFE_PN0P__1137  (.L_HI(net1137));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[20]$_SDFFE_PN0P__1138  (.L_HI(net1138));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[21]$_SDFFE_PN0P__1139  (.L_HI(net1139));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[22]$_SDFFE_PN0P__1140  (.L_HI(net1140));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[23]$_SDFFE_PN0P__1141  (.L_HI(net1141));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[2]$_SDFFE_PN0P__1142  (.L_HI(net1142));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[3]$_SDFFE_PN0P__1143  (.L_HI(net1143));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[4]$_SDFFE_PN0P__1144  (.L_HI(net1144));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[5]$_SDFFE_PN0P__1145  (.L_HI(net1145));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[6]$_SDFFE_PN0P__1146  (.L_HI(net1146));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[7]$_SDFFE_PN0P__1147  (.L_HI(net1147));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[8]$_SDFFE_PN0P__1148  (.L_HI(net1148));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd0[9]$_SDFFE_PN0P__1149  (.L_HI(net1149));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[0]$_SDFFE_PN0P__1150  (.L_HI(net1150));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[10]$_SDFFE_PN0P__1151  (.L_HI(net1151));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[11]$_SDFFE_PN0P__1152  (.L_HI(net1152));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[12]$_SDFFE_PN0P__1153  (.L_HI(net1153));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[13]$_SDFFE_PN0P__1154  (.L_HI(net1154));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[14]$_SDFFE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[15]$_SDFFE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[16]$_SDFFE_PN0P__1157  (.L_HI(net1157));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[17]$_SDFFE_PN0P__1158  (.L_HI(net1158));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[18]$_SDFFE_PN0P__1159  (.L_HI(net1159));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[19]$_SDFFE_PN0P__1160  (.L_HI(net1160));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[1]$_SDFFE_PN0P__1161  (.L_HI(net1161));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[20]$_SDFFE_PN0P__1162  (.L_HI(net1162));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[21]$_SDFFE_PN0P__1163  (.L_HI(net1163));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[22]$_SDFFE_PN0P__1164  (.L_HI(net1164));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[23]$_SDFFE_PN0P__1165  (.L_HI(net1165));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[2]$_SDFFE_PN0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[3]$_SDFFE_PN0P__1167  (.L_HI(net1167));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[4]$_SDFFE_PN0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[5]$_SDFFE_PN0P__1169  (.L_HI(net1169));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[6]$_SDFFE_PN0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[7]$_SDFFE_PN0P__1171  (.L_HI(net1171));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[8]$_SDFFE_PN0P__1172  (.L_HI(net1172));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd1[9]$_SDFFE_PN0P__1173  (.L_HI(net1173));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[0]$_SDFFE_PN0P__1174  (.L_HI(net1174));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[10]$_SDFFE_PN0P__1175  (.L_HI(net1175));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[11]$_SDFFE_PN0P__1176  (.L_HI(net1176));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[12]$_SDFFE_PN0P__1177  (.L_HI(net1177));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[13]$_SDFFE_PN0P__1178  (.L_HI(net1178));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[14]$_SDFFE_PN0P__1179  (.L_HI(net1179));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[15]$_SDFFE_PN0P__1180  (.L_HI(net1180));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[16]$_SDFFE_PN0P__1181  (.L_HI(net1181));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[17]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[18]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[19]$_SDFFE_PN0P__1184  (.L_HI(net1184));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[1]$_SDFFE_PN0P__1185  (.L_HI(net1185));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[20]$_SDFFE_PN0P__1186  (.L_HI(net1186));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[21]$_SDFFE_PN0P__1187  (.L_HI(net1187));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[22]$_SDFFE_PN0P__1188  (.L_HI(net1188));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[23]$_SDFFE_PN0P__1189  (.L_HI(net1189));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[2]$_SDFFE_PN0P__1190  (.L_HI(net1190));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[3]$_SDFFE_PN0P__1191  (.L_HI(net1191));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[4]$_SDFFE_PN0P__1192  (.L_HI(net1192));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[5]$_SDFFE_PN0P__1193  (.L_HI(net1193));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[6]$_SDFFE_PN0P__1194  (.L_HI(net1194));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[7]$_SDFFE_PN0P__1195  (.L_HI(net1195));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[8]$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd2[9]$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[0]$_SDFFE_PN0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[10]$_SDFFE_PN0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[11]$_SDFFE_PN0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[12]$_SDFFE_PN0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[13]$_SDFFE_PN0P__1202  (.L_HI(net1202));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[14]$_SDFFE_PN0P__1203  (.L_HI(net1203));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[15]$_SDFFE_PN0P__1204  (.L_HI(net1204));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[16]$_SDFFE_PN0P__1205  (.L_HI(net1205));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[17]$_SDFFE_PN0P__1206  (.L_HI(net1206));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[18]$_SDFFE_PN0P__1207  (.L_HI(net1207));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[19]$_SDFFE_PN0P__1208  (.L_HI(net1208));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[1]$_SDFFE_PN0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[20]$_SDFFE_PN0P__1210  (.L_HI(net1210));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[21]$_SDFFE_PN0P__1211  (.L_HI(net1211));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[22]$_SDFFE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[23]$_SDFFE_PN0P__1213  (.L_HI(net1213));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[2]$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[3]$_SDFFE_PN0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[4]$_SDFFE_PN0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[5]$_SDFFE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[6]$_SDFFE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[7]$_SDFFE_PN0P__1219  (.L_HI(net1219));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[8]$_SDFFE_PN0P__1220  (.L_HI(net1220));
 sg13g2_tiehi \rbzero.spi_registers.buf_texadd3[9]$_SDFFE_PN0P__1221  (.L_HI(net1221));
 sg13g2_tiehi \rbzero.spi_registers.buf_vinf$_SDFFE_PN0P__1222  (.L_HI(net1222));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[0]$_SDFFE_PN0P__1223  (.L_HI(net1223));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[1]$_SDFFE_PN0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[2]$_SDFFE_PN0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[3]$_SDFFE_PN0P__1226  (.L_HI(net1226));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[4]$_SDFFE_PN0P__1227  (.L_HI(net1227));
 sg13g2_tiehi \rbzero.spi_registers.buf_vshift[5]$_SDFFE_PN0P__1228  (.L_HI(net1228));
 sg13g2_tiehi \rbzero.spi_registers.floor[0]$_SDFFE_PN0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \rbzero.spi_registers.floor[1]$_SDFFE_PN1P__1230  (.L_HI(net1230));
 sg13g2_tiehi \rbzero.spi_registers.floor[2]$_SDFFE_PN0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \rbzero.spi_registers.floor[3]$_SDFFE_PN1P__1232  (.L_HI(net1232));
 sg13g2_tiehi \rbzero.spi_registers.floor[4]$_SDFFE_PN0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \rbzero.spi_registers.floor[5]$_SDFFE_PN1P__1234  (.L_HI(net1234));
 sg13g2_tiehi \rbzero.spi_registers.leak[0]$_SDFFE_PN0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \rbzero.spi_registers.leak[1]$_SDFFE_PN0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \rbzero.spi_registers.leak[2]$_SDFFE_PN0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \rbzero.spi_registers.leak[3]$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \rbzero.spi_registers.leak[4]$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \rbzero.spi_registers.leak[5]$_SDFFE_PN0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \rbzero.spi_registers.mapdx[0]$_SDFFE_PN0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \rbzero.spi_registers.mapdx[1]$_SDFFE_PN0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \rbzero.spi_registers.mapdx[2]$_SDFFE_PN0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \rbzero.spi_registers.mapdx[3]$_SDFFE_PN0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \rbzero.spi_registers.mapdx[4]$_SDFFE_PN0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \rbzero.spi_registers.mapdxw[0]$_SDFFE_PN0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \rbzero.spi_registers.mapdxw[1]$_SDFFE_PN0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \rbzero.spi_registers.mapdy[0]$_SDFFE_PN0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \rbzero.spi_registers.mapdy[1]$_SDFFE_PN0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \rbzero.spi_registers.mapdy[2]$_SDFFE_PN0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \rbzero.spi_registers.mapdy[3]$_SDFFE_PN0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \rbzero.spi_registers.mapdy[4]$_SDFFE_PN0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \rbzero.spi_registers.mapdyw[0]$_SDFFE_PN0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \rbzero.spi_registers.mapdyw[1]$_SDFFE_PN0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \rbzero.spi_registers.mosi_buffer[0]$_SDFF_PN0__1255  (.L_HI(net1255));
 sg13g2_tiehi \rbzero.spi_registers.mosi_buffer[1]$_SDFF_PN0__1256  (.L_HI(net1256));
 sg13g2_tiehi \rbzero.spi_registers.otherx[0]$_SDFFE_PN0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \rbzero.spi_registers.otherx[1]$_SDFFE_PN0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \rbzero.spi_registers.otherx[2]$_SDFFE_PN0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \rbzero.spi_registers.otherx[3]$_SDFFE_PN0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \rbzero.spi_registers.otherx[4]$_SDFFE_PN0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \rbzero.spi_registers.othery[0]$_SDFFE_PN0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \rbzero.spi_registers.othery[1]$_SDFFE_PN0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \rbzero.spi_registers.othery[2]$_SDFFE_PN0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \rbzero.spi_registers.othery[3]$_SDFFE_PN0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \rbzero.spi_registers.othery[4]$_SDFFE_PN0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \rbzero.spi_registers.sclk_buffer[0]$_SDFF_PN0__1267  (.L_HI(net1267));
 sg13g2_tiehi \rbzero.spi_registers.sclk_buffer[1]$_SDFF_PN0__1268  (.L_HI(net1268));
 sg13g2_tiehi \rbzero.spi_registers.sclk_buffer[2]$_SDFF_PN0__1269  (.L_HI(net1269));
 sg13g2_tiehi \rbzero.spi_registers.sky[0]$_SDFFE_PN1P__1270  (.L_HI(net1270));
 sg13g2_tiehi \rbzero.spi_registers.sky[1]$_SDFFE_PN0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \rbzero.spi_registers.sky[2]$_SDFFE_PN1P__1272  (.L_HI(net1272));
 sg13g2_tiehi \rbzero.spi_registers.sky[3]$_SDFFE_PN0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \rbzero.spi_registers.sky[4]$_SDFFE_PN1P__1274  (.L_HI(net1274));
 sg13g2_tiehi \rbzero.spi_registers.sky[5]$_SDFFE_PN0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[0]$_SDFFE_PN0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[10]$_SDFFE_PN0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[11]$_SDFFE_PN0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[12]$_SDFFE_PN0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[13]$_SDFFE_PN0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[14]$_SDFFE_PN0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[15]$_SDFFE_PN0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[16]$_SDFFE_PN0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[17]$_SDFFE_PN0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[18]$_SDFFE_PN0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[19]$_SDFFE_PN0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[1]$_SDFFE_PN0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[20]$_SDFFE_PN0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[21]$_SDFFE_PN0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[22]$_SDFFE_PN0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[23]$_SDFFE_PN0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[2]$_SDFFE_PN0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[3]$_SDFFE_PN0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[4]$_SDFFE_PN0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[5]$_SDFFE_PN0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[6]$_SDFFE_PN0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[7]$_SDFFE_PN0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[8]$_SDFFE_PN0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \rbzero.spi_registers.spi_buffer[9]$_SDFFE_PN0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \rbzero.spi_registers.spi_cmd[0]$_SDFFE_PP0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \rbzero.spi_registers.spi_cmd[1]$_SDFFE_PP0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \rbzero.spi_registers.spi_cmd[2]$_SDFFE_PP0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \rbzero.spi_registers.spi_cmd[3]$_SDFFE_PP0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[0]$_SDFFE_PP0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[1]$_SDFFE_PP0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[2]$_SDFFE_PP0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[3]$_SDFFE_PP0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[4]$_SDFFE_PP0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[5]$_SDFFE_PP0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \rbzero.spi_registers.spi_counter[6]$_SDFFE_PP0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \rbzero.spi_registers.spi_done$_SDFF_PP0__1311  (.L_HI(net1311));
 sg13g2_tiehi \rbzero.spi_registers.ss_buffer[0]$_SDFF_PN0__1312  (.L_HI(net1312));
 sg13g2_tiehi \rbzero.spi_registers.ss_buffer[1]$_SDFF_PN0__1313  (.L_HI(net1313));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[0]$_SDFFE_PN0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[10]$_SDFFE_PN0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[11]$_SDFFE_PN0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[12]$_SDFFE_PN0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[13]$_SDFFE_PN0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[14]$_SDFFE_PN0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[15]$_SDFFE_PN0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[16]$_SDFFE_PN0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[17]$_SDFFE_PN0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[18]$_SDFFE_PN0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[19]$_SDFFE_PN0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[1]$_SDFFE_PN0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[20]$_SDFFE_PN0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[21]$_SDFFE_PN0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[22]$_SDFFE_PN0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[23]$_SDFFE_PN0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[2]$_SDFFE_PN0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[3]$_SDFFE_PN0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[4]$_SDFFE_PN0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[5]$_SDFFE_PN0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[6]$_SDFFE_PN0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[7]$_SDFFE_PN0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[8]$_SDFFE_PN0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \rbzero.spi_registers.texadd0[9]$_SDFFE_PN0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[0]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[10]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[11]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[12]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[13]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[14]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[15]$_SDFFE_PN0P__1344  (.L_HI(net1344));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[16]$_SDFFE_PN0P__1345  (.L_HI(net1345));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[17]$_SDFFE_PN0P__1346  (.L_HI(net1346));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[18]$_SDFFE_PN0P__1347  (.L_HI(net1347));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[19]$_SDFFE_PN0P__1348  (.L_HI(net1348));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[1]$_SDFFE_PN0P__1349  (.L_HI(net1349));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[20]$_SDFFE_PN0P__1350  (.L_HI(net1350));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[21]$_SDFFE_PN0P__1351  (.L_HI(net1351));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[22]$_SDFFE_PN0P__1352  (.L_HI(net1352));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[23]$_SDFFE_PN0P__1353  (.L_HI(net1353));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[2]$_SDFFE_PN0P__1354  (.L_HI(net1354));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[3]$_SDFFE_PN0P__1355  (.L_HI(net1355));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[4]$_SDFFE_PN0P__1356  (.L_HI(net1356));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[5]$_SDFFE_PN0P__1357  (.L_HI(net1357));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[6]$_SDFFE_PN0P__1358  (.L_HI(net1358));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[7]$_SDFFE_PN0P__1359  (.L_HI(net1359));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[8]$_SDFFE_PN0P__1360  (.L_HI(net1360));
 sg13g2_tiehi \rbzero.spi_registers.texadd1[9]$_SDFFE_PN0P__1361  (.L_HI(net1361));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[0]$_SDFFE_PN0P__1362  (.L_HI(net1362));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[10]$_SDFFE_PN0P__1363  (.L_HI(net1363));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[11]$_SDFFE_PN0P__1364  (.L_HI(net1364));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[12]$_SDFFE_PN0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[13]$_SDFFE_PN0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[14]$_SDFFE_PN0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[15]$_SDFFE_PN0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[16]$_SDFFE_PN0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[17]$_SDFFE_PN0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[18]$_SDFFE_PN0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[19]$_SDFFE_PN0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[1]$_SDFFE_PN0P__1373  (.L_HI(net1373));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[20]$_SDFFE_PN0P__1374  (.L_HI(net1374));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[21]$_SDFFE_PN0P__1375  (.L_HI(net1375));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[22]$_SDFFE_PN0P__1376  (.L_HI(net1376));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[23]$_SDFFE_PN0P__1377  (.L_HI(net1377));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[2]$_SDFFE_PN0P__1378  (.L_HI(net1378));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[3]$_SDFFE_PN0P__1379  (.L_HI(net1379));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[4]$_SDFFE_PN0P__1380  (.L_HI(net1380));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[5]$_SDFFE_PN0P__1381  (.L_HI(net1381));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[6]$_SDFFE_PN0P__1382  (.L_HI(net1382));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[7]$_SDFFE_PN0P__1383  (.L_HI(net1383));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[8]$_SDFFE_PN0P__1384  (.L_HI(net1384));
 sg13g2_tiehi \rbzero.spi_registers.texadd2[9]$_SDFFE_PN0P__1385  (.L_HI(net1385));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[0]$_SDFFE_PN0P__1386  (.L_HI(net1386));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[10]$_SDFFE_PN0P__1387  (.L_HI(net1387));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[11]$_SDFFE_PN0P__1388  (.L_HI(net1388));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[12]$_SDFFE_PN0P__1389  (.L_HI(net1389));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[13]$_SDFFE_PN0P__1390  (.L_HI(net1390));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[14]$_SDFFE_PN0P__1391  (.L_HI(net1391));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[15]$_SDFFE_PN0P__1392  (.L_HI(net1392));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[16]$_SDFFE_PN0P__1393  (.L_HI(net1393));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[17]$_SDFFE_PN0P__1394  (.L_HI(net1394));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[18]$_SDFFE_PN0P__1395  (.L_HI(net1395));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[19]$_SDFFE_PN0P__1396  (.L_HI(net1396));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[1]$_SDFFE_PN0P__1397  (.L_HI(net1397));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[20]$_SDFFE_PN0P__1398  (.L_HI(net1398));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[21]$_SDFFE_PN0P__1399  (.L_HI(net1399));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[22]$_SDFFE_PN0P__1400  (.L_HI(net1400));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[23]$_SDFFE_PN0P__1401  (.L_HI(net1401));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[2]$_SDFFE_PN0P__1402  (.L_HI(net1402));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[3]$_SDFFE_PN0P__1403  (.L_HI(net1403));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[4]$_SDFFE_PN0P__1404  (.L_HI(net1404));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[5]$_SDFFE_PN0P__1405  (.L_HI(net1405));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[6]$_SDFFE_PN0P__1406  (.L_HI(net1406));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[7]$_SDFFE_PN0P__1407  (.L_HI(net1407));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[8]$_SDFFE_PN0P__1408  (.L_HI(net1408));
 sg13g2_tiehi \rbzero.spi_registers.texadd3[9]$_SDFFE_PN0P__1409  (.L_HI(net1409));
 sg13g2_tiehi \rbzero.spi_registers.vinf$_SDFFE_PN0P__1410  (.L_HI(net1410));
 sg13g2_tiehi \rbzero.spi_registers.vshift[0]$_SDFFE_PN0P__1411  (.L_HI(net1411));
 sg13g2_tiehi \rbzero.spi_registers.vshift[1]$_SDFFE_PN0P__1412  (.L_HI(net1412));
 sg13g2_tiehi \rbzero.spi_registers.vshift[2]$_SDFFE_PN0P__1413  (.L_HI(net1413));
 sg13g2_tiehi \rbzero.spi_registers.vshift[3]$_SDFFE_PN0P__1414  (.L_HI(net1414));
 sg13g2_tiehi \rbzero.spi_registers.vshift[4]$_SDFFE_PN0P__1415  (.L_HI(net1415));
 sg13g2_tiehi \rbzero.spi_registers.vshift[5]$_SDFFE_PN0P__1416  (.L_HI(net1416));
 sg13g2_tiehi \rbzero.texV[0]$_SDFF_PP0__1417  (.L_HI(net1417));
 sg13g2_tiehi \rbzero.texV[10]$_SDFF_PP0__1418  (.L_HI(net1418));
 sg13g2_tiehi \rbzero.texV[11]$_SDFF_PP0__1419  (.L_HI(net1419));
 sg13g2_tiehi \rbzero.texV[12]$_SDFF_PP0__1420  (.L_HI(net1420));
 sg13g2_tiehi \rbzero.texV[13]$_SDFF_PP0__1421  (.L_HI(net1421));
 sg13g2_tiehi \rbzero.texV[14]$_SDFF_PP0__1422  (.L_HI(net1422));
 sg13g2_tiehi \rbzero.texV[15]$_SDFF_PP0__1423  (.L_HI(net1423));
 sg13g2_tiehi \rbzero.texV[16]$_SDFF_PP0__1424  (.L_HI(net1424));
 sg13g2_tiehi \rbzero.texV[17]$_SDFF_PP0__1425  (.L_HI(net1425));
 sg13g2_tiehi \rbzero.texV[18]$_SDFF_PP0__1426  (.L_HI(net1426));
 sg13g2_tiehi \rbzero.texV[19]$_SDFF_PP0__1427  (.L_HI(net1427));
 sg13g2_tiehi \rbzero.texV[1]$_SDFF_PP0__1428  (.L_HI(net1428));
 sg13g2_tiehi \rbzero.texV[20]$_SDFF_PP0__1429  (.L_HI(net1429));
 sg13g2_tiehi \rbzero.texV[21]$_SDFF_PP0__1430  (.L_HI(net1430));
 sg13g2_tiehi \rbzero.texV[2]$_SDFF_PP0__1431  (.L_HI(net1431));
 sg13g2_tiehi \rbzero.texV[3]$_SDFF_PP0__1432  (.L_HI(net1432));
 sg13g2_tiehi \rbzero.texV[4]$_SDFF_PP0__1433  (.L_HI(net1433));
 sg13g2_tiehi \rbzero.texV[5]$_SDFF_PP0__1434  (.L_HI(net1434));
 sg13g2_tiehi \rbzero.texV[6]$_SDFF_PP0__1435  (.L_HI(net1435));
 sg13g2_tiehi \rbzero.texV[7]$_SDFF_PP0__1436  (.L_HI(net1436));
 sg13g2_tiehi \rbzero.texV[8]$_SDFF_PP0__1437  (.L_HI(net1437));
 sg13g2_tiehi \rbzero.texV[9]$_SDFF_PP0__1438  (.L_HI(net1438));
 sg13g2_tiehi \rbzero.tex_b0[0]$_DFFE_NP__1439  (.L_HI(net1439));
 sg13g2_tiehi \rbzero.tex_b0[10]$_DFFE_NP__1440  (.L_HI(net1440));
 sg13g2_tiehi \rbzero.tex_b0[11]$_DFFE_NP__1441  (.L_HI(net1441));
 sg13g2_tiehi \rbzero.tex_b0[12]$_DFFE_NP__1442  (.L_HI(net1442));
 sg13g2_tiehi \rbzero.tex_b0[13]$_DFFE_NP__1443  (.L_HI(net1443));
 sg13g2_tiehi \rbzero.tex_b0[14]$_DFFE_NP__1444  (.L_HI(net1444));
 sg13g2_tiehi \rbzero.tex_b0[15]$_DFFE_NP__1445  (.L_HI(net1445));
 sg13g2_tiehi \rbzero.tex_b0[16]$_DFFE_NP__1446  (.L_HI(net1446));
 sg13g2_tiehi \rbzero.tex_b0[17]$_DFFE_NP__1447  (.L_HI(net1447));
 sg13g2_tiehi \rbzero.tex_b0[18]$_DFFE_NP__1448  (.L_HI(net1448));
 sg13g2_tiehi \rbzero.tex_b0[19]$_DFFE_NP__1449  (.L_HI(net1449));
 sg13g2_tiehi \rbzero.tex_b0[1]$_DFFE_NP__1450  (.L_HI(net1450));
 sg13g2_tiehi \rbzero.tex_b0[20]$_DFFE_NP__1451  (.L_HI(net1451));
 sg13g2_tiehi \rbzero.tex_b0[21]$_DFFE_NP__1452  (.L_HI(net1452));
 sg13g2_tiehi \rbzero.tex_b0[22]$_DFFE_NP__1453  (.L_HI(net1453));
 sg13g2_tiehi \rbzero.tex_b0[23]$_DFFE_NP__1454  (.L_HI(net1454));
 sg13g2_tiehi \rbzero.tex_b0[24]$_DFFE_NP__1455  (.L_HI(net1455));
 sg13g2_tiehi \rbzero.tex_b0[25]$_DFFE_NP__1456  (.L_HI(net1456));
 sg13g2_tiehi \rbzero.tex_b0[26]$_DFFE_NP__1457  (.L_HI(net1457));
 sg13g2_tiehi \rbzero.tex_b0[27]$_DFFE_NP__1458  (.L_HI(net1458));
 sg13g2_tiehi \rbzero.tex_b0[28]$_DFFE_NP__1459  (.L_HI(net1459));
 sg13g2_tiehi \rbzero.tex_b0[29]$_DFFE_NP__1460  (.L_HI(net1460));
 sg13g2_tiehi \rbzero.tex_b0[2]$_DFFE_NP__1461  (.L_HI(net1461));
 sg13g2_tiehi \rbzero.tex_b0[30]$_DFFE_NP__1462  (.L_HI(net1462));
 sg13g2_tiehi \rbzero.tex_b0[31]$_DFFE_NP__1463  (.L_HI(net1463));
 sg13g2_tiehi \rbzero.tex_b0[32]$_DFFE_NP__1464  (.L_HI(net1464));
 sg13g2_tiehi \rbzero.tex_b0[33]$_DFFE_NP__1465  (.L_HI(net1465));
 sg13g2_tiehi \rbzero.tex_b0[34]$_DFFE_NP__1466  (.L_HI(net1466));
 sg13g2_tiehi \rbzero.tex_b0[35]$_DFFE_NP__1467  (.L_HI(net1467));
 sg13g2_tiehi \rbzero.tex_b0[36]$_DFFE_NP__1468  (.L_HI(net1468));
 sg13g2_tiehi \rbzero.tex_b0[37]$_DFFE_NP__1469  (.L_HI(net1469));
 sg13g2_tiehi \rbzero.tex_b0[38]$_DFFE_NP__1470  (.L_HI(net1470));
 sg13g2_tiehi \rbzero.tex_b0[39]$_DFFE_NP__1471  (.L_HI(net1471));
 sg13g2_tiehi \rbzero.tex_b0[3]$_DFFE_NP__1472  (.L_HI(net1472));
 sg13g2_tiehi \rbzero.tex_b0[40]$_DFFE_NP__1473  (.L_HI(net1473));
 sg13g2_tiehi \rbzero.tex_b0[41]$_DFFE_NP__1474  (.L_HI(net1474));
 sg13g2_tiehi \rbzero.tex_b0[42]$_DFFE_NP__1475  (.L_HI(net1475));
 sg13g2_tiehi \rbzero.tex_b0[43]$_DFFE_NP__1476  (.L_HI(net1476));
 sg13g2_tiehi \rbzero.tex_b0[44]$_DFFE_NP__1477  (.L_HI(net1477));
 sg13g2_tiehi \rbzero.tex_b0[45]$_DFFE_NP__1478  (.L_HI(net1478));
 sg13g2_tiehi \rbzero.tex_b0[46]$_DFFE_NP__1479  (.L_HI(net1479));
 sg13g2_tiehi \rbzero.tex_b0[47]$_DFFE_NP__1480  (.L_HI(net1480));
 sg13g2_tiehi \rbzero.tex_b0[48]$_DFFE_NP__1481  (.L_HI(net1481));
 sg13g2_tiehi \rbzero.tex_b0[49]$_DFFE_NP__1482  (.L_HI(net1482));
 sg13g2_tiehi \rbzero.tex_b0[4]$_DFFE_NP__1483  (.L_HI(net1483));
 sg13g2_tiehi \rbzero.tex_b0[50]$_DFFE_NP__1484  (.L_HI(net1484));
 sg13g2_tiehi \rbzero.tex_b0[51]$_DFFE_NP__1485  (.L_HI(net1485));
 sg13g2_tiehi \rbzero.tex_b0[52]$_DFFE_NP__1486  (.L_HI(net1486));
 sg13g2_tiehi \rbzero.tex_b0[53]$_DFFE_NP__1487  (.L_HI(net1487));
 sg13g2_tiehi \rbzero.tex_b0[54]$_DFFE_NP__1488  (.L_HI(net1488));
 sg13g2_tiehi \rbzero.tex_b0[55]$_DFFE_NP__1489  (.L_HI(net1489));
 sg13g2_tiehi \rbzero.tex_b0[56]$_DFFE_NP__1490  (.L_HI(net1490));
 sg13g2_tiehi \rbzero.tex_b0[57]$_DFFE_NP__1491  (.L_HI(net1491));
 sg13g2_tiehi \rbzero.tex_b0[58]$_DFFE_NP__1492  (.L_HI(net1492));
 sg13g2_tiehi \rbzero.tex_b0[59]$_DFFE_NP__1493  (.L_HI(net1493));
 sg13g2_tiehi \rbzero.tex_b0[5]$_DFFE_NP__1494  (.L_HI(net1494));
 sg13g2_tiehi \rbzero.tex_b0[60]$_DFFE_NP__1495  (.L_HI(net1495));
 sg13g2_tiehi \rbzero.tex_b0[61]$_DFFE_NP__1496  (.L_HI(net1496));
 sg13g2_tiehi \rbzero.tex_b0[62]$_DFFE_NP__1497  (.L_HI(net1497));
 sg13g2_tiehi \rbzero.tex_b0[63]$_DFFE_NP__1498  (.L_HI(net1498));
 sg13g2_tiehi \rbzero.tex_b0[6]$_DFFE_NP__1499  (.L_HI(net1499));
 sg13g2_tiehi \rbzero.tex_b0[7]$_DFFE_NP__1500  (.L_HI(net1500));
 sg13g2_tiehi \rbzero.tex_b0[8]$_DFFE_NP__1501  (.L_HI(net1501));
 sg13g2_tiehi \rbzero.tex_b0[9]$_DFFE_NP__1502  (.L_HI(net1502));
 sg13g2_tiehi \rbzero.tex_b1[0]$_DFFE_NP__1503  (.L_HI(net1503));
 sg13g2_tiehi \rbzero.tex_b1[10]$_DFFE_NP__1504  (.L_HI(net1504));
 sg13g2_tiehi \rbzero.tex_b1[11]$_DFFE_NP__1505  (.L_HI(net1505));
 sg13g2_tiehi \rbzero.tex_b1[12]$_DFFE_NP__1506  (.L_HI(net1506));
 sg13g2_tiehi \rbzero.tex_b1[13]$_DFFE_NP__1507  (.L_HI(net1507));
 sg13g2_tiehi \rbzero.tex_b1[14]$_DFFE_NP__1508  (.L_HI(net1508));
 sg13g2_tiehi \rbzero.tex_b1[15]$_DFFE_NP__1509  (.L_HI(net1509));
 sg13g2_tiehi \rbzero.tex_b1[16]$_DFFE_NP__1510  (.L_HI(net1510));
 sg13g2_tiehi \rbzero.tex_b1[17]$_DFFE_NP__1511  (.L_HI(net1511));
 sg13g2_tiehi \rbzero.tex_b1[18]$_DFFE_NP__1512  (.L_HI(net1512));
 sg13g2_tiehi \rbzero.tex_b1[19]$_DFFE_NP__1513  (.L_HI(net1513));
 sg13g2_tiehi \rbzero.tex_b1[1]$_DFFE_NP__1514  (.L_HI(net1514));
 sg13g2_tiehi \rbzero.tex_b1[20]$_DFFE_NP__1515  (.L_HI(net1515));
 sg13g2_tiehi \rbzero.tex_b1[21]$_DFFE_NP__1516  (.L_HI(net1516));
 sg13g2_tiehi \rbzero.tex_b1[22]$_DFFE_NP__1517  (.L_HI(net1517));
 sg13g2_tiehi \rbzero.tex_b1[23]$_DFFE_NP__1518  (.L_HI(net1518));
 sg13g2_tiehi \rbzero.tex_b1[24]$_DFFE_NP__1519  (.L_HI(net1519));
 sg13g2_tiehi \rbzero.tex_b1[25]$_DFFE_NP__1520  (.L_HI(net1520));
 sg13g2_tiehi \rbzero.tex_b1[26]$_DFFE_NP__1521  (.L_HI(net1521));
 sg13g2_tiehi \rbzero.tex_b1[27]$_DFFE_NP__1522  (.L_HI(net1522));
 sg13g2_tiehi \rbzero.tex_b1[28]$_DFFE_NP__1523  (.L_HI(net1523));
 sg13g2_tiehi \rbzero.tex_b1[29]$_DFFE_NP__1524  (.L_HI(net1524));
 sg13g2_tiehi \rbzero.tex_b1[2]$_DFFE_NP__1525  (.L_HI(net1525));
 sg13g2_tiehi \rbzero.tex_b1[30]$_DFFE_NP__1526  (.L_HI(net1526));
 sg13g2_tiehi \rbzero.tex_b1[31]$_DFFE_NP__1527  (.L_HI(net1527));
 sg13g2_tiehi \rbzero.tex_b1[32]$_DFFE_NP__1528  (.L_HI(net1528));
 sg13g2_tiehi \rbzero.tex_b1[33]$_DFFE_NP__1529  (.L_HI(net1529));
 sg13g2_tiehi \rbzero.tex_b1[34]$_DFFE_NP__1530  (.L_HI(net1530));
 sg13g2_tiehi \rbzero.tex_b1[35]$_DFFE_NP__1531  (.L_HI(net1531));
 sg13g2_tiehi \rbzero.tex_b1[36]$_DFFE_NP__1532  (.L_HI(net1532));
 sg13g2_tiehi \rbzero.tex_b1[37]$_DFFE_NP__1533  (.L_HI(net1533));
 sg13g2_tiehi \rbzero.tex_b1[38]$_DFFE_NP__1534  (.L_HI(net1534));
 sg13g2_tiehi \rbzero.tex_b1[39]$_DFFE_NP__1535  (.L_HI(net1535));
 sg13g2_tiehi \rbzero.tex_b1[3]$_DFFE_NP__1536  (.L_HI(net1536));
 sg13g2_tiehi \rbzero.tex_b1[40]$_DFFE_NP__1537  (.L_HI(net1537));
 sg13g2_tiehi \rbzero.tex_b1[41]$_DFFE_NP__1538  (.L_HI(net1538));
 sg13g2_tiehi \rbzero.tex_b1[42]$_DFFE_NP__1539  (.L_HI(net1539));
 sg13g2_tiehi \rbzero.tex_b1[43]$_DFFE_NP__1540  (.L_HI(net1540));
 sg13g2_tiehi \rbzero.tex_b1[44]$_DFFE_NP__1541  (.L_HI(net1541));
 sg13g2_tiehi \rbzero.tex_b1[45]$_DFFE_NP__1542  (.L_HI(net1542));
 sg13g2_tiehi \rbzero.tex_b1[46]$_DFFE_NP__1543  (.L_HI(net1543));
 sg13g2_tiehi \rbzero.tex_b1[47]$_DFFE_NP__1544  (.L_HI(net1544));
 sg13g2_tiehi \rbzero.tex_b1[48]$_DFFE_NP__1545  (.L_HI(net1545));
 sg13g2_tiehi \rbzero.tex_b1[49]$_DFFE_NP__1546  (.L_HI(net1546));
 sg13g2_tiehi \rbzero.tex_b1[4]$_DFFE_NP__1547  (.L_HI(net1547));
 sg13g2_tiehi \rbzero.tex_b1[50]$_DFFE_NP__1548  (.L_HI(net1548));
 sg13g2_tiehi \rbzero.tex_b1[51]$_DFFE_NP__1549  (.L_HI(net1549));
 sg13g2_tiehi \rbzero.tex_b1[52]$_DFFE_NP__1550  (.L_HI(net1550));
 sg13g2_tiehi \rbzero.tex_b1[53]$_DFFE_NP__1551  (.L_HI(net1551));
 sg13g2_tiehi \rbzero.tex_b1[54]$_DFFE_NP__1552  (.L_HI(net1552));
 sg13g2_tiehi \rbzero.tex_b1[55]$_DFFE_NP__1553  (.L_HI(net1553));
 sg13g2_tiehi \rbzero.tex_b1[56]$_DFFE_NP__1554  (.L_HI(net1554));
 sg13g2_tiehi \rbzero.tex_b1[57]$_DFFE_NP__1555  (.L_HI(net1555));
 sg13g2_tiehi \rbzero.tex_b1[58]$_DFFE_NP__1556  (.L_HI(net1556));
 sg13g2_tiehi \rbzero.tex_b1[59]$_DFFE_NP__1557  (.L_HI(net1557));
 sg13g2_tiehi \rbzero.tex_b1[5]$_DFFE_NP__1558  (.L_HI(net1558));
 sg13g2_tiehi \rbzero.tex_b1[60]$_DFFE_NP__1559  (.L_HI(net1559));
 sg13g2_tiehi \rbzero.tex_b1[61]$_DFFE_NP__1560  (.L_HI(net1560));
 sg13g2_tiehi \rbzero.tex_b1[62]$_DFFE_NP__1561  (.L_HI(net1561));
 sg13g2_tiehi \rbzero.tex_b1[63]$_DFFE_NP__1562  (.L_HI(net1562));
 sg13g2_tiehi \rbzero.tex_b1[6]$_DFFE_NP__1563  (.L_HI(net1563));
 sg13g2_tiehi \rbzero.tex_b1[7]$_DFFE_NP__1564  (.L_HI(net1564));
 sg13g2_tiehi \rbzero.tex_b1[8]$_DFFE_NP__1565  (.L_HI(net1565));
 sg13g2_tiehi \rbzero.tex_b1[9]$_DFFE_NP__1566  (.L_HI(net1566));
 sg13g2_tiehi \rbzero.tex_g0[0]$_DFFE_NP__1567  (.L_HI(net1567));
 sg13g2_tiehi \rbzero.tex_g0[10]$_DFFE_NP__1568  (.L_HI(net1568));
 sg13g2_tiehi \rbzero.tex_g0[11]$_DFFE_NP__1569  (.L_HI(net1569));
 sg13g2_tiehi \rbzero.tex_g0[12]$_DFFE_NP__1570  (.L_HI(net1570));
 sg13g2_tiehi \rbzero.tex_g0[13]$_DFFE_NP__1571  (.L_HI(net1571));
 sg13g2_tiehi \rbzero.tex_g0[14]$_DFFE_NP__1572  (.L_HI(net1572));
 sg13g2_tiehi \rbzero.tex_g0[15]$_DFFE_NP__1573  (.L_HI(net1573));
 sg13g2_tiehi \rbzero.tex_g0[16]$_DFFE_NP__1574  (.L_HI(net1574));
 sg13g2_tiehi \rbzero.tex_g0[17]$_DFFE_NP__1575  (.L_HI(net1575));
 sg13g2_tiehi \rbzero.tex_g0[18]$_DFFE_NP__1576  (.L_HI(net1576));
 sg13g2_tiehi \rbzero.tex_g0[19]$_DFFE_NP__1577  (.L_HI(net1577));
 sg13g2_tiehi \rbzero.tex_g0[1]$_DFFE_NP__1578  (.L_HI(net1578));
 sg13g2_tiehi \rbzero.tex_g0[20]$_DFFE_NP__1579  (.L_HI(net1579));
 sg13g2_tiehi \rbzero.tex_g0[21]$_DFFE_NP__1580  (.L_HI(net1580));
 sg13g2_tiehi \rbzero.tex_g0[22]$_DFFE_NP__1581  (.L_HI(net1581));
 sg13g2_tiehi \rbzero.tex_g0[23]$_DFFE_NP__1582  (.L_HI(net1582));
 sg13g2_tiehi \rbzero.tex_g0[24]$_DFFE_NP__1583  (.L_HI(net1583));
 sg13g2_tiehi \rbzero.tex_g0[25]$_DFFE_NP__1584  (.L_HI(net1584));
 sg13g2_tiehi \rbzero.tex_g0[26]$_DFFE_NP__1585  (.L_HI(net1585));
 sg13g2_tiehi \rbzero.tex_g0[27]$_DFFE_NP__1586  (.L_HI(net1586));
 sg13g2_tiehi \rbzero.tex_g0[28]$_DFFE_NP__1587  (.L_HI(net1587));
 sg13g2_tiehi \rbzero.tex_g0[29]$_DFFE_NP__1588  (.L_HI(net1588));
 sg13g2_tiehi \rbzero.tex_g0[2]$_DFFE_NP__1589  (.L_HI(net1589));
 sg13g2_tiehi \rbzero.tex_g0[30]$_DFFE_NP__1590  (.L_HI(net1590));
 sg13g2_tiehi \rbzero.tex_g0[31]$_DFFE_NP__1591  (.L_HI(net1591));
 sg13g2_tiehi \rbzero.tex_g0[32]$_DFFE_NP__1592  (.L_HI(net1592));
 sg13g2_tiehi \rbzero.tex_g0[33]$_DFFE_NP__1593  (.L_HI(net1593));
 sg13g2_tiehi \rbzero.tex_g0[34]$_DFFE_NP__1594  (.L_HI(net1594));
 sg13g2_tiehi \rbzero.tex_g0[35]$_DFFE_NP__1595  (.L_HI(net1595));
 sg13g2_tiehi \rbzero.tex_g0[36]$_DFFE_NP__1596  (.L_HI(net1596));
 sg13g2_tiehi \rbzero.tex_g0[37]$_DFFE_NP__1597  (.L_HI(net1597));
 sg13g2_tiehi \rbzero.tex_g0[38]$_DFFE_NP__1598  (.L_HI(net1598));
 sg13g2_tiehi \rbzero.tex_g0[39]$_DFFE_NP__1599  (.L_HI(net1599));
 sg13g2_tiehi \rbzero.tex_g0[3]$_DFFE_NP__1600  (.L_HI(net1600));
 sg13g2_tiehi \rbzero.tex_g0[40]$_DFFE_NP__1601  (.L_HI(net1601));
 sg13g2_tiehi \rbzero.tex_g0[41]$_DFFE_NP__1602  (.L_HI(net1602));
 sg13g2_tiehi \rbzero.tex_g0[42]$_DFFE_NP__1603  (.L_HI(net1603));
 sg13g2_tiehi \rbzero.tex_g0[43]$_DFFE_NP__1604  (.L_HI(net1604));
 sg13g2_tiehi \rbzero.tex_g0[44]$_DFFE_NP__1605  (.L_HI(net1605));
 sg13g2_tiehi \rbzero.tex_g0[45]$_DFFE_NP__1606  (.L_HI(net1606));
 sg13g2_tiehi \rbzero.tex_g0[46]$_DFFE_NP__1607  (.L_HI(net1607));
 sg13g2_tiehi \rbzero.tex_g0[47]$_DFFE_NP__1608  (.L_HI(net1608));
 sg13g2_tiehi \rbzero.tex_g0[48]$_DFFE_NP__1609  (.L_HI(net1609));
 sg13g2_tiehi \rbzero.tex_g0[49]$_DFFE_NP__1610  (.L_HI(net1610));
 sg13g2_tiehi \rbzero.tex_g0[4]$_DFFE_NP__1611  (.L_HI(net1611));
 sg13g2_tiehi \rbzero.tex_g0[50]$_DFFE_NP__1612  (.L_HI(net1612));
 sg13g2_tiehi \rbzero.tex_g0[51]$_DFFE_NP__1613  (.L_HI(net1613));
 sg13g2_tiehi \rbzero.tex_g0[52]$_DFFE_NP__1614  (.L_HI(net1614));
 sg13g2_tiehi \rbzero.tex_g0[53]$_DFFE_NP__1615  (.L_HI(net1615));
 sg13g2_tiehi \rbzero.tex_g0[54]$_DFFE_NP__1616  (.L_HI(net1616));
 sg13g2_tiehi \rbzero.tex_g0[55]$_DFFE_NP__1617  (.L_HI(net1617));
 sg13g2_tiehi \rbzero.tex_g0[56]$_DFFE_NP__1618  (.L_HI(net1618));
 sg13g2_tiehi \rbzero.tex_g0[57]$_DFFE_NP__1619  (.L_HI(net1619));
 sg13g2_tiehi \rbzero.tex_g0[58]$_DFFE_NP__1620  (.L_HI(net1620));
 sg13g2_tiehi \rbzero.tex_g0[59]$_DFFE_NP__1621  (.L_HI(net1621));
 sg13g2_tiehi \rbzero.tex_g0[5]$_DFFE_NP__1622  (.L_HI(net1622));
 sg13g2_tiehi \rbzero.tex_g0[60]$_DFFE_NP__1623  (.L_HI(net1623));
 sg13g2_tiehi \rbzero.tex_g0[61]$_DFFE_NP__1624  (.L_HI(net1624));
 sg13g2_tiehi \rbzero.tex_g0[62]$_DFFE_NP__1625  (.L_HI(net1625));
 sg13g2_tiehi \rbzero.tex_g0[63]$_DFFE_NP__1626  (.L_HI(net1626));
 sg13g2_tiehi \rbzero.tex_g0[6]$_DFFE_NP__1627  (.L_HI(net1627));
 sg13g2_tiehi \rbzero.tex_g0[7]$_DFFE_NP__1628  (.L_HI(net1628));
 sg13g2_tiehi \rbzero.tex_g0[8]$_DFFE_NP__1629  (.L_HI(net1629));
 sg13g2_tiehi \rbzero.tex_g0[9]$_DFFE_NP__1630  (.L_HI(net1630));
 sg13g2_tiehi \rbzero.tex_g1[0]$_DFFE_NP__1631  (.L_HI(net1631));
 sg13g2_tiehi \rbzero.tex_g1[10]$_DFFE_NP__1632  (.L_HI(net1632));
 sg13g2_tiehi \rbzero.tex_g1[11]$_DFFE_NP__1633  (.L_HI(net1633));
 sg13g2_tiehi \rbzero.tex_g1[12]$_DFFE_NP__1634  (.L_HI(net1634));
 sg13g2_tiehi \rbzero.tex_g1[13]$_DFFE_NP__1635  (.L_HI(net1635));
 sg13g2_tiehi \rbzero.tex_g1[14]$_DFFE_NP__1636  (.L_HI(net1636));
 sg13g2_tiehi \rbzero.tex_g1[15]$_DFFE_NP__1637  (.L_HI(net1637));
 sg13g2_tiehi \rbzero.tex_g1[16]$_DFFE_NP__1638  (.L_HI(net1638));
 sg13g2_tiehi \rbzero.tex_g1[17]$_DFFE_NP__1639  (.L_HI(net1639));
 sg13g2_tiehi \rbzero.tex_g1[18]$_DFFE_NP__1640  (.L_HI(net1640));
 sg13g2_tiehi \rbzero.tex_g1[19]$_DFFE_NP__1641  (.L_HI(net1641));
 sg13g2_tiehi \rbzero.tex_g1[1]$_DFFE_NP__1642  (.L_HI(net1642));
 sg13g2_tiehi \rbzero.tex_g1[20]$_DFFE_NP__1643  (.L_HI(net1643));
 sg13g2_tiehi \rbzero.tex_g1[21]$_DFFE_NP__1644  (.L_HI(net1644));
 sg13g2_tiehi \rbzero.tex_g1[22]$_DFFE_NP__1645  (.L_HI(net1645));
 sg13g2_tiehi \rbzero.tex_g1[23]$_DFFE_NP__1646  (.L_HI(net1646));
 sg13g2_tiehi \rbzero.tex_g1[24]$_DFFE_NP__1647  (.L_HI(net1647));
 sg13g2_tiehi \rbzero.tex_g1[25]$_DFFE_NP__1648  (.L_HI(net1648));
 sg13g2_tiehi \rbzero.tex_g1[26]$_DFFE_NP__1649  (.L_HI(net1649));
 sg13g2_tiehi \rbzero.tex_g1[27]$_DFFE_NP__1650  (.L_HI(net1650));
 sg13g2_tiehi \rbzero.tex_g1[28]$_DFFE_NP__1651  (.L_HI(net1651));
 sg13g2_tiehi \rbzero.tex_g1[29]$_DFFE_NP__1652  (.L_HI(net1652));
 sg13g2_tiehi \rbzero.tex_g1[2]$_DFFE_NP__1653  (.L_HI(net1653));
 sg13g2_tiehi \rbzero.tex_g1[30]$_DFFE_NP__1654  (.L_HI(net1654));
 sg13g2_tiehi \rbzero.tex_g1[31]$_DFFE_NP__1655  (.L_HI(net1655));
 sg13g2_tiehi \rbzero.tex_g1[32]$_DFFE_NP__1656  (.L_HI(net1656));
 sg13g2_tiehi \rbzero.tex_g1[33]$_DFFE_NP__1657  (.L_HI(net1657));
 sg13g2_tiehi \rbzero.tex_g1[34]$_DFFE_NP__1658  (.L_HI(net1658));
 sg13g2_tiehi \rbzero.tex_g1[35]$_DFFE_NP__1659  (.L_HI(net1659));
 sg13g2_tiehi \rbzero.tex_g1[36]$_DFFE_NP__1660  (.L_HI(net1660));
 sg13g2_tiehi \rbzero.tex_g1[37]$_DFFE_NP__1661  (.L_HI(net1661));
 sg13g2_tiehi \rbzero.tex_g1[38]$_DFFE_NP__1662  (.L_HI(net1662));
 sg13g2_tiehi \rbzero.tex_g1[39]$_DFFE_NP__1663  (.L_HI(net1663));
 sg13g2_tiehi \rbzero.tex_g1[3]$_DFFE_NP__1664  (.L_HI(net1664));
 sg13g2_tiehi \rbzero.tex_g1[40]$_DFFE_NP__1665  (.L_HI(net1665));
 sg13g2_tiehi \rbzero.tex_g1[41]$_DFFE_NP__1666  (.L_HI(net1666));
 sg13g2_tiehi \rbzero.tex_g1[42]$_DFFE_NP__1667  (.L_HI(net1667));
 sg13g2_tiehi \rbzero.tex_g1[43]$_DFFE_NP__1668  (.L_HI(net1668));
 sg13g2_tiehi \rbzero.tex_g1[44]$_DFFE_NP__1669  (.L_HI(net1669));
 sg13g2_tiehi \rbzero.tex_g1[45]$_DFFE_NP__1670  (.L_HI(net1670));
 sg13g2_tiehi \rbzero.tex_g1[46]$_DFFE_NP__1671  (.L_HI(net1671));
 sg13g2_tiehi \rbzero.tex_g1[47]$_DFFE_NP__1672  (.L_HI(net1672));
 sg13g2_tiehi \rbzero.tex_g1[48]$_DFFE_NP__1673  (.L_HI(net1673));
 sg13g2_tiehi \rbzero.tex_g1[49]$_DFFE_NP__1674  (.L_HI(net1674));
 sg13g2_tiehi \rbzero.tex_g1[4]$_DFFE_NP__1675  (.L_HI(net1675));
 sg13g2_tiehi \rbzero.tex_g1[50]$_DFFE_NP__1676  (.L_HI(net1676));
 sg13g2_tiehi \rbzero.tex_g1[51]$_DFFE_NP__1677  (.L_HI(net1677));
 sg13g2_tiehi \rbzero.tex_g1[52]$_DFFE_NP__1678  (.L_HI(net1678));
 sg13g2_tiehi \rbzero.tex_g1[53]$_DFFE_NP__1679  (.L_HI(net1679));
 sg13g2_tiehi \rbzero.tex_g1[54]$_DFFE_NP__1680  (.L_HI(net1680));
 sg13g2_tiehi \rbzero.tex_g1[55]$_DFFE_NP__1681  (.L_HI(net1681));
 sg13g2_tiehi \rbzero.tex_g1[56]$_DFFE_NP__1682  (.L_HI(net1682));
 sg13g2_tiehi \rbzero.tex_g1[57]$_DFFE_NP__1683  (.L_HI(net1683));
 sg13g2_tiehi \rbzero.tex_g1[58]$_DFFE_NP__1684  (.L_HI(net1684));
 sg13g2_tiehi \rbzero.tex_g1[59]$_DFFE_NP__1685  (.L_HI(net1685));
 sg13g2_tiehi \rbzero.tex_g1[5]$_DFFE_NP__1686  (.L_HI(net1686));
 sg13g2_tiehi \rbzero.tex_g1[60]$_DFFE_NP__1687  (.L_HI(net1687));
 sg13g2_tiehi \rbzero.tex_g1[61]$_DFFE_NP__1688  (.L_HI(net1688));
 sg13g2_tiehi \rbzero.tex_g1[62]$_DFFE_NP__1689  (.L_HI(net1689));
 sg13g2_tiehi \rbzero.tex_g1[63]$_DFFE_NP__1690  (.L_HI(net1690));
 sg13g2_tiehi \rbzero.tex_g1[6]$_DFFE_NP__1691  (.L_HI(net1691));
 sg13g2_tiehi \rbzero.tex_g1[7]$_DFFE_NP__1692  (.L_HI(net1692));
 sg13g2_tiehi \rbzero.tex_g1[8]$_DFFE_NP__1693  (.L_HI(net1693));
 sg13g2_tiehi \rbzero.tex_g1[9]$_DFFE_NP__1694  (.L_HI(net1694));
 sg13g2_tiehi \rbzero.tex_r0[0]$_DFFE_NP__1695  (.L_HI(net1695));
 sg13g2_tiehi \rbzero.tex_r0[10]$_DFFE_NP__1696  (.L_HI(net1696));
 sg13g2_tiehi \rbzero.tex_r0[11]$_DFFE_NP__1697  (.L_HI(net1697));
 sg13g2_tiehi \rbzero.tex_r0[12]$_DFFE_NP__1698  (.L_HI(net1698));
 sg13g2_tiehi \rbzero.tex_r0[13]$_DFFE_NP__1699  (.L_HI(net1699));
 sg13g2_tiehi \rbzero.tex_r0[14]$_DFFE_NP__1700  (.L_HI(net1700));
 sg13g2_tiehi \rbzero.tex_r0[15]$_DFFE_NP__1701  (.L_HI(net1701));
 sg13g2_tiehi \rbzero.tex_r0[16]$_DFFE_NP__1702  (.L_HI(net1702));
 sg13g2_tiehi \rbzero.tex_r0[17]$_DFFE_NP__1703  (.L_HI(net1703));
 sg13g2_tiehi \rbzero.tex_r0[18]$_DFFE_NP__1704  (.L_HI(net1704));
 sg13g2_tiehi \rbzero.tex_r0[19]$_DFFE_NP__1705  (.L_HI(net1705));
 sg13g2_tiehi \rbzero.tex_r0[1]$_DFFE_NP__1706  (.L_HI(net1706));
 sg13g2_tiehi \rbzero.tex_r0[20]$_DFFE_NP__1707  (.L_HI(net1707));
 sg13g2_tiehi \rbzero.tex_r0[21]$_DFFE_NP__1708  (.L_HI(net1708));
 sg13g2_tiehi \rbzero.tex_r0[22]$_DFFE_NP__1709  (.L_HI(net1709));
 sg13g2_tiehi \rbzero.tex_r0[23]$_DFFE_NP__1710  (.L_HI(net1710));
 sg13g2_tiehi \rbzero.tex_r0[24]$_DFFE_NP__1711  (.L_HI(net1711));
 sg13g2_tiehi \rbzero.tex_r0[25]$_DFFE_NP__1712  (.L_HI(net1712));
 sg13g2_tiehi \rbzero.tex_r0[26]$_DFFE_NP__1713  (.L_HI(net1713));
 sg13g2_tiehi \rbzero.tex_r0[27]$_DFFE_NP__1714  (.L_HI(net1714));
 sg13g2_tiehi \rbzero.tex_r0[28]$_DFFE_NP__1715  (.L_HI(net1715));
 sg13g2_tiehi \rbzero.tex_r0[29]$_DFFE_NP__1716  (.L_HI(net1716));
 sg13g2_tiehi \rbzero.tex_r0[2]$_DFFE_NP__1717  (.L_HI(net1717));
 sg13g2_tiehi \rbzero.tex_r0[30]$_DFFE_NP__1718  (.L_HI(net1718));
 sg13g2_tiehi \rbzero.tex_r0[31]$_DFFE_NP__1719  (.L_HI(net1719));
 sg13g2_tiehi \rbzero.tex_r0[32]$_DFFE_NP__1720  (.L_HI(net1720));
 sg13g2_tiehi \rbzero.tex_r0[33]$_DFFE_NP__1721  (.L_HI(net1721));
 sg13g2_tiehi \rbzero.tex_r0[34]$_DFFE_NP__1722  (.L_HI(net1722));
 sg13g2_tiehi \rbzero.tex_r0[35]$_DFFE_NP__1723  (.L_HI(net1723));
 sg13g2_tiehi \rbzero.tex_r0[36]$_DFFE_NP__1724  (.L_HI(net1724));
 sg13g2_tiehi \rbzero.tex_r0[37]$_DFFE_NP__1725  (.L_HI(net1725));
 sg13g2_tiehi \rbzero.tex_r0[38]$_DFFE_NP__1726  (.L_HI(net1726));
 sg13g2_tiehi \rbzero.tex_r0[39]$_DFFE_NP__1727  (.L_HI(net1727));
 sg13g2_tiehi \rbzero.tex_r0[3]$_DFFE_NP__1728  (.L_HI(net1728));
 sg13g2_tiehi \rbzero.tex_r0[40]$_DFFE_NP__1729  (.L_HI(net1729));
 sg13g2_tiehi \rbzero.tex_r0[41]$_DFFE_NP__1730  (.L_HI(net1730));
 sg13g2_tiehi \rbzero.tex_r0[42]$_DFFE_NP__1731  (.L_HI(net1731));
 sg13g2_tiehi \rbzero.tex_r0[43]$_DFFE_NP__1732  (.L_HI(net1732));
 sg13g2_tiehi \rbzero.tex_r0[44]$_DFFE_NP__1733  (.L_HI(net1733));
 sg13g2_tiehi \rbzero.tex_r0[45]$_DFFE_NP__1734  (.L_HI(net1734));
 sg13g2_tiehi \rbzero.tex_r0[46]$_DFFE_NP__1735  (.L_HI(net1735));
 sg13g2_tiehi \rbzero.tex_r0[47]$_DFFE_NP__1736  (.L_HI(net1736));
 sg13g2_tiehi \rbzero.tex_r0[48]$_DFFE_NP__1737  (.L_HI(net1737));
 sg13g2_tiehi \rbzero.tex_r0[49]$_DFFE_NP__1738  (.L_HI(net1738));
 sg13g2_tiehi \rbzero.tex_r0[4]$_DFFE_NP__1739  (.L_HI(net1739));
 sg13g2_tiehi \rbzero.tex_r0[50]$_DFFE_NP__1740  (.L_HI(net1740));
 sg13g2_tiehi \rbzero.tex_r0[51]$_DFFE_NP__1741  (.L_HI(net1741));
 sg13g2_tiehi \rbzero.tex_r0[52]$_DFFE_NP__1742  (.L_HI(net1742));
 sg13g2_tiehi \rbzero.tex_r0[53]$_DFFE_NP__1743  (.L_HI(net1743));
 sg13g2_tiehi \rbzero.tex_r0[54]$_DFFE_NP__1744  (.L_HI(net1744));
 sg13g2_tiehi \rbzero.tex_r0[55]$_DFFE_NP__1745  (.L_HI(net1745));
 sg13g2_tiehi \rbzero.tex_r0[56]$_DFFE_NP__1746  (.L_HI(net1746));
 sg13g2_tiehi \rbzero.tex_r0[57]$_DFFE_NP__1747  (.L_HI(net1747));
 sg13g2_tiehi \rbzero.tex_r0[58]$_DFFE_NP__1748  (.L_HI(net1748));
 sg13g2_tiehi \rbzero.tex_r0[59]$_DFFE_NP__1749  (.L_HI(net1749));
 sg13g2_tiehi \rbzero.tex_r0[5]$_DFFE_NP__1750  (.L_HI(net1750));
 sg13g2_tiehi \rbzero.tex_r0[60]$_DFFE_NP__1751  (.L_HI(net1751));
 sg13g2_tiehi \rbzero.tex_r0[61]$_DFFE_NP__1752  (.L_HI(net1752));
 sg13g2_tiehi \rbzero.tex_r0[62]$_DFFE_NP__1753  (.L_HI(net1753));
 sg13g2_tiehi \rbzero.tex_r0[63]$_DFFE_NP__1754  (.L_HI(net1754));
 sg13g2_tiehi \rbzero.tex_r0[6]$_DFFE_NP__1755  (.L_HI(net1755));
 sg13g2_tiehi \rbzero.tex_r0[7]$_DFFE_NP__1756  (.L_HI(net1756));
 sg13g2_tiehi \rbzero.tex_r0[8]$_DFFE_NP__1757  (.L_HI(net1757));
 sg13g2_tiehi \rbzero.tex_r0[9]$_DFFE_NP__1758  (.L_HI(net1758));
 sg13g2_tiehi \rbzero.tex_r1[0]$_DFFE_NP__1759  (.L_HI(net1759));
 sg13g2_tiehi \rbzero.tex_r1[10]$_DFFE_NP__1760  (.L_HI(net1760));
 sg13g2_tiehi \rbzero.tex_r1[11]$_DFFE_NP__1761  (.L_HI(net1761));
 sg13g2_tiehi \rbzero.tex_r1[12]$_DFFE_NP__1762  (.L_HI(net1762));
 sg13g2_tiehi \rbzero.tex_r1[13]$_DFFE_NP__1763  (.L_HI(net1763));
 sg13g2_tiehi \rbzero.tex_r1[14]$_DFFE_NP__1764  (.L_HI(net1764));
 sg13g2_tiehi \rbzero.tex_r1[15]$_DFFE_NP__1765  (.L_HI(net1765));
 sg13g2_tiehi \rbzero.tex_r1[16]$_DFFE_NP__1766  (.L_HI(net1766));
 sg13g2_tiehi \rbzero.tex_r1[17]$_DFFE_NP__1767  (.L_HI(net1767));
 sg13g2_tiehi \rbzero.tex_r1[18]$_DFFE_NP__1768  (.L_HI(net1768));
 sg13g2_tiehi \rbzero.tex_r1[19]$_DFFE_NP__1769  (.L_HI(net1769));
 sg13g2_tiehi \rbzero.tex_r1[1]$_DFFE_NP__1770  (.L_HI(net1770));
 sg13g2_tiehi \rbzero.tex_r1[20]$_DFFE_NP__1771  (.L_HI(net1771));
 sg13g2_tiehi \rbzero.tex_r1[21]$_DFFE_NP__1772  (.L_HI(net1772));
 sg13g2_tiehi \rbzero.tex_r1[22]$_DFFE_NP__1773  (.L_HI(net1773));
 sg13g2_tiehi \rbzero.tex_r1[23]$_DFFE_NP__1774  (.L_HI(net1774));
 sg13g2_tiehi \rbzero.tex_r1[24]$_DFFE_NP__1775  (.L_HI(net1775));
 sg13g2_tiehi \rbzero.tex_r1[25]$_DFFE_NP__1776  (.L_HI(net1776));
 sg13g2_tiehi \rbzero.tex_r1[26]$_DFFE_NP__1777  (.L_HI(net1777));
 sg13g2_tiehi \rbzero.tex_r1[27]$_DFFE_NP__1778  (.L_HI(net1778));
 sg13g2_tiehi \rbzero.tex_r1[28]$_DFFE_NP__1779  (.L_HI(net1779));
 sg13g2_tiehi \rbzero.tex_r1[29]$_DFFE_NP__1780  (.L_HI(net1780));
 sg13g2_tiehi \rbzero.tex_r1[2]$_DFFE_NP__1781  (.L_HI(net1781));
 sg13g2_tiehi \rbzero.tex_r1[30]$_DFFE_NP__1782  (.L_HI(net1782));
 sg13g2_tiehi \rbzero.tex_r1[31]$_DFFE_NP__1783  (.L_HI(net1783));
 sg13g2_tiehi \rbzero.tex_r1[32]$_DFFE_NP__1784  (.L_HI(net1784));
 sg13g2_tiehi \rbzero.tex_r1[33]$_DFFE_NP__1785  (.L_HI(net1785));
 sg13g2_tiehi \rbzero.tex_r1[34]$_DFFE_NP__1786  (.L_HI(net1786));
 sg13g2_tiehi \rbzero.tex_r1[35]$_DFFE_NP__1787  (.L_HI(net1787));
 sg13g2_tiehi \rbzero.tex_r1[36]$_DFFE_NP__1788  (.L_HI(net1788));
 sg13g2_tiehi \rbzero.tex_r1[37]$_DFFE_NP__1789  (.L_HI(net1789));
 sg13g2_tiehi \rbzero.tex_r1[38]$_DFFE_NP__1790  (.L_HI(net1790));
 sg13g2_tiehi \rbzero.tex_r1[39]$_DFFE_NP__1791  (.L_HI(net1791));
 sg13g2_tiehi \rbzero.tex_r1[3]$_DFFE_NP__1792  (.L_HI(net1792));
 sg13g2_tiehi \rbzero.tex_r1[40]$_DFFE_NP__1793  (.L_HI(net1793));
 sg13g2_tiehi \rbzero.tex_r1[41]$_DFFE_NP__1794  (.L_HI(net1794));
 sg13g2_tiehi \rbzero.tex_r1[42]$_DFFE_NP__1795  (.L_HI(net1795));
 sg13g2_tiehi \rbzero.tex_r1[43]$_DFFE_NP__1796  (.L_HI(net1796));
 sg13g2_tiehi \rbzero.tex_r1[44]$_DFFE_NP__1797  (.L_HI(net1797));
 sg13g2_tiehi \rbzero.tex_r1[45]$_DFFE_NP__1798  (.L_HI(net1798));
 sg13g2_tiehi \rbzero.tex_r1[46]$_DFFE_NP__1799  (.L_HI(net1799));
 sg13g2_tiehi \rbzero.tex_r1[47]$_DFFE_NP__1800  (.L_HI(net1800));
 sg13g2_tiehi \rbzero.tex_r1[48]$_DFFE_NP__1801  (.L_HI(net1801));
 sg13g2_tiehi \rbzero.tex_r1[49]$_DFFE_NP__1802  (.L_HI(net1802));
 sg13g2_tiehi \rbzero.tex_r1[4]$_DFFE_NP__1803  (.L_HI(net1803));
 sg13g2_tiehi \rbzero.tex_r1[50]$_DFFE_NP__1804  (.L_HI(net1804));
 sg13g2_tiehi \rbzero.tex_r1[51]$_DFFE_NP__1805  (.L_HI(net1805));
 sg13g2_tiehi \rbzero.tex_r1[52]$_DFFE_NP__1806  (.L_HI(net1806));
 sg13g2_tiehi \rbzero.tex_r1[53]$_DFFE_NP__1807  (.L_HI(net1807));
 sg13g2_tiehi \rbzero.tex_r1[54]$_DFFE_NP__1808  (.L_HI(net1808));
 sg13g2_tiehi \rbzero.tex_r1[55]$_DFFE_NP__1809  (.L_HI(net1809));
 sg13g2_tiehi \rbzero.tex_r1[56]$_DFFE_NP__1810  (.L_HI(net1810));
 sg13g2_tiehi \rbzero.tex_r1[57]$_DFFE_NP__1811  (.L_HI(net1811));
 sg13g2_tiehi \rbzero.tex_r1[58]$_DFFE_NP__1812  (.L_HI(net1812));
 sg13g2_tiehi \rbzero.tex_r1[59]$_DFFE_NP__1813  (.L_HI(net1813));
 sg13g2_tiehi \rbzero.tex_r1[5]$_DFFE_NP__1814  (.L_HI(net1814));
 sg13g2_tiehi \rbzero.tex_r1[60]$_DFFE_NP__1815  (.L_HI(net1815));
 sg13g2_tiehi \rbzero.tex_r1[61]$_DFFE_NP__1816  (.L_HI(net1816));
 sg13g2_tiehi \rbzero.tex_r1[62]$_DFFE_NP__1817  (.L_HI(net1817));
 sg13g2_tiehi \rbzero.tex_r1[63]$_DFFE_NP__1818  (.L_HI(net1818));
 sg13g2_tiehi \rbzero.tex_r1[6]$_DFFE_NP__1819  (.L_HI(net1819));
 sg13g2_tiehi \rbzero.tex_r1[7]$_DFFE_NP__1820  (.L_HI(net1820));
 sg13g2_tiehi \rbzero.tex_r1[8]$_DFFE_NP__1821  (.L_HI(net1821));
 sg13g2_tiehi \rbzero.tex_r1[9]$_DFFE_NP__1822  (.L_HI(net1822));
 sg13g2_tiehi \rbzero.vga_sync.hpos[0]$_SDFF_PP0__1823  (.L_HI(net1823));
 sg13g2_tiehi \rbzero.vga_sync.hpos[1]$_SDFF_PP0__1824  (.L_HI(net1824));
 sg13g2_tiehi \rbzero.vga_sync.hpos[2]$_SDFF_PP0__1825  (.L_HI(net1825));
 sg13g2_tiehi \rbzero.vga_sync.hpos[3]$_SDFF_PP0__1826  (.L_HI(net1826));
 sg13g2_tiehi \rbzero.vga_sync.hpos[4]$_SDFF_PP0__1827  (.L_HI(net1827));
 sg13g2_tiehi \rbzero.vga_sync.hpos[5]$_SDFF_PP0__1828  (.L_HI(net1828));
 sg13g2_tiehi \rbzero.vga_sync.hpos[6]$_SDFF_PP0__1829  (.L_HI(net1829));
 sg13g2_tiehi \rbzero.vga_sync.hpos[7]$_SDFF_PP0__1830  (.L_HI(net1830));
 sg13g2_tiehi \rbzero.vga_sync.hpos[8]$_SDFF_PP0__1831  (.L_HI(net1831));
 sg13g2_tiehi \rbzero.vga_sync.hpos[9]$_SDFF_PP0__1832  (.L_HI(net1832));
 sg13g2_tiehi \rbzero.vga_sync.hsync$_SDFFE_PP0N__1833  (.L_HI(net1833));
 sg13g2_tiehi \rbzero.vga_sync.vpos[0]$_SDFFE_PN0P__1834  (.L_HI(net1834));
 sg13g2_tiehi \rbzero.vga_sync.vpos[1]$_SDFFE_PN0P__1835  (.L_HI(net1835));
 sg13g2_tiehi \rbzero.vga_sync.vpos[2]$_SDFFE_PN0P__1836  (.L_HI(net1836));
 sg13g2_tiehi \rbzero.vga_sync.vpos[3]$_SDFFE_PN0P__1837  (.L_HI(net1837));
 sg13g2_tiehi \rbzero.vga_sync.vpos[4]$_SDFFE_PN0P__1838  (.L_HI(net1838));
 sg13g2_tiehi \rbzero.vga_sync.vpos[5]$_SDFFE_PN0P__1839  (.L_HI(net1839));
 sg13g2_tiehi \rbzero.vga_sync.vpos[6]$_SDFFE_PN0P__1840  (.L_HI(net1840));
 sg13g2_tiehi \rbzero.vga_sync.vpos[7]$_SDFFE_PN0P__1841  (.L_HI(net1841));
 sg13g2_tiehi \rbzero.vga_sync.vpos[8]$_SDFFE_PN0P__1842  (.L_HI(net1842));
 sg13g2_tiehi \rbzero.vga_sync.vpos[9]$_SDFFE_PN0P__1843  (.L_HI(net1843));
 sg13g2_tiehi \rbzero.vga_sync.vsync$_SDFFE_PP0N__1844  (.L_HI(net1844));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[0]$_SDFFE_PN0P__1845  (.L_HI(net1845));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[10]$_SDFFE_PN0P__1846  (.L_HI(net1846));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[1]$_SDFFE_PN0P__1847  (.L_HI(net1847));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[2]$_SDFFE_PN0P__1848  (.L_HI(net1848));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[3]$_SDFFE_PN0P__1849  (.L_HI(net1849));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[4]$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[5]$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[6]$_SDFFE_PN0P__1852  (.L_HI(net1852));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[7]$_SDFFE_PN0P__1853  (.L_HI(net1853));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[8]$_SDFFE_PN0P__1854  (.L_HI(net1854));
 sg13g2_tiehi \rbzero.wall_tracer.mapX[9]$_SDFFE_PN0P__1855  (.L_HI(net1855));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[0]$_SDFFE_PN0P__1856  (.L_HI(net1856));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[10]$_SDFFE_PN0P__1857  (.L_HI(net1857));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[1]$_SDFFE_PN0P__1858  (.L_HI(net1858));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[2]$_SDFFE_PN0P__1859  (.L_HI(net1859));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[3]$_SDFFE_PN0P__1860  (.L_HI(net1860));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[4]$_SDFFE_PN0P__1861  (.L_HI(net1861));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[5]$_SDFFE_PN0P__1862  (.L_HI(net1862));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[6]$_SDFFE_PN0P__1863  (.L_HI(net1863));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[7]$_SDFFE_PN0P__1864  (.L_HI(net1864));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[8]$_SDFFE_PN0P__1865  (.L_HI(net1865));
 sg13g2_tiehi \rbzero.wall_tracer.mapY[9]$_SDFFE_PN0P__1866  (.L_HI(net1866));
 sg13g2_tiehi \rbzero.wall_tracer.o_side$_SDFFE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \rbzero.wall_tracer.o_side_hot$_SDFFE_PN0P__1868  (.L_HI(net1868));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[0]$_SDFFE_PN0P__1869  (.L_HI(net1869));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[10]$_SDFFE_PN0P__1870  (.L_HI(net1870));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[1]$_SDFFE_PN0P__1871  (.L_HI(net1871));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[2]$_SDFFE_PN0P__1872  (.L_HI(net1872));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[3]$_SDFFE_PN0P__1873  (.L_HI(net1873));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[4]$_SDFFE_PN0P__1874  (.L_HI(net1874));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[5]$_SDFFE_PN0P__1875  (.L_HI(net1875));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[6]$_SDFFE_PN0P__1876  (.L_HI(net1876));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[7]$_SDFFE_PN0P__1877  (.L_HI(net1877));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[8]$_SDFFE_PN0P__1878  (.L_HI(net1878));
 sg13g2_tiehi \rbzero.wall_tracer.o_size[9]$_SDFFE_PN0P__1879  (.L_HI(net1879));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[11]$_SDFFE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[12]$_SDFFE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[13]$_SDFFE_PN0P__1882  (.L_HI(net1882));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[14]$_SDFFE_PN0P__1883  (.L_HI(net1883));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[15]$_SDFFE_PN0P__1884  (.L_HI(net1884));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[16]$_SDFFE_PN0P__1885  (.L_HI(net1885));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[17]$_SDFFE_PN0P__1886  (.L_HI(net1886));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[18]$_SDFFE_PN0P__1887  (.L_HI(net1887));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[19]$_SDFFE_PN0P__1888  (.L_HI(net1888));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[20]$_SDFFE_PN0P__1889  (.L_HI(net1889));
 sg13g2_tiehi \rbzero.wall_tracer.o_texVinit[21]$_SDFFE_PN0P__1890  (.L_HI(net1890));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[0]$_SDFFE_PN0P__1891  (.L_HI(net1891));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[10]$_SDFFE_PN0P__1892  (.L_HI(net1892));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[11]$_SDFFE_PN0P__1893  (.L_HI(net1893));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[12]$_SDFFE_PN0P__1894  (.L_HI(net1894));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[13]$_SDFFE_PN0P__1895  (.L_HI(net1895));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[14]$_SDFFE_PN0P__1896  (.L_HI(net1896));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[15]$_SDFFE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[16]$_SDFFE_PN0P__1898  (.L_HI(net1898));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[17]$_SDFFE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[18]$_SDFFE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[19]$_SDFFE_PN0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[1]$_SDFFE_PN0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[20]$_SDFFE_PN0P__1903  (.L_HI(net1903));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[21]$_SDFFE_PN0P__1904  (.L_HI(net1904));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[2]$_SDFFE_PN0P__1905  (.L_HI(net1905));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[3]$_SDFFE_PN0P__1906  (.L_HI(net1906));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[4]$_SDFFE_PN0P__1907  (.L_HI(net1907));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[5]$_SDFFE_PN0P__1908  (.L_HI(net1908));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[6]$_SDFFE_PN0P__1909  (.L_HI(net1909));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[7]$_SDFFE_PN0P__1910  (.L_HI(net1910));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[8]$_SDFFE_PN0P__1911  (.L_HI(net1911));
 sg13g2_tiehi \rbzero.wall_tracer.o_texa[9]$_SDFFE_PN0P__1912  (.L_HI(net1912));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu[0]$_SDFFE_PN0P__1913  (.L_HI(net1913));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu[1]$_SDFFE_PN0P__1914  (.L_HI(net1914));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu[2]$_SDFFE_PN0P__1915  (.L_HI(net1915));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu[3]$_SDFFE_PN0P__1916  (.L_HI(net1916));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu[4]$_SDFFE_PN0P__1917  (.L_HI(net1917));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[0]$_SDFFE_PN0P__1918  (.L_HI(net1918));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[1]$_SDFFE_PN0P__1919  (.L_HI(net1919));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[2]$_SDFFE_PN0P__1920  (.L_HI(net1920));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[3]$_SDFFE_PN0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[4]$_SDFFE_PN0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \rbzero.wall_tracer.o_texu_hot[5]$_SDFFE_PN0P__1923  (.L_HI(net1923));
 sg13g2_tiehi \rbzero.wall_tracer.o_wall[0]$_SDFFE_PN0P__1924  (.L_HI(net1924));
 sg13g2_tiehi \rbzero.wall_tracer.o_wall[1]$_SDFFE_PN0P__1925  (.L_HI(net1925));
 sg13g2_tiehi \rbzero.wall_tracer.o_wall_hot[0]$_SDFFE_PN0P__1926  (.L_HI(net1926));
 sg13g2_tiehi \rbzero.wall_tracer.o_wall_hot[1]$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[10]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[11]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[12]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[13]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[14]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[15]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[16]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[17]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[18]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[19]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[20]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[21]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[2]$_SDFFCE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[3]$_SDFFCE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[4]$_SDFFCE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[5]$_SDFFCE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[6]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[7]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[8]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendX[9]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[10]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[11]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[12]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[13]$_DFFE_PP__1951  (.L_HI(net1951));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[14]$_DFFE_PP__1952  (.L_HI(net1952));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[15]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[16]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[17]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[18]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[19]$_DFFE_PP__1957  (.L_HI(net1957));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[20]$_DFFE_PP__1958  (.L_HI(net1958));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[21]$_DFFE_PP__1959  (.L_HI(net1959));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[2]$_SDFFCE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[3]$_SDFFCE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[4]$_SDFFCE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[5]$_SDFFCE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[6]$_DFFE_PP__1964  (.L_HI(net1964));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[7]$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[8]$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \rbzero.wall_tracer.rayAddendY[9]$_DFFE_PP__1967  (.L_HI(net1967));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[0]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[10]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[11]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[12]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[13]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[14]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[15]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[16]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[17]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[18]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[19]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[1]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[20]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[21]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[2]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[3]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[4]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[5]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[6]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[7]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[8]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_data[9]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.o_done$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[0]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[10]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[11]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[12]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[13]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[14]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[15]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[16]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[17]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[18]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[19]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[1]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[20]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[21]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[2]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[3]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[4]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[5]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[6]$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[7]$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[8]$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.operand[9]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.state[0]$_DFF_P__2013  (.L_HI(net2013));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.state[1]$_DFF_P__2014  (.L_HI(net2014));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.state[2]$_DFF_P__2015  (.L_HI(net2015));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.state[3]$_DFF_P__2016  (.L_HI(net2016));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_fsm.state[4]$_DFF_P__2017  (.L_HI(net2017));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[0]$_SDFFE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[10]$_SDFFE_PN0P__2019  (.L_HI(net2019));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[11]$_SDFFE_PN0P__2020  (.L_HI(net2020));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[12]$_SDFFE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[13]$_SDFFE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[14]$_SDFFE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[15]$_SDFFE_PN0P__2024  (.L_HI(net2024));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[16]$_SDFFE_PN0P__2025  (.L_HI(net2025));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[17]$_SDFFE_PN0P__2026  (.L_HI(net2026));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[18]$_SDFFE_PN0P__2027  (.L_HI(net2027));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[19]$_SDFFE_PN0P__2028  (.L_HI(net2028));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[1]$_SDFFE_PN0P__2029  (.L_HI(net2029));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[20]$_SDFFE_PN0P__2030  (.L_HI(net2030));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[21]$_SDFFE_PN0P__2031  (.L_HI(net2031));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[2]$_SDFFE_PN0P__2032  (.L_HI(net2032));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[3]$_SDFFE_PN0P__2033  (.L_HI(net2033));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[4]$_SDFFE_PN0P__2034  (.L_HI(net2034));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[5]$_SDFFE_PN0P__2035  (.L_HI(net2035));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[6]$_SDFFE_PN0P__2036  (.L_HI(net2036));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[7]$_SDFFE_PN0P__2037  (.L_HI(net2037));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[8]$_SDFFE_PN0P__2038  (.L_HI(net2038));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_in[9]$_SDFFE_PN0P__2039  (.L_HI(net2039));
 sg13g2_tiehi \rbzero.wall_tracer.rcp_start$_SDFFE_PN0P__2040  (.L_HI(net2040));
 sg13g2_tiehi \rbzero.wall_tracer.side$_SDFFE_PN0P__2041  (.L_HI(net2041));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[0]$_SDFFE_PN0P__2042  (.L_HI(net2042));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[10]$_SDFFE_PN0P__2043  (.L_HI(net2043));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[11]$_SDFFE_PN0P__2044  (.L_HI(net2044));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[12]$_SDFFE_PN0P__2045  (.L_HI(net2045));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[13]$_SDFFE_PN0P__2046  (.L_HI(net2046));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[14]$_SDFFE_PN0P__2047  (.L_HI(net2047));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[15]$_SDFFE_PN0P__2048  (.L_HI(net2048));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[16]$_SDFFE_PN0P__2049  (.L_HI(net2049));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[17]$_SDFFE_PN0P__2050  (.L_HI(net2050));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[18]$_SDFFE_PN0P__2051  (.L_HI(net2051));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[19]$_SDFFE_PN0P__2052  (.L_HI(net2052));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[1]$_SDFFE_PN0P__2053  (.L_HI(net2053));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[20]$_SDFFE_PN0P__2054  (.L_HI(net2054));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[21]$_SDFFE_PN0P__2055  (.L_HI(net2055));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[2]$_SDFFE_PN0P__2056  (.L_HI(net2056));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[3]$_SDFFE_PN0P__2057  (.L_HI(net2057));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[4]$_SDFFE_PN0P__2058  (.L_HI(net2058));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[5]$_SDFFE_PN0P__2059  (.L_HI(net2059));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[6]$_SDFFE_PN0P__2060  (.L_HI(net2060));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[7]$_SDFFE_PN0P__2061  (.L_HI(net2061));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[8]$_SDFFE_PN0P__2062  (.L_HI(net2062));
 sg13g2_tiehi \rbzero.wall_tracer.size_full[9]$_SDFFE_PN0P__2063  (.L_HI(net2063));
 sg13g2_tiehi \rbzero.wall_tracer.state[0]$_DFF_P__2064  (.L_HI(net2064));
 sg13g2_tiehi \rbzero.wall_tracer.state[1]$_DFF_P__2065  (.L_HI(net2065));
 sg13g2_tiehi \rbzero.wall_tracer.state[2]$_DFF_P__2066  (.L_HI(net2066));
 sg13g2_tiehi \rbzero.wall_tracer.state[3]$_DFF_P__2067  (.L_HI(net2067));
 sg13g2_tiehi \rbzero.wall_tracer.state[4]$_DFF_P__2068  (.L_HI(net2068));
 sg13g2_tiehi \rbzero.wall_tracer.state[5]$_DFF_P__2069  (.L_HI(net2069));
 sg13g2_tiehi \rbzero.wall_tracer.state[6]$_DFF_P__2070  (.L_HI(net2070));
 sg13g2_tiehi \rbzero.wall_tracer.state[7]$_DFF_P__2071  (.L_HI(net2071));
 sg13g2_tiehi \rbzero.wall_tracer.state[8]$_DFF_P__2072  (.L_HI(net2072));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[0]$_SDFFE_PN0P__2073  (.L_HI(net2073));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[10]$_SDFFE_PN0P__2074  (.L_HI(net2074));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[11]$_SDFFE_PN0P__2075  (.L_HI(net2075));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[12]$_SDFFE_PN0P__2076  (.L_HI(net2076));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[13]$_SDFFE_PN0P__2077  (.L_HI(net2077));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[14]$_SDFFE_PN0P__2078  (.L_HI(net2078));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[15]$_SDFFE_PN0P__2079  (.L_HI(net2079));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[16]$_SDFFE_PN0P__2080  (.L_HI(net2080));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[17]$_SDFFE_PN0P__2081  (.L_HI(net2081));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[18]$_SDFFE_PN0P__2082  (.L_HI(net2082));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[19]$_SDFFE_PN0P__2083  (.L_HI(net2083));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[1]$_SDFFE_PN0P__2084  (.L_HI(net2084));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[20]$_SDFFE_PN0P__2085  (.L_HI(net2085));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[21]$_SDFFE_PN0P__2086  (.L_HI(net2086));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[2]$_SDFFE_PN0P__2087  (.L_HI(net2087));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[3]$_SDFFE_PN0P__2088  (.L_HI(net2088));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[4]$_SDFFE_PN0P__2089  (.L_HI(net2089));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[5]$_SDFFE_PN0P__2090  (.L_HI(net2090));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[6]$_SDFFE_PN0P__2091  (.L_HI(net2091));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[7]$_SDFFE_PN0P__2092  (.L_HI(net2092));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[8]$_SDFFE_PN0P__2093  (.L_HI(net2093));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistX[9]$_SDFFE_PN0P__2094  (.L_HI(net2094));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[0]$_SDFFE_PN0P__2095  (.L_HI(net2095));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[10]$_SDFFE_PN0P__2096  (.L_HI(net2096));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[11]$_SDFFE_PN0P__2097  (.L_HI(net2097));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[12]$_SDFFE_PN0P__2098  (.L_HI(net2098));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[13]$_SDFFE_PN0P__2099  (.L_HI(net2099));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[14]$_SDFFE_PN0P__2100  (.L_HI(net2100));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[15]$_SDFFE_PN0P__2101  (.L_HI(net2101));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[16]$_SDFFE_PN0P__2102  (.L_HI(net2102));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[17]$_SDFFE_PN0P__2103  (.L_HI(net2103));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[18]$_SDFFE_PN0P__2104  (.L_HI(net2104));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[19]$_SDFFE_PN0P__2105  (.L_HI(net2105));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[1]$_SDFFE_PN0P__2106  (.L_HI(net2106));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[20]$_SDFFE_PN0P__2107  (.L_HI(net2107));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[21]$_SDFFE_PN0P__2108  (.L_HI(net2108));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[2]$_SDFFE_PN0P__2109  (.L_HI(net2109));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[3]$_SDFFE_PN0P__2110  (.L_HI(net2110));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[4]$_SDFFE_PN0P__2111  (.L_HI(net2111));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[5]$_SDFFE_PN0P__2112  (.L_HI(net2112));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[6]$_SDFFE_PN0P__2113  (.L_HI(net2113));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[7]$_SDFFE_PN0P__2114  (.L_HI(net2114));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[8]$_SDFFE_PN0P__2115  (.L_HI(net2115));
 sg13g2_tiehi \rbzero.wall_tracer.stepDistY[9]$_SDFFE_PN0P__2116  (.L_HI(net2116));
 sg13g2_tiehi \rbzero.wall_tracer.texu[0]$_SDFFE_PN0P__2117  (.L_HI(net2117));
 sg13g2_tiehi \rbzero.wall_tracer.texu[1]$_SDFFE_PN0P__2118  (.L_HI(net2118));
 sg13g2_tiehi \rbzero.wall_tracer.texu[2]$_SDFFE_PN0P__2119  (.L_HI(net2119));
 sg13g2_tiehi \rbzero.wall_tracer.texu[3]$_SDFFE_PN0P__2120  (.L_HI(net2120));
 sg13g2_tiehi \rbzero.wall_tracer.texu[4]$_SDFFE_PN0P__2121  (.L_HI(net2121));
 sg13g2_tiehi \rbzero.wall_tracer.texu[5]$_SDFFE_PN0P__2122  (.L_HI(net2122));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[0]$_SDFFE_PN0P__2123  (.L_HI(net2123));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[10]$_SDFFE_PN0P__2124  (.L_HI(net2124));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[11]$_SDFFE_PN0P__2125  (.L_HI(net2125));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[12]$_SDFFE_PN0P__2126  (.L_HI(net2126));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[13]$_SDFFE_PN0P__2127  (.L_HI(net2127));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[14]$_SDFFE_PN0P__2128  (.L_HI(net2128));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[15]$_SDFFE_PN0P__2129  (.L_HI(net2129));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[16]$_SDFFE_PN0P__2130  (.L_HI(net2130));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[17]$_SDFFE_PN0P__2131  (.L_HI(net2131));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[18]$_SDFFE_PN0P__2132  (.L_HI(net2132));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[19]$_SDFFE_PN0P__2133  (.L_HI(net2133));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[1]$_SDFFE_PN0P__2134  (.L_HI(net2134));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[20]$_SDFFE_PN0P__2135  (.L_HI(net2135));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[21]$_SDFFE_PN0P__2136  (.L_HI(net2136));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[2]$_SDFFE_PN0P__2137  (.L_HI(net2137));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[3]$_SDFFE_PN0P__2138  (.L_HI(net2138));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[4]$_SDFFE_PN0P__2139  (.L_HI(net2139));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[5]$_SDFFE_PN0P__2140  (.L_HI(net2140));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[6]$_SDFFE_PN0P__2141  (.L_HI(net2141));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[7]$_SDFFE_PN0P__2142  (.L_HI(net2142));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[8]$_SDFFE_PN0P__2143  (.L_HI(net2143));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistX[9]$_SDFFE_PN0P__2144  (.L_HI(net2144));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[0]$_SDFFE_PN0P__2145  (.L_HI(net2145));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[10]$_SDFFE_PN0P__2146  (.L_HI(net2146));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[11]$_SDFFE_PN0P__2147  (.L_HI(net2147));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[12]$_SDFFE_PN0P__2148  (.L_HI(net2148));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[13]$_SDFFE_PN0P__2149  (.L_HI(net2149));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[14]$_SDFFE_PN0P__2150  (.L_HI(net2150));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[15]$_SDFFE_PN0P__2151  (.L_HI(net2151));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[16]$_SDFFE_PN0P__2152  (.L_HI(net2152));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[17]$_SDFFE_PN0P__2153  (.L_HI(net2153));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[18]$_SDFFE_PN0P__2154  (.L_HI(net2154));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[19]$_SDFFE_PN0P__2155  (.L_HI(net2155));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[1]$_SDFFE_PN0P__2156  (.L_HI(net2156));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[20]$_SDFFE_PN0P__2157  (.L_HI(net2157));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[21]$_SDFFE_PN0P__2158  (.L_HI(net2158));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[2]$_SDFFE_PN0P__2159  (.L_HI(net2159));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[3]$_SDFFE_PN0P__2160  (.L_HI(net2160));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[4]$_SDFFE_PN0P__2161  (.L_HI(net2161));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[5]$_SDFFE_PN0P__2162  (.L_HI(net2162));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[6]$_SDFFE_PN0P__2163  (.L_HI(net2163));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[7]$_SDFFE_PN0P__2164  (.L_HI(net2164));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[8]$_SDFFE_PN0P__2165  (.L_HI(net2165));
 sg13g2_tiehi \rbzero.wall_tracer.trackDistY[9]$_SDFFE_PN0P__2166  (.L_HI(net2166));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[0]$_SDFFE_PN0P__2167  (.L_HI(net2167));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[10]$_SDFFE_PN0P__2168  (.L_HI(net2168));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[11]$_SDFFE_PN0P__2169  (.L_HI(net2169));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[12]$_SDFFE_PN0P__2170  (.L_HI(net2170));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[13]$_SDFFE_PN0P__2171  (.L_HI(net2171));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[14]$_SDFFE_PN0P__2172  (.L_HI(net2172));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[15]$_SDFFE_PN0P__2173  (.L_HI(net2173));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[16]$_SDFFE_PN0P__2174  (.L_HI(net2174));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[17]$_SDFFE_PN0P__2175  (.L_HI(net2175));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[18]$_SDFFE_PN0P__2176  (.L_HI(net2176));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[19]$_SDFFE_PN0P__2177  (.L_HI(net2177));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[1]$_SDFFE_PN0P__2178  (.L_HI(net2178));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[20]$_SDFFE_PN0P__2179  (.L_HI(net2179));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[21]$_SDFFE_PN0P__2180  (.L_HI(net2180));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[2]$_SDFFE_PN0P__2181  (.L_HI(net2181));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[3]$_SDFFE_PN0P__2182  (.L_HI(net2182));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[4]$_SDFFE_PN0P__2183  (.L_HI(net2183));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[5]$_SDFFE_PN0P__2184  (.L_HI(net2184));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[6]$_SDFFE_PN0P__2185  (.L_HI(net2185));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[7]$_SDFFE_PN0P__2186  (.L_HI(net2186));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[8]$_SDFFE_PN0P__2187  (.L_HI(net2187));
 sg13g2_tiehi \rbzero.wall_tracer.visualWallDist[9]$_SDFFE_PN0P__2188  (.L_HI(net2188));
 sg13g2_tiehi \rbzero.wall_tracer.w[0]$_SDFFE_PN0P__2189  (.L_HI(net2189));
 sg13g2_tiehi \rbzero.wall_tracer.w[1]$_SDFFE_PN0P__2190  (.L_HI(net2190));
 sg13g2_tiehi \rbzero.wall_tracer.w[2]$_SDFFE_PN0P__2191  (.L_HI(net2191));
 sg13g2_tiehi \rbzero.wall_tracer.wall[0]$_SDFFE_PN0P__2192  (.L_HI(net2192));
 sg13g2_tiehi \rbzero.wall_tracer.wall[1]$_SDFFE_PN0P__2193  (.L_HI(net2193));
 sg13g2_tiehi \registered_vga_output[0]$_DFF_P__2194  (.L_HI(net2194));
 sg13g2_tiehi \registered_vga_output[1]$_DFF_P__2195  (.L_HI(net2195));
 sg13g2_tiehi \registered_vga_output[2]$_DFF_P__2196  (.L_HI(net2196));
 sg13g2_tiehi \registered_vga_output[3]$_DFF_P__2197  (.L_HI(net2197));
 sg13g2_tiehi \registered_vga_output[4]$_DFF_P__2198  (.L_HI(net2198));
 sg13g2_tiehi \registered_vga_output[5]$_DFF_P__2199  (.L_HI(net2199));
 sg13g2_tiehi \registered_vga_output[6]$_DFF_P__2200  (.L_HI(net2200));
 sg13g2_tiehi \registered_vga_output[7]$_DFF_P__2201  (.L_HI(net2201));
 sg13g2_inv_1 net2047_2 (.Y(net2203),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 net2047_3 (.Y(net2204),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 net2047_4 (.Y(net2205),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_5 (.Y(net2206),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 net2047_6 (.Y(net2207),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 net2047_7 (.Y(net2208),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 net2047_8 (.Y(net2209),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 net2047_9 (.Y(net2210),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_10 (.Y(net2211),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 net2047_11 (.Y(net2212),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 net2047_12 (.Y(net2213),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_13 (.Y(net2214),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_14 (.Y(net2215),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 net2047_15 (.Y(net2216),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_16 (.Y(net2217),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 net2047_17 (.Y(net2218),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_18 (.Y(net2219),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_19 (.Y(net2220),
    .A(clknet_leaf_95_clk));
 sg13g2_inv_1 net2047_20 (.Y(net2221),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_21 (.Y(net2222),
    .A(clknet_leaf_95_clk));
 sg13g2_inv_1 net2047_22 (.Y(net2223),
    .A(clknet_leaf_96_clk));
 sg13g2_inv_1 net2047_23 (.Y(net2224),
    .A(clknet_leaf_95_clk));
 sg13g2_inv_1 net2047_24 (.Y(net2225),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_25 (.Y(net2226),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_26 (.Y(net2227),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_27 (.Y(net2228),
    .A(clknet_leaf_95_clk));
 sg13g2_inv_1 net2047_28 (.Y(net2229),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_29 (.Y(net2230),
    .A(clknet_leaf_89_clk));
 sg13g2_inv_1 net2047_30 (.Y(net2231),
    .A(clknet_leaf_85_clk));
 sg13g2_inv_1 net2047_31 (.Y(net2232),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_32 (.Y(net2233),
    .A(clknet_leaf_85_clk));
 sg13g2_inv_1 net2047_33 (.Y(net2234),
    .A(clknet_leaf_85_clk));
 sg13g2_inv_1 net2047_34 (.Y(net2235),
    .A(clknet_leaf_85_clk));
 sg13g2_inv_1 net2047_35 (.Y(net2236),
    .A(clknet_leaf_85_clk));
 sg13g2_inv_1 net2047_36 (.Y(net2237),
    .A(clknet_leaf_84_clk));
 sg13g2_inv_1 net2047_37 (.Y(net2238),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_38 (.Y(net2239),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_39 (.Y(net2240),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_40 (.Y(net2241),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_41 (.Y(net2242),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_42 (.Y(net2243),
    .A(clknet_leaf_78_clk));
 sg13g2_inv_1 net2047_43 (.Y(net2244),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 net2047_44 (.Y(net2245),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 net2047_45 (.Y(net2246),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 net2047_46 (.Y(net2247),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 net2047_47 (.Y(net2248),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 net2047_48 (.Y(net2249),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 net2047_49 (.Y(net2250),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 net2047_50 (.Y(net2251),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 net2047_51 (.Y(net2252),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 _52 (.Y(net2253),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 _52_53 (.Y(net2254),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_54 (.Y(net2255),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_55 (.Y(net2256),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 _52_56 (.Y(net2257),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 _52_57 (.Y(net2258),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 _52_58 (.Y(net2259),
    .A(clknet_leaf_79_clk));
 sg13g2_inv_1 _52_59 (.Y(net2260),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_60 (.Y(net2261),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_61 (.Y(net2262),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_62 (.Y(net2263),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_63 (.Y(net2264),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 _52_64 (.Y(net2265),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _52_65 (.Y(net2266),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_66 (.Y(net2267),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_67 (.Y(net2268),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_68 (.Y(net2269),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_69 (.Y(net2270),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_70 (.Y(net2271),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_71 (.Y(net2272),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_72 (.Y(net2273),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_73 (.Y(net2274),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_74 (.Y(net2275),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_75 (.Y(net2276),
    .A(clknet_leaf_105_clk));
 sg13g2_inv_1 _52_76 (.Y(net2277),
    .A(clknet_leaf_105_clk));
 sg13g2_inv_1 _52_77 (.Y(net2278),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_78 (.Y(net2279),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_79 (.Y(net2280),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_80 (.Y(net2281),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_81 (.Y(net2282),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_82 (.Y(net2283),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_83 (.Y(net2284),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_84 (.Y(net2285),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_85 (.Y(net2286),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_86 (.Y(net2287),
    .A(clknet_leaf_103_clk));
 sg13g2_inv_1 _52_87 (.Y(net2288),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_88 (.Y(net2289),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_89 (.Y(net2290),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_90 (.Y(net2291),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_91 (.Y(net2292),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_92 (.Y(net2293),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_93 (.Y(net2294),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_94 (.Y(net2295),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_95 (.Y(net2296),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_96 (.Y(net2297),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_97 (.Y(net2298),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_98 (.Y(net2299),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_99 (.Y(net2300),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _52_100 (.Y(net2301),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 _52_101 (.Y(net2302),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 _52_102 (.Y(net2303),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 _52_103 (.Y(net2304),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_104 (.Y(net2305),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_105 (.Y(net2306),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_106 (.Y(net2307),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_107 (.Y(net2308),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_108 (.Y(net2309),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_109 (.Y(net2310),
    .A(clknet_leaf_105_clk));
 sg13g2_inv_1 _52_110 (.Y(net2311),
    .A(clknet_leaf_105_clk));
 sg13g2_inv_1 _52_111 (.Y(net2312),
    .A(clknet_leaf_105_clk));
 sg13g2_inv_1 _52_112 (.Y(net2313),
    .A(clknet_leaf_104_clk));
 sg13g2_inv_1 _52_113 (.Y(net2314),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_114 (.Y(net2315),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_115 (.Y(net2316),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_116 (.Y(net2317),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_117 (.Y(net2318),
    .A(clknet_leaf_100_clk));
 sg13g2_inv_1 _52_118 (.Y(net2319),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_119 (.Y(net2320),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_120 (.Y(net2321),
    .A(clknet_leaf_98_clk));
 sg13g2_inv_1 _52_121 (.Y(net2322),
    .A(clknet_leaf_102_clk));
 sg13g2_inv_1 _52_122 (.Y(net2323),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_123 (.Y(net2324),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_124 (.Y(net2325),
    .A(clknet_leaf_94_clk));
 sg13g2_inv_1 _52_125 (.Y(net2326),
    .A(clknet_leaf_94_clk));
 sg13g2_inv_1 _52_126 (.Y(net2327),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_127 (.Y(net2328),
    .A(clknet_leaf_97_clk));
 sg13g2_inv_1 _52_128 (.Y(net2329),
    .A(clknet_leaf_101_clk));
 sg13g2_inv_1 _52_129 (.Y(net2330),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _52_130 (.Y(net2331),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _52_131 (.Y(net2332),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_132 (.Y(net2333),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_133 (.Y(net2334),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _52_134 (.Y(net2335),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _52_135 (.Y(net2336),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _52_136 (.Y(net2337),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _52_137 (.Y(net2338),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_138 (.Y(net2339),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _52_139 (.Y(net2340),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _52_140 (.Y(net2341),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _52_141 (.Y(net2342),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _52_142 (.Y(net2343),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_143 (.Y(net2344),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _52_144 (.Y(net2345),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _52_145 (.Y(net2346),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _52_146 (.Y(net2347),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_147 (.Y(net2348),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_148 (.Y(net2349),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_149 (.Y(net2350),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_150 (.Y(net2351),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_151 (.Y(net2352),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_152 (.Y(net2353),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _52_153 (.Y(net2354),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _52_154 (.Y(net2355),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _52_155 (.Y(net2356),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_156 (.Y(net2357),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_157 (.Y(net2358),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _52_158 (.Y(net2359),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_159 (.Y(net2360),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_160 (.Y(net2361),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_161 (.Y(net2362),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_162 (.Y(net2363),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_163 (.Y(net2364),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_164 (.Y(net2365),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_165 (.Y(net2366),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_166 (.Y(net2367),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_167 (.Y(net2368),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_168 (.Y(net2369),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_169 (.Y(net2370),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _52_170 (.Y(net2371),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _52_171 (.Y(net2372),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_172 (.Y(net2373),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_173 (.Y(net2374),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_174 (.Y(net2375),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_175 (.Y(net2376),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_176 (.Y(net2377),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _52_177 (.Y(net2378),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _52_178 (.Y(net2379),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _52_179 (.Y(net2380),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _180 (.Y(net2381),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _180_181 (.Y(net2382),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _180_182 (.Y(net2383),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _180_183 (.Y(net2384),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _180_184 (.Y(net2385),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _180_185 (.Y(net2386),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _180_186 (.Y(net2387),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_187 (.Y(net2388),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_188 (.Y(net2389),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_189 (.Y(net2390),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_190 (.Y(net2391),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_191 (.Y(net2392),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _180_192 (.Y(net2393),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _180_193 (.Y(net2394),
    .A(clknet_leaf_77_clk));
 sg13g2_inv_1 _180_194 (.Y(net2395),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 _180_195 (.Y(net2396),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_196 (.Y(net2397),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_197 (.Y(net2398),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_198 (.Y(net2399),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_199 (.Y(net2400),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_200 (.Y(net2401),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_201 (.Y(net2402),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_202 (.Y(net2403),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_203 (.Y(net2404),
    .A(clknet_leaf_99_clk));
 sg13g2_inv_1 _180_204 (.Y(net2405),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_205 (.Y(net2406),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_206 (.Y(net2407),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_207 (.Y(net2408),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_208 (.Y(net2409),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_209 (.Y(net2410),
    .A(clknet_leaf_75_clk));
 sg13g2_inv_1 _180_210 (.Y(net2411),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 _180_211 (.Y(net2412),
    .A(clknet_leaf_76_clk));
 sg13g2_inv_1 _180_212 (.Y(net2413),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_213 (.Y(net2414),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_214 (.Y(net2415),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_215 (.Y(net2416),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_216 (.Y(net2417),
    .A(clknet_leaf_74_clk));
 sg13g2_inv_1 _180_217 (.Y(net2418),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_218 (.Y(net2419),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_219 (.Y(net2420),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_220 (.Y(net2421),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_221 (.Y(net2422),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_222 (.Y(net2423),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_223 (.Y(net2424),
    .A(clknet_leaf_73_clk));
 sg13g2_inv_1 _180_224 (.Y(net2425),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_225 (.Y(net2426),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_226 (.Y(net2427),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_227 (.Y(net2428),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_228 (.Y(net2429),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_229 (.Y(net2430),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_230 (.Y(net2431),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_231 (.Y(net2432),
    .A(clknet_leaf_71_clk));
 sg13g2_inv_1 _180_232 (.Y(net2433),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_233 (.Y(net2434),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_234 (.Y(net2435),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_235 (.Y(net2436),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_236 (.Y(net2437),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_237 (.Y(net2438),
    .A(clknet_leaf_70_clk));
 sg13g2_inv_1 _180_238 (.Y(net2439),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _180_239 (.Y(net2440),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_240 (.Y(net2441),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_241 (.Y(net2442),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _180_242 (.Y(net2443),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _180_243 (.Y(net2444),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _180_244 (.Y(net2445),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _180_245 (.Y(net2446),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_246 (.Y(net2447),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_247 (.Y(net2448),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_248 (.Y(net2449),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_249 (.Y(net2450),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 _180_250 (.Y(net2451),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _180_251 (.Y(net2452),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 _180_252 (.Y(net2453),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_253 (.Y(net2454),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 _180_254 (.Y(net2455),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_255 (.Y(net2456),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_256 (.Y(net2457),
    .A(clknet_leaf_72_clk));
 sg13g2_inv_1 _180_257 (.Y(net2458),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _180_258 (.Y(net2459),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _180_259 (.Y(net2460),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _180_260 (.Y(net2461),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _180_261 (.Y(net2462),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_262 (.Y(net2463),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_263 (.Y(net2464),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_264 (.Y(net2465),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _180_265 (.Y(net2466),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _180_266 (.Y(net2467),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _180_267 (.Y(net2468),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _180_268 (.Y(net2469),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_269 (.Y(net2470),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_270 (.Y(net2471),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_271 (.Y(net2472),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_272 (.Y(net2473),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_273 (.Y(net2474),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_274 (.Y(net2475),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_275 (.Y(net2476),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_276 (.Y(net2477),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _180_277 (.Y(net2478),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_278 (.Y(net2479),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_279 (.Y(net2480),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_280 (.Y(net2481),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _180_281 (.Y(net2482),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_282 (.Y(net2483),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_283 (.Y(net2484),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_284 (.Y(net2485),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_285 (.Y(net2486),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_286 (.Y(net2487),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_287 (.Y(net2488),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _180_288 (.Y(net2489),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_289 (.Y(net2490),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _180_290 (.Y(net2491),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _180_291 (.Y(net2492),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_292 (.Y(net2493),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_293 (.Y(net2494),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_294 (.Y(net2495),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _180_295 (.Y(net2496),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _180_296 (.Y(net2497),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _180_297 (.Y(net2498),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _180_298 (.Y(net2499),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _180_299 (.Y(net2500),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _180_300 (.Y(net2501),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _180_301 (.Y(net2502),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_302 (.Y(net2503),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_303 (.Y(net2504),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _180_304 (.Y(net2505),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _180_305 (.Y(net2506),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _180_306 (.Y(net2507),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _180_307 (.Y(net2508),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _308 (.Y(net2509),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _308_309 (.Y(net2510),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _308_310 (.Y(net2511),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _308_311 (.Y(net2512),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _308_312 (.Y(net2513),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _308_313 (.Y(net2514),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _308_314 (.Y(net2515),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_315 (.Y(net2516),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _308_316 (.Y(net2517),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _308_317 (.Y(net2518),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_318 (.Y(net2519),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_319 (.Y(net2520),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _308_320 (.Y(net2521),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _308_321 (.Y(net2522),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_322 (.Y(net2523),
    .A(clknet_leaf_68_clk));
 sg13g2_inv_1 _308_323 (.Y(net2524),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_324 (.Y(net2525),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_325 (.Y(net2526),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_326 (.Y(net2527),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_327 (.Y(net2528),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_328 (.Y(net2529),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 _308_329 (.Y(net2530),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_330 (.Y(net2531),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_331 (.Y(net2532),
    .A(clknet_leaf_80_clk));
 sg13g2_inv_1 _308_332 (.Y(net2533),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_333 (.Y(net2534),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_334 (.Y(net2535),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_335 (.Y(net2536),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_336 (.Y(net2537),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_337 (.Y(net2538),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_338 (.Y(net2539),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_339 (.Y(net2540),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_340 (.Y(net2541),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_341 (.Y(net2542),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _308_342 (.Y(net2543),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_343 (.Y(net2544),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_344 (.Y(net2545),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_345 (.Y(net2546),
    .A(clknet_leaf_82_clk));
 sg13g2_inv_1 _308_346 (.Y(net2547),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_347 (.Y(net2548),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_348 (.Y(net2549),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_349 (.Y(net2550),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_350 (.Y(net2551),
    .A(clknet_leaf_83_clk));
 sg13g2_inv_1 _308_351 (.Y(net2552),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_352 (.Y(net2553),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _308_353 (.Y(net2554),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _308_354 (.Y(net2555),
    .A(clknet_leaf_81_clk));
 sg13g2_inv_1 _308_355 (.Y(net2556),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _308_356 (.Y(net2557),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_357 (.Y(net2558),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_358 (.Y(net2559),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_359 (.Y(net2560),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_360 (.Y(net2561),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _308_361 (.Y(net2562),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _308_362 (.Y(net2563),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_363 (.Y(net2564),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_364 (.Y(net2565),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _308_365 (.Y(net2566),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _308_366 (.Y(net2567),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _308_367 (.Y(net2568),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_368 (.Y(net2569),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_369 (.Y(net2570),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _308_370 (.Y(net2571),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_371 (.Y(net2572),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_372 (.Y(net2573),
    .A(clknet_leaf_66_clk));
 sg13g2_inv_1 _308_373 (.Y(net2574),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_374 (.Y(net2575),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_375 (.Y(net2576),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_376 (.Y(net2577),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_377 (.Y(net2578),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _308_378 (.Y(net2579),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _308_379 (.Y(net2580),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_380 (.Y(net2581),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _308_381 (.Y(net2582),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _308_382 (.Y(net2583),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_383 (.Y(net2584),
    .A(clknet_leaf_69_clk));
 sg13g2_inv_1 _308_384 (.Y(net2585),
    .A(clknet_leaf_67_clk));
 sg13g2_inv_1 _308_385 (.Y(net2586),
    .A(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_5_0__f_clk (.X(clknet_5_0__leaf_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_5_1__f_clk (.X(clknet_5_1__leaf_clk),
    .A(clknet_4_0_0_clk));
 sg13g2_buf_4 clkbuf_5_2__f_clk (.X(clknet_5_2__leaf_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_5_3__f_clk (.X(clknet_5_3__leaf_clk),
    .A(clknet_4_1_0_clk));
 sg13g2_buf_4 clkbuf_5_4__f_clk (.X(clknet_5_4__leaf_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_5_5__f_clk (.X(clknet_5_5__leaf_clk),
    .A(clknet_4_2_0_clk));
 sg13g2_buf_4 clkbuf_5_6__f_clk (.X(clknet_5_6__leaf_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_5_7__f_clk (.X(clknet_5_7__leaf_clk),
    .A(clknet_4_3_0_clk));
 sg13g2_buf_4 clkbuf_5_8__f_clk (.X(clknet_5_8__leaf_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_5_9__f_clk (.X(clknet_5_9__leaf_clk),
    .A(clknet_4_4_0_clk));
 sg13g2_buf_4 clkbuf_5_10__f_clk (.X(clknet_5_10__leaf_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_5_11__f_clk (.X(clknet_5_11__leaf_clk),
    .A(clknet_4_5_0_clk));
 sg13g2_buf_4 clkbuf_5_12__f_clk (.X(clknet_5_12__leaf_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_5_13__f_clk (.X(clknet_5_13__leaf_clk),
    .A(clknet_4_6_0_clk));
 sg13g2_buf_4 clkbuf_5_14__f_clk (.X(clknet_5_14__leaf_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_5_15__f_clk (.X(clknet_5_15__leaf_clk),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_4 clkbuf_5_16__f_clk (.X(clknet_5_16__leaf_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_5_17__f_clk (.X(clknet_5_17__leaf_clk),
    .A(clknet_4_8_0_clk));
 sg13g2_buf_4 clkbuf_5_18__f_clk (.X(clknet_5_18__leaf_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_5_19__f_clk (.X(clknet_5_19__leaf_clk),
    .A(clknet_4_9_0_clk));
 sg13g2_buf_4 clkbuf_5_20__f_clk (.X(clknet_5_20__leaf_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_5_21__f_clk (.X(clknet_5_21__leaf_clk),
    .A(clknet_4_10_0_clk));
 sg13g2_buf_4 clkbuf_5_22__f_clk (.X(clknet_5_22__leaf_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_5_23__f_clk (.X(clknet_5_23__leaf_clk),
    .A(clknet_4_11_0_clk));
 sg13g2_buf_4 clkbuf_5_24__f_clk (.X(clknet_5_24__leaf_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_5_25__f_clk (.X(clknet_5_25__leaf_clk),
    .A(clknet_4_12_0_clk));
 sg13g2_buf_4 clkbuf_5_26__f_clk (.X(clknet_5_26__leaf_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_5_27__f_clk (.X(clknet_5_27__leaf_clk),
    .A(clknet_4_13_0_clk));
 sg13g2_buf_4 clkbuf_5_28__f_clk (.X(clknet_5_28__leaf_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_5_29__f_clk (.X(clknet_5_29__leaf_clk),
    .A(clknet_4_14_0_clk));
 sg13g2_buf_4 clkbuf_5_30__f_clk (.X(clknet_5_30__leaf_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_4 clkbuf_5_31__f_clk (.X(clknet_5_31__leaf_clk),
    .A(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_169_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00000_));
 sg13g2_antennanp ANTENNA_2 (.A(_00499_));
 sg13g2_antennanp ANTENNA_3 (.A(_07956_));
 sg13g2_antennanp ANTENNA_4 (.A(_07956_));
 sg13g2_antennanp ANTENNA_5 (.A(_07956_));
 sg13g2_antennanp ANTENNA_6 (.A(_08542_));
 sg13g2_antennanp ANTENNA_7 (.A(_08542_));
 sg13g2_antennanp ANTENNA_8 (.A(_08542_));
 sg13g2_antennanp ANTENNA_9 (.A(_08542_));
 sg13g2_antennanp ANTENNA_10 (.A(_08542_));
 sg13g2_antennanp ANTENNA_11 (.A(_08542_));
 sg13g2_antennanp ANTENNA_12 (.A(_08542_));
 sg13g2_antennanp ANTENNA_13 (.A(_08542_));
 sg13g2_antennanp ANTENNA_14 (.A(_08542_));
 sg13g2_antennanp ANTENNA_15 (.A(_08542_));
 sg13g2_antennanp ANTENNA_16 (.A(_08542_));
 sg13g2_antennanp ANTENNA_17 (.A(_08543_));
 sg13g2_antennanp ANTENNA_18 (.A(_08543_));
 sg13g2_antennanp ANTENNA_19 (.A(_08543_));
 sg13g2_antennanp ANTENNA_20 (.A(_08543_));
 sg13g2_antennanp ANTENNA_21 (.A(_08543_));
 sg13g2_antennanp ANTENNA_22 (.A(_08639_));
 sg13g2_antennanp ANTENNA_23 (.A(_08639_));
 sg13g2_antennanp ANTENNA_24 (.A(_10379_));
 sg13g2_antennanp ANTENNA_25 (.A(_10379_));
 sg13g2_antennanp ANTENNA_26 (.A(_10379_));
 sg13g2_antennanp ANTENNA_27 (.A(_11353_));
 sg13g2_antennanp ANTENNA_28 (.A(_11353_));
 sg13g2_antennanp ANTENNA_29 (.A(_11353_));
 sg13g2_antennanp ANTENNA_30 (.A(_11353_));
 sg13g2_antennanp ANTENNA_31 (.A(_13629_));
 sg13g2_antennanp ANTENNA_32 (.A(_13724_));
 sg13g2_antennanp ANTENNA_33 (.A(_13724_));
 sg13g2_antennanp ANTENNA_34 (.A(_13724_));
 sg13g2_antennanp ANTENNA_35 (.A(_13724_));
 sg13g2_antennanp ANTENNA_36 (.A(_13724_));
 sg13g2_antennanp ANTENNA_37 (.A(\rbzero.spi_registers.vshift[3] ));
 sg13g2_antennanp ANTENNA_38 (.A(\rbzero.spi_registers.vshift[3] ));
 sg13g2_antennanp ANTENNA_39 (.A(\rbzero.spi_registers.vshift[3] ));
 sg13g2_antennanp ANTENNA_40 (.A(net9));
 sg13g2_antennanp ANTENNA_41 (.A(net10));
 sg13g2_antennanp ANTENNA_42 (.A(net10));
 sg13g2_antennanp ANTENNA_43 (.A(net10));
 sg13g2_antennanp ANTENNA_44 (.A(net562));
 sg13g2_antennanp ANTENNA_45 (.A(net562));
 sg13g2_antennanp ANTENNA_46 (.A(net562));
 sg13g2_antennanp ANTENNA_47 (.A(net562));
 sg13g2_antennanp ANTENNA_48 (.A(net562));
 sg13g2_antennanp ANTENNA_49 (.A(net562));
 sg13g2_antennanp ANTENNA_50 (.A(net562));
 sg13g2_antennanp ANTENNA_51 (.A(net562));
 sg13g2_antennanp ANTENNA_52 (.A(net562));
 sg13g2_antennanp ANTENNA_53 (.A(net700));
 sg13g2_antennanp ANTENNA_54 (.A(net700));
 sg13g2_antennanp ANTENNA_55 (.A(net700));
 sg13g2_antennanp ANTENNA_56 (.A(net700));
 sg13g2_antennanp ANTENNA_57 (.A(net700));
 sg13g2_antennanp ANTENNA_58 (.A(net700));
 sg13g2_antennanp ANTENNA_59 (.A(net700));
 sg13g2_antennanp ANTENNA_60 (.A(net700));
 sg13g2_antennanp ANTENNA_61 (.A(net700));
 sg13g2_antennanp ANTENNA_62 (.A(net700));
 sg13g2_antennanp ANTENNA_63 (.A(net700));
 sg13g2_antennanp ANTENNA_64 (.A(net700));
 sg13g2_antennanp ANTENNA_65 (.A(net700));
 sg13g2_antennanp ANTENNA_66 (.A(_00499_));
 sg13g2_antennanp ANTENNA_67 (.A(_07956_));
 sg13g2_antennanp ANTENNA_68 (.A(_07956_));
 sg13g2_antennanp ANTENNA_69 (.A(_07956_));
 sg13g2_antennanp ANTENNA_70 (.A(_08543_));
 sg13g2_antennanp ANTENNA_71 (.A(_08543_));
 sg13g2_antennanp ANTENNA_72 (.A(_08543_));
 sg13g2_antennanp ANTENNA_73 (.A(_08543_));
 sg13g2_antennanp ANTENNA_74 (.A(_08543_));
 sg13g2_antennanp ANTENNA_75 (.A(_08543_));
 sg13g2_antennanp ANTENNA_76 (.A(_08543_));
 sg13g2_antennanp ANTENNA_77 (.A(_08543_));
 sg13g2_antennanp ANTENNA_78 (.A(_08639_));
 sg13g2_antennanp ANTENNA_79 (.A(_08639_));
 sg13g2_antennanp ANTENNA_80 (.A(_10379_));
 sg13g2_antennanp ANTENNA_81 (.A(_10379_));
 sg13g2_antennanp ANTENNA_82 (.A(_10379_));
 sg13g2_antennanp ANTENNA_83 (.A(_13724_));
 sg13g2_antennanp ANTENNA_84 (.A(_13724_));
 sg13g2_antennanp ANTENNA_85 (.A(_13724_));
 sg13g2_antennanp ANTENNA_86 (.A(_13724_));
 sg13g2_antennanp ANTENNA_87 (.A(_13724_));
 sg13g2_antennanp ANTENNA_88 (.A(_13724_));
 sg13g2_antennanp ANTENNA_89 (.A(_13724_));
 sg13g2_antennanp ANTENNA_90 (.A(_13724_));
 sg13g2_antennanp ANTENNA_91 (.A(net9));
 sg13g2_antennanp ANTENNA_92 (.A(net2347));
 sg13g2_antennanp ANTENNA_93 (.A(_00499_));
 sg13g2_antennanp ANTENNA_94 (.A(_07956_));
 sg13g2_antennanp ANTENNA_95 (.A(_07956_));
 sg13g2_antennanp ANTENNA_96 (.A(_07956_));
 sg13g2_antennanp ANTENNA_97 (.A(_07956_));
 sg13g2_antennanp ANTENNA_98 (.A(_10379_));
 sg13g2_antennanp ANTENNA_99 (.A(_10379_));
 sg13g2_antennanp ANTENNA_100 (.A(_10379_));
 sg13g2_antennanp ANTENNA_101 (.A(_13724_));
 sg13g2_antennanp ANTENNA_102 (.A(_13724_));
 sg13g2_antennanp ANTENNA_103 (.A(_13724_));
 sg13g2_antennanp ANTENNA_104 (.A(_13724_));
 sg13g2_antennanp ANTENNA_105 (.A(_13724_));
 sg13g2_antennanp ANTENNA_106 (.A(net9));
 sg13g2_antennanp ANTENNA_107 (.A(net2336));
 sg13g2_antennanp ANTENNA_108 (.A(net2337));
 sg13g2_antennanp ANTENNA_109 (.A(_00499_));
 sg13g2_antennanp ANTENNA_110 (.A(_10379_));
 sg13g2_antennanp ANTENNA_111 (.A(_10379_));
 sg13g2_antennanp ANTENNA_112 (.A(_10379_));
 sg13g2_antennanp ANTENNA_113 (.A(_13724_));
 sg13g2_antennanp ANTENNA_114 (.A(_13724_));
 sg13g2_antennanp ANTENNA_115 (.A(_13724_));
 sg13g2_antennanp ANTENNA_116 (.A(_13724_));
 sg13g2_antennanp ANTENNA_117 (.A(_13724_));
 sg13g2_antennanp ANTENNA_118 (.A(_13724_));
 sg13g2_antennanp ANTENNA_119 (.A(_13724_));
 sg13g2_antennanp ANTENNA_120 (.A(net9));
 sg13g2_antennanp ANTENNA_121 (.A(_00499_));
 sg13g2_antennanp ANTENNA_122 (.A(_10379_));
 sg13g2_antennanp ANTENNA_123 (.A(_10379_));
 sg13g2_antennanp ANTENNA_124 (.A(_10379_));
 sg13g2_antennanp ANTENNA_125 (.A(_10379_));
 sg13g2_antennanp ANTENNA_126 (.A(_10379_));
 sg13g2_antennanp ANTENNA_127 (.A(_10379_));
 sg13g2_antennanp ANTENNA_128 (.A(_13724_));
 sg13g2_antennanp ANTENNA_129 (.A(_13724_));
 sg13g2_antennanp ANTENNA_130 (.A(_13724_));
 sg13g2_antennanp ANTENNA_131 (.A(_13724_));
 sg13g2_antennanp ANTENNA_132 (.A(_13724_));
 sg13g2_antennanp ANTENNA_133 (.A(_13724_));
 sg13g2_antennanp ANTENNA_134 (.A(_13724_));
 sg13g2_antennanp ANTENNA_135 (.A(_13724_));
 sg13g2_antennanp ANTENNA_136 (.A(net9));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_42 ();
 sg13g2_fill_1 FILLER_0_46 ();
 sg13g2_decap_8 FILLER_0_51 ();
 sg13g2_decap_8 FILLER_0_58 ();
 sg13g2_decap_8 FILLER_0_65 ();
 sg13g2_decap_8 FILLER_0_72 ();
 sg13g2_decap_8 FILLER_0_79 ();
 sg13g2_decap_8 FILLER_0_86 ();
 sg13g2_decap_8 FILLER_0_93 ();
 sg13g2_decap_8 FILLER_0_100 ();
 sg13g2_decap_8 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_142 ();
 sg13g2_decap_8 FILLER_0_149 ();
 sg13g2_decap_8 FILLER_0_156 ();
 sg13g2_decap_8 FILLER_0_163 ();
 sg13g2_fill_1 FILLER_0_170 ();
 sg13g2_decap_4 FILLER_0_176 ();
 sg13g2_fill_1 FILLER_0_180 ();
 sg13g2_fill_2 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_217 ();
 sg13g2_fill_2 FILLER_0_244 ();
 sg13g2_fill_1 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_281 ();
 sg13g2_fill_1 FILLER_0_288 ();
 sg13g2_fill_2 FILLER_0_323 ();
 sg13g2_fill_1 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_fill_1 FILLER_0_392 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_fill_2 FILLER_0_478 ();
 sg13g2_fill_2 FILLER_0_577 ();
 sg13g2_fill_1 FILLER_0_579 ();
 sg13g2_fill_1 FILLER_0_607 ();
 sg13g2_fill_2 FILLER_0_616 ();
 sg13g2_fill_1 FILLER_0_618 ();
 sg13g2_fill_2 FILLER_0_628 ();
 sg13g2_fill_1 FILLER_0_630 ();
 sg13g2_fill_1 FILLER_0_665 ();
 sg13g2_fill_1 FILLER_0_675 ();
 sg13g2_fill_2 FILLER_0_702 ();
 sg13g2_fill_1 FILLER_0_708 ();
 sg13g2_fill_1 FILLER_0_718 ();
 sg13g2_fill_2 FILLER_0_723 ();
 sg13g2_fill_2 FILLER_0_729 ();
 sg13g2_decap_4 FILLER_0_761 ();
 sg13g2_fill_2 FILLER_0_770 ();
 sg13g2_fill_2 FILLER_0_786 ();
 sg13g2_fill_1 FILLER_0_799 ();
 sg13g2_fill_2 FILLER_0_809 ();
 sg13g2_fill_1 FILLER_0_811 ();
 sg13g2_fill_2 FILLER_0_816 ();
 sg13g2_fill_2 FILLER_0_822 ();
 sg13g2_fill_2 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_834 ();
 sg13g2_fill_1 FILLER_0_841 ();
 sg13g2_decap_8 FILLER_0_846 ();
 sg13g2_fill_2 FILLER_0_853 ();
 sg13g2_fill_1 FILLER_0_855 ();
 sg13g2_decap_8 FILLER_0_872 ();
 sg13g2_fill_1 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_900 ();
 sg13g2_decap_8 FILLER_0_907 ();
 sg13g2_decap_8 FILLER_0_914 ();
 sg13g2_decap_8 FILLER_0_921 ();
 sg13g2_decap_8 FILLER_0_928 ();
 sg13g2_decap_8 FILLER_0_935 ();
 sg13g2_decap_8 FILLER_0_942 ();
 sg13g2_decap_8 FILLER_0_949 ();
 sg13g2_decap_8 FILLER_0_956 ();
 sg13g2_decap_8 FILLER_0_963 ();
 sg13g2_decap_8 FILLER_0_970 ();
 sg13g2_decap_8 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_984 ();
 sg13g2_decap_8 FILLER_0_991 ();
 sg13g2_decap_8 FILLER_0_998 ();
 sg13g2_decap_8 FILLER_0_1005 ();
 sg13g2_decap_8 FILLER_0_1012 ();
 sg13g2_decap_8 FILLER_0_1019 ();
 sg13g2_decap_8 FILLER_0_1026 ();
 sg13g2_decap_8 FILLER_0_1033 ();
 sg13g2_decap_8 FILLER_0_1040 ();
 sg13g2_decap_8 FILLER_0_1047 ();
 sg13g2_decap_8 FILLER_0_1054 ();
 sg13g2_decap_8 FILLER_0_1061 ();
 sg13g2_decap_8 FILLER_0_1068 ();
 sg13g2_decap_8 FILLER_0_1075 ();
 sg13g2_decap_8 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1089 ();
 sg13g2_decap_8 FILLER_0_1096 ();
 sg13g2_decap_8 FILLER_0_1103 ();
 sg13g2_decap_8 FILLER_0_1110 ();
 sg13g2_decap_8 FILLER_0_1117 ();
 sg13g2_decap_8 FILLER_0_1124 ();
 sg13g2_decap_8 FILLER_0_1131 ();
 sg13g2_decap_8 FILLER_0_1138 ();
 sg13g2_decap_8 FILLER_0_1145 ();
 sg13g2_decap_8 FILLER_0_1152 ();
 sg13g2_decap_8 FILLER_0_1159 ();
 sg13g2_decap_8 FILLER_0_1166 ();
 sg13g2_decap_8 FILLER_0_1173 ();
 sg13g2_decap_8 FILLER_0_1180 ();
 sg13g2_decap_8 FILLER_0_1187 ();
 sg13g2_decap_8 FILLER_0_1194 ();
 sg13g2_decap_8 FILLER_0_1201 ();
 sg13g2_decap_8 FILLER_0_1208 ();
 sg13g2_decap_8 FILLER_0_1215 ();
 sg13g2_decap_8 FILLER_0_1222 ();
 sg13g2_decap_8 FILLER_0_1229 ();
 sg13g2_fill_2 FILLER_0_1236 ();
 sg13g2_fill_1 FILLER_0_1238 ();
 sg13g2_fill_2 FILLER_0_1243 ();
 sg13g2_decap_8 FILLER_0_1250 ();
 sg13g2_decap_8 FILLER_0_1257 ();
 sg13g2_decap_8 FILLER_0_1264 ();
 sg13g2_decap_8 FILLER_0_1271 ();
 sg13g2_decap_8 FILLER_0_1278 ();
 sg13g2_decap_4 FILLER_0_1285 ();
 sg13g2_fill_1 FILLER_0_1289 ();
 sg13g2_decap_8 FILLER_0_1303 ();
 sg13g2_fill_1 FILLER_0_1310 ();
 sg13g2_decap_4 FILLER_0_1335 ();
 sg13g2_fill_2 FILLER_0_1339 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_4 FILLER_0_1365 ();
 sg13g2_decap_8 FILLER_0_1374 ();
 sg13g2_decap_4 FILLER_0_1410 ();
 sg13g2_fill_1 FILLER_0_1414 ();
 sg13g2_fill_2 FILLER_0_1419 ();
 sg13g2_fill_1 FILLER_0_1442 ();
 sg13g2_fill_2 FILLER_0_1456 ();
 sg13g2_fill_2 FILLER_0_1485 ();
 sg13g2_fill_1 FILLER_0_1487 ();
 sg13g2_decap_4 FILLER_0_1495 ();
 sg13g2_fill_2 FILLER_0_1499 ();
 sg13g2_decap_4 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_fill_2 FILLER_0_1576 ();
 sg13g2_fill_1 FILLER_0_1578 ();
 sg13g2_decap_4 FILLER_0_1584 ();
 sg13g2_fill_1 FILLER_0_1597 ();
 sg13g2_fill_1 FILLER_0_1607 ();
 sg13g2_fill_1 FILLER_0_1613 ();
 sg13g2_fill_1 FILLER_0_1618 ();
 sg13g2_fill_1 FILLER_0_1623 ();
 sg13g2_decap_8 FILLER_0_1632 ();
 sg13g2_decap_4 FILLER_0_1639 ();
 sg13g2_fill_1 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1649 ();
 sg13g2_decap_8 FILLER_0_1656 ();
 sg13g2_fill_2 FILLER_0_1663 ();
 sg13g2_fill_1 FILLER_0_1665 ();
 sg13g2_decap_4 FILLER_0_1675 ();
 sg13g2_fill_1 FILLER_0_1684 ();
 sg13g2_decap_8 FILLER_0_1697 ();
 sg13g2_decap_8 FILLER_0_1704 ();
 sg13g2_decap_8 FILLER_0_1711 ();
 sg13g2_decap_8 FILLER_0_1718 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_decap_8 FILLER_0_1739 ();
 sg13g2_decap_8 FILLER_0_1746 ();
 sg13g2_decap_8 FILLER_0_1753 ();
 sg13g2_decap_8 FILLER_0_1760 ();
 sg13g2_decap_8 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_4 FILLER_1_35 ();
 sg13g2_fill_1 FILLER_1_39 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_fill_1 FILLER_1_203 ();
 sg13g2_decap_4 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_212 ();
 sg13g2_fill_2 FILLER_1_235 ();
 sg13g2_decap_8 FILLER_1_264 ();
 sg13g2_decap_8 FILLER_1_271 ();
 sg13g2_fill_1 FILLER_1_278 ();
 sg13g2_fill_2 FILLER_1_309 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_341 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_fill_1 FILLER_1_355 ();
 sg13g2_fill_1 FILLER_1_360 ();
 sg13g2_fill_1 FILLER_1_364 ();
 sg13g2_fill_1 FILLER_1_369 ();
 sg13g2_fill_2 FILLER_1_374 ();
 sg13g2_fill_2 FILLER_1_380 ();
 sg13g2_fill_2 FILLER_1_410 ();
 sg13g2_fill_1 FILLER_1_499 ();
 sg13g2_fill_2 FILLER_1_526 ();
 sg13g2_fill_2 FILLER_1_537 ();
 sg13g2_fill_2 FILLER_1_544 ();
 sg13g2_fill_1 FILLER_1_551 ();
 sg13g2_fill_1 FILLER_1_560 ();
 sg13g2_fill_2 FILLER_1_566 ();
 sg13g2_fill_1 FILLER_1_568 ();
 sg13g2_fill_1 FILLER_1_595 ();
 sg13g2_fill_1 FILLER_1_622 ();
 sg13g2_fill_1 FILLER_1_654 ();
 sg13g2_fill_2 FILLER_1_660 ();
 sg13g2_fill_1 FILLER_1_662 ();
 sg13g2_fill_2 FILLER_1_710 ();
 sg13g2_fill_1 FILLER_1_753 ();
 sg13g2_fill_2 FILLER_1_758 ();
 sg13g2_fill_1 FILLER_1_760 ();
 sg13g2_fill_1 FILLER_1_774 ();
 sg13g2_fill_1 FILLER_1_780 ();
 sg13g2_fill_2 FILLER_1_789 ();
 sg13g2_fill_1 FILLER_1_795 ();
 sg13g2_fill_1 FILLER_1_806 ();
 sg13g2_fill_1 FILLER_1_812 ();
 sg13g2_fill_1 FILLER_1_817 ();
 sg13g2_fill_2 FILLER_1_823 ();
 sg13g2_fill_2 FILLER_1_845 ();
 sg13g2_fill_1 FILLER_1_855 ();
 sg13g2_fill_2 FILLER_1_871 ();
 sg13g2_fill_2 FILLER_1_891 ();
 sg13g2_decap_8 FILLER_1_901 ();
 sg13g2_decap_8 FILLER_1_908 ();
 sg13g2_fill_1 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_920 ();
 sg13g2_decap_8 FILLER_1_927 ();
 sg13g2_decap_8 FILLER_1_934 ();
 sg13g2_decap_8 FILLER_1_941 ();
 sg13g2_decap_8 FILLER_1_948 ();
 sg13g2_decap_8 FILLER_1_955 ();
 sg13g2_decap_8 FILLER_1_962 ();
 sg13g2_decap_8 FILLER_1_969 ();
 sg13g2_decap_8 FILLER_1_976 ();
 sg13g2_decap_8 FILLER_1_983 ();
 sg13g2_decap_8 FILLER_1_990 ();
 sg13g2_decap_8 FILLER_1_997 ();
 sg13g2_decap_8 FILLER_1_1004 ();
 sg13g2_decap_8 FILLER_1_1011 ();
 sg13g2_decap_8 FILLER_1_1018 ();
 sg13g2_decap_8 FILLER_1_1025 ();
 sg13g2_decap_8 FILLER_1_1032 ();
 sg13g2_decap_8 FILLER_1_1039 ();
 sg13g2_decap_4 FILLER_1_1046 ();
 sg13g2_decap_8 FILLER_1_1054 ();
 sg13g2_decap_4 FILLER_1_1061 ();
 sg13g2_decap_8 FILLER_1_1070 ();
 sg13g2_decap_8 FILLER_1_1077 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_8 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_fill_1 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1110 ();
 sg13g2_decap_8 FILLER_1_1117 ();
 sg13g2_decap_8 FILLER_1_1124 ();
 sg13g2_decap_8 FILLER_1_1131 ();
 sg13g2_decap_8 FILLER_1_1138 ();
 sg13g2_decap_8 FILLER_1_1145 ();
 sg13g2_decap_8 FILLER_1_1152 ();
 sg13g2_decap_8 FILLER_1_1159 ();
 sg13g2_decap_8 FILLER_1_1166 ();
 sg13g2_decap_8 FILLER_1_1173 ();
 sg13g2_decap_4 FILLER_1_1180 ();
 sg13g2_decap_8 FILLER_1_1192 ();
 sg13g2_decap_8 FILLER_1_1199 ();
 sg13g2_decap_8 FILLER_1_1206 ();
 sg13g2_decap_8 FILLER_1_1213 ();
 sg13g2_fill_1 FILLER_1_1220 ();
 sg13g2_fill_2 FILLER_1_1234 ();
 sg13g2_fill_1 FILLER_1_1247 ();
 sg13g2_fill_1 FILLER_1_1252 ();
 sg13g2_decap_8 FILLER_1_1258 ();
 sg13g2_decap_8 FILLER_1_1265 ();
 sg13g2_decap_4 FILLER_1_1272 ();
 sg13g2_fill_1 FILLER_1_1276 ();
 sg13g2_fill_2 FILLER_1_1281 ();
 sg13g2_fill_1 FILLER_1_1283 ();
 sg13g2_fill_1 FILLER_1_1308 ();
 sg13g2_decap_4 FILLER_1_1323 ();
 sg13g2_fill_2 FILLER_1_1327 ();
 sg13g2_fill_2 FILLER_1_1334 ();
 sg13g2_fill_1 FILLER_1_1342 ();
 sg13g2_fill_1 FILLER_1_1351 ();
 sg13g2_fill_2 FILLER_1_1358 ();
 sg13g2_fill_2 FILLER_1_1373 ();
 sg13g2_fill_2 FILLER_1_1398 ();
 sg13g2_fill_1 FILLER_1_1400 ();
 sg13g2_decap_4 FILLER_1_1409 ();
 sg13g2_fill_1 FILLER_1_1452 ();
 sg13g2_fill_2 FILLER_1_1463 ();
 sg13g2_fill_1 FILLER_1_1469 ();
 sg13g2_fill_1 FILLER_1_1474 ();
 sg13g2_fill_1 FILLER_1_1486 ();
 sg13g2_fill_2 FILLER_1_1520 ();
 sg13g2_fill_1 FILLER_1_1522 ();
 sg13g2_fill_2 FILLER_1_1551 ();
 sg13g2_fill_1 FILLER_1_1553 ();
 sg13g2_decap_8 FILLER_1_1575 ();
 sg13g2_decap_4 FILLER_1_1582 ();
 sg13g2_fill_2 FILLER_1_1614 ();
 sg13g2_fill_2 FILLER_1_1621 ();
 sg13g2_fill_1 FILLER_1_1623 ();
 sg13g2_decap_8 FILLER_1_1632 ();
 sg13g2_decap_8 FILLER_1_1639 ();
 sg13g2_fill_1 FILLER_1_1646 ();
 sg13g2_fill_1 FILLER_1_1651 ();
 sg13g2_decap_8 FILLER_1_1656 ();
 sg13g2_decap_4 FILLER_1_1663 ();
 sg13g2_fill_2 FILLER_1_1672 ();
 sg13g2_fill_1 FILLER_1_1705 ();
 sg13g2_decap_8 FILLER_1_1710 ();
 sg13g2_decap_8 FILLER_1_1717 ();
 sg13g2_decap_8 FILLER_1_1724 ();
 sg13g2_decap_8 FILLER_1_1731 ();
 sg13g2_decap_8 FILLER_1_1738 ();
 sg13g2_decap_8 FILLER_1_1745 ();
 sg13g2_decap_8 FILLER_1_1752 ();
 sg13g2_decap_8 FILLER_1_1759 ();
 sg13g2_decap_8 FILLER_1_1766 ();
 sg13g2_fill_1 FILLER_1_1773 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_7 ();
 sg13g2_fill_2 FILLER_2_11 ();
 sg13g2_fill_1 FILLER_2_18 ();
 sg13g2_fill_1 FILLER_2_29 ();
 sg13g2_fill_2 FILLER_2_40 ();
 sg13g2_fill_2 FILLER_2_57 ();
 sg13g2_fill_1 FILLER_2_59 ();
 sg13g2_fill_2 FILLER_2_64 ();
 sg13g2_decap_4 FILLER_2_74 ();
 sg13g2_fill_2 FILLER_2_78 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_101 ();
 sg13g2_fill_2 FILLER_2_108 ();
 sg13g2_fill_1 FILLER_2_110 ();
 sg13g2_decap_8 FILLER_2_120 ();
 sg13g2_fill_2 FILLER_2_132 ();
 sg13g2_decap_8 FILLER_2_139 ();
 sg13g2_fill_2 FILLER_2_146 ();
 sg13g2_fill_1 FILLER_2_148 ();
 sg13g2_fill_1 FILLER_2_180 ();
 sg13g2_fill_2 FILLER_2_248 ();
 sg13g2_fill_1 FILLER_2_285 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_decap_4 FILLER_2_297 ();
 sg13g2_fill_2 FILLER_2_305 ();
 sg13g2_fill_2 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_450 ();
 sg13g2_fill_1 FILLER_2_465 ();
 sg13g2_fill_2 FILLER_2_471 ();
 sg13g2_fill_2 FILLER_2_504 ();
 sg13g2_fill_2 FILLER_2_531 ();
 sg13g2_fill_1 FILLER_2_533 ();
 sg13g2_fill_2 FILLER_2_570 ();
 sg13g2_fill_1 FILLER_2_572 ();
 sg13g2_fill_2 FILLER_2_582 ();
 sg13g2_fill_1 FILLER_2_584 ();
 sg13g2_fill_2 FILLER_2_608 ();
 sg13g2_fill_2 FILLER_2_644 ();
 sg13g2_fill_1 FILLER_2_694 ();
 sg13g2_fill_2 FILLER_2_699 ();
 sg13g2_fill_1 FILLER_2_701 ();
 sg13g2_fill_1 FILLER_2_706 ();
 sg13g2_fill_2 FILLER_2_793 ();
 sg13g2_decap_4 FILLER_2_812 ();
 sg13g2_fill_2 FILLER_2_816 ();
 sg13g2_fill_2 FILLER_2_867 ();
 sg13g2_fill_1 FILLER_2_891 ();
 sg13g2_fill_2 FILLER_2_900 ();
 sg13g2_fill_2 FILLER_2_906 ();
 sg13g2_fill_1 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_940 ();
 sg13g2_decap_8 FILLER_2_947 ();
 sg13g2_decap_8 FILLER_2_954 ();
 sg13g2_decap_8 FILLER_2_961 ();
 sg13g2_fill_1 FILLER_2_968 ();
 sg13g2_decap_8 FILLER_2_973 ();
 sg13g2_fill_1 FILLER_2_980 ();
 sg13g2_decap_4 FILLER_2_991 ();
 sg13g2_fill_1 FILLER_2_995 ();
 sg13g2_fill_2 FILLER_2_1000 ();
 sg13g2_fill_2 FILLER_2_1007 ();
 sg13g2_fill_2 FILLER_2_1016 ();
 sg13g2_fill_1 FILLER_2_1018 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_fill_1 FILLER_2_1033 ();
 sg13g2_fill_1 FILLER_2_1038 ();
 sg13g2_fill_2 FILLER_2_1052 ();
 sg13g2_fill_2 FILLER_2_1061 ();
 sg13g2_fill_1 FILLER_2_1063 ();
 sg13g2_decap_8 FILLER_2_1079 ();
 sg13g2_fill_2 FILLER_2_1086 ();
 sg13g2_fill_1 FILLER_2_1088 ();
 sg13g2_decap_4 FILLER_2_1093 ();
 sg13g2_fill_1 FILLER_2_1097 ();
 sg13g2_fill_2 FILLER_2_1118 ();
 sg13g2_decap_8 FILLER_2_1128 ();
 sg13g2_decap_8 FILLER_2_1135 ();
 sg13g2_fill_2 FILLER_2_1151 ();
 sg13g2_fill_1 FILLER_2_1153 ();
 sg13g2_decap_8 FILLER_2_1158 ();
 sg13g2_fill_2 FILLER_2_1178 ();
 sg13g2_fill_2 FILLER_2_1193 ();
 sg13g2_fill_1 FILLER_2_1195 ();
 sg13g2_fill_2 FILLER_2_1209 ();
 sg13g2_fill_1 FILLER_2_1211 ();
 sg13g2_fill_2 FILLER_2_1225 ();
 sg13g2_decap_4 FILLER_2_1237 ();
 sg13g2_fill_2 FILLER_2_1278 ();
 sg13g2_fill_1 FILLER_2_1302 ();
 sg13g2_fill_1 FILLER_2_1308 ();
 sg13g2_fill_2 FILLER_2_1313 ();
 sg13g2_fill_1 FILLER_2_1320 ();
 sg13g2_fill_1 FILLER_2_1326 ();
 sg13g2_fill_1 FILLER_2_1334 ();
 sg13g2_fill_2 FILLER_2_1353 ();
 sg13g2_fill_1 FILLER_2_1355 ();
 sg13g2_fill_1 FILLER_2_1364 ();
 sg13g2_fill_2 FILLER_2_1387 ();
 sg13g2_fill_2 FILLER_2_1398 ();
 sg13g2_fill_2 FILLER_2_1420 ();
 sg13g2_decap_8 FILLER_2_1449 ();
 sg13g2_fill_2 FILLER_2_1461 ();
 sg13g2_fill_2 FILLER_2_1476 ();
 sg13g2_decap_4 FILLER_2_1482 ();
 sg13g2_fill_2 FILLER_2_1491 ();
 sg13g2_fill_2 FILLER_2_1497 ();
 sg13g2_fill_1 FILLER_2_1499 ();
 sg13g2_fill_1 FILLER_2_1505 ();
 sg13g2_fill_1 FILLER_2_1510 ();
 sg13g2_fill_1 FILLER_2_1517 ();
 sg13g2_fill_2 FILLER_2_1522 ();
 sg13g2_fill_2 FILLER_2_1531 ();
 sg13g2_fill_2 FILLER_2_1538 ();
 sg13g2_fill_1 FILLER_2_1540 ();
 sg13g2_fill_2 FILLER_2_1545 ();
 sg13g2_fill_1 FILLER_2_1551 ();
 sg13g2_fill_1 FILLER_2_1557 ();
 sg13g2_fill_1 FILLER_2_1563 ();
 sg13g2_decap_8 FILLER_2_1573 ();
 sg13g2_fill_1 FILLER_2_1580 ();
 sg13g2_fill_2 FILLER_2_1586 ();
 sg13g2_fill_1 FILLER_2_1588 ();
 sg13g2_fill_2 FILLER_2_1633 ();
 sg13g2_decap_8 FILLER_2_1653 ();
 sg13g2_decap_4 FILLER_2_1660 ();
 sg13g2_fill_1 FILLER_2_1680 ();
 sg13g2_fill_1 FILLER_2_1686 ();
 sg13g2_fill_1 FILLER_2_1696 ();
 sg13g2_fill_2 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1713 ();
 sg13g2_decap_8 FILLER_2_1720 ();
 sg13g2_decap_8 FILLER_2_1727 ();
 sg13g2_decap_8 FILLER_2_1734 ();
 sg13g2_decap_8 FILLER_2_1741 ();
 sg13g2_decap_8 FILLER_2_1748 ();
 sg13g2_decap_8 FILLER_2_1755 ();
 sg13g2_decap_8 FILLER_2_1762 ();
 sg13g2_decap_4 FILLER_2_1769 ();
 sg13g2_fill_1 FILLER_2_1773 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_219 ();
 sg13g2_fill_2 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_237 ();
 sg13g2_decap_4 FILLER_3_244 ();
 sg13g2_decap_4 FILLER_3_279 ();
 sg13g2_fill_2 FILLER_3_283 ();
 sg13g2_fill_2 FILLER_3_350 ();
 sg13g2_fill_2 FILLER_3_405 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_1 FILLER_3_499 ();
 sg13g2_fill_1 FILLER_3_526 ();
 sg13g2_decap_4 FILLER_3_535 ();
 sg13g2_fill_2 FILLER_3_544 ();
 sg13g2_fill_1 FILLER_3_546 ();
 sg13g2_fill_2 FILLER_3_552 ();
 sg13g2_fill_1 FILLER_3_554 ();
 sg13g2_fill_1 FILLER_3_590 ();
 sg13g2_fill_2 FILLER_3_634 ();
 sg13g2_fill_2 FILLER_3_662 ();
 sg13g2_fill_2 FILLER_3_728 ();
 sg13g2_fill_1 FILLER_3_746 ();
 sg13g2_fill_1 FILLER_3_761 ();
 sg13g2_fill_1 FILLER_3_767 ();
 sg13g2_decap_4 FILLER_3_795 ();
 sg13g2_fill_1 FILLER_3_799 ();
 sg13g2_decap_4 FILLER_3_805 ();
 sg13g2_fill_1 FILLER_3_809 ();
 sg13g2_fill_1 FILLER_3_840 ();
 sg13g2_fill_2 FILLER_3_845 ();
 sg13g2_fill_2 FILLER_3_852 ();
 sg13g2_fill_2 FILLER_3_858 ();
 sg13g2_fill_1 FILLER_3_860 ();
 sg13g2_fill_1 FILLER_3_865 ();
 sg13g2_fill_1 FILLER_3_871 ();
 sg13g2_fill_1 FILLER_3_877 ();
 sg13g2_fill_1 FILLER_3_886 ();
 sg13g2_fill_1 FILLER_3_895 ();
 sg13g2_fill_2 FILLER_3_900 ();
 sg13g2_decap_4 FILLER_3_907 ();
 sg13g2_fill_2 FILLER_3_942 ();
 sg13g2_fill_1 FILLER_3_944 ();
 sg13g2_decap_4 FILLER_3_949 ();
 sg13g2_decap_4 FILLER_3_958 ();
 sg13g2_fill_2 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1030 ();
 sg13g2_fill_1 FILLER_3_1042 ();
 sg13g2_fill_1 FILLER_3_1058 ();
 sg13g2_fill_1 FILLER_3_1085 ();
 sg13g2_fill_1 FILLER_3_1099 ();
 sg13g2_fill_1 FILLER_3_1124 ();
 sg13g2_fill_2 FILLER_3_1135 ();
 sg13g2_fill_1 FILLER_3_1154 ();
 sg13g2_decap_4 FILLER_3_1196 ();
 sg13g2_fill_1 FILLER_3_1200 ();
 sg13g2_decap_4 FILLER_3_1253 ();
 sg13g2_fill_1 FILLER_3_1257 ();
 sg13g2_fill_1 FILLER_3_1262 ();
 sg13g2_fill_1 FILLER_3_1267 ();
 sg13g2_fill_1 FILLER_3_1276 ();
 sg13g2_fill_2 FILLER_3_1281 ();
 sg13g2_fill_1 FILLER_3_1293 ();
 sg13g2_fill_1 FILLER_3_1306 ();
 sg13g2_fill_2 FILLER_3_1316 ();
 sg13g2_fill_2 FILLER_3_1323 ();
 sg13g2_decap_8 FILLER_3_1332 ();
 sg13g2_decap_8 FILLER_3_1339 ();
 sg13g2_fill_2 FILLER_3_1346 ();
 sg13g2_fill_1 FILLER_3_1348 ();
 sg13g2_fill_2 FILLER_3_1367 ();
 sg13g2_fill_1 FILLER_3_1369 ();
 sg13g2_decap_8 FILLER_3_1375 ();
 sg13g2_fill_2 FILLER_3_1382 ();
 sg13g2_decap_4 FILLER_3_1399 ();
 sg13g2_fill_1 FILLER_3_1403 ();
 sg13g2_fill_1 FILLER_3_1409 ();
 sg13g2_fill_1 FILLER_3_1415 ();
 sg13g2_fill_1 FILLER_3_1428 ();
 sg13g2_fill_1 FILLER_3_1434 ();
 sg13g2_fill_1 FILLER_3_1439 ();
 sg13g2_fill_1 FILLER_3_1447 ();
 sg13g2_fill_1 FILLER_3_1458 ();
 sg13g2_fill_1 FILLER_3_1464 ();
 sg13g2_fill_2 FILLER_3_1469 ();
 sg13g2_fill_1 FILLER_3_1484 ();
 sg13g2_fill_2 FILLER_3_1503 ();
 sg13g2_fill_1 FILLER_3_1509 ();
 sg13g2_fill_1 FILLER_3_1543 ();
 sg13g2_fill_2 FILLER_3_1554 ();
 sg13g2_fill_1 FILLER_3_1556 ();
 sg13g2_fill_1 FILLER_3_1562 ();
 sg13g2_fill_2 FILLER_3_1571 ();
 sg13g2_fill_1 FILLER_3_1573 ();
 sg13g2_fill_1 FILLER_3_1582 ();
 sg13g2_fill_1 FILLER_3_1587 ();
 sg13g2_fill_1 FILLER_3_1596 ();
 sg13g2_fill_1 FILLER_3_1601 ();
 sg13g2_fill_2 FILLER_3_1631 ();
 sg13g2_fill_2 FILLER_3_1638 ();
 sg13g2_fill_2 FILLER_3_1647 ();
 sg13g2_decap_8 FILLER_3_1657 ();
 sg13g2_fill_2 FILLER_3_1664 ();
 sg13g2_fill_2 FILLER_3_1705 ();
 sg13g2_decap_8 FILLER_3_1716 ();
 sg13g2_decap_8 FILLER_3_1723 ();
 sg13g2_decap_8 FILLER_3_1730 ();
 sg13g2_decap_8 FILLER_3_1737 ();
 sg13g2_decap_8 FILLER_3_1744 ();
 sg13g2_decap_8 FILLER_3_1751 ();
 sg13g2_decap_8 FILLER_3_1758 ();
 sg13g2_decap_8 FILLER_3_1765 ();
 sg13g2_fill_2 FILLER_3_1772 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_2 FILLER_4_5 ();
 sg13g2_fill_1 FILLER_4_7 ();
 sg13g2_fill_1 FILLER_4_45 ();
 sg13g2_fill_1 FILLER_4_76 ();
 sg13g2_fill_2 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_fill_1 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_fill_2 FILLER_4_171 ();
 sg13g2_decap_8 FILLER_4_190 ();
 sg13g2_decap_4 FILLER_4_197 ();
 sg13g2_decap_4 FILLER_4_205 ();
 sg13g2_fill_1 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_257 ();
 sg13g2_fill_1 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_275 ();
 sg13g2_fill_1 FILLER_4_311 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_fill_1 FILLER_4_322 ();
 sg13g2_fill_1 FILLER_4_327 ();
 sg13g2_fill_1 FILLER_4_332 ();
 sg13g2_fill_1 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_364 ();
 sg13g2_fill_1 FILLER_4_370 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_1 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_440 ();
 sg13g2_fill_1 FILLER_4_442 ();
 sg13g2_fill_2 FILLER_4_451 ();
 sg13g2_fill_2 FILLER_4_458 ();
 sg13g2_fill_1 FILLER_4_460 ();
 sg13g2_fill_2 FILLER_4_466 ();
 sg13g2_fill_2 FILLER_4_472 ();
 sg13g2_fill_1 FILLER_4_474 ();
 sg13g2_fill_2 FILLER_4_515 ();
 sg13g2_fill_2 FILLER_4_614 ();
 sg13g2_fill_1 FILLER_4_616 ();
 sg13g2_fill_2 FILLER_4_683 ();
 sg13g2_fill_2 FILLER_4_689 ();
 sg13g2_fill_1 FILLER_4_696 ();
 sg13g2_fill_2 FILLER_4_706 ();
 sg13g2_fill_2 FILLER_4_712 ();
 sg13g2_fill_1 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_fill_1 FILLER_4_734 ();
 sg13g2_fill_2 FILLER_4_740 ();
 sg13g2_fill_2 FILLER_4_746 ();
 sg13g2_fill_1 FILLER_4_752 ();
 sg13g2_fill_2 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_813 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_fill_2 FILLER_4_864 ();
 sg13g2_fill_1 FILLER_4_915 ();
 sg13g2_decap_8 FILLER_4_985 ();
 sg13g2_fill_2 FILLER_4_992 ();
 sg13g2_fill_2 FILLER_4_999 ();
 sg13g2_fill_1 FILLER_4_1001 ();
 sg13g2_fill_1 FILLER_4_1014 ();
 sg13g2_fill_2 FILLER_4_1027 ();
 sg13g2_fill_1 FILLER_4_1034 ();
 sg13g2_fill_2 FILLER_4_1039 ();
 sg13g2_fill_2 FILLER_4_1054 ();
 sg13g2_fill_1 FILLER_4_1064 ();
 sg13g2_fill_2 FILLER_4_1070 ();
 sg13g2_fill_1 FILLER_4_1072 ();
 sg13g2_fill_2 FILLER_4_1085 ();
 sg13g2_fill_1 FILLER_4_1092 ();
 sg13g2_fill_2 FILLER_4_1117 ();
 sg13g2_fill_1 FILLER_4_1119 ();
 sg13g2_decap_8 FILLER_4_1125 ();
 sg13g2_fill_1 FILLER_4_1132 ();
 sg13g2_fill_2 FILLER_4_1137 ();
 sg13g2_decap_4 FILLER_4_1147 ();
 sg13g2_decap_4 FILLER_4_1161 ();
 sg13g2_fill_2 FILLER_4_1175 ();
 sg13g2_fill_1 FILLER_4_1177 ();
 sg13g2_fill_2 FILLER_4_1214 ();
 sg13g2_decap_8 FILLER_4_1220 ();
 sg13g2_fill_2 FILLER_4_1227 ();
 sg13g2_decap_4 FILLER_4_1233 ();
 sg13g2_decap_4 FILLER_4_1247 ();
 sg13g2_fill_1 FILLER_4_1251 ();
 sg13g2_fill_2 FILLER_4_1257 ();
 sg13g2_decap_8 FILLER_4_1268 ();
 sg13g2_fill_2 FILLER_4_1275 ();
 sg13g2_fill_1 FILLER_4_1277 ();
 sg13g2_decap_4 FILLER_4_1283 ();
 sg13g2_fill_2 FILLER_4_1287 ();
 sg13g2_fill_1 FILLER_4_1293 ();
 sg13g2_fill_2 FILLER_4_1298 ();
 sg13g2_fill_1 FILLER_4_1305 ();
 sg13g2_fill_1 FILLER_4_1311 ();
 sg13g2_fill_1 FILLER_4_1324 ();
 sg13g2_fill_2 FILLER_4_1329 ();
 sg13g2_fill_2 FILLER_4_1344 ();
 sg13g2_fill_1 FILLER_4_1346 ();
 sg13g2_fill_2 FILLER_4_1351 ();
 sg13g2_fill_1 FILLER_4_1353 ();
 sg13g2_fill_2 FILLER_4_1359 ();
 sg13g2_fill_2 FILLER_4_1412 ();
 sg13g2_fill_1 FILLER_4_1428 ();
 sg13g2_fill_1 FILLER_4_1434 ();
 sg13g2_fill_1 FILLER_4_1444 ();
 sg13g2_decap_8 FILLER_4_1449 ();
 sg13g2_fill_2 FILLER_4_1456 ();
 sg13g2_fill_2 FILLER_4_1462 ();
 sg13g2_fill_1 FILLER_4_1464 ();
 sg13g2_fill_2 FILLER_4_1493 ();
 sg13g2_fill_2 FILLER_4_1500 ();
 sg13g2_fill_2 FILLER_4_1507 ();
 sg13g2_fill_2 FILLER_4_1517 ();
 sg13g2_fill_1 FILLER_4_1519 ();
 sg13g2_fill_1 FILLER_4_1550 ();
 sg13g2_fill_2 FILLER_4_1555 ();
 sg13g2_fill_2 FILLER_4_1562 ();
 sg13g2_fill_2 FILLER_4_1568 ();
 sg13g2_fill_1 FILLER_4_1578 ();
 sg13g2_fill_1 FILLER_4_1589 ();
 sg13g2_fill_1 FILLER_4_1598 ();
 sg13g2_fill_1 FILLER_4_1615 ();
 sg13g2_fill_1 FILLER_4_1621 ();
 sg13g2_decap_8 FILLER_4_1643 ();
 sg13g2_decap_4 FILLER_4_1663 ();
 sg13g2_fill_1 FILLER_4_1698 ();
 sg13g2_decap_8 FILLER_4_1732 ();
 sg13g2_decap_8 FILLER_4_1739 ();
 sg13g2_decap_8 FILLER_4_1746 ();
 sg13g2_decap_8 FILLER_4_1753 ();
 sg13g2_decap_8 FILLER_4_1760 ();
 sg13g2_decap_8 FILLER_4_1767 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_31 ();
 sg13g2_fill_2 FILLER_5_67 ();
 sg13g2_fill_1 FILLER_5_82 ();
 sg13g2_fill_2 FILLER_5_127 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_2 FILLER_5_165 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_294 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_4 FILLER_5_347 ();
 sg13g2_fill_2 FILLER_5_351 ();
 sg13g2_fill_2 FILLER_5_424 ();
 sg13g2_fill_1 FILLER_5_426 ();
 sg13g2_fill_1 FILLER_5_445 ();
 sg13g2_fill_2 FILLER_5_450 ();
 sg13g2_fill_1 FILLER_5_473 ();
 sg13g2_fill_2 FILLER_5_478 ();
 sg13g2_fill_1 FILLER_5_484 ();
 sg13g2_fill_2 FILLER_5_490 ();
 sg13g2_decap_4 FILLER_5_500 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_2 FILLER_5_558 ();
 sg13g2_fill_1 FILLER_5_565 ();
 sg13g2_fill_1 FILLER_5_574 ();
 sg13g2_fill_2 FILLER_5_606 ();
 sg13g2_fill_1 FILLER_5_608 ();
 sg13g2_fill_1 FILLER_5_626 ();
 sg13g2_fill_1 FILLER_5_631 ();
 sg13g2_fill_2 FILLER_5_645 ();
 sg13g2_fill_2 FILLER_5_659 ();
 sg13g2_fill_1 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_696 ();
 sg13g2_fill_2 FILLER_5_701 ();
 sg13g2_fill_1 FILLER_5_707 ();
 sg13g2_fill_2 FILLER_5_712 ();
 sg13g2_fill_1 FILLER_5_768 ();
 sg13g2_fill_2 FILLER_5_773 ();
 sg13g2_fill_1 FILLER_5_780 ();
 sg13g2_fill_2 FILLER_5_786 ();
 sg13g2_fill_1 FILLER_5_803 ();
 sg13g2_fill_1 FILLER_5_812 ();
 sg13g2_fill_1 FILLER_5_821 ();
 sg13g2_fill_2 FILLER_5_826 ();
 sg13g2_fill_1 FILLER_5_849 ();
 sg13g2_fill_1 FILLER_5_860 ();
 sg13g2_fill_1 FILLER_5_866 ();
 sg13g2_fill_1 FILLER_5_872 ();
 sg13g2_fill_1 FILLER_5_878 ();
 sg13g2_fill_1 FILLER_5_887 ();
 sg13g2_fill_1 FILLER_5_893 ();
 sg13g2_fill_1 FILLER_5_897 ();
 sg13g2_fill_2 FILLER_5_906 ();
 sg13g2_fill_1 FILLER_5_908 ();
 sg13g2_fill_1 FILLER_5_914 ();
 sg13g2_fill_2 FILLER_5_963 ();
 sg13g2_fill_1 FILLER_5_965 ();
 sg13g2_fill_1 FILLER_5_970 ();
 sg13g2_fill_2 FILLER_5_979 ();
 sg13g2_fill_2 FILLER_5_987 ();
 sg13g2_fill_1 FILLER_5_993 ();
 sg13g2_fill_1 FILLER_5_1000 ();
 sg13g2_fill_1 FILLER_5_1006 ();
 sg13g2_fill_1 FILLER_5_1023 ();
 sg13g2_fill_1 FILLER_5_1032 ();
 sg13g2_fill_2 FILLER_5_1041 ();
 sg13g2_fill_2 FILLER_5_1063 ();
 sg13g2_fill_1 FILLER_5_1070 ();
 sg13g2_fill_1 FILLER_5_1104 ();
 sg13g2_fill_2 FILLER_5_1124 ();
 sg13g2_fill_2 FILLER_5_1130 ();
 sg13g2_fill_1 FILLER_5_1132 ();
 sg13g2_fill_2 FILLER_5_1137 ();
 sg13g2_fill_1 FILLER_5_1139 ();
 sg13g2_fill_2 FILLER_5_1144 ();
 sg13g2_fill_1 FILLER_5_1167 ();
 sg13g2_fill_1 FILLER_5_1189 ();
 sg13g2_fill_1 FILLER_5_1194 ();
 sg13g2_fill_2 FILLER_5_1202 ();
 sg13g2_fill_1 FILLER_5_1209 ();
 sg13g2_fill_1 FILLER_5_1227 ();
 sg13g2_fill_2 FILLER_5_1260 ();
 sg13g2_fill_2 FILLER_5_1293 ();
 sg13g2_fill_1 FILLER_5_1335 ();
 sg13g2_fill_1 FILLER_5_1355 ();
 sg13g2_fill_1 FILLER_5_1376 ();
 sg13g2_fill_1 FILLER_5_1397 ();
 sg13g2_fill_1 FILLER_5_1402 ();
 sg13g2_fill_1 FILLER_5_1427 ();
 sg13g2_fill_2 FILLER_5_1433 ();
 sg13g2_fill_2 FILLER_5_1450 ();
 sg13g2_fill_1 FILLER_5_1469 ();
 sg13g2_fill_1 FILLER_5_1476 ();
 sg13g2_fill_1 FILLER_5_1488 ();
 sg13g2_fill_2 FILLER_5_1493 ();
 sg13g2_fill_2 FILLER_5_1504 ();
 sg13g2_decap_4 FILLER_5_1521 ();
 sg13g2_fill_1 FILLER_5_1539 ();
 sg13g2_fill_2 FILLER_5_1549 ();
 sg13g2_fill_2 FILLER_5_1558 ();
 sg13g2_decap_8 FILLER_5_1586 ();
 sg13g2_fill_2 FILLER_5_1593 ();
 sg13g2_fill_1 FILLER_5_1595 ();
 sg13g2_decap_8 FILLER_5_1600 ();
 sg13g2_decap_8 FILLER_5_1607 ();
 sg13g2_fill_2 FILLER_5_1614 ();
 sg13g2_fill_1 FILLER_5_1616 ();
 sg13g2_decap_8 FILLER_5_1621 ();
 sg13g2_fill_1 FILLER_5_1628 ();
 sg13g2_decap_4 FILLER_5_1641 ();
 sg13g2_fill_1 FILLER_5_1645 ();
 sg13g2_decap_4 FILLER_5_1660 ();
 sg13g2_fill_1 FILLER_5_1664 ();
 sg13g2_fill_1 FILLER_5_1670 ();
 sg13g2_decap_8 FILLER_5_1684 ();
 sg13g2_decap_8 FILLER_5_1691 ();
 sg13g2_fill_2 FILLER_5_1698 ();
 sg13g2_decap_4 FILLER_5_1717 ();
 sg13g2_decap_8 FILLER_5_1740 ();
 sg13g2_decap_8 FILLER_5_1747 ();
 sg13g2_decap_8 FILLER_5_1754 ();
 sg13g2_decap_8 FILLER_5_1761 ();
 sg13g2_decap_4 FILLER_5_1768 ();
 sg13g2_fill_2 FILLER_5_1772 ();
 sg13g2_fill_2 FILLER_6_51 ();
 sg13g2_fill_1 FILLER_6_53 ();
 sg13g2_fill_2 FILLER_6_89 ();
 sg13g2_fill_2 FILLER_6_95 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_1 FILLER_6_213 ();
 sg13g2_fill_2 FILLER_6_254 ();
 sg13g2_fill_2 FILLER_6_309 ();
 sg13g2_fill_2 FILLER_6_336 ();
 sg13g2_fill_2 FILLER_6_343 ();
 sg13g2_fill_2 FILLER_6_349 ();
 sg13g2_fill_1 FILLER_6_351 ();
 sg13g2_decap_4 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_364 ();
 sg13g2_fill_2 FILLER_6_436 ();
 sg13g2_fill_1 FILLER_6_455 ();
 sg13g2_fill_2 FILLER_6_482 ();
 sg13g2_fill_2 FILLER_6_515 ();
 sg13g2_fill_2 FILLER_6_569 ();
 sg13g2_fill_1 FILLER_6_580 ();
 sg13g2_fill_2 FILLER_6_586 ();
 sg13g2_fill_1 FILLER_6_619 ();
 sg13g2_fill_1 FILLER_6_651 ();
 sg13g2_fill_1 FILLER_6_670 ();
 sg13g2_fill_1 FILLER_6_692 ();
 sg13g2_fill_1 FILLER_6_701 ();
 sg13g2_decap_4 FILLER_6_737 ();
 sg13g2_fill_2 FILLER_6_741 ();
 sg13g2_fill_1 FILLER_6_752 ();
 sg13g2_fill_1 FILLER_6_756 ();
 sg13g2_fill_2 FILLER_6_762 ();
 sg13g2_fill_1 FILLER_6_769 ();
 sg13g2_fill_2 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_811 ();
 sg13g2_fill_1 FILLER_6_819 ();
 sg13g2_fill_1 FILLER_6_833 ();
 sg13g2_fill_2 FILLER_6_844 ();
 sg13g2_fill_2 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_856 ();
 sg13g2_fill_1 FILLER_6_868 ();
 sg13g2_fill_2 FILLER_6_903 ();
 sg13g2_fill_1 FILLER_6_905 ();
 sg13g2_decap_4 FILLER_6_914 ();
 sg13g2_fill_2 FILLER_6_918 ();
 sg13g2_fill_2 FILLER_6_927 ();
 sg13g2_fill_1 FILLER_6_929 ();
 sg13g2_fill_1 FILLER_6_972 ();
 sg13g2_fill_1 FILLER_6_977 ();
 sg13g2_fill_1 FILLER_6_982 ();
 sg13g2_fill_1 FILLER_6_1005 ();
 sg13g2_fill_2 FILLER_6_1023 ();
 sg13g2_fill_1 FILLER_6_1025 ();
 sg13g2_fill_2 FILLER_6_1040 ();
 sg13g2_fill_2 FILLER_6_1066 ();
 sg13g2_fill_1 FILLER_6_1068 ();
 sg13g2_fill_1 FILLER_6_1074 ();
 sg13g2_fill_1 FILLER_6_1079 ();
 sg13g2_fill_2 FILLER_6_1085 ();
 sg13g2_fill_1 FILLER_6_1087 ();
 sg13g2_fill_2 FILLER_6_1092 ();
 sg13g2_fill_1 FILLER_6_1094 ();
 sg13g2_decap_4 FILLER_6_1106 ();
 sg13g2_fill_1 FILLER_6_1110 ();
 sg13g2_fill_2 FILLER_6_1121 ();
 sg13g2_decap_8 FILLER_6_1143 ();
 sg13g2_decap_8 FILLER_6_1150 ();
 sg13g2_decap_4 FILLER_6_1157 ();
 sg13g2_fill_1 FILLER_6_1174 ();
 sg13g2_fill_1 FILLER_6_1204 ();
 sg13g2_fill_1 FILLER_6_1210 ();
 sg13g2_fill_1 FILLER_6_1215 ();
 sg13g2_fill_1 FILLER_6_1221 ();
 sg13g2_fill_1 FILLER_6_1236 ();
 sg13g2_fill_1 FILLER_6_1253 ();
 sg13g2_fill_2 FILLER_6_1262 ();
 sg13g2_decap_8 FILLER_6_1274 ();
 sg13g2_decap_4 FILLER_6_1285 ();
 sg13g2_fill_2 FILLER_6_1289 ();
 sg13g2_decap_8 FILLER_6_1295 ();
 sg13g2_fill_2 FILLER_6_1302 ();
 sg13g2_decap_8 FILLER_6_1312 ();
 sg13g2_decap_8 FILLER_6_1319 ();
 sg13g2_fill_2 FILLER_6_1335 ();
 sg13g2_fill_1 FILLER_6_1337 ();
 sg13g2_fill_1 FILLER_6_1352 ();
 sg13g2_fill_1 FILLER_6_1360 ();
 sg13g2_fill_1 FILLER_6_1382 ();
 sg13g2_fill_2 FILLER_6_1400 ();
 sg13g2_fill_2 FILLER_6_1418 ();
 sg13g2_fill_1 FILLER_6_1420 ();
 sg13g2_fill_1 FILLER_6_1448 ();
 sg13g2_fill_2 FILLER_6_1454 ();
 sg13g2_fill_2 FILLER_6_1514 ();
 sg13g2_fill_1 FILLER_6_1521 ();
 sg13g2_fill_1 FILLER_6_1527 ();
 sg13g2_fill_2 FILLER_6_1540 ();
 sg13g2_fill_1 FILLER_6_1542 ();
 sg13g2_fill_2 FILLER_6_1567 ();
 sg13g2_fill_2 FILLER_6_1573 ();
 sg13g2_fill_1 FILLER_6_1575 ();
 sg13g2_decap_8 FILLER_6_1583 ();
 sg13g2_fill_1 FILLER_6_1594 ();
 sg13g2_fill_1 FILLER_6_1603 ();
 sg13g2_decap_8 FILLER_6_1612 ();
 sg13g2_fill_1 FILLER_6_1619 ();
 sg13g2_decap_4 FILLER_6_1639 ();
 sg13g2_fill_1 FILLER_6_1659 ();
 sg13g2_fill_1 FILLER_6_1677 ();
 sg13g2_fill_2 FILLER_6_1682 ();
 sg13g2_fill_1 FILLER_6_1692 ();
 sg13g2_fill_1 FILLER_6_1714 ();
 sg13g2_fill_1 FILLER_6_1733 ();
 sg13g2_decap_8 FILLER_6_1739 ();
 sg13g2_decap_8 FILLER_6_1759 ();
 sg13g2_decap_8 FILLER_6_1766 ();
 sg13g2_fill_1 FILLER_6_1773 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_2 ();
 sg13g2_fill_1 FILLER_7_33 ();
 sg13g2_fill_2 FILLER_7_39 ();
 sg13g2_fill_2 FILLER_7_55 ();
 sg13g2_fill_1 FILLER_7_57 ();
 sg13g2_fill_2 FILLER_7_62 ();
 sg13g2_fill_1 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_236 ();
 sg13g2_fill_1 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_289 ();
 sg13g2_decap_4 FILLER_7_316 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_fill_2 FILLER_7_339 ();
 sg13g2_fill_1 FILLER_7_351 ();
 sg13g2_decap_4 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_366 ();
 sg13g2_fill_1 FILLER_7_372 ();
 sg13g2_fill_1 FILLER_7_421 ();
 sg13g2_fill_1 FILLER_7_448 ();
 sg13g2_fill_1 FILLER_7_462 ();
 sg13g2_fill_1 FILLER_7_489 ();
 sg13g2_fill_2 FILLER_7_500 ();
 sg13g2_fill_1 FILLER_7_502 ();
 sg13g2_fill_2 FILLER_7_507 ();
 sg13g2_fill_2 FILLER_7_540 ();
 sg13g2_fill_1 FILLER_7_547 ();
 sg13g2_fill_2 FILLER_7_575 ();
 sg13g2_fill_1 FILLER_7_577 ();
 sg13g2_fill_2 FILLER_7_610 ();
 sg13g2_fill_1 FILLER_7_625 ();
 sg13g2_fill_2 FILLER_7_630 ();
 sg13g2_fill_1 FILLER_7_636 ();
 sg13g2_fill_1 FILLER_7_653 ();
 sg13g2_fill_2 FILLER_7_715 ();
 sg13g2_fill_1 FILLER_7_717 ();
 sg13g2_fill_1 FILLER_7_723 ();
 sg13g2_fill_2 FILLER_7_762 ();
 sg13g2_fill_1 FILLER_7_764 ();
 sg13g2_decap_8 FILLER_7_832 ();
 sg13g2_decap_4 FILLER_7_847 ();
 sg13g2_fill_2 FILLER_7_851 ();
 sg13g2_fill_2 FILLER_7_858 ();
 sg13g2_fill_1 FILLER_7_860 ();
 sg13g2_fill_2 FILLER_7_886 ();
 sg13g2_fill_2 FILLER_7_893 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_fill_1 FILLER_7_980 ();
 sg13g2_fill_1 FILLER_7_1005 ();
 sg13g2_fill_2 FILLER_7_1019 ();
 sg13g2_fill_2 FILLER_7_1026 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_fill_2 FILLER_7_1046 ();
 sg13g2_fill_2 FILLER_7_1059 ();
 sg13g2_fill_2 FILLER_7_1069 ();
 sg13g2_fill_1 FILLER_7_1071 ();
 sg13g2_fill_2 FILLER_7_1102 ();
 sg13g2_fill_1 FILLER_7_1114 ();
 sg13g2_decap_8 FILLER_7_1128 ();
 sg13g2_fill_1 FILLER_7_1135 ();
 sg13g2_decap_4 FILLER_7_1141 ();
 sg13g2_fill_2 FILLER_7_1145 ();
 sg13g2_fill_1 FILLER_7_1159 ();
 sg13g2_fill_2 FILLER_7_1201 ();
 sg13g2_fill_1 FILLER_7_1250 ();
 sg13g2_decap_8 FILLER_7_1264 ();
 sg13g2_decap_8 FILLER_7_1271 ();
 sg13g2_fill_1 FILLER_7_1301 ();
 sg13g2_fill_2 FILLER_7_1307 ();
 sg13g2_decap_8 FILLER_7_1317 ();
 sg13g2_decap_4 FILLER_7_1324 ();
 sg13g2_fill_2 FILLER_7_1336 ();
 sg13g2_fill_1 FILLER_7_1338 ();
 sg13g2_fill_1 FILLER_7_1344 ();
 sg13g2_fill_1 FILLER_7_1350 ();
 sg13g2_fill_1 FILLER_7_1376 ();
 sg13g2_fill_2 FILLER_7_1383 ();
 sg13g2_fill_1 FILLER_7_1390 ();
 sg13g2_fill_2 FILLER_7_1396 ();
 sg13g2_fill_2 FILLER_7_1416 ();
 sg13g2_fill_1 FILLER_7_1422 ();
 sg13g2_fill_2 FILLER_7_1431 ();
 sg13g2_fill_1 FILLER_7_1437 ();
 sg13g2_fill_1 FILLER_7_1443 ();
 sg13g2_fill_1 FILLER_7_1454 ();
 sg13g2_fill_2 FILLER_7_1461 ();
 sg13g2_fill_1 FILLER_7_1463 ();
 sg13g2_decap_4 FILLER_7_1513 ();
 sg13g2_decap_4 FILLER_7_1563 ();
 sg13g2_fill_1 FILLER_7_1575 ();
 sg13g2_fill_2 FILLER_7_1596 ();
 sg13g2_fill_1 FILLER_7_1608 ();
 sg13g2_fill_1 FILLER_7_1614 ();
 sg13g2_fill_1 FILLER_7_1620 ();
 sg13g2_fill_2 FILLER_7_1626 ();
 sg13g2_fill_2 FILLER_7_1650 ();
 sg13g2_fill_1 FILLER_7_1657 ();
 sg13g2_fill_1 FILLER_7_1665 ();
 sg13g2_fill_2 FILLER_7_1671 ();
 sg13g2_fill_2 FILLER_7_1681 ();
 sg13g2_fill_1 FILLER_7_1683 ();
 sg13g2_fill_1 FILLER_7_1689 ();
 sg13g2_fill_2 FILLER_7_1722 ();
 sg13g2_fill_1 FILLER_7_1724 ();
 sg13g2_fill_2 FILLER_7_1729 ();
 sg13g2_fill_1 FILLER_7_1731 ();
 sg13g2_fill_1 FILLER_7_1740 ();
 sg13g2_fill_2 FILLER_7_1763 ();
 sg13g2_fill_2 FILLER_7_1771 ();
 sg13g2_fill_1 FILLER_7_1773 ();
 sg13g2_fill_2 FILLER_8_5 ();
 sg13g2_fill_1 FILLER_8_11 ();
 sg13g2_fill_1 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_132 ();
 sg13g2_fill_2 FILLER_8_141 ();
 sg13g2_fill_1 FILLER_8_169 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_decap_4 FILLER_8_227 ();
 sg13g2_fill_1 FILLER_8_231 ();
 sg13g2_fill_2 FILLER_8_271 ();
 sg13g2_fill_1 FILLER_8_303 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_1 FILLER_8_402 ();
 sg13g2_fill_2 FILLER_8_412 ();
 sg13g2_fill_2 FILLER_8_423 ();
 sg13g2_fill_1 FILLER_8_437 ();
 sg13g2_fill_1 FILLER_8_453 ();
 sg13g2_fill_2 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_478 ();
 sg13g2_fill_1 FILLER_8_485 ();
 sg13g2_fill_2 FILLER_8_552 ();
 sg13g2_fill_1 FILLER_8_559 ();
 sg13g2_fill_2 FILLER_8_612 ();
 sg13g2_fill_1 FILLER_8_614 ();
 sg13g2_fill_1 FILLER_8_628 ();
 sg13g2_fill_1 FILLER_8_655 ();
 sg13g2_fill_2 FILLER_8_661 ();
 sg13g2_fill_1 FILLER_8_663 ();
 sg13g2_fill_2 FILLER_8_690 ();
 sg13g2_fill_2 FILLER_8_727 ();
 sg13g2_decap_4 FILLER_8_741 ();
 sg13g2_fill_2 FILLER_8_745 ();
 sg13g2_decap_8 FILLER_8_751 ();
 sg13g2_fill_2 FILLER_8_758 ();
 sg13g2_fill_1 FILLER_8_760 ();
 sg13g2_decap_4 FILLER_8_773 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_fill_2 FILLER_8_788 ();
 sg13g2_fill_1 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_800 ();
 sg13g2_fill_2 FILLER_8_813 ();
 sg13g2_fill_2 FILLER_8_823 ();
 sg13g2_fill_2 FILLER_8_830 ();
 sg13g2_fill_1 FILLER_8_872 ();
 sg13g2_fill_1 FILLER_8_881 ();
 sg13g2_fill_1 FILLER_8_896 ();
 sg13g2_fill_1 FILLER_8_901 ();
 sg13g2_fill_1 FILLER_8_910 ();
 sg13g2_fill_2 FILLER_8_915 ();
 sg13g2_fill_2 FILLER_8_961 ();
 sg13g2_decap_8 FILLER_8_968 ();
 sg13g2_decap_8 FILLER_8_975 ();
 sg13g2_fill_1 FILLER_8_994 ();
 sg13g2_decap_4 FILLER_8_1005 ();
 sg13g2_fill_2 FILLER_8_1013 ();
 sg13g2_fill_1 FILLER_8_1023 ();
 sg13g2_fill_1 FILLER_8_1032 ();
 sg13g2_fill_1 FILLER_8_1046 ();
 sg13g2_fill_1 FILLER_8_1061 ();
 sg13g2_fill_1 FILLER_8_1072 ();
 sg13g2_fill_2 FILLER_8_1083 ();
 sg13g2_decap_4 FILLER_8_1089 ();
 sg13g2_fill_1 FILLER_8_1110 ();
 sg13g2_fill_2 FILLER_8_1116 ();
 sg13g2_fill_2 FILLER_8_1126 ();
 sg13g2_fill_2 FILLER_8_1136 ();
 sg13g2_fill_1 FILLER_8_1138 ();
 sg13g2_fill_2 FILLER_8_1144 ();
 sg13g2_decap_4 FILLER_8_1155 ();
 sg13g2_fill_2 FILLER_8_1180 ();
 sg13g2_fill_1 FILLER_8_1182 ();
 sg13g2_fill_2 FILLER_8_1204 ();
 sg13g2_fill_1 FILLER_8_1242 ();
 sg13g2_fill_2 FILLER_8_1262 ();
 sg13g2_fill_1 FILLER_8_1280 ();
 sg13g2_fill_1 FILLER_8_1313 ();
 sg13g2_fill_1 FILLER_8_1327 ();
 sg13g2_fill_1 FILLER_8_1332 ();
 sg13g2_fill_1 FILLER_8_1363 ();
 sg13g2_fill_1 FILLER_8_1369 ();
 sg13g2_fill_1 FILLER_8_1388 ();
 sg13g2_fill_1 FILLER_8_1393 ();
 sg13g2_decap_8 FILLER_8_1412 ();
 sg13g2_decap_4 FILLER_8_1419 ();
 sg13g2_fill_1 FILLER_8_1423 ();
 sg13g2_decap_4 FILLER_8_1429 ();
 sg13g2_fill_1 FILLER_8_1468 ();
 sg13g2_fill_1 FILLER_8_1474 ();
 sg13g2_fill_1 FILLER_8_1480 ();
 sg13g2_fill_2 FILLER_8_1486 ();
 sg13g2_fill_2 FILLER_8_1492 ();
 sg13g2_fill_2 FILLER_8_1504 ();
 sg13g2_decap_8 FILLER_8_1526 ();
 sg13g2_fill_1 FILLER_8_1542 ();
 sg13g2_fill_1 FILLER_8_1547 ();
 sg13g2_fill_1 FILLER_8_1554 ();
 sg13g2_fill_1 FILLER_8_1567 ();
 sg13g2_fill_2 FILLER_8_1581 ();
 sg13g2_decap_8 FILLER_8_1592 ();
 sg13g2_fill_1 FILLER_8_1599 ();
 sg13g2_decap_8 FILLER_8_1604 ();
 sg13g2_fill_2 FILLER_8_1611 ();
 sg13g2_fill_1 FILLER_8_1613 ();
 sg13g2_decap_4 FILLER_8_1624 ();
 sg13g2_fill_2 FILLER_8_1628 ();
 sg13g2_fill_1 FILLER_8_1644 ();
 sg13g2_fill_1 FILLER_8_1658 ();
 sg13g2_fill_1 FILLER_8_1675 ();
 sg13g2_fill_2 FILLER_8_1689 ();
 sg13g2_fill_1 FILLER_8_1705 ();
 sg13g2_decap_8 FILLER_8_1717 ();
 sg13g2_decap_4 FILLER_8_1724 ();
 sg13g2_fill_2 FILLER_8_1728 ();
 sg13g2_fill_1 FILLER_8_1741 ();
 sg13g2_fill_1 FILLER_8_1747 ();
 sg13g2_fill_1 FILLER_8_1757 ();
 sg13g2_fill_2 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_34 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_2 FILLER_9_63 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_70 ();
 sg13g2_fill_1 FILLER_9_72 ();
 sg13g2_fill_1 FILLER_9_85 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_fill_2 FILLER_9_135 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_2 FILLER_9_143 ();
 sg13g2_fill_2 FILLER_9_149 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_decap_4 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_219 ();
 sg13g2_fill_1 FILLER_9_285 ();
 sg13g2_fill_2 FILLER_9_307 ();
 sg13g2_fill_2 FILLER_9_348 ();
 sg13g2_decap_4 FILLER_9_368 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_fill_1 FILLER_9_412 ();
 sg13g2_fill_2 FILLER_9_539 ();
 sg13g2_fill_2 FILLER_9_575 ();
 sg13g2_fill_1 FILLER_9_582 ();
 sg13g2_fill_2 FILLER_9_649 ();
 sg13g2_fill_2 FILLER_9_693 ();
 sg13g2_decap_4 FILLER_9_703 ();
 sg13g2_fill_1 FILLER_9_707 ();
 sg13g2_fill_2 FILLER_9_716 ();
 sg13g2_fill_1 FILLER_9_800 ();
 sg13g2_decap_4 FILLER_9_805 ();
 sg13g2_fill_1 FILLER_9_826 ();
 sg13g2_fill_1 FILLER_9_831 ();
 sg13g2_fill_1 FILLER_9_840 ();
 sg13g2_fill_1 FILLER_9_848 ();
 sg13g2_fill_2 FILLER_9_853 ();
 sg13g2_fill_2 FILLER_9_859 ();
 sg13g2_fill_2 FILLER_9_866 ();
 sg13g2_fill_1 FILLER_9_872 ();
 sg13g2_fill_2 FILLER_9_878 ();
 sg13g2_fill_1 FILLER_9_880 ();
 sg13g2_fill_1 FILLER_9_886 ();
 sg13g2_fill_2 FILLER_9_892 ();
 sg13g2_fill_1 FILLER_9_894 ();
 sg13g2_decap_4 FILLER_9_899 ();
 sg13g2_decap_4 FILLER_9_980 ();
 sg13g2_fill_1 FILLER_9_984 ();
 sg13g2_fill_2 FILLER_9_995 ();
 sg13g2_fill_2 FILLER_9_1002 ();
 sg13g2_fill_1 FILLER_9_1004 ();
 sg13g2_fill_2 FILLER_9_1010 ();
 sg13g2_fill_1 FILLER_9_1012 ();
 sg13g2_fill_2 FILLER_9_1029 ();
 sg13g2_fill_2 FILLER_9_1041 ();
 sg13g2_fill_1 FILLER_9_1053 ();
 sg13g2_fill_1 FILLER_9_1058 ();
 sg13g2_fill_1 FILLER_9_1095 ();
 sg13g2_decap_4 FILLER_9_1130 ();
 sg13g2_fill_2 FILLER_9_1140 ();
 sg13g2_decap_4 FILLER_9_1146 ();
 sg13g2_fill_1 FILLER_9_1150 ();
 sg13g2_fill_2 FILLER_9_1160 ();
 sg13g2_fill_1 FILLER_9_1167 ();
 sg13g2_fill_2 FILLER_9_1194 ();
 sg13g2_fill_2 FILLER_9_1202 ();
 sg13g2_fill_1 FILLER_9_1204 ();
 sg13g2_fill_2 FILLER_9_1210 ();
 sg13g2_fill_1 FILLER_9_1212 ();
 sg13g2_fill_2 FILLER_9_1219 ();
 sg13g2_decap_4 FILLER_9_1226 ();
 sg13g2_fill_2 FILLER_9_1248 ();
 sg13g2_decap_4 FILLER_9_1254 ();
 sg13g2_fill_1 FILLER_9_1262 ();
 sg13g2_decap_4 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1280 ();
 sg13g2_decap_4 FILLER_9_1287 ();
 sg13g2_fill_2 FILLER_9_1291 ();
 sg13g2_fill_2 FILLER_9_1297 ();
 sg13g2_fill_1 FILLER_9_1299 ();
 sg13g2_decap_4 FILLER_9_1311 ();
 sg13g2_decap_4 FILLER_9_1319 ();
 sg13g2_fill_1 FILLER_9_1345 ();
 sg13g2_fill_1 FILLER_9_1383 ();
 sg13g2_decap_4 FILLER_9_1392 ();
 sg13g2_fill_1 FILLER_9_1396 ();
 sg13g2_fill_2 FILLER_9_1402 ();
 sg13g2_fill_1 FILLER_9_1431 ();
 sg13g2_fill_2 FILLER_9_1437 ();
 sg13g2_fill_2 FILLER_9_1444 ();
 sg13g2_fill_1 FILLER_9_1446 ();
 sg13g2_fill_2 FILLER_9_1451 ();
 sg13g2_fill_1 FILLER_9_1453 ();
 sg13g2_fill_1 FILLER_9_1458 ();
 sg13g2_fill_2 FILLER_9_1475 ();
 sg13g2_fill_1 FILLER_9_1487 ();
 sg13g2_fill_2 FILLER_9_1506 ();
 sg13g2_fill_1 FILLER_9_1514 ();
 sg13g2_fill_1 FILLER_9_1522 ();
 sg13g2_fill_2 FILLER_9_1528 ();
 sg13g2_fill_1 FILLER_9_1541 ();
 sg13g2_fill_2 FILLER_9_1565 ();
 sg13g2_fill_1 FILLER_9_1567 ();
 sg13g2_decap_8 FILLER_9_1574 ();
 sg13g2_fill_2 FILLER_9_1581 ();
 sg13g2_fill_1 FILLER_9_1583 ();
 sg13g2_fill_1 FILLER_9_1593 ();
 sg13g2_fill_2 FILLER_9_1599 ();
 sg13g2_fill_1 FILLER_9_1606 ();
 sg13g2_fill_2 FILLER_9_1616 ();
 sg13g2_fill_1 FILLER_9_1618 ();
 sg13g2_decap_4 FILLER_9_1630 ();
 sg13g2_fill_1 FILLER_9_1634 ();
 sg13g2_decap_8 FILLER_9_1655 ();
 sg13g2_fill_2 FILLER_9_1662 ();
 sg13g2_fill_2 FILLER_9_1672 ();
 sg13g2_fill_2 FILLER_9_1682 ();
 sg13g2_fill_2 FILLER_9_1700 ();
 sg13g2_fill_1 FILLER_9_1714 ();
 sg13g2_fill_1 FILLER_9_1733 ();
 sg13g2_fill_2 FILLER_9_1746 ();
 sg13g2_decap_4 FILLER_9_1765 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_fill_2 FILLER_10_15 ();
 sg13g2_fill_1 FILLER_10_17 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_fill_1 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_216 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_235 ();
 sg13g2_fill_1 FILLER_10_237 ();
 sg13g2_decap_4 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_328 ();
 sg13g2_fill_1 FILLER_10_333 ();
 sg13g2_fill_2 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_344 ();
 sg13g2_fill_1 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_354 ();
 sg13g2_fill_2 FILLER_10_360 ();
 sg13g2_fill_2 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_407 ();
 sg13g2_fill_2 FILLER_10_413 ();
 sg13g2_fill_1 FILLER_10_415 ();
 sg13g2_fill_1 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_427 ();
 sg13g2_fill_2 FILLER_10_470 ();
 sg13g2_fill_1 FILLER_10_472 ();
 sg13g2_fill_1 FILLER_10_495 ();
 sg13g2_fill_2 FILLER_10_500 ();
 sg13g2_fill_1 FILLER_10_506 ();
 sg13g2_fill_1 FILLER_10_538 ();
 sg13g2_fill_1 FILLER_10_544 ();
 sg13g2_fill_1 FILLER_10_549 ();
 sg13g2_fill_1 FILLER_10_555 ();
 sg13g2_fill_1 FILLER_10_591 ();
 sg13g2_fill_1 FILLER_10_597 ();
 sg13g2_fill_1 FILLER_10_602 ();
 sg13g2_fill_1 FILLER_10_607 ();
 sg13g2_fill_1 FILLER_10_613 ();
 sg13g2_fill_1 FILLER_10_635 ();
 sg13g2_fill_2 FILLER_10_640 ();
 sg13g2_fill_1 FILLER_10_647 ();
 sg13g2_fill_2 FILLER_10_722 ();
 sg13g2_decap_8 FILLER_10_736 ();
 sg13g2_fill_1 FILLER_10_743 ();
 sg13g2_decap_4 FILLER_10_748 ();
 sg13g2_fill_2 FILLER_10_752 ();
 sg13g2_fill_2 FILLER_10_778 ();
 sg13g2_fill_1 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_789 ();
 sg13g2_decap_4 FILLER_10_796 ();
 sg13g2_decap_4 FILLER_10_848 ();
 sg13g2_fill_2 FILLER_10_852 ();
 sg13g2_fill_2 FILLER_10_866 ();
 sg13g2_fill_1 FILLER_10_868 ();
 sg13g2_fill_2 FILLER_10_897 ();
 sg13g2_fill_2 FILLER_10_903 ();
 sg13g2_fill_2 FILLER_10_910 ();
 sg13g2_fill_1 FILLER_10_912 ();
 sg13g2_fill_1 FILLER_10_931 ();
 sg13g2_fill_2 FILLER_10_961 ();
 sg13g2_decap_8 FILLER_10_967 ();
 sg13g2_decap_8 FILLER_10_974 ();
 sg13g2_fill_2 FILLER_10_981 ();
 sg13g2_fill_1 FILLER_10_983 ();
 sg13g2_decap_4 FILLER_10_994 ();
 sg13g2_fill_1 FILLER_10_998 ();
 sg13g2_fill_2 FILLER_10_1008 ();
 sg13g2_fill_1 FILLER_10_1010 ();
 sg13g2_fill_2 FILLER_10_1077 ();
 sg13g2_fill_1 FILLER_10_1079 ();
 sg13g2_decap_4 FILLER_10_1084 ();
 sg13g2_fill_2 FILLER_10_1088 ();
 sg13g2_decap_8 FILLER_10_1103 ();
 sg13g2_fill_1 FILLER_10_1110 ();
 sg13g2_decap_4 FILLER_10_1115 ();
 sg13g2_decap_4 FILLER_10_1124 ();
 sg13g2_fill_1 FILLER_10_1140 ();
 sg13g2_decap_4 FILLER_10_1145 ();
 sg13g2_fill_2 FILLER_10_1153 ();
 sg13g2_fill_2 FILLER_10_1224 ();
 sg13g2_fill_1 FILLER_10_1226 ();
 sg13g2_fill_1 FILLER_10_1232 ();
 sg13g2_decap_4 FILLER_10_1247 ();
 sg13g2_decap_8 FILLER_10_1266 ();
 sg13g2_fill_1 FILLER_10_1324 ();
 sg13g2_fill_1 FILLER_10_1343 ();
 sg13g2_fill_2 FILLER_10_1349 ();
 sg13g2_fill_2 FILLER_10_1355 ();
 sg13g2_fill_1 FILLER_10_1357 ();
 sg13g2_fill_1 FILLER_10_1371 ();
 sg13g2_decap_4 FILLER_10_1387 ();
 sg13g2_fill_1 FILLER_10_1405 ();
 sg13g2_fill_1 FILLER_10_1411 ();
 sg13g2_fill_1 FILLER_10_1441 ();
 sg13g2_fill_2 FILLER_10_1448 ();
 sg13g2_fill_2 FILLER_10_1460 ();
 sg13g2_fill_2 FILLER_10_1496 ();
 sg13g2_fill_1 FILLER_10_1503 ();
 sg13g2_fill_1 FILLER_10_1524 ();
 sg13g2_fill_1 FILLER_10_1542 ();
 sg13g2_fill_1 FILLER_10_1547 ();
 sg13g2_decap_4 FILLER_10_1568 ();
 sg13g2_fill_1 FILLER_10_1598 ();
 sg13g2_fill_1 FILLER_10_1604 ();
 sg13g2_fill_1 FILLER_10_1613 ();
 sg13g2_fill_1 FILLER_10_1619 ();
 sg13g2_decap_4 FILLER_10_1629 ();
 sg13g2_fill_1 FILLER_10_1638 ();
 sg13g2_fill_2 FILLER_10_1644 ();
 sg13g2_fill_2 FILLER_10_1651 ();
 sg13g2_decap_8 FILLER_10_1658 ();
 sg13g2_decap_4 FILLER_10_1690 ();
 sg13g2_fill_2 FILLER_10_1699 ();
 sg13g2_fill_2 FILLER_10_1735 ();
 sg13g2_fill_2 FILLER_10_1764 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_43 ();
 sg13g2_fill_1 FILLER_11_53 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_1 FILLER_11_95 ();
 sg13g2_fill_2 FILLER_11_110 ();
 sg13g2_fill_1 FILLER_11_112 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_fill_2 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_323 ();
 sg13g2_fill_2 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_485 ();
 sg13g2_fill_2 FILLER_11_538 ();
 sg13g2_fill_2 FILLER_11_566 ();
 sg13g2_fill_1 FILLER_11_568 ();
 sg13g2_fill_1 FILLER_11_573 ();
 sg13g2_fill_2 FILLER_11_634 ();
 sg13g2_fill_1 FILLER_11_640 ();
 sg13g2_fill_1 FILLER_11_650 ();
 sg13g2_fill_1 FILLER_11_659 ();
 sg13g2_fill_2 FILLER_11_673 ();
 sg13g2_fill_1 FILLER_11_675 ();
 sg13g2_fill_1 FILLER_11_696 ();
 sg13g2_fill_2 FILLER_11_739 ();
 sg13g2_fill_1 FILLER_11_749 ();
 sg13g2_fill_1 FILLER_11_754 ();
 sg13g2_fill_1 FILLER_11_763 ();
 sg13g2_fill_1 FILLER_11_772 ();
 sg13g2_fill_1 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_814 ();
 sg13g2_fill_1 FILLER_11_825 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_4 FILLER_11_875 ();
 sg13g2_fill_1 FILLER_11_892 ();
 sg13g2_fill_2 FILLER_11_901 ();
 sg13g2_fill_1 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_926 ();
 sg13g2_decap_4 FILLER_11_933 ();
 sg13g2_fill_2 FILLER_11_937 ();
 sg13g2_fill_2 FILLER_11_1024 ();
 sg13g2_fill_1 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1032 ();
 sg13g2_fill_1 FILLER_11_1044 ();
 sg13g2_fill_1 FILLER_11_1076 ();
 sg13g2_fill_1 FILLER_11_1086 ();
 sg13g2_fill_2 FILLER_11_1091 ();
 sg13g2_fill_2 FILLER_11_1103 ();
 sg13g2_decap_8 FILLER_11_1109 ();
 sg13g2_fill_1 FILLER_11_1116 ();
 sg13g2_fill_2 FILLER_11_1132 ();
 sg13g2_decap_8 FILLER_11_1147 ();
 sg13g2_decap_8 FILLER_11_1158 ();
 sg13g2_decap_8 FILLER_11_1165 ();
 sg13g2_decap_8 FILLER_11_1172 ();
 sg13g2_fill_1 FILLER_11_1179 ();
 sg13g2_fill_2 FILLER_11_1229 ();
 sg13g2_fill_1 FILLER_11_1231 ();
 sg13g2_decap_4 FILLER_11_1236 ();
 sg13g2_fill_1 FILLER_11_1240 ();
 sg13g2_fill_2 FILLER_11_1248 ();
 sg13g2_fill_1 FILLER_11_1250 ();
 sg13g2_fill_2 FILLER_11_1263 ();
 sg13g2_fill_1 FILLER_11_1265 ();
 sg13g2_fill_2 FILLER_11_1271 ();
 sg13g2_fill_1 FILLER_11_1273 ();
 sg13g2_decap_8 FILLER_11_1284 ();
 sg13g2_fill_2 FILLER_11_1291 ();
 sg13g2_fill_1 FILLER_11_1293 ();
 sg13g2_decap_4 FILLER_11_1330 ();
 sg13g2_decap_4 FILLER_11_1338 ();
 sg13g2_fill_1 FILLER_11_1342 ();
 sg13g2_fill_2 FILLER_11_1355 ();
 sg13g2_fill_1 FILLER_11_1385 ();
 sg13g2_fill_1 FILLER_11_1394 ();
 sg13g2_fill_1 FILLER_11_1403 ();
 sg13g2_fill_1 FILLER_11_1439 ();
 sg13g2_fill_1 FILLER_11_1445 ();
 sg13g2_fill_1 FILLER_11_1451 ();
 sg13g2_fill_1 FILLER_11_1459 ();
 sg13g2_fill_1 FILLER_11_1468 ();
 sg13g2_fill_1 FILLER_11_1474 ();
 sg13g2_fill_1 FILLER_11_1478 ();
 sg13g2_fill_1 FILLER_11_1499 ();
 sg13g2_fill_2 FILLER_11_1514 ();
 sg13g2_fill_2 FILLER_11_1521 ();
 sg13g2_decap_4 FILLER_11_1568 ();
 sg13g2_fill_1 FILLER_11_1572 ();
 sg13g2_fill_2 FILLER_11_1577 ();
 sg13g2_fill_1 FILLER_11_1595 ();
 sg13g2_fill_1 FILLER_11_1623 ();
 sg13g2_fill_1 FILLER_11_1638 ();
 sg13g2_fill_2 FILLER_11_1644 ();
 sg13g2_fill_1 FILLER_11_1651 ();
 sg13g2_decap_8 FILLER_11_1656 ();
 sg13g2_fill_1 FILLER_11_1663 ();
 sg13g2_fill_2 FILLER_11_1688 ();
 sg13g2_fill_2 FILLER_11_1697 ();
 sg13g2_fill_2 FILLER_11_1704 ();
 sg13g2_decap_4 FILLER_11_1710 ();
 sg13g2_fill_1 FILLER_11_1714 ();
 sg13g2_fill_2 FILLER_11_1723 ();
 sg13g2_fill_1 FILLER_11_1725 ();
 sg13g2_fill_1 FILLER_11_1746 ();
 sg13g2_decap_4 FILLER_11_1768 ();
 sg13g2_fill_2 FILLER_11_1772 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_6 ();
 sg13g2_fill_1 FILLER_12_22 ();
 sg13g2_fill_1 FILLER_12_53 ();
 sg13g2_fill_2 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_fill_2 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_275 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_357 ();
 sg13g2_fill_2 FILLER_12_363 ();
 sg13g2_fill_2 FILLER_12_386 ();
 sg13g2_fill_1 FILLER_12_410 ();
 sg13g2_fill_2 FILLER_12_469 ();
 sg13g2_fill_1 FILLER_12_476 ();
 sg13g2_fill_1 FILLER_12_481 ();
 sg13g2_fill_1 FILLER_12_486 ();
 sg13g2_fill_1 FILLER_12_491 ();
 sg13g2_fill_1 FILLER_12_496 ();
 sg13g2_fill_1 FILLER_12_501 ();
 sg13g2_fill_1 FILLER_12_507 ();
 sg13g2_fill_2 FILLER_12_512 ();
 sg13g2_fill_1 FILLER_12_518 ();
 sg13g2_fill_2 FILLER_12_524 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_fill_1 FILLER_12_536 ();
 sg13g2_fill_1 FILLER_12_563 ();
 sg13g2_fill_1 FILLER_12_568 ();
 sg13g2_fill_1 FILLER_12_574 ();
 sg13g2_fill_1 FILLER_12_672 ();
 sg13g2_fill_1 FILLER_12_677 ();
 sg13g2_fill_1 FILLER_12_685 ();
 sg13g2_fill_1 FILLER_12_696 ();
 sg13g2_fill_2 FILLER_12_706 ();
 sg13g2_fill_1 FILLER_12_741 ();
 sg13g2_fill_1 FILLER_12_745 ();
 sg13g2_fill_1 FILLER_12_751 ();
 sg13g2_decap_4 FILLER_12_760 ();
 sg13g2_fill_2 FILLER_12_764 ();
 sg13g2_fill_1 FILLER_12_798 ();
 sg13g2_fill_1 FILLER_12_803 ();
 sg13g2_fill_1 FILLER_12_842 ();
 sg13g2_fill_2 FILLER_12_847 ();
 sg13g2_fill_2 FILLER_12_853 ();
 sg13g2_decap_8 FILLER_12_859 ();
 sg13g2_fill_2 FILLER_12_866 ();
 sg13g2_decap_4 FILLER_12_872 ();
 sg13g2_fill_2 FILLER_12_881 ();
 sg13g2_fill_1 FILLER_12_883 ();
 sg13g2_fill_1 FILLER_12_887 ();
 sg13g2_fill_1 FILLER_12_893 ();
 sg13g2_fill_1 FILLER_12_946 ();
 sg13g2_fill_2 FILLER_12_986 ();
 sg13g2_fill_2 FILLER_12_993 ();
 sg13g2_fill_1 FILLER_12_995 ();
 sg13g2_fill_2 FILLER_12_1014 ();
 sg13g2_fill_2 FILLER_12_1035 ();
 sg13g2_fill_2 FILLER_12_1057 ();
 sg13g2_fill_1 FILLER_12_1072 ();
 sg13g2_fill_2 FILLER_12_1083 ();
 sg13g2_fill_1 FILLER_12_1105 ();
 sg13g2_fill_2 FILLER_12_1111 ();
 sg13g2_fill_1 FILLER_12_1113 ();
 sg13g2_fill_2 FILLER_12_1151 ();
 sg13g2_fill_1 FILLER_12_1153 ();
 sg13g2_fill_1 FILLER_12_1235 ();
 sg13g2_fill_1 FILLER_12_1244 ();
 sg13g2_fill_2 FILLER_12_1254 ();
 sg13g2_fill_1 FILLER_12_1256 ();
 sg13g2_fill_1 FILLER_12_1262 ();
 sg13g2_fill_2 FILLER_12_1268 ();
 sg13g2_fill_2 FILLER_12_1275 ();
 sg13g2_fill_2 FILLER_12_1283 ();
 sg13g2_decap_8 FILLER_12_1294 ();
 sg13g2_decap_8 FILLER_12_1318 ();
 sg13g2_decap_4 FILLER_12_1325 ();
 sg13g2_fill_1 FILLER_12_1329 ();
 sg13g2_decap_4 FILLER_12_1343 ();
 sg13g2_fill_2 FILLER_12_1347 ();
 sg13g2_fill_2 FILLER_12_1370 ();
 sg13g2_fill_1 FILLER_12_1372 ();
 sg13g2_fill_2 FILLER_12_1383 ();
 sg13g2_fill_2 FILLER_12_1390 ();
 sg13g2_decap_8 FILLER_12_1412 ();
 sg13g2_fill_1 FILLER_12_1419 ();
 sg13g2_fill_2 FILLER_12_1434 ();
 sg13g2_fill_1 FILLER_12_1472 ();
 sg13g2_fill_1 FILLER_12_1477 ();
 sg13g2_decap_8 FILLER_12_1483 ();
 sg13g2_decap_4 FILLER_12_1495 ();
 sg13g2_fill_2 FILLER_12_1499 ();
 sg13g2_fill_2 FILLER_12_1511 ();
 sg13g2_fill_1 FILLER_12_1513 ();
 sg13g2_fill_2 FILLER_12_1519 ();
 sg13g2_fill_2 FILLER_12_1559 ();
 sg13g2_fill_2 FILLER_12_1573 ();
 sg13g2_fill_1 FILLER_12_1575 ();
 sg13g2_fill_2 FILLER_12_1580 ();
 sg13g2_fill_1 FILLER_12_1582 ();
 sg13g2_fill_1 FILLER_12_1588 ();
 sg13g2_fill_1 FILLER_12_1594 ();
 sg13g2_fill_1 FILLER_12_1603 ();
 sg13g2_fill_1 FILLER_12_1609 ();
 sg13g2_fill_1 FILLER_12_1615 ();
 sg13g2_fill_2 FILLER_12_1621 ();
 sg13g2_fill_1 FILLER_12_1623 ();
 sg13g2_fill_2 FILLER_12_1628 ();
 sg13g2_fill_1 FILLER_12_1630 ();
 sg13g2_fill_2 FILLER_12_1636 ();
 sg13g2_fill_2 FILLER_12_1667 ();
 sg13g2_fill_1 FILLER_12_1669 ();
 sg13g2_decap_8 FILLER_12_1681 ();
 sg13g2_decap_4 FILLER_12_1688 ();
 sg13g2_fill_2 FILLER_12_1692 ();
 sg13g2_decap_4 FILLER_12_1712 ();
 sg13g2_fill_1 FILLER_12_1719 ();
 sg13g2_fill_1 FILLER_12_1724 ();
 sg13g2_fill_1 FILLER_12_1729 ();
 sg13g2_fill_1 FILLER_12_1745 ();
 sg13g2_fill_2 FILLER_12_1771 ();
 sg13g2_fill_1 FILLER_12_1773 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_27 ();
 sg13g2_fill_2 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_158 ();
 sg13g2_fill_1 FILLER_13_213 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_fill_1 FILLER_13_276 ();
 sg13g2_fill_2 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_337 ();
 sg13g2_fill_1 FILLER_13_364 ();
 sg13g2_fill_1 FILLER_13_370 ();
 sg13g2_fill_1 FILLER_13_402 ();
 sg13g2_fill_2 FILLER_13_426 ();
 sg13g2_fill_1 FILLER_13_476 ();
 sg13g2_fill_2 FILLER_13_508 ();
 sg13g2_fill_2 FILLER_13_541 ();
 sg13g2_fill_1 FILLER_13_543 ();
 sg13g2_fill_1 FILLER_13_548 ();
 sg13g2_fill_1 FILLER_13_557 ();
 sg13g2_fill_1 FILLER_13_580 ();
 sg13g2_fill_1 FILLER_13_585 ();
 sg13g2_fill_1 FILLER_13_595 ();
 sg13g2_fill_1 FILLER_13_601 ();
 sg13g2_fill_1 FILLER_13_610 ();
 sg13g2_fill_1 FILLER_13_646 ();
 sg13g2_fill_2 FILLER_13_658 ();
 sg13g2_fill_1 FILLER_13_660 ();
 sg13g2_decap_4 FILLER_13_665 ();
 sg13g2_fill_1 FILLER_13_674 ();
 sg13g2_fill_1 FILLER_13_679 ();
 sg13g2_fill_2 FILLER_13_688 ();
 sg13g2_fill_2 FILLER_13_694 ();
 sg13g2_fill_1 FILLER_13_706 ();
 sg13g2_fill_2 FILLER_13_712 ();
 sg13g2_decap_4 FILLER_13_718 ();
 sg13g2_decap_4 FILLER_13_727 ();
 sg13g2_fill_2 FILLER_13_736 ();
 sg13g2_fill_2 FILLER_13_743 ();
 sg13g2_fill_1 FILLER_13_745 ();
 sg13g2_decap_4 FILLER_13_760 ();
 sg13g2_fill_2 FILLER_13_764 ();
 sg13g2_decap_8 FILLER_13_779 ();
 sg13g2_fill_1 FILLER_13_797 ();
 sg13g2_fill_2 FILLER_13_802 ();
 sg13g2_fill_1 FILLER_13_830 ();
 sg13g2_fill_2 FILLER_13_877 ();
 sg13g2_fill_1 FILLER_13_879 ();
 sg13g2_fill_1 FILLER_13_888 ();
 sg13g2_fill_2 FILLER_13_902 ();
 sg13g2_fill_1 FILLER_13_904 ();
 sg13g2_fill_2 FILLER_13_908 ();
 sg13g2_fill_1 FILLER_13_910 ();
 sg13g2_fill_1 FILLER_13_915 ();
 sg13g2_fill_2 FILLER_13_940 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_fill_1 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_967 ();
 sg13g2_fill_2 FILLER_13_974 ();
 sg13g2_fill_1 FILLER_13_1006 ();
 sg13g2_fill_1 FILLER_13_1012 ();
 sg13g2_decap_4 FILLER_13_1034 ();
 sg13g2_fill_2 FILLER_13_1054 ();
 sg13g2_fill_1 FILLER_13_1056 ();
 sg13g2_fill_2 FILLER_13_1064 ();
 sg13g2_decap_4 FILLER_13_1074 ();
 sg13g2_fill_2 FILLER_13_1078 ();
 sg13g2_fill_1 FILLER_13_1085 ();
 sg13g2_fill_1 FILLER_13_1090 ();
 sg13g2_fill_2 FILLER_13_1095 ();
 sg13g2_fill_1 FILLER_13_1107 ();
 sg13g2_fill_1 FILLER_13_1132 ();
 sg13g2_fill_2 FILLER_13_1141 ();
 sg13g2_decap_4 FILLER_13_1156 ();
 sg13g2_fill_1 FILLER_13_1160 ();
 sg13g2_fill_2 FILLER_13_1182 ();
 sg13g2_fill_1 FILLER_13_1192 ();
 sg13g2_fill_1 FILLER_13_1214 ();
 sg13g2_fill_1 FILLER_13_1219 ();
 sg13g2_fill_1 FILLER_13_1236 ();
 sg13g2_decap_4 FILLER_13_1242 ();
 sg13g2_fill_2 FILLER_13_1267 ();
 sg13g2_fill_1 FILLER_13_1269 ();
 sg13g2_fill_1 FILLER_13_1277 ();
 sg13g2_fill_1 FILLER_13_1282 ();
 sg13g2_fill_1 FILLER_13_1287 ();
 sg13g2_fill_2 FILLER_13_1292 ();
 sg13g2_decap_8 FILLER_13_1298 ();
 sg13g2_decap_8 FILLER_13_1305 ();
 sg13g2_decap_8 FILLER_13_1312 ();
 sg13g2_decap_4 FILLER_13_1324 ();
 sg13g2_fill_2 FILLER_13_1346 ();
 sg13g2_fill_1 FILLER_13_1348 ();
 sg13g2_fill_1 FILLER_13_1374 ();
 sg13g2_fill_1 FILLER_13_1394 ();
 sg13g2_fill_2 FILLER_13_1400 ();
 sg13g2_fill_1 FILLER_13_1407 ();
 sg13g2_fill_1 FILLER_13_1414 ();
 sg13g2_fill_2 FILLER_13_1424 ();
 sg13g2_fill_1 FILLER_13_1431 ();
 sg13g2_fill_1 FILLER_13_1443 ();
 sg13g2_fill_1 FILLER_13_1448 ();
 sg13g2_fill_1 FILLER_13_1459 ();
 sg13g2_fill_1 FILLER_13_1464 ();
 sg13g2_fill_1 FILLER_13_1483 ();
 sg13g2_fill_1 FILLER_13_1489 ();
 sg13g2_fill_1 FILLER_13_1494 ();
 sg13g2_fill_1 FILLER_13_1500 ();
 sg13g2_fill_1 FILLER_13_1507 ();
 sg13g2_fill_2 FILLER_13_1513 ();
 sg13g2_fill_1 FILLER_13_1520 ();
 sg13g2_fill_2 FILLER_13_1526 ();
 sg13g2_fill_2 FILLER_13_1538 ();
 sg13g2_decap_8 FILLER_13_1548 ();
 sg13g2_fill_1 FILLER_13_1555 ();
 sg13g2_fill_1 FILLER_13_1560 ();
 sg13g2_fill_1 FILLER_13_1566 ();
 sg13g2_fill_1 FILLER_13_1583 ();
 sg13g2_fill_1 FILLER_13_1610 ();
 sg13g2_fill_1 FILLER_13_1616 ();
 sg13g2_decap_8 FILLER_13_1625 ();
 sg13g2_fill_2 FILLER_13_1643 ();
 sg13g2_fill_1 FILLER_13_1650 ();
 sg13g2_fill_1 FILLER_13_1663 ();
 sg13g2_fill_1 FILLER_13_1669 ();
 sg13g2_fill_2 FILLER_13_1676 ();
 sg13g2_fill_1 FILLER_13_1678 ();
 sg13g2_fill_2 FILLER_13_1692 ();
 sg13g2_fill_1 FILLER_13_1708 ();
 sg13g2_fill_1 FILLER_13_1734 ();
 sg13g2_decap_4 FILLER_13_1740 ();
 sg13g2_fill_2 FILLER_13_1744 ();
 sg13g2_decap_4 FILLER_13_1770 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_2 ();
 sg13g2_fill_2 FILLER_14_18 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_80 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_fill_1 FILLER_14_113 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_fill_2 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_2 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_287 ();
 sg13g2_fill_2 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_303 ();
 sg13g2_fill_2 FILLER_14_343 ();
 sg13g2_fill_1 FILLER_14_345 ();
 sg13g2_fill_2 FILLER_14_374 ();
 sg13g2_fill_1 FILLER_14_442 ();
 sg13g2_fill_1 FILLER_14_456 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_fill_2 FILLER_14_504 ();
 sg13g2_fill_1 FILLER_14_506 ();
 sg13g2_fill_1 FILLER_14_554 ();
 sg13g2_fill_1 FILLER_14_560 ();
 sg13g2_fill_1 FILLER_14_587 ();
 sg13g2_fill_1 FILLER_14_592 ();
 sg13g2_fill_2 FILLER_14_619 ();
 sg13g2_fill_1 FILLER_14_631 ();
 sg13g2_fill_2 FILLER_14_644 ();
 sg13g2_fill_2 FILLER_14_672 ();
 sg13g2_fill_1 FILLER_14_674 ();
 sg13g2_fill_1 FILLER_14_758 ();
 sg13g2_fill_1 FILLER_14_764 ();
 sg13g2_fill_2 FILLER_14_782 ();
 sg13g2_fill_1 FILLER_14_784 ();
 sg13g2_fill_1 FILLER_14_790 ();
 sg13g2_fill_1 FILLER_14_797 ();
 sg13g2_fill_2 FILLER_14_838 ();
 sg13g2_fill_1 FILLER_14_850 ();
 sg13g2_decap_4 FILLER_14_875 ();
 sg13g2_fill_2 FILLER_14_891 ();
 sg13g2_fill_2 FILLER_14_904 ();
 sg13g2_fill_1 FILLER_14_906 ();
 sg13g2_fill_2 FILLER_14_912 ();
 sg13g2_decap_8 FILLER_14_923 ();
 sg13g2_fill_2 FILLER_14_930 ();
 sg13g2_fill_1 FILLER_14_932 ();
 sg13g2_decap_4 FILLER_14_964 ();
 sg13g2_decap_4 FILLER_14_972 ();
 sg13g2_fill_1 FILLER_14_976 ();
 sg13g2_decap_4 FILLER_14_982 ();
 sg13g2_decap_4 FILLER_14_990 ();
 sg13g2_fill_1 FILLER_14_998 ();
 sg13g2_fill_1 FILLER_14_1012 ();
 sg13g2_fill_1 FILLER_14_1018 ();
 sg13g2_fill_2 FILLER_14_1055 ();
 sg13g2_fill_1 FILLER_14_1057 ();
 sg13g2_fill_2 FILLER_14_1073 ();
 sg13g2_fill_1 FILLER_14_1075 ();
 sg13g2_decap_4 FILLER_14_1081 ();
 sg13g2_decap_8 FILLER_14_1095 ();
 sg13g2_fill_1 FILLER_14_1109 ();
 sg13g2_fill_2 FILLER_14_1123 ();
 sg13g2_decap_8 FILLER_14_1129 ();
 sg13g2_fill_2 FILLER_14_1136 ();
 sg13g2_fill_1 FILLER_14_1138 ();
 sg13g2_fill_2 FILLER_14_1154 ();
 sg13g2_fill_1 FILLER_14_1156 ();
 sg13g2_fill_1 FILLER_14_1170 ();
 sg13g2_fill_2 FILLER_14_1191 ();
 sg13g2_fill_2 FILLER_14_1201 ();
 sg13g2_decap_4 FILLER_14_1207 ();
 sg13g2_fill_1 FILLER_14_1215 ();
 sg13g2_fill_2 FILLER_14_1224 ();
 sg13g2_fill_1 FILLER_14_1233 ();
 sg13g2_decap_8 FILLER_14_1268 ();
 sg13g2_fill_2 FILLER_14_1275 ();
 sg13g2_fill_1 FILLER_14_1277 ();
 sg13g2_fill_2 FILLER_14_1289 ();
 sg13g2_fill_1 FILLER_14_1298 ();
 sg13g2_fill_2 FILLER_14_1304 ();
 sg13g2_fill_1 FILLER_14_1306 ();
 sg13g2_decap_8 FILLER_14_1316 ();
 sg13g2_fill_2 FILLER_14_1328 ();
 sg13g2_fill_2 FILLER_14_1347 ();
 sg13g2_fill_1 FILLER_14_1364 ();
 sg13g2_fill_1 FILLER_14_1420 ();
 sg13g2_fill_2 FILLER_14_1472 ();
 sg13g2_fill_1 FILLER_14_1479 ();
 sg13g2_fill_1 FILLER_14_1484 ();
 sg13g2_fill_1 FILLER_14_1499 ();
 sg13g2_fill_1 FILLER_14_1528 ();
 sg13g2_fill_1 FILLER_14_1537 ();
 sg13g2_fill_1 FILLER_14_1561 ();
 sg13g2_fill_1 FILLER_14_1567 ();
 sg13g2_fill_2 FILLER_14_1576 ();
 sg13g2_decap_8 FILLER_14_1591 ();
 sg13g2_decap_8 FILLER_14_1598 ();
 sg13g2_decap_8 FILLER_14_1637 ();
 sg13g2_decap_8 FILLER_14_1644 ();
 sg13g2_fill_1 FILLER_14_1655 ();
 sg13g2_fill_1 FILLER_14_1675 ();
 sg13g2_decap_4 FILLER_14_1696 ();
 sg13g2_decap_8 FILLER_14_1710 ();
 sg13g2_fill_2 FILLER_14_1717 ();
 sg13g2_fill_1 FILLER_14_1719 ();
 sg13g2_decap_4 FILLER_14_1732 ();
 sg13g2_fill_2 FILLER_14_1736 ();
 sg13g2_fill_2 FILLER_14_1764 ();
 sg13g2_fill_2 FILLER_14_1771 ();
 sg13g2_fill_1 FILLER_14_1773 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_6 ();
 sg13g2_fill_2 FILLER_15_22 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_78 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_149 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_fill_2 FILLER_15_239 ();
 sg13g2_fill_2 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_261 ();
 sg13g2_fill_1 FILLER_15_263 ();
 sg13g2_fill_2 FILLER_15_276 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_fill_2 FILLER_15_314 ();
 sg13g2_fill_2 FILLER_15_410 ();
 sg13g2_fill_1 FILLER_15_412 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_15_461 ();
 sg13g2_fill_1 FILLER_15_463 ();
 sg13g2_fill_2 FILLER_15_469 ();
 sg13g2_fill_1 FILLER_15_471 ();
 sg13g2_fill_1 FILLER_15_477 ();
 sg13g2_fill_1 FILLER_15_483 ();
 sg13g2_fill_1 FILLER_15_489 ();
 sg13g2_fill_2 FILLER_15_516 ();
 sg13g2_fill_1 FILLER_15_579 ();
 sg13g2_fill_2 FILLER_15_606 ();
 sg13g2_fill_1 FILLER_15_624 ();
 sg13g2_fill_2 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_656 ();
 sg13g2_fill_2 FILLER_15_681 ();
 sg13g2_fill_1 FILLER_15_683 ();
 sg13g2_fill_2 FILLER_15_702 ();
 sg13g2_fill_1 FILLER_15_704 ();
 sg13g2_fill_2 FILLER_15_736 ();
 sg13g2_decap_4 FILLER_15_753 ();
 sg13g2_fill_1 FILLER_15_757 ();
 sg13g2_decap_4 FILLER_15_764 ();
 sg13g2_fill_2 FILLER_15_798 ();
 sg13g2_fill_1 FILLER_15_825 ();
 sg13g2_decap_4 FILLER_15_848 ();
 sg13g2_fill_2 FILLER_15_852 ();
 sg13g2_fill_2 FILLER_15_862 ();
 sg13g2_decap_4 FILLER_15_868 ();
 sg13g2_fill_1 FILLER_15_872 ();
 sg13g2_fill_2 FILLER_15_881 ();
 sg13g2_fill_1 FILLER_15_887 ();
 sg13g2_fill_2 FILLER_15_893 ();
 sg13g2_fill_1 FILLER_15_927 ();
 sg13g2_fill_1 FILLER_15_936 ();
 sg13g2_fill_2 FILLER_15_941 ();
 sg13g2_fill_1 FILLER_15_943 ();
 sg13g2_fill_1 FILLER_15_948 ();
 sg13g2_decap_8 FILLER_15_953 ();
 sg13g2_fill_1 FILLER_15_960 ();
 sg13g2_fill_2 FILLER_15_987 ();
 sg13g2_fill_1 FILLER_15_989 ();
 sg13g2_fill_2 FILLER_15_1008 ();
 sg13g2_fill_1 FILLER_15_1019 ();
 sg13g2_decap_4 FILLER_15_1025 ();
 sg13g2_fill_1 FILLER_15_1029 ();
 sg13g2_decap_4 FILLER_15_1035 ();
 sg13g2_fill_1 FILLER_15_1049 ();
 sg13g2_fill_1 FILLER_15_1055 ();
 sg13g2_fill_1 FILLER_15_1077 ();
 sg13g2_fill_2 FILLER_15_1097 ();
 sg13g2_fill_1 FILLER_15_1099 ();
 sg13g2_fill_1 FILLER_15_1104 ();
 sg13g2_fill_1 FILLER_15_1110 ();
 sg13g2_fill_2 FILLER_15_1115 ();
 sg13g2_decap_8 FILLER_15_1131 ();
 sg13g2_decap_8 FILLER_15_1138 ();
 sg13g2_decap_4 FILLER_15_1145 ();
 sg13g2_fill_2 FILLER_15_1149 ();
 sg13g2_fill_1 FILLER_15_1164 ();
 sg13g2_fill_1 FILLER_15_1170 ();
 sg13g2_decap_4 FILLER_15_1183 ();
 sg13g2_fill_2 FILLER_15_1227 ();
 sg13g2_decap_4 FILLER_15_1274 ();
 sg13g2_decap_4 FILLER_15_1296 ();
 sg13g2_decap_8 FILLER_15_1326 ();
 sg13g2_fill_1 FILLER_15_1363 ();
 sg13g2_fill_2 FILLER_15_1388 ();
 sg13g2_fill_1 FILLER_15_1394 ();
 sg13g2_fill_1 FILLER_15_1413 ();
 sg13g2_fill_2 FILLER_15_1431 ();
 sg13g2_fill_1 FILLER_15_1433 ();
 sg13g2_fill_2 FILLER_15_1449 ();
 sg13g2_fill_1 FILLER_15_1451 ();
 sg13g2_fill_2 FILLER_15_1456 ();
 sg13g2_fill_1 FILLER_15_1458 ();
 sg13g2_fill_1 FILLER_15_1465 ();
 sg13g2_fill_1 FILLER_15_1479 ();
 sg13g2_fill_1 FILLER_15_1485 ();
 sg13g2_fill_1 FILLER_15_1502 ();
 sg13g2_fill_2 FILLER_15_1517 ();
 sg13g2_fill_1 FILLER_15_1527 ();
 sg13g2_fill_2 FILLER_15_1544 ();
 sg13g2_fill_1 FILLER_15_1546 ();
 sg13g2_fill_1 FILLER_15_1576 ();
 sg13g2_fill_2 FILLER_15_1583 ();
 sg13g2_fill_1 FILLER_15_1585 ();
 sg13g2_fill_2 FILLER_15_1594 ();
 sg13g2_fill_1 FILLER_15_1616 ();
 sg13g2_fill_2 FILLER_15_1622 ();
 sg13g2_decap_4 FILLER_15_1637 ();
 sg13g2_fill_2 FILLER_15_1641 ();
 sg13g2_decap_4 FILLER_15_1646 ();
 sg13g2_fill_1 FILLER_15_1650 ();
 sg13g2_decap_8 FILLER_15_1668 ();
 sg13g2_fill_2 FILLER_15_1675 ();
 sg13g2_fill_2 FILLER_15_1701 ();
 sg13g2_fill_1 FILLER_15_1703 ();
 sg13g2_fill_1 FILLER_15_1709 ();
 sg13g2_fill_2 FILLER_15_1719 ();
 sg13g2_fill_1 FILLER_15_1725 ();
 sg13g2_fill_2 FILLER_15_1734 ();
 sg13g2_fill_2 FILLER_15_1772 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_66 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_377 ();
 sg13g2_fill_2 FILLER_16_435 ();
 sg13g2_fill_1 FILLER_16_437 ();
 sg13g2_fill_2 FILLER_16_503 ();
 sg13g2_fill_1 FILLER_16_510 ();
 sg13g2_fill_2 FILLER_16_516 ();
 sg13g2_fill_1 FILLER_16_569 ();
 sg13g2_fill_2 FILLER_16_583 ();
 sg13g2_fill_1 FILLER_16_610 ();
 sg13g2_fill_1 FILLER_16_646 ();
 sg13g2_fill_1 FILLER_16_672 ();
 sg13g2_fill_2 FILLER_16_679 ();
 sg13g2_fill_2 FILLER_16_687 ();
 sg13g2_fill_1 FILLER_16_689 ();
 sg13g2_fill_2 FILLER_16_701 ();
 sg13g2_fill_2 FILLER_16_758 ();
 sg13g2_fill_2 FILLER_16_773 ();
 sg13g2_fill_1 FILLER_16_775 ();
 sg13g2_fill_2 FILLER_16_781 ();
 sg13g2_fill_2 FILLER_16_793 ();
 sg13g2_fill_1 FILLER_16_795 ();
 sg13g2_fill_1 FILLER_16_805 ();
 sg13g2_fill_1 FILLER_16_838 ();
 sg13g2_fill_2 FILLER_16_855 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_fill_2 FILLER_16_870 ();
 sg13g2_fill_2 FILLER_16_919 ();
 sg13g2_fill_2 FILLER_16_929 ();
 sg13g2_fill_1 FILLER_16_943 ();
 sg13g2_fill_1 FILLER_16_952 ();
 sg13g2_fill_2 FILLER_16_967 ();
 sg13g2_fill_2 FILLER_16_1002 ();
 sg13g2_fill_1 FILLER_16_1013 ();
 sg13g2_fill_1 FILLER_16_1023 ();
 sg13g2_fill_1 FILLER_16_1050 ();
 sg13g2_fill_2 FILLER_16_1056 ();
 sg13g2_fill_1 FILLER_16_1058 ();
 sg13g2_fill_1 FILLER_16_1095 ();
 sg13g2_fill_2 FILLER_16_1117 ();
 sg13g2_fill_1 FILLER_16_1119 ();
 sg13g2_decap_8 FILLER_16_1125 ();
 sg13g2_fill_1 FILLER_16_1132 ();
 sg13g2_fill_2 FILLER_16_1137 ();
 sg13g2_fill_1 FILLER_16_1139 ();
 sg13g2_fill_1 FILLER_16_1148 ();
 sg13g2_fill_1 FILLER_16_1157 ();
 sg13g2_fill_1 FILLER_16_1162 ();
 sg13g2_fill_2 FILLER_16_1166 ();
 sg13g2_fill_1 FILLER_16_1176 ();
 sg13g2_fill_1 FILLER_16_1182 ();
 sg13g2_fill_1 FILLER_16_1188 ();
 sg13g2_fill_1 FILLER_16_1194 ();
 sg13g2_fill_2 FILLER_16_1210 ();
 sg13g2_fill_1 FILLER_16_1212 ();
 sg13g2_decap_8 FILLER_16_1217 ();
 sg13g2_fill_1 FILLER_16_1234 ();
 sg13g2_fill_2 FILLER_16_1243 ();
 sg13g2_fill_1 FILLER_16_1249 ();
 sg13g2_fill_2 FILLER_16_1255 ();
 sg13g2_fill_1 FILLER_16_1261 ();
 sg13g2_fill_1 FILLER_16_1269 ();
 sg13g2_fill_1 FILLER_16_1275 ();
 sg13g2_fill_1 FILLER_16_1280 ();
 sg13g2_fill_1 FILLER_16_1294 ();
 sg13g2_decap_4 FILLER_16_1300 ();
 sg13g2_fill_2 FILLER_16_1304 ();
 sg13g2_decap_4 FILLER_16_1326 ();
 sg13g2_decap_4 FILLER_16_1335 ();
 sg13g2_decap_4 FILLER_16_1380 ();
 sg13g2_fill_1 FILLER_16_1393 ();
 sg13g2_fill_2 FILLER_16_1413 ();
 sg13g2_fill_1 FILLER_16_1415 ();
 sg13g2_fill_2 FILLER_16_1442 ();
 sg13g2_fill_1 FILLER_16_1492 ();
 sg13g2_fill_1 FILLER_16_1541 ();
 sg13g2_fill_1 FILLER_16_1550 ();
 sg13g2_fill_2 FILLER_16_1563 ();
 sg13g2_fill_2 FILLER_16_1573 ();
 sg13g2_fill_1 FILLER_16_1588 ();
 sg13g2_fill_2 FILLER_16_1597 ();
 sg13g2_decap_8 FILLER_16_1612 ();
 sg13g2_decap_4 FILLER_16_1619 ();
 sg13g2_decap_4 FILLER_16_1628 ();
 sg13g2_fill_2 FILLER_16_1632 ();
 sg13g2_fill_2 FILLER_16_1649 ();
 sg13g2_decap_8 FILLER_16_1674 ();
 sg13g2_fill_1 FILLER_16_1681 ();
 sg13g2_fill_1 FILLER_16_1691 ();
 sg13g2_fill_1 FILLER_16_1697 ();
 sg13g2_fill_2 FILLER_16_1727 ();
 sg13g2_fill_2 FILLER_16_1733 ();
 sg13g2_decap_4 FILLER_16_1738 ();
 sg13g2_fill_1 FILLER_16_1753 ();
 sg13g2_fill_2 FILLER_16_1767 ();
 sg13g2_fill_1 FILLER_16_1769 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_fill_2 FILLER_17_130 ();
 sg13g2_fill_2 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_297 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_1 FILLER_17_351 ();
 sg13g2_decap_4 FILLER_17_366 ();
 sg13g2_fill_1 FILLER_17_370 ();
 sg13g2_decap_4 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_419 ();
 sg13g2_fill_1 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_431 ();
 sg13g2_fill_2 FILLER_17_456 ();
 sg13g2_fill_2 FILLER_17_467 ();
 sg13g2_fill_1 FILLER_17_469 ();
 sg13g2_fill_2 FILLER_17_592 ();
 sg13g2_fill_1 FILLER_17_620 ();
 sg13g2_fill_2 FILLER_17_628 ();
 sg13g2_fill_1 FILLER_17_639 ();
 sg13g2_fill_2 FILLER_17_671 ();
 sg13g2_fill_2 FILLER_17_685 ();
 sg13g2_fill_2 FILLER_17_693 ();
 sg13g2_fill_2 FILLER_17_699 ();
 sg13g2_fill_1 FILLER_17_725 ();
 sg13g2_fill_1 FILLER_17_730 ();
 sg13g2_fill_1 FILLER_17_743 ();
 sg13g2_decap_4 FILLER_17_776 ();
 sg13g2_fill_2 FILLER_17_780 ();
 sg13g2_fill_2 FILLER_17_798 ();
 sg13g2_fill_1 FILLER_17_800 ();
 sg13g2_fill_1 FILLER_17_811 ();
 sg13g2_fill_1 FILLER_17_835 ();
 sg13g2_fill_2 FILLER_17_841 ();
 sg13g2_fill_2 FILLER_17_851 ();
 sg13g2_fill_2 FILLER_17_857 ();
 sg13g2_fill_2 FILLER_17_864 ();
 sg13g2_fill_1 FILLER_17_866 ();
 sg13g2_fill_2 FILLER_17_892 ();
 sg13g2_fill_1 FILLER_17_922 ();
 sg13g2_fill_1 FILLER_17_931 ();
 sg13g2_fill_2 FILLER_17_966 ();
 sg13g2_fill_1 FILLER_17_968 ();
 sg13g2_decap_4 FILLER_17_983 ();
 sg13g2_fill_1 FILLER_17_995 ();
 sg13g2_fill_1 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1009 ();
 sg13g2_decap_4 FILLER_17_1021 ();
 sg13g2_fill_2 FILLER_17_1025 ();
 sg13g2_decap_8 FILLER_17_1040 ();
 sg13g2_decap_4 FILLER_17_1047 ();
 sg13g2_fill_1 FILLER_17_1051 ();
 sg13g2_fill_2 FILLER_17_1062 ();
 sg13g2_fill_1 FILLER_17_1068 ();
 sg13g2_fill_2 FILLER_17_1077 ();
 sg13g2_fill_1 FILLER_17_1093 ();
 sg13g2_fill_1 FILLER_17_1105 ();
 sg13g2_decap_4 FILLER_17_1116 ();
 sg13g2_fill_2 FILLER_17_1120 ();
 sg13g2_fill_2 FILLER_17_1131 ();
 sg13g2_fill_1 FILLER_17_1133 ();
 sg13g2_fill_1 FILLER_17_1138 ();
 sg13g2_fill_1 FILLER_17_1160 ();
 sg13g2_fill_2 FILLER_17_1166 ();
 sg13g2_fill_1 FILLER_17_1168 ();
 sg13g2_fill_1 FILLER_17_1174 ();
 sg13g2_fill_2 FILLER_17_1180 ();
 sg13g2_fill_2 FILLER_17_1194 ();
 sg13g2_fill_1 FILLER_17_1201 ();
 sg13g2_fill_1 FILLER_17_1211 ();
 sg13g2_fill_1 FILLER_17_1217 ();
 sg13g2_fill_1 FILLER_17_1222 ();
 sg13g2_decap_4 FILLER_17_1255 ();
 sg13g2_fill_1 FILLER_17_1264 ();
 sg13g2_fill_1 FILLER_17_1270 ();
 sg13g2_fill_2 FILLER_17_1275 ();
 sg13g2_fill_1 FILLER_17_1281 ();
 sg13g2_fill_2 FILLER_17_1291 ();
 sg13g2_decap_8 FILLER_17_1297 ();
 sg13g2_decap_4 FILLER_17_1304 ();
 sg13g2_decap_4 FILLER_17_1313 ();
 sg13g2_decap_4 FILLER_17_1335 ();
 sg13g2_fill_1 FILLER_17_1363 ();
 sg13g2_fill_1 FILLER_17_1384 ();
 sg13g2_fill_1 FILLER_17_1391 ();
 sg13g2_fill_1 FILLER_17_1397 ();
 sg13g2_fill_2 FILLER_17_1403 ();
 sg13g2_fill_2 FILLER_17_1415 ();
 sg13g2_decap_4 FILLER_17_1434 ();
 sg13g2_fill_1 FILLER_17_1438 ();
 sg13g2_fill_1 FILLER_17_1444 ();
 sg13g2_fill_2 FILLER_17_1454 ();
 sg13g2_fill_1 FILLER_17_1456 ();
 sg13g2_decap_4 FILLER_17_1542 ();
 sg13g2_fill_1 FILLER_17_1546 ();
 sg13g2_fill_2 FILLER_17_1570 ();
 sg13g2_decap_8 FILLER_17_1585 ();
 sg13g2_fill_1 FILLER_17_1592 ();
 sg13g2_fill_2 FILLER_17_1603 ();
 sg13g2_fill_1 FILLER_17_1605 ();
 sg13g2_fill_1 FILLER_17_1629 ();
 sg13g2_fill_1 FILLER_17_1638 ();
 sg13g2_fill_1 FILLER_17_1649 ();
 sg13g2_fill_2 FILLER_17_1660 ();
 sg13g2_fill_1 FILLER_17_1662 ();
 sg13g2_fill_1 FILLER_17_1668 ();
 sg13g2_fill_1 FILLER_17_1707 ();
 sg13g2_fill_2 FILLER_17_1713 ();
 sg13g2_fill_2 FILLER_17_1720 ();
 sg13g2_fill_1 FILLER_17_1736 ();
 sg13g2_fill_2 FILLER_17_1764 ();
 sg13g2_fill_1 FILLER_17_1773 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_fill_2 FILLER_18_95 ();
 sg13g2_fill_2 FILLER_18_122 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_173 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_1 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_268 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_320 ();
 sg13g2_fill_2 FILLER_18_326 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_348 ();
 sg13g2_fill_2 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_413 ();
 sg13g2_fill_2 FILLER_18_420 ();
 sg13g2_fill_2 FILLER_18_448 ();
 sg13g2_fill_1 FILLER_18_510 ();
 sg13g2_fill_2 FILLER_18_520 ();
 sg13g2_fill_2 FILLER_18_531 ();
 sg13g2_fill_1 FILLER_18_533 ();
 sg13g2_fill_2 FILLER_18_547 ();
 sg13g2_fill_1 FILLER_18_549 ();
 sg13g2_fill_2 FILLER_18_571 ();
 sg13g2_fill_1 FILLER_18_578 ();
 sg13g2_fill_1 FILLER_18_609 ();
 sg13g2_fill_2 FILLER_18_691 ();
 sg13g2_fill_2 FILLER_18_698 ();
 sg13g2_fill_1 FILLER_18_700 ();
 sg13g2_fill_2 FILLER_18_709 ();
 sg13g2_fill_1 FILLER_18_711 ();
 sg13g2_fill_2 FILLER_18_725 ();
 sg13g2_fill_2 FILLER_18_764 ();
 sg13g2_fill_1 FILLER_18_766 ();
 sg13g2_fill_2 FILLER_18_771 ();
 sg13g2_fill_1 FILLER_18_773 ();
 sg13g2_fill_1 FILLER_18_783 ();
 sg13g2_fill_2 FILLER_18_788 ();
 sg13g2_fill_1 FILLER_18_794 ();
 sg13g2_fill_2 FILLER_18_811 ();
 sg13g2_fill_1 FILLER_18_822 ();
 sg13g2_fill_2 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_892 ();
 sg13g2_fill_2 FILLER_18_898 ();
 sg13g2_fill_1 FILLER_18_900 ();
 sg13g2_fill_1 FILLER_18_909 ();
 sg13g2_fill_1 FILLER_18_918 ();
 sg13g2_fill_2 FILLER_18_927 ();
 sg13g2_fill_2 FILLER_18_934 ();
 sg13g2_fill_1 FILLER_18_957 ();
 sg13g2_fill_1 FILLER_18_963 ();
 sg13g2_fill_1 FILLER_18_1024 ();
 sg13g2_fill_2 FILLER_18_1068 ();
 sg13g2_decap_8 FILLER_18_1074 ();
 sg13g2_fill_1 FILLER_18_1090 ();
 sg13g2_fill_1 FILLER_18_1099 ();
 sg13g2_fill_1 FILLER_18_1110 ();
 sg13g2_fill_1 FILLER_18_1114 ();
 sg13g2_fill_2 FILLER_18_1123 ();
 sg13g2_fill_2 FILLER_18_1130 ();
 sg13g2_fill_1 FILLER_18_1132 ();
 sg13g2_fill_2 FILLER_18_1147 ();
 sg13g2_fill_1 FILLER_18_1149 ();
 sg13g2_fill_1 FILLER_18_1168 ();
 sg13g2_fill_1 FILLER_18_1173 ();
 sg13g2_fill_2 FILLER_18_1185 ();
 sg13g2_fill_1 FILLER_18_1187 ();
 sg13g2_decap_8 FILLER_18_1193 ();
 sg13g2_fill_2 FILLER_18_1207 ();
 sg13g2_decap_4 FILLER_18_1214 ();
 sg13g2_decap_4 FILLER_18_1222 ();
 sg13g2_fill_2 FILLER_18_1226 ();
 sg13g2_fill_1 FILLER_18_1233 ();
 sg13g2_fill_1 FILLER_18_1239 ();
 sg13g2_fill_1 FILLER_18_1245 ();
 sg13g2_fill_1 FILLER_18_1251 ();
 sg13g2_fill_2 FILLER_18_1256 ();
 sg13g2_fill_1 FILLER_18_1262 ();
 sg13g2_fill_1 FILLER_18_1267 ();
 sg13g2_fill_2 FILLER_18_1274 ();
 sg13g2_fill_1 FILLER_18_1281 ();
 sg13g2_fill_1 FILLER_18_1292 ();
 sg13g2_fill_1 FILLER_18_1297 ();
 sg13g2_fill_2 FILLER_18_1305 ();
 sg13g2_fill_2 FILLER_18_1311 ();
 sg13g2_fill_2 FILLER_18_1330 ();
 sg13g2_decap_4 FILLER_18_1345 ();
 sg13g2_fill_2 FILLER_18_1349 ();
 sg13g2_fill_2 FILLER_18_1360 ();
 sg13g2_fill_1 FILLER_18_1362 ();
 sg13g2_fill_1 FILLER_18_1367 ();
 sg13g2_fill_1 FILLER_18_1373 ();
 sg13g2_fill_1 FILLER_18_1409 ();
 sg13g2_fill_1 FILLER_18_1425 ();
 sg13g2_fill_1 FILLER_18_1438 ();
 sg13g2_decap_8 FILLER_18_1443 ();
 sg13g2_fill_2 FILLER_18_1508 ();
 sg13g2_fill_1 FILLER_18_1525 ();
 sg13g2_fill_1 FILLER_18_1530 ();
 sg13g2_fill_1 FILLER_18_1546 ();
 sg13g2_fill_1 FILLER_18_1551 ();
 sg13g2_fill_2 FILLER_18_1556 ();
 sg13g2_fill_2 FILLER_18_1562 ();
 sg13g2_fill_1 FILLER_18_1564 ();
 sg13g2_fill_2 FILLER_18_1602 ();
 sg13g2_fill_1 FILLER_18_1609 ();
 sg13g2_fill_2 FILLER_18_1614 ();
 sg13g2_fill_2 FILLER_18_1620 ();
 sg13g2_fill_2 FILLER_18_1627 ();
 sg13g2_fill_2 FILLER_18_1633 ();
 sg13g2_fill_2 FILLER_18_1639 ();
 sg13g2_fill_2 FILLER_18_1650 ();
 sg13g2_fill_1 FILLER_18_1661 ();
 sg13g2_fill_1 FILLER_18_1667 ();
 sg13g2_decap_4 FILLER_18_1676 ();
 sg13g2_fill_2 FILLER_18_1729 ();
 sg13g2_decap_8 FILLER_18_1739 ();
 sg13g2_decap_4 FILLER_18_1746 ();
 sg13g2_fill_1 FILLER_18_1750 ();
 sg13g2_fill_2 FILLER_18_1756 ();
 sg13g2_fill_2 FILLER_18_1771 ();
 sg13g2_fill_1 FILLER_18_1773 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_fill_1 FILLER_19_42 ();
 sg13g2_fill_1 FILLER_19_48 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_fill_1 FILLER_19_91 ();
 sg13g2_fill_2 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_232 ();
 sg13g2_fill_2 FILLER_19_241 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_343 ();
 sg13g2_fill_1 FILLER_19_345 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_353 ();
 sg13g2_fill_2 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_361 ();
 sg13g2_fill_2 FILLER_19_381 ();
 sg13g2_fill_1 FILLER_19_383 ();
 sg13g2_fill_1 FILLER_19_431 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_1 FILLER_19_468 ();
 sg13g2_fill_2 FILLER_19_487 ();
 sg13g2_fill_1 FILLER_19_489 ();
 sg13g2_fill_1 FILLER_19_503 ();
 sg13g2_fill_2 FILLER_19_526 ();
 sg13g2_fill_1 FILLER_19_559 ();
 sg13g2_fill_1 FILLER_19_565 ();
 sg13g2_fill_1 FILLER_19_571 ();
 sg13g2_fill_1 FILLER_19_576 ();
 sg13g2_fill_2 FILLER_19_581 ();
 sg13g2_fill_1 FILLER_19_583 ();
 sg13g2_fill_1 FILLER_19_631 ();
 sg13g2_fill_2 FILLER_19_641 ();
 sg13g2_fill_1 FILLER_19_648 ();
 sg13g2_fill_1 FILLER_19_654 ();
 sg13g2_fill_1 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_702 ();
 sg13g2_fill_1 FILLER_19_718 ();
 sg13g2_fill_1 FILLER_19_763 ();
 sg13g2_fill_2 FILLER_19_769 ();
 sg13g2_fill_1 FILLER_19_771 ();
 sg13g2_fill_1 FILLER_19_810 ();
 sg13g2_decap_4 FILLER_19_815 ();
 sg13g2_decap_8 FILLER_19_894 ();
 sg13g2_decap_4 FILLER_19_901 ();
 sg13g2_fill_2 FILLER_19_905 ();
 sg13g2_fill_1 FILLER_19_944 ();
 sg13g2_fill_2 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_962 ();
 sg13g2_fill_2 FILLER_19_969 ();
 sg13g2_fill_2 FILLER_19_980 ();
 sg13g2_fill_1 FILLER_19_982 ();
 sg13g2_fill_2 FILLER_19_987 ();
 sg13g2_fill_1 FILLER_19_989 ();
 sg13g2_fill_2 FILLER_19_994 ();
 sg13g2_fill_1 FILLER_19_996 ();
 sg13g2_fill_2 FILLER_19_1023 ();
 sg13g2_fill_1 FILLER_19_1025 ();
 sg13g2_fill_1 FILLER_19_1087 ();
 sg13g2_fill_2 FILLER_19_1092 ();
 sg13g2_fill_2 FILLER_19_1098 ();
 sg13g2_decap_4 FILLER_19_1120 ();
 sg13g2_decap_4 FILLER_19_1132 ();
 sg13g2_fill_2 FILLER_19_1136 ();
 sg13g2_fill_2 FILLER_19_1143 ();
 sg13g2_fill_1 FILLER_19_1145 ();
 sg13g2_decap_4 FILLER_19_1150 ();
 sg13g2_fill_2 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1159 ();
 sg13g2_decap_8 FILLER_19_1166 ();
 sg13g2_fill_1 FILLER_19_1173 ();
 sg13g2_fill_2 FILLER_19_1187 ();
 sg13g2_fill_1 FILLER_19_1189 ();
 sg13g2_fill_2 FILLER_19_1213 ();
 sg13g2_decap_8 FILLER_19_1228 ();
 sg13g2_decap_4 FILLER_19_1235 ();
 sg13g2_fill_2 FILLER_19_1253 ();
 sg13g2_fill_1 FILLER_19_1286 ();
 sg13g2_fill_1 FILLER_19_1291 ();
 sg13g2_fill_1 FILLER_19_1297 ();
 sg13g2_fill_1 FILLER_19_1306 ();
 sg13g2_fill_1 FILLER_19_1312 ();
 sg13g2_fill_2 FILLER_19_1329 ();
 sg13g2_fill_1 FILLER_19_1331 ();
 sg13g2_fill_2 FILLER_19_1336 ();
 sg13g2_fill_1 FILLER_19_1338 ();
 sg13g2_fill_1 FILLER_19_1344 ();
 sg13g2_fill_1 FILLER_19_1357 ();
 sg13g2_decap_4 FILLER_19_1363 ();
 sg13g2_fill_2 FILLER_19_1367 ();
 sg13g2_decap_8 FILLER_19_1373 ();
 sg13g2_fill_1 FILLER_19_1380 ();
 sg13g2_fill_2 FILLER_19_1385 ();
 sg13g2_fill_1 FILLER_19_1405 ();
 sg13g2_decap_8 FILLER_19_1410 ();
 sg13g2_fill_2 FILLER_19_1422 ();
 sg13g2_fill_2 FILLER_19_1433 ();
 sg13g2_decap_4 FILLER_19_1440 ();
 sg13g2_fill_1 FILLER_19_1444 ();
 sg13g2_decap_4 FILLER_19_1468 ();
 sg13g2_decap_4 FILLER_19_1506 ();
 sg13g2_fill_2 FILLER_19_1519 ();
 sg13g2_fill_1 FILLER_19_1572 ();
 sg13g2_decap_8 FILLER_19_1594 ();
 sg13g2_fill_1 FILLER_19_1606 ();
 sg13g2_fill_2 FILLER_19_1615 ();
 sg13g2_fill_1 FILLER_19_1617 ();
 sg13g2_fill_2 FILLER_19_1627 ();
 sg13g2_fill_1 FILLER_19_1629 ();
 sg13g2_fill_2 FILLER_19_1645 ();
 sg13g2_fill_1 FILLER_19_1647 ();
 sg13g2_decap_4 FILLER_19_1652 ();
 sg13g2_fill_1 FILLER_19_1664 ();
 sg13g2_fill_2 FILLER_19_1678 ();
 sg13g2_fill_1 FILLER_19_1680 ();
 sg13g2_fill_2 FILLER_19_1696 ();
 sg13g2_fill_1 FILLER_19_1698 ();
 sg13g2_fill_1 FILLER_19_1739 ();
 sg13g2_fill_2 FILLER_19_1748 ();
 sg13g2_decap_8 FILLER_19_1755 ();
 sg13g2_fill_1 FILLER_19_1762 ();
 sg13g2_decap_8 FILLER_19_1767 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_2 FILLER_20_153 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_fill_1 FILLER_20_170 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_188 ();
 sg13g2_decap_4 FILLER_20_225 ();
 sg13g2_decap_4 FILLER_20_234 ();
 sg13g2_fill_2 FILLER_20_242 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_321 ();
 sg13g2_fill_1 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_362 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_394 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_fill_1 FILLER_20_402 ();
 sg13g2_fill_2 FILLER_20_412 ();
 sg13g2_fill_1 FILLER_20_414 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_fill_1 FILLER_20_430 ();
 sg13g2_fill_2 FILLER_20_436 ();
 sg13g2_fill_1 FILLER_20_438 ();
 sg13g2_fill_1 FILLER_20_473 ();
 sg13g2_fill_2 FILLER_20_534 ();
 sg13g2_fill_2 FILLER_20_566 ();
 sg13g2_fill_1 FILLER_20_730 ();
 sg13g2_fill_2 FILLER_20_736 ();
 sg13g2_fill_2 FILLER_20_746 ();
 sg13g2_decap_4 FILLER_20_774 ();
 sg13g2_fill_2 FILLER_20_790 ();
 sg13g2_fill_1 FILLER_20_804 ();
 sg13g2_fill_1 FILLER_20_815 ();
 sg13g2_fill_2 FILLER_20_877 ();
 sg13g2_fill_1 FILLER_20_883 ();
 sg13g2_decap_8 FILLER_20_892 ();
 sg13g2_decap_4 FILLER_20_899 ();
 sg13g2_fill_1 FILLER_20_923 ();
 sg13g2_fill_2 FILLER_20_929 ();
 sg13g2_fill_1 FILLER_20_959 ();
 sg13g2_fill_2 FILLER_20_968 ();
 sg13g2_fill_1 FILLER_20_978 ();
 sg13g2_fill_1 FILLER_20_1016 ();
 sg13g2_fill_2 FILLER_20_1021 ();
 sg13g2_fill_2 FILLER_20_1031 ();
 sg13g2_fill_2 FILLER_20_1076 ();
 sg13g2_fill_1 FILLER_20_1113 ();
 sg13g2_fill_1 FILLER_20_1148 ();
 sg13g2_fill_2 FILLER_20_1153 ();
 sg13g2_fill_1 FILLER_20_1155 ();
 sg13g2_decap_8 FILLER_20_1182 ();
 sg13g2_fill_2 FILLER_20_1189 ();
 sg13g2_fill_1 FILLER_20_1209 ();
 sg13g2_decap_4 FILLER_20_1225 ();
 sg13g2_fill_1 FILLER_20_1239 ();
 sg13g2_fill_1 FILLER_20_1246 ();
 sg13g2_fill_1 FILLER_20_1255 ();
 sg13g2_fill_1 FILLER_20_1260 ();
 sg13g2_fill_2 FILLER_20_1266 ();
 sg13g2_decap_4 FILLER_20_1276 ();
 sg13g2_fill_1 FILLER_20_1280 ();
 sg13g2_decap_4 FILLER_20_1311 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_fill_2 FILLER_20_1358 ();
 sg13g2_fill_2 FILLER_20_1365 ();
 sg13g2_decap_8 FILLER_20_1372 ();
 sg13g2_decap_8 FILLER_20_1379 ();
 sg13g2_fill_1 FILLER_20_1386 ();
 sg13g2_fill_1 FILLER_20_1395 ();
 sg13g2_fill_1 FILLER_20_1410 ();
 sg13g2_fill_1 FILLER_20_1416 ();
 sg13g2_fill_1 FILLER_20_1422 ();
 sg13g2_fill_2 FILLER_20_1443 ();
 sg13g2_decap_8 FILLER_20_1463 ();
 sg13g2_fill_1 FILLER_20_1470 ();
 sg13g2_fill_1 FILLER_20_1480 ();
 sg13g2_fill_1 FILLER_20_1486 ();
 sg13g2_fill_1 FILLER_20_1491 ();
 sg13g2_fill_1 FILLER_20_1497 ();
 sg13g2_fill_1 FILLER_20_1503 ();
 sg13g2_fill_1 FILLER_20_1510 ();
 sg13g2_decap_4 FILLER_20_1515 ();
 sg13g2_fill_2 FILLER_20_1546 ();
 sg13g2_fill_2 FILLER_20_1573 ();
 sg13g2_fill_1 FILLER_20_1587 ();
 sg13g2_fill_2 FILLER_20_1600 ();
 sg13g2_fill_1 FILLER_20_1602 ();
 sg13g2_decap_4 FILLER_20_1633 ();
 sg13g2_fill_1 FILLER_20_1637 ();
 sg13g2_fill_1 FILLER_20_1647 ();
 sg13g2_fill_2 FILLER_20_1680 ();
 sg13g2_fill_2 FILLER_20_1691 ();
 sg13g2_fill_1 FILLER_20_1702 ();
 sg13g2_fill_1 FILLER_20_1725 ();
 sg13g2_decap_8 FILLER_20_1736 ();
 sg13g2_fill_2 FILLER_20_1743 ();
 sg13g2_decap_4 FILLER_20_1770 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_139 ();
 sg13g2_fill_2 FILLER_21_201 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_fill_2 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_225 ();
 sg13g2_fill_1 FILLER_21_257 ();
 sg13g2_fill_2 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_425 ();
 sg13g2_fill_2 FILLER_21_475 ();
 sg13g2_fill_2 FILLER_21_482 ();
 sg13g2_fill_1 FILLER_21_488 ();
 sg13g2_fill_1 FILLER_21_533 ();
 sg13g2_fill_2 FILLER_21_557 ();
 sg13g2_fill_1 FILLER_21_564 ();
 sg13g2_fill_2 FILLER_21_570 ();
 sg13g2_fill_1 FILLER_21_576 ();
 sg13g2_fill_1 FILLER_21_647 ();
 sg13g2_fill_1 FILLER_21_652 ();
 sg13g2_fill_1 FILLER_21_658 ();
 sg13g2_fill_1 FILLER_21_663 ();
 sg13g2_fill_1 FILLER_21_690 ();
 sg13g2_fill_1 FILLER_21_696 ();
 sg13g2_fill_1 FILLER_21_701 ();
 sg13g2_fill_2 FILLER_21_706 ();
 sg13g2_fill_1 FILLER_21_712 ();
 sg13g2_fill_1 FILLER_21_718 ();
 sg13g2_fill_1 FILLER_21_724 ();
 sg13g2_fill_1 FILLER_21_732 ();
 sg13g2_fill_1 FILLER_21_738 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_fill_2 FILLER_21_754 ();
 sg13g2_fill_2 FILLER_21_769 ();
 sg13g2_fill_1 FILLER_21_771 ();
 sg13g2_decap_4 FILLER_21_780 ();
 sg13g2_fill_1 FILLER_21_845 ();
 sg13g2_fill_1 FILLER_21_871 ();
 sg13g2_decap_8 FILLER_21_898 ();
 sg13g2_fill_2 FILLER_21_905 ();
 sg13g2_decap_4 FILLER_21_922 ();
 sg13g2_decap_8 FILLER_21_931 ();
 sg13g2_decap_4 FILLER_21_938 ();
 sg13g2_fill_2 FILLER_21_942 ();
 sg13g2_fill_1 FILLER_21_954 ();
 sg13g2_fill_2 FILLER_21_960 ();
 sg13g2_decap_8 FILLER_21_966 ();
 sg13g2_fill_2 FILLER_21_978 ();
 sg13g2_decap_4 FILLER_21_993 ();
 sg13g2_fill_2 FILLER_21_1002 ();
 sg13g2_fill_1 FILLER_21_1004 ();
 sg13g2_fill_2 FILLER_21_1083 ();
 sg13g2_fill_1 FILLER_21_1102 ();
 sg13g2_fill_2 FILLER_21_1113 ();
 sg13g2_fill_1 FILLER_21_1115 ();
 sg13g2_fill_1 FILLER_21_1172 ();
 sg13g2_fill_2 FILLER_21_1177 ();
 sg13g2_fill_2 FILLER_21_1183 ();
 sg13g2_fill_1 FILLER_21_1189 ();
 sg13g2_fill_1 FILLER_21_1195 ();
 sg13g2_fill_1 FILLER_21_1244 ();
 sg13g2_fill_1 FILLER_21_1248 ();
 sg13g2_fill_2 FILLER_21_1269 ();
 sg13g2_decap_4 FILLER_21_1276 ();
 sg13g2_fill_1 FILLER_21_1280 ();
 sg13g2_fill_1 FILLER_21_1308 ();
 sg13g2_decap_8 FILLER_21_1377 ();
 sg13g2_fill_2 FILLER_21_1384 ();
 sg13g2_fill_1 FILLER_21_1386 ();
 sg13g2_decap_4 FILLER_21_1402 ();
 sg13g2_fill_2 FILLER_21_1410 ();
 sg13g2_fill_1 FILLER_21_1412 ();
 sg13g2_fill_2 FILLER_21_1435 ();
 sg13g2_fill_2 FILLER_21_1462 ();
 sg13g2_fill_1 FILLER_21_1464 ();
 sg13g2_decap_8 FILLER_21_1469 ();
 sg13g2_fill_1 FILLER_21_1476 ();
 sg13g2_fill_1 FILLER_21_1481 ();
 sg13g2_fill_2 FILLER_21_1513 ();
 sg13g2_decap_8 FILLER_21_1520 ();
 sg13g2_fill_2 FILLER_21_1531 ();
 sg13g2_fill_1 FILLER_21_1542 ();
 sg13g2_fill_2 FILLER_21_1547 ();
 sg13g2_fill_1 FILLER_21_1549 ();
 sg13g2_decap_4 FILLER_21_1578 ();
 sg13g2_fill_2 FILLER_21_1582 ();
 sg13g2_fill_2 FILLER_21_1619 ();
 sg13g2_fill_1 FILLER_21_1638 ();
 sg13g2_decap_8 FILLER_21_1671 ();
 sg13g2_fill_1 FILLER_21_1682 ();
 sg13g2_fill_1 FILLER_21_1692 ();
 sg13g2_fill_2 FILLER_21_1701 ();
 sg13g2_fill_1 FILLER_21_1709 ();
 sg13g2_fill_2 FILLER_21_1716 ();
 sg13g2_decap_4 FILLER_21_1723 ();
 sg13g2_fill_1 FILLER_21_1727 ();
 sg13g2_fill_1 FILLER_21_1740 ();
 sg13g2_fill_1 FILLER_21_1745 ();
 sg13g2_fill_1 FILLER_21_1750 ();
 sg13g2_fill_1 FILLER_21_1762 ();
 sg13g2_decap_4 FILLER_21_1768 ();
 sg13g2_fill_2 FILLER_21_1772 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_45 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_fill_1 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_79 ();
 sg13g2_fill_1 FILLER_22_81 ();
 sg13g2_fill_1 FILLER_22_118 ();
 sg13g2_fill_1 FILLER_22_124 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_290 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_361 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_378 ();
 sg13g2_fill_1 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_420 ();
 sg13g2_fill_1 FILLER_22_455 ();
 sg13g2_fill_1 FILLER_22_474 ();
 sg13g2_fill_2 FILLER_22_484 ();
 sg13g2_fill_1 FILLER_22_486 ();
 sg13g2_fill_1 FILLER_22_509 ();
 sg13g2_fill_1 FILLER_22_514 ();
 sg13g2_fill_2 FILLER_22_519 ();
 sg13g2_fill_1 FILLER_22_529 ();
 sg13g2_fill_1 FILLER_22_561 ();
 sg13g2_fill_2 FILLER_22_597 ();
 sg13g2_fill_1 FILLER_22_599 ();
 sg13g2_fill_2 FILLER_22_610 ();
 sg13g2_fill_2 FILLER_22_666 ();
 sg13g2_fill_1 FILLER_22_668 ();
 sg13g2_fill_2 FILLER_22_690 ();
 sg13g2_decap_4 FILLER_22_723 ();
 sg13g2_fill_1 FILLER_22_732 ();
 sg13g2_fill_2 FILLER_22_784 ();
 sg13g2_fill_1 FILLER_22_786 ();
 sg13g2_fill_1 FILLER_22_792 ();
 sg13g2_fill_2 FILLER_22_816 ();
 sg13g2_fill_2 FILLER_22_836 ();
 sg13g2_fill_1 FILLER_22_842 ();
 sg13g2_fill_1 FILLER_22_848 ();
 sg13g2_fill_1 FILLER_22_872 ();
 sg13g2_decap_4 FILLER_22_878 ();
 sg13g2_decap_4 FILLER_22_886 ();
 sg13g2_fill_2 FILLER_22_890 ();
 sg13g2_fill_2 FILLER_22_897 ();
 sg13g2_fill_1 FILLER_22_899 ();
 sg13g2_fill_2 FILLER_22_916 ();
 sg13g2_fill_1 FILLER_22_918 ();
 sg13g2_decap_8 FILLER_22_997 ();
 sg13g2_fill_2 FILLER_22_1019 ();
 sg13g2_fill_1 FILLER_22_1021 ();
 sg13g2_fill_1 FILLER_22_1026 ();
 sg13g2_fill_2 FILLER_22_1058 ();
 sg13g2_fill_1 FILLER_22_1060 ();
 sg13g2_fill_1 FILLER_22_1092 ();
 sg13g2_fill_1 FILLER_22_1105 ();
 sg13g2_fill_1 FILLER_22_1111 ();
 sg13g2_fill_2 FILLER_22_1117 ();
 sg13g2_fill_1 FILLER_22_1119 ();
 sg13g2_fill_1 FILLER_22_1190 ();
 sg13g2_fill_1 FILLER_22_1195 ();
 sg13g2_fill_2 FILLER_22_1222 ();
 sg13g2_fill_1 FILLER_22_1229 ();
 sg13g2_fill_1 FILLER_22_1234 ();
 sg13g2_fill_2 FILLER_22_1240 ();
 sg13g2_fill_1 FILLER_22_1247 ();
 sg13g2_fill_2 FILLER_22_1253 ();
 sg13g2_fill_1 FILLER_22_1255 ();
 sg13g2_decap_4 FILLER_22_1263 ();
 sg13g2_decap_4 FILLER_22_1272 ();
 sg13g2_decap_4 FILLER_22_1283 ();
 sg13g2_decap_4 FILLER_22_1304 ();
 sg13g2_fill_1 FILLER_22_1308 ();
 sg13g2_fill_1 FILLER_22_1314 ();
 sg13g2_fill_1 FILLER_22_1324 ();
 sg13g2_fill_1 FILLER_22_1330 ();
 sg13g2_fill_2 FILLER_22_1335 ();
 sg13g2_fill_1 FILLER_22_1340 ();
 sg13g2_fill_1 FILLER_22_1349 ();
 sg13g2_fill_1 FILLER_22_1380 ();
 sg13g2_fill_2 FILLER_22_1386 ();
 sg13g2_fill_1 FILLER_22_1388 ();
 sg13g2_fill_1 FILLER_22_1394 ();
 sg13g2_fill_2 FILLER_22_1403 ();
 sg13g2_decap_4 FILLER_22_1413 ();
 sg13g2_fill_1 FILLER_22_1417 ();
 sg13g2_fill_2 FILLER_22_1431 ();
 sg13g2_fill_1 FILLER_22_1433 ();
 sg13g2_decap_8 FILLER_22_1451 ();
 sg13g2_decap_8 FILLER_22_1458 ();
 sg13g2_fill_2 FILLER_22_1465 ();
 sg13g2_fill_2 FILLER_22_1471 ();
 sg13g2_fill_2 FILLER_22_1493 ();
 sg13g2_fill_1 FILLER_22_1505 ();
 sg13g2_fill_2 FILLER_22_1511 ();
 sg13g2_fill_1 FILLER_22_1513 ();
 sg13g2_decap_4 FILLER_22_1519 ();
 sg13g2_decap_4 FILLER_22_1535 ();
 sg13g2_fill_1 FILLER_22_1539 ();
 sg13g2_fill_2 FILLER_22_1544 ();
 sg13g2_fill_1 FILLER_22_1546 ();
 sg13g2_fill_2 FILLER_22_1581 ();
 sg13g2_fill_1 FILLER_22_1646 ();
 sg13g2_fill_1 FILLER_22_1656 ();
 sg13g2_fill_2 FILLER_22_1665 ();
 sg13g2_fill_1 FILLER_22_1685 ();
 sg13g2_fill_1 FILLER_22_1703 ();
 sg13g2_fill_1 FILLER_22_1708 ();
 sg13g2_fill_1 FILLER_22_1714 ();
 sg13g2_fill_2 FILLER_22_1732 ();
 sg13g2_fill_1 FILLER_22_1734 ();
 sg13g2_fill_1 FILLER_22_1745 ();
 sg13g2_fill_1 FILLER_22_1751 ();
 sg13g2_fill_2 FILLER_22_1757 ();
 sg13g2_fill_2 FILLER_22_1763 ();
 sg13g2_fill_1 FILLER_22_1773 ();
 sg13g2_fill_2 FILLER_23_26 ();
 sg13g2_fill_1 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_fill_2 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_88 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_259 ();
 sg13g2_fill_2 FILLER_23_265 ();
 sg13g2_fill_1 FILLER_23_267 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_2 FILLER_23_355 ();
 sg13g2_fill_2 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_396 ();
 sg13g2_fill_1 FILLER_23_415 ();
 sg13g2_fill_1 FILLER_23_420 ();
 sg13g2_fill_1 FILLER_23_426 ();
 sg13g2_fill_2 FILLER_23_432 ();
 sg13g2_fill_1 FILLER_23_490 ();
 sg13g2_fill_1 FILLER_23_532 ();
 sg13g2_fill_1 FILLER_23_564 ();
 sg13g2_fill_1 FILLER_23_570 ();
 sg13g2_fill_1 FILLER_23_623 ();
 sg13g2_fill_2 FILLER_23_629 ();
 sg13g2_fill_2 FILLER_23_640 ();
 sg13g2_fill_2 FILLER_23_651 ();
 sg13g2_fill_1 FILLER_23_653 ();
 sg13g2_fill_1 FILLER_23_659 ();
 sg13g2_fill_1 FILLER_23_704 ();
 sg13g2_decap_4 FILLER_23_709 ();
 sg13g2_fill_1 FILLER_23_713 ();
 sg13g2_fill_2 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_737 ();
 sg13g2_decap_4 FILLER_23_751 ();
 sg13g2_fill_1 FILLER_23_755 ();
 sg13g2_fill_1 FILLER_23_767 ();
 sg13g2_fill_1 FILLER_23_803 ();
 sg13g2_fill_2 FILLER_23_812 ();
 sg13g2_fill_1 FILLER_23_822 ();
 sg13g2_fill_1 FILLER_23_859 ();
 sg13g2_fill_1 FILLER_23_863 ();
 sg13g2_fill_1 FILLER_23_870 ();
 sg13g2_fill_1 FILLER_23_874 ();
 sg13g2_fill_2 FILLER_23_901 ();
 sg13g2_fill_1 FILLER_23_903 ();
 sg13g2_fill_1 FILLER_23_910 ();
 sg13g2_fill_1 FILLER_23_917 ();
 sg13g2_decap_4 FILLER_23_932 ();
 sg13g2_fill_1 FILLER_23_936 ();
 sg13g2_fill_2 FILLER_23_942 ();
 sg13g2_fill_2 FILLER_23_953 ();
 sg13g2_fill_1 FILLER_23_995 ();
 sg13g2_fill_2 FILLER_23_1001 ();
 sg13g2_fill_2 FILLER_23_1013 ();
 sg13g2_fill_1 FILLER_23_1015 ();
 sg13g2_decap_4 FILLER_23_1086 ();
 sg13g2_fill_1 FILLER_23_1151 ();
 sg13g2_fill_1 FILLER_23_1160 ();
 sg13g2_fill_1 FILLER_23_1165 ();
 sg13g2_fill_2 FILLER_23_1171 ();
 sg13g2_fill_1 FILLER_23_1173 ();
 sg13g2_fill_2 FILLER_23_1197 ();
 sg13g2_fill_1 FILLER_23_1199 ();
 sg13g2_fill_2 FILLER_23_1205 ();
 sg13g2_fill_1 FILLER_23_1228 ();
 sg13g2_fill_1 FILLER_23_1234 ();
 sg13g2_fill_1 FILLER_23_1247 ();
 sg13g2_fill_1 FILLER_23_1257 ();
 sg13g2_decap_4 FILLER_23_1281 ();
 sg13g2_fill_1 FILLER_23_1285 ();
 sg13g2_fill_1 FILLER_23_1295 ();
 sg13g2_fill_1 FILLER_23_1357 ();
 sg13g2_decap_8 FILLER_23_1367 ();
 sg13g2_decap_4 FILLER_23_1374 ();
 sg13g2_fill_2 FILLER_23_1378 ();
 sg13g2_fill_1 FILLER_23_1385 ();
 sg13g2_fill_1 FILLER_23_1389 ();
 sg13g2_decap_8 FILLER_23_1410 ();
 sg13g2_decap_4 FILLER_23_1417 ();
 sg13g2_fill_1 FILLER_23_1421 ();
 sg13g2_decap_8 FILLER_23_1426 ();
 sg13g2_fill_1 FILLER_23_1442 ();
 sg13g2_fill_2 FILLER_23_1460 ();
 sg13g2_decap_8 FILLER_23_1471 ();
 sg13g2_decap_8 FILLER_23_1478 ();
 sg13g2_fill_2 FILLER_23_1485 ();
 sg13g2_decap_4 FILLER_23_1494 ();
 sg13g2_fill_2 FILLER_23_1548 ();
 sg13g2_fill_1 FILLER_23_1566 ();
 sg13g2_fill_1 FILLER_23_1571 ();
 sg13g2_fill_1 FILLER_23_1578 ();
 sg13g2_fill_1 FILLER_23_1583 ();
 sg13g2_fill_1 FILLER_23_1601 ();
 sg13g2_fill_2 FILLER_23_1606 ();
 sg13g2_fill_1 FILLER_23_1662 ();
 sg13g2_fill_2 FILLER_23_1673 ();
 sg13g2_fill_1 FILLER_23_1675 ();
 sg13g2_fill_1 FILLER_23_1681 ();
 sg13g2_fill_2 FILLER_23_1687 ();
 sg13g2_fill_1 FILLER_23_1689 ();
 sg13g2_fill_1 FILLER_23_1693 ();
 sg13g2_fill_1 FILLER_23_1699 ();
 sg13g2_fill_1 FILLER_23_1710 ();
 sg13g2_fill_1 FILLER_23_1716 ();
 sg13g2_fill_2 FILLER_23_1726 ();
 sg13g2_fill_1 FILLER_23_1735 ();
 sg13g2_decap_8 FILLER_23_1740 ();
 sg13g2_fill_2 FILLER_23_1755 ();
 sg13g2_fill_2 FILLER_23_1771 ();
 sg13g2_fill_1 FILLER_23_1773 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_68 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_80 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_234 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_fill_1 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_411 ();
 sg13g2_fill_1 FILLER_24_438 ();
 sg13g2_fill_2 FILLER_24_465 ();
 sg13g2_fill_1 FILLER_24_467 ();
 sg13g2_fill_1 FILLER_24_493 ();
 sg13g2_fill_1 FILLER_24_546 ();
 sg13g2_fill_1 FILLER_24_551 ();
 sg13g2_fill_1 FILLER_24_556 ();
 sg13g2_decap_8 FILLER_24_562 ();
 sg13g2_fill_2 FILLER_24_573 ();
 sg13g2_fill_2 FILLER_24_579 ();
 sg13g2_fill_1 FILLER_24_581 ();
 sg13g2_fill_1 FILLER_24_586 ();
 sg13g2_fill_2 FILLER_24_669 ();
 sg13g2_fill_2 FILLER_24_688 ();
 sg13g2_fill_2 FILLER_24_696 ();
 sg13g2_decap_4 FILLER_24_707 ();
 sg13g2_fill_1 FILLER_24_715 ();
 sg13g2_fill_1 FILLER_24_724 ();
 sg13g2_fill_1 FILLER_24_729 ();
 sg13g2_fill_1 FILLER_24_738 ();
 sg13g2_fill_2 FILLER_24_756 ();
 sg13g2_fill_1 FILLER_24_774 ();
 sg13g2_fill_1 FILLER_24_821 ();
 sg13g2_fill_1 FILLER_24_834 ();
 sg13g2_fill_1 FILLER_24_840 ();
 sg13g2_fill_1 FILLER_24_845 ();
 sg13g2_fill_1 FILLER_24_850 ();
 sg13g2_fill_1 FILLER_24_854 ();
 sg13g2_fill_2 FILLER_24_867 ();
 sg13g2_fill_1 FILLER_24_869 ();
 sg13g2_decap_4 FILLER_24_886 ();
 sg13g2_fill_2 FILLER_24_890 ();
 sg13g2_fill_1 FILLER_24_898 ();
 sg13g2_fill_2 FILLER_24_924 ();
 sg13g2_fill_1 FILLER_24_926 ();
 sg13g2_fill_1 FILLER_24_958 ();
 sg13g2_fill_2 FILLER_24_986 ();
 sg13g2_fill_2 FILLER_24_1032 ();
 sg13g2_fill_2 FILLER_24_1052 ();
 sg13g2_fill_1 FILLER_24_1054 ();
 sg13g2_fill_2 FILLER_24_1060 ();
 sg13g2_fill_1 FILLER_24_1067 ();
 sg13g2_fill_1 FILLER_24_1094 ();
 sg13g2_fill_2 FILLER_24_1134 ();
 sg13g2_fill_2 FILLER_24_1175 ();
 sg13g2_fill_2 FILLER_24_1189 ();
 sg13g2_fill_1 FILLER_24_1191 ();
 sg13g2_decap_8 FILLER_24_1210 ();
 sg13g2_fill_2 FILLER_24_1217 ();
 sg13g2_fill_1 FILLER_24_1236 ();
 sg13g2_fill_1 FILLER_24_1257 ();
 sg13g2_fill_2 FILLER_24_1276 ();
 sg13g2_fill_1 FILLER_24_1283 ();
 sg13g2_decap_4 FILLER_24_1291 ();
 sg13g2_fill_2 FILLER_24_1295 ();
 sg13g2_fill_1 FILLER_24_1302 ();
 sg13g2_fill_1 FILLER_24_1317 ();
 sg13g2_fill_2 FILLER_24_1412 ();
 sg13g2_fill_2 FILLER_24_1432 ();
 sg13g2_fill_1 FILLER_24_1434 ();
 sg13g2_fill_2 FILLER_24_1443 ();
 sg13g2_fill_1 FILLER_24_1445 ();
 sg13g2_fill_1 FILLER_24_1485 ();
 sg13g2_fill_2 FILLER_24_1490 ();
 sg13g2_decap_4 FILLER_24_1528 ();
 sg13g2_fill_2 FILLER_24_1540 ();
 sg13g2_fill_2 FILLER_24_1557 ();
 sg13g2_fill_1 FILLER_24_1597 ();
 sg13g2_fill_1 FILLER_24_1603 ();
 sg13g2_fill_1 FILLER_24_1609 ();
 sg13g2_fill_1 FILLER_24_1615 ();
 sg13g2_fill_1 FILLER_24_1620 ();
 sg13g2_fill_1 FILLER_24_1629 ();
 sg13g2_decap_8 FILLER_24_1638 ();
 sg13g2_fill_1 FILLER_24_1660 ();
 sg13g2_fill_2 FILLER_24_1665 ();
 sg13g2_fill_1 FILLER_24_1671 ();
 sg13g2_fill_1 FILLER_24_1704 ();
 sg13g2_decap_4 FILLER_24_1710 ();
 sg13g2_fill_2 FILLER_24_1714 ();
 sg13g2_fill_1 FILLER_24_1761 ();
 sg13g2_fill_2 FILLER_24_1766 ();
 sg13g2_fill_2 FILLER_24_1772 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_43 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_fill_2 FILLER_25_104 ();
 sg13g2_fill_1 FILLER_25_106 ();
 sg13g2_fill_1 FILLER_25_111 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_decap_4 FILLER_25_319 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_331 ();
 sg13g2_decap_8 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_415 ();
 sg13g2_fill_1 FILLER_25_426 ();
 sg13g2_fill_2 FILLER_25_436 ();
 sg13g2_fill_1 FILLER_25_438 ();
 sg13g2_fill_1 FILLER_25_452 ();
 sg13g2_fill_2 FILLER_25_471 ();
 sg13g2_fill_2 FILLER_25_477 ();
 sg13g2_fill_1 FILLER_25_484 ();
 sg13g2_fill_2 FILLER_25_511 ();
 sg13g2_fill_1 FILLER_25_513 ();
 sg13g2_fill_1 FILLER_25_518 ();
 sg13g2_fill_1 FILLER_25_523 ();
 sg13g2_fill_2 FILLER_25_528 ();
 sg13g2_fill_2 FILLER_25_534 ();
 sg13g2_fill_1 FILLER_25_536 ();
 sg13g2_fill_2 FILLER_25_576 ();
 sg13g2_fill_1 FILLER_25_586 ();
 sg13g2_fill_1 FILLER_25_592 ();
 sg13g2_decap_4 FILLER_25_619 ();
 sg13g2_decap_4 FILLER_25_631 ();
 sg13g2_decap_4 FILLER_25_640 ();
 sg13g2_fill_2 FILLER_25_661 ();
 sg13g2_fill_2 FILLER_25_701 ();
 sg13g2_fill_2 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_738 ();
 sg13g2_fill_1 FILLER_25_745 ();
 sg13g2_fill_2 FILLER_25_775 ();
 sg13g2_fill_1 FILLER_25_851 ();
 sg13g2_fill_1 FILLER_25_879 ();
 sg13g2_fill_1 FILLER_25_888 ();
 sg13g2_fill_1 FILLER_25_899 ();
 sg13g2_fill_1 FILLER_25_909 ();
 sg13g2_fill_1 FILLER_25_916 ();
 sg13g2_decap_4 FILLER_25_932 ();
 sg13g2_fill_2 FILLER_25_950 ();
 sg13g2_fill_1 FILLER_25_982 ();
 sg13g2_fill_1 FILLER_25_1066 ();
 sg13g2_fill_1 FILLER_25_1077 ();
 sg13g2_fill_2 FILLER_25_1087 ();
 sg13g2_fill_2 FILLER_25_1124 ();
 sg13g2_fill_1 FILLER_25_1170 ();
 sg13g2_fill_1 FILLER_25_1199 ();
 sg13g2_fill_2 FILLER_25_1204 ();
 sg13g2_fill_1 FILLER_25_1211 ();
 sg13g2_fill_2 FILLER_25_1216 ();
 sg13g2_fill_2 FILLER_25_1222 ();
 sg13g2_fill_1 FILLER_25_1259 ();
 sg13g2_decap_4 FILLER_25_1292 ();
 sg13g2_decap_4 FILLER_25_1301 ();
 sg13g2_fill_1 FILLER_25_1305 ();
 sg13g2_fill_1 FILLER_25_1320 ();
 sg13g2_fill_1 FILLER_25_1328 ();
 sg13g2_fill_1 FILLER_25_1336 ();
 sg13g2_fill_2 FILLER_25_1341 ();
 sg13g2_decap_4 FILLER_25_1353 ();
 sg13g2_fill_1 FILLER_25_1357 ();
 sg13g2_fill_2 FILLER_25_1400 ();
 sg13g2_fill_1 FILLER_25_1402 ();
 sg13g2_decap_8 FILLER_25_1411 ();
 sg13g2_decap_4 FILLER_25_1418 ();
 sg13g2_fill_1 FILLER_25_1422 ();
 sg13g2_fill_2 FILLER_25_1460 ();
 sg13g2_decap_4 FILLER_25_1475 ();
 sg13g2_fill_1 FILLER_25_1492 ();
 sg13g2_decap_4 FILLER_25_1497 ();
 sg13g2_fill_2 FILLER_25_1501 ();
 sg13g2_fill_2 FILLER_25_1508 ();
 sg13g2_fill_2 FILLER_25_1527 ();
 sg13g2_decap_8 FILLER_25_1537 ();
 sg13g2_decap_8 FILLER_25_1544 ();
 sg13g2_fill_1 FILLER_25_1551 ();
 sg13g2_fill_2 FILLER_25_1571 ();
 sg13g2_fill_1 FILLER_25_1573 ();
 sg13g2_fill_1 FILLER_25_1584 ();
 sg13g2_fill_2 FILLER_25_1621 ();
 sg13g2_fill_1 FILLER_25_1629 ();
 sg13g2_fill_1 FILLER_25_1641 ();
 sg13g2_decap_4 FILLER_25_1646 ();
 sg13g2_fill_2 FILLER_25_1650 ();
 sg13g2_decap_8 FILLER_25_1660 ();
 sg13g2_fill_1 FILLER_25_1667 ();
 sg13g2_fill_2 FILLER_25_1717 ();
 sg13g2_fill_1 FILLER_25_1723 ();
 sg13g2_fill_1 FILLER_25_1729 ();
 sg13g2_fill_1 FILLER_25_1734 ();
 sg13g2_fill_1 FILLER_25_1739 ();
 sg13g2_fill_1 FILLER_25_1747 ();
 sg13g2_fill_2 FILLER_25_1757 ();
 sg13g2_fill_1 FILLER_25_1759 ();
 sg13g2_fill_2 FILLER_25_1772 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_101 ();
 sg13g2_fill_1 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_165 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_fill_2 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_235 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_263 ();
 sg13g2_fill_1 FILLER_26_265 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_fill_1 FILLER_26_349 ();
 sg13g2_fill_1 FILLER_26_354 ();
 sg13g2_fill_2 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_407 ();
 sg13g2_fill_2 FILLER_26_438 ();
 sg13g2_fill_1 FILLER_26_444 ();
 sg13g2_fill_1 FILLER_26_450 ();
 sg13g2_fill_1 FILLER_26_456 ();
 sg13g2_fill_2 FILLER_26_488 ();
 sg13g2_fill_2 FILLER_26_494 ();
 sg13g2_fill_1 FILLER_26_496 ();
 sg13g2_fill_1 FILLER_26_546 ();
 sg13g2_fill_1 FILLER_26_552 ();
 sg13g2_fill_1 FILLER_26_558 ();
 sg13g2_fill_1 FILLER_26_564 ();
 sg13g2_fill_1 FILLER_26_570 ();
 sg13g2_fill_2 FILLER_26_575 ();
 sg13g2_decap_4 FILLER_26_582 ();
 sg13g2_fill_1 FILLER_26_591 ();
 sg13g2_fill_1 FILLER_26_602 ();
 sg13g2_fill_2 FILLER_26_607 ();
 sg13g2_fill_2 FILLER_26_635 ();
 sg13g2_fill_2 FILLER_26_663 ();
 sg13g2_fill_1 FILLER_26_696 ();
 sg13g2_fill_1 FILLER_26_723 ();
 sg13g2_fill_1 FILLER_26_729 ();
 sg13g2_decap_4 FILLER_26_756 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_fill_2 FILLER_26_772 ();
 sg13g2_decap_8 FILLER_26_778 ();
 sg13g2_decap_4 FILLER_26_785 ();
 sg13g2_fill_1 FILLER_26_789 ();
 sg13g2_fill_1 FILLER_26_807 ();
 sg13g2_fill_1 FILLER_26_816 ();
 sg13g2_fill_2 FILLER_26_837 ();
 sg13g2_decap_4 FILLER_26_850 ();
 sg13g2_fill_1 FILLER_26_854 ();
 sg13g2_fill_2 FILLER_26_862 ();
 sg13g2_fill_2 FILLER_26_868 ();
 sg13g2_fill_2 FILLER_26_891 ();
 sg13g2_fill_1 FILLER_26_893 ();
 sg13g2_fill_1 FILLER_26_897 ();
 sg13g2_fill_2 FILLER_26_902 ();
 sg13g2_fill_1 FILLER_26_904 ();
 sg13g2_fill_1 FILLER_26_924 ();
 sg13g2_fill_2 FILLER_26_930 ();
 sg13g2_fill_1 FILLER_26_936 ();
 sg13g2_fill_1 FILLER_26_981 ();
 sg13g2_decap_4 FILLER_26_987 ();
 sg13g2_fill_1 FILLER_26_996 ();
 sg13g2_fill_1 FILLER_26_1001 ();
 sg13g2_fill_1 FILLER_26_1006 ();
 sg13g2_decap_4 FILLER_26_1016 ();
 sg13g2_fill_2 FILLER_26_1036 ();
 sg13g2_fill_1 FILLER_26_1038 ();
 sg13g2_fill_2 FILLER_26_1056 ();
 sg13g2_fill_2 FILLER_26_1067 ();
 sg13g2_fill_1 FILLER_26_1095 ();
 sg13g2_fill_1 FILLER_26_1101 ();
 sg13g2_decap_8 FILLER_26_1115 ();
 sg13g2_decap_4 FILLER_26_1122 ();
 sg13g2_fill_1 FILLER_26_1126 ();
 sg13g2_fill_1 FILLER_26_1162 ();
 sg13g2_fill_2 FILLER_26_1194 ();
 sg13g2_fill_2 FILLER_26_1227 ();
 sg13g2_decap_4 FILLER_26_1237 ();
 sg13g2_fill_1 FILLER_26_1241 ();
 sg13g2_fill_2 FILLER_26_1260 ();
 sg13g2_fill_1 FILLER_26_1272 ();
 sg13g2_fill_1 FILLER_26_1277 ();
 sg13g2_decap_8 FILLER_26_1285 ();
 sg13g2_decap_8 FILLER_26_1292 ();
 sg13g2_decap_8 FILLER_26_1304 ();
 sg13g2_fill_2 FILLER_26_1311 ();
 sg13g2_fill_2 FILLER_26_1323 ();
 sg13g2_decap_8 FILLER_26_1334 ();
 sg13g2_fill_2 FILLER_26_1341 ();
 sg13g2_fill_1 FILLER_26_1343 ();
 sg13g2_decap_8 FILLER_26_1348 ();
 sg13g2_decap_8 FILLER_26_1355 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_fill_2 FILLER_26_1369 ();
 sg13g2_fill_1 FILLER_26_1388 ();
 sg13g2_fill_1 FILLER_26_1397 ();
 sg13g2_fill_2 FILLER_26_1420 ();
 sg13g2_fill_1 FILLER_26_1427 ();
 sg13g2_fill_1 FILLER_26_1432 ();
 sg13g2_fill_1 FILLER_26_1472 ();
 sg13g2_decap_4 FILLER_26_1477 ();
 sg13g2_fill_1 FILLER_26_1506 ();
 sg13g2_decap_4 FILLER_26_1518 ();
 sg13g2_fill_1 FILLER_26_1543 ();
 sg13g2_fill_2 FILLER_26_1549 ();
 sg13g2_fill_1 FILLER_26_1618 ();
 sg13g2_fill_1 FILLER_26_1649 ();
 sg13g2_fill_1 FILLER_26_1663 ();
 sg13g2_fill_2 FILLER_26_1668 ();
 sg13g2_fill_1 FILLER_26_1670 ();
 sg13g2_fill_1 FILLER_26_1675 ();
 sg13g2_fill_1 FILLER_26_1686 ();
 sg13g2_fill_1 FILLER_26_1691 ();
 sg13g2_fill_1 FILLER_26_1701 ();
 sg13g2_fill_1 FILLER_26_1708 ();
 sg13g2_fill_2 FILLER_26_1763 ();
 sg13g2_decap_4 FILLER_26_1770 ();
 sg13g2_fill_2 FILLER_27_26 ();
 sg13g2_fill_2 FILLER_27_47 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_1 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_162 ();
 sg13g2_fill_2 FILLER_27_167 ();
 sg13g2_fill_1 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_175 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_380 ();
 sg13g2_fill_2 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_388 ();
 sg13g2_fill_1 FILLER_27_398 ();
 sg13g2_fill_2 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_433 ();
 sg13g2_fill_1 FILLER_27_442 ();
 sg13g2_fill_1 FILLER_27_527 ();
 sg13g2_fill_1 FILLER_27_592 ();
 sg13g2_decap_4 FILLER_27_597 ();
 sg13g2_fill_2 FILLER_27_616 ();
 sg13g2_fill_2 FILLER_27_622 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_decap_4 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_633 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_fill_2 FILLER_27_657 ();
 sg13g2_fill_1 FILLER_27_664 ();
 sg13g2_fill_2 FILLER_27_670 ();
 sg13g2_fill_1 FILLER_27_718 ();
 sg13g2_fill_1 FILLER_27_729 ();
 sg13g2_fill_1 FILLER_27_734 ();
 sg13g2_decap_4 FILLER_27_787 ();
 sg13g2_fill_2 FILLER_27_791 ();
 sg13g2_fill_2 FILLER_27_819 ();
 sg13g2_fill_1 FILLER_27_831 ();
 sg13g2_decap_4 FILLER_27_855 ();
 sg13g2_fill_1 FILLER_27_864 ();
 sg13g2_fill_2 FILLER_27_875 ();
 sg13g2_fill_2 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_901 ();
 sg13g2_fill_1 FILLER_27_908 ();
 sg13g2_fill_1 FILLER_27_932 ();
 sg13g2_fill_1 FILLER_27_937 ();
 sg13g2_fill_1 FILLER_27_943 ();
 sg13g2_fill_1 FILLER_27_956 ();
 sg13g2_fill_1 FILLER_27_965 ();
 sg13g2_fill_1 FILLER_27_970 ();
 sg13g2_fill_1 FILLER_27_989 ();
 sg13g2_decap_4 FILLER_27_1025 ();
 sg13g2_fill_1 FILLER_27_1034 ();
 sg13g2_fill_1 FILLER_27_1051 ();
 sg13g2_fill_1 FILLER_27_1061 ();
 sg13g2_fill_2 FILLER_27_1131 ();
 sg13g2_fill_2 FILLER_27_1149 ();
 sg13g2_fill_1 FILLER_27_1156 ();
 sg13g2_fill_2 FILLER_27_1162 ();
 sg13g2_fill_2 FILLER_27_1181 ();
 sg13g2_fill_2 FILLER_27_1204 ();
 sg13g2_fill_1 FILLER_27_1210 ();
 sg13g2_fill_2 FILLER_27_1215 ();
 sg13g2_fill_1 FILLER_27_1221 ();
 sg13g2_fill_2 FILLER_27_1227 ();
 sg13g2_fill_2 FILLER_27_1246 ();
 sg13g2_fill_1 FILLER_27_1248 ();
 sg13g2_decap_4 FILLER_27_1254 ();
 sg13g2_fill_2 FILLER_27_1276 ();
 sg13g2_fill_1 FILLER_27_1278 ();
 sg13g2_fill_2 FILLER_27_1309 ();
 sg13g2_decap_4 FILLER_27_1315 ();
 sg13g2_decap_8 FILLER_27_1322 ();
 sg13g2_decap_8 FILLER_27_1329 ();
 sg13g2_decap_8 FILLER_27_1336 ();
 sg13g2_decap_8 FILLER_27_1343 ();
 sg13g2_decap_4 FILLER_27_1355 ();
 sg13g2_fill_1 FILLER_27_1363 ();
 sg13g2_fill_1 FILLER_27_1371 ();
 sg13g2_fill_1 FILLER_27_1382 ();
 sg13g2_fill_1 FILLER_27_1391 ();
 sg13g2_fill_1 FILLER_27_1403 ();
 sg13g2_fill_1 FILLER_27_1417 ();
 sg13g2_fill_1 FILLER_27_1439 ();
 sg13g2_fill_1 FILLER_27_1448 ();
 sg13g2_fill_1 FILLER_27_1458 ();
 sg13g2_fill_2 FILLER_27_1467 ();
 sg13g2_fill_1 FILLER_27_1469 ();
 sg13g2_decap_4 FILLER_27_1474 ();
 sg13g2_fill_1 FILLER_27_1478 ();
 sg13g2_fill_1 FILLER_27_1491 ();
 sg13g2_fill_1 FILLER_27_1506 ();
 sg13g2_fill_2 FILLER_27_1518 ();
 sg13g2_fill_2 FILLER_27_1543 ();
 sg13g2_decap_4 FILLER_27_1550 ();
 sg13g2_fill_2 FILLER_27_1554 ();
 sg13g2_fill_1 FILLER_27_1566 ();
 sg13g2_fill_1 FILLER_27_1576 ();
 sg13g2_fill_2 FILLER_27_1592 ();
 sg13g2_fill_1 FILLER_27_1594 ();
 sg13g2_fill_1 FILLER_27_1614 ();
 sg13g2_decap_4 FILLER_27_1620 ();
 sg13g2_fill_1 FILLER_27_1629 ();
 sg13g2_fill_1 FILLER_27_1634 ();
 sg13g2_fill_2 FILLER_27_1660 ();
 sg13g2_fill_2 FILLER_27_1667 ();
 sg13g2_fill_1 FILLER_27_1680 ();
 sg13g2_fill_2 FILLER_27_1686 ();
 sg13g2_fill_1 FILLER_27_1688 ();
 sg13g2_fill_2 FILLER_27_1693 ();
 sg13g2_fill_1 FILLER_27_1695 ();
 sg13g2_fill_1 FILLER_27_1701 ();
 sg13g2_fill_1 FILLER_27_1709 ();
 sg13g2_fill_1 FILLER_27_1714 ();
 sg13g2_fill_1 FILLER_27_1719 ();
 sg13g2_fill_2 FILLER_27_1725 ();
 sg13g2_fill_1 FILLER_27_1732 ();
 sg13g2_fill_1 FILLER_27_1737 ();
 sg13g2_fill_2 FILLER_27_1743 ();
 sg13g2_fill_2 FILLER_27_1772 ();
 sg13g2_fill_1 FILLER_28_12 ();
 sg13g2_fill_1 FILLER_28_49 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_130 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_140 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_195 ();
 sg13g2_fill_1 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_250 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_340 ();
 sg13g2_decap_4 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_351 ();
 sg13g2_fill_1 FILLER_28_357 ();
 sg13g2_fill_2 FILLER_28_419 ();
 sg13g2_fill_1 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_426 ();
 sg13g2_fill_1 FILLER_28_454 ();
 sg13g2_fill_1 FILLER_28_460 ();
 sg13g2_fill_2 FILLER_28_487 ();
 sg13g2_decap_4 FILLER_28_493 ();
 sg13g2_fill_2 FILLER_28_497 ();
 sg13g2_fill_2 FILLER_28_504 ();
 sg13g2_fill_2 FILLER_28_555 ();
 sg13g2_fill_1 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_4 FILLER_28_616 ();
 sg13g2_fill_1 FILLER_28_660 ();
 sg13g2_fill_2 FILLER_28_666 ();
 sg13g2_decap_4 FILLER_28_672 ();
 sg13g2_fill_1 FILLER_28_681 ();
 sg13g2_fill_2 FILLER_28_691 ();
 sg13g2_fill_2 FILLER_28_742 ();
 sg13g2_fill_2 FILLER_28_748 ();
 sg13g2_fill_1 FILLER_28_817 ();
 sg13g2_fill_2 FILLER_28_822 ();
 sg13g2_fill_1 FILLER_28_824 ();
 sg13g2_fill_2 FILLER_28_830 ();
 sg13g2_fill_2 FILLER_28_835 ();
 sg13g2_fill_2 FILLER_28_847 ();
 sg13g2_fill_1 FILLER_28_849 ();
 sg13g2_decap_8 FILLER_28_879 ();
 sg13g2_decap_4 FILLER_28_894 ();
 sg13g2_fill_1 FILLER_28_898 ();
 sg13g2_fill_1 FILLER_28_975 ();
 sg13g2_fill_2 FILLER_28_980 ();
 sg13g2_fill_1 FILLER_28_982 ();
 sg13g2_fill_2 FILLER_28_988 ();
 sg13g2_fill_2 FILLER_28_995 ();
 sg13g2_fill_2 FILLER_28_1002 ();
 sg13g2_fill_1 FILLER_28_1081 ();
 sg13g2_fill_1 FILLER_28_1098 ();
 sg13g2_fill_1 FILLER_28_1112 ();
 sg13g2_fill_2 FILLER_28_1117 ();
 sg13g2_fill_2 FILLER_28_1192 ();
 sg13g2_decap_8 FILLER_28_1341 ();
 sg13g2_decap_4 FILLER_28_1348 ();
 sg13g2_fill_2 FILLER_28_1352 ();
 sg13g2_fill_1 FILLER_28_1394 ();
 sg13g2_decap_4 FILLER_28_1405 ();
 sg13g2_fill_1 FILLER_28_1409 ();
 sg13g2_fill_1 FILLER_28_1428 ();
 sg13g2_decap_8 FILLER_28_1438 ();
 sg13g2_decap_4 FILLER_28_1445 ();
 sg13g2_fill_2 FILLER_28_1449 ();
 sg13g2_decap_8 FILLER_28_1463 ();
 sg13g2_fill_2 FILLER_28_1470 ();
 sg13g2_fill_1 FILLER_28_1496 ();
 sg13g2_fill_1 FILLER_28_1502 ();
 sg13g2_fill_1 FILLER_28_1508 ();
 sg13g2_fill_1 FILLER_28_1514 ();
 sg13g2_fill_2 FILLER_28_1527 ();
 sg13g2_fill_1 FILLER_28_1529 ();
 sg13g2_fill_1 FILLER_28_1560 ();
 sg13g2_fill_1 FILLER_28_1571 ();
 sg13g2_fill_1 FILLER_28_1580 ();
 sg13g2_fill_1 FILLER_28_1586 ();
 sg13g2_fill_1 FILLER_28_1597 ();
 sg13g2_fill_1 FILLER_28_1606 ();
 sg13g2_fill_1 FILLER_28_1615 ();
 sg13g2_decap_4 FILLER_28_1620 ();
 sg13g2_fill_2 FILLER_28_1624 ();
 sg13g2_fill_1 FILLER_28_1630 ();
 sg13g2_fill_1 FILLER_28_1636 ();
 sg13g2_fill_1 FILLER_28_1657 ();
 sg13g2_fill_2 FILLER_28_1677 ();
 sg13g2_fill_1 FILLER_28_1684 ();
 sg13g2_fill_1 FILLER_28_1690 ();
 sg13g2_fill_2 FILLER_28_1697 ();
 sg13g2_decap_4 FILLER_28_1712 ();
 sg13g2_fill_1 FILLER_28_1726 ();
 sg13g2_fill_2 FILLER_28_1731 ();
 sg13g2_fill_2 FILLER_28_1748 ();
 sg13g2_decap_4 FILLER_28_1754 ();
 sg13g2_fill_2 FILLER_28_1771 ();
 sg13g2_fill_1 FILLER_28_1773 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_1 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_173 ();
 sg13g2_fill_1 FILLER_29_179 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_fill_2 FILLER_29_222 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_fill_2 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_403 ();
 sg13g2_fill_1 FILLER_29_405 ();
 sg13g2_fill_1 FILLER_29_410 ();
 sg13g2_fill_2 FILLER_29_421 ();
 sg13g2_fill_1 FILLER_29_441 ();
 sg13g2_fill_2 FILLER_29_456 ();
 sg13g2_decap_4 FILLER_29_493 ();
 sg13g2_fill_2 FILLER_29_524 ();
 sg13g2_fill_1 FILLER_29_526 ();
 sg13g2_decap_4 FILLER_29_563 ();
 sg13g2_fill_1 FILLER_29_567 ();
 sg13g2_fill_2 FILLER_29_586 ();
 sg13g2_fill_1 FILLER_29_592 ();
 sg13g2_fill_1 FILLER_29_623 ();
 sg13g2_fill_1 FILLER_29_629 ();
 sg13g2_fill_1 FILLER_29_634 ();
 sg13g2_decap_4 FILLER_29_700 ();
 sg13g2_fill_1 FILLER_29_730 ();
 sg13g2_fill_1 FILLER_29_736 ();
 sg13g2_fill_2 FILLER_29_768 ();
 sg13g2_fill_2 FILLER_29_796 ();
 sg13g2_decap_4 FILLER_29_824 ();
 sg13g2_fill_2 FILLER_29_828 ();
 sg13g2_fill_2 FILLER_29_834 ();
 sg13g2_fill_1 FILLER_29_836 ();
 sg13g2_decap_4 FILLER_29_841 ();
 sg13g2_fill_1 FILLER_29_845 ();
 sg13g2_fill_1 FILLER_29_863 ();
 sg13g2_fill_1 FILLER_29_869 ();
 sg13g2_fill_1 FILLER_29_879 ();
 sg13g2_fill_2 FILLER_29_885 ();
 sg13g2_fill_2 FILLER_29_922 ();
 sg13g2_fill_1 FILLER_29_975 ();
 sg13g2_fill_2 FILLER_29_981 ();
 sg13g2_fill_1 FILLER_29_983 ();
 sg13g2_fill_2 FILLER_29_998 ();
 sg13g2_fill_1 FILLER_29_1000 ();
 sg13g2_fill_2 FILLER_29_1010 ();
 sg13g2_fill_1 FILLER_29_1016 ();
 sg13g2_fill_2 FILLER_29_1021 ();
 sg13g2_fill_1 FILLER_29_1027 ();
 sg13g2_fill_1 FILLER_29_1032 ();
 sg13g2_fill_1 FILLER_29_1038 ();
 sg13g2_fill_2 FILLER_29_1049 ();
 sg13g2_fill_1 FILLER_29_1051 ();
 sg13g2_fill_2 FILLER_29_1122 ();
 sg13g2_fill_1 FILLER_29_1132 ();
 sg13g2_fill_2 FILLER_29_1180 ();
 sg13g2_fill_1 FILLER_29_1182 ();
 sg13g2_fill_2 FILLER_29_1203 ();
 sg13g2_fill_1 FILLER_29_1205 ();
 sg13g2_fill_1 FILLER_29_1223 ();
 sg13g2_fill_2 FILLER_29_1259 ();
 sg13g2_fill_1 FILLER_29_1265 ();
 sg13g2_fill_1 FILLER_29_1271 ();
 sg13g2_fill_1 FILLER_29_1276 ();
 sg13g2_fill_1 FILLER_29_1282 ();
 sg13g2_fill_1 FILLER_29_1287 ();
 sg13g2_fill_2 FILLER_29_1303 ();
 sg13g2_fill_1 FILLER_29_1305 ();
 sg13g2_fill_2 FILLER_29_1310 ();
 sg13g2_decap_8 FILLER_29_1342 ();
 sg13g2_decap_8 FILLER_29_1349 ();
 sg13g2_fill_2 FILLER_29_1377 ();
 sg13g2_fill_1 FILLER_29_1399 ();
 sg13g2_fill_1 FILLER_29_1415 ();
 sg13g2_fill_1 FILLER_29_1421 ();
 sg13g2_fill_2 FILLER_29_1430 ();
 sg13g2_decap_4 FILLER_29_1442 ();
 sg13g2_fill_2 FILLER_29_1459 ();
 sg13g2_decap_8 FILLER_29_1465 ();
 sg13g2_fill_2 FILLER_29_1472 ();
 sg13g2_fill_1 FILLER_29_1490 ();
 sg13g2_fill_1 FILLER_29_1513 ();
 sg13g2_fill_1 FILLER_29_1526 ();
 sg13g2_fill_1 FILLER_29_1532 ();
 sg13g2_fill_1 FILLER_29_1538 ();
 sg13g2_fill_1 FILLER_29_1543 ();
 sg13g2_fill_2 FILLER_29_1551 ();
 sg13g2_fill_1 FILLER_29_1559 ();
 sg13g2_fill_2 FILLER_29_1564 ();
 sg13g2_fill_2 FILLER_29_1571 ();
 sg13g2_fill_1 FILLER_29_1578 ();
 sg13g2_fill_2 FILLER_29_1614 ();
 sg13g2_decap_4 FILLER_29_1644 ();
 sg13g2_fill_2 FILLER_29_1698 ();
 sg13g2_fill_1 FILLER_29_1700 ();
 sg13g2_fill_2 FILLER_29_1721 ();
 sg13g2_fill_2 FILLER_29_1737 ();
 sg13g2_fill_2 FILLER_29_1771 ();
 sg13g2_fill_1 FILLER_29_1773 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_79 ();
 sg13g2_fill_2 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_fill_2 FILLER_30_246 ();
 sg13g2_decap_4 FILLER_30_261 ();
 sg13g2_decap_4 FILLER_30_269 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_decap_4 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_fill_2 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_1 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_359 ();
 sg13g2_fill_2 FILLER_30_365 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_4 FILLER_30_386 ();
 sg13g2_fill_1 FILLER_30_390 ();
 sg13g2_fill_1 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_2 FILLER_30_434 ();
 sg13g2_fill_1 FILLER_30_436 ();
 sg13g2_fill_2 FILLER_30_454 ();
 sg13g2_fill_2 FILLER_30_473 ();
 sg13g2_decap_4 FILLER_30_575 ();
 sg13g2_fill_1 FILLER_30_579 ();
 sg13g2_fill_1 FILLER_30_589 ();
 sg13g2_fill_2 FILLER_30_595 ();
 sg13g2_fill_1 FILLER_30_610 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_1 FILLER_30_650 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_fill_1 FILLER_30_662 ();
 sg13g2_fill_2 FILLER_30_720 ();
 sg13g2_fill_1 FILLER_30_748 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_fill_1 FILLER_30_760 ();
 sg13g2_fill_2 FILLER_30_798 ();
 sg13g2_fill_2 FILLER_30_808 ();
 sg13g2_fill_1 FILLER_30_810 ();
 sg13g2_decap_8 FILLER_30_853 ();
 sg13g2_fill_2 FILLER_30_860 ();
 sg13g2_fill_2 FILLER_30_867 ();
 sg13g2_fill_2 FILLER_30_873 ();
 sg13g2_decap_8 FILLER_30_879 ();
 sg13g2_fill_2 FILLER_30_961 ();
 sg13g2_fill_1 FILLER_30_981 ();
 sg13g2_fill_2 FILLER_30_1063 ();
 sg13g2_fill_1 FILLER_30_1065 ();
 sg13g2_fill_1 FILLER_30_1077 ();
 sg13g2_fill_1 FILLER_30_1085 ();
 sg13g2_fill_1 FILLER_30_1090 ();
 sg13g2_fill_1 FILLER_30_1095 ();
 sg13g2_fill_1 FILLER_30_1157 ();
 sg13g2_fill_2 FILLER_30_1263 ();
 sg13g2_fill_1 FILLER_30_1265 ();
 sg13g2_fill_2 FILLER_30_1296 ();
 sg13g2_fill_1 FILLER_30_1328 ();
 sg13g2_fill_2 FILLER_30_1359 ();
 sg13g2_decap_4 FILLER_30_1369 ();
 sg13g2_fill_1 FILLER_30_1373 ();
 sg13g2_fill_2 FILLER_30_1383 ();
 sg13g2_fill_1 FILLER_30_1385 ();
 sg13g2_fill_1 FILLER_30_1396 ();
 sg13g2_fill_2 FILLER_30_1402 ();
 sg13g2_fill_2 FILLER_30_1408 ();
 sg13g2_fill_2 FILLER_30_1415 ();
 sg13g2_decap_4 FILLER_30_1421 ();
 sg13g2_fill_1 FILLER_30_1425 ();
 sg13g2_fill_2 FILLER_30_1433 ();
 sg13g2_fill_1 FILLER_30_1435 ();
 sg13g2_fill_1 FILLER_30_1459 ();
 sg13g2_fill_2 FILLER_30_1468 ();
 sg13g2_fill_1 FILLER_30_1470 ();
 sg13g2_fill_1 FILLER_30_1496 ();
 sg13g2_fill_1 FILLER_30_1512 ();
 sg13g2_fill_1 FILLER_30_1521 ();
 sg13g2_fill_2 FILLER_30_1600 ();
 sg13g2_fill_1 FILLER_30_1606 ();
 sg13g2_fill_1 FILLER_30_1616 ();
 sg13g2_fill_1 FILLER_30_1620 ();
 sg13g2_fill_1 FILLER_30_1627 ();
 sg13g2_fill_1 FILLER_30_1650 ();
 sg13g2_fill_1 FILLER_30_1657 ();
 sg13g2_fill_1 FILLER_30_1684 ();
 sg13g2_fill_1 FILLER_30_1690 ();
 sg13g2_fill_1 FILLER_30_1704 ();
 sg13g2_fill_1 FILLER_30_1711 ();
 sg13g2_fill_2 FILLER_30_1720 ();
 sg13g2_fill_1 FILLER_30_1722 ();
 sg13g2_fill_2 FILLER_30_1742 ();
 sg13g2_fill_1 FILLER_30_1752 ();
 sg13g2_fill_1 FILLER_30_1758 ();
 sg13g2_decap_8 FILLER_30_1767 ();
 sg13g2_fill_1 FILLER_31_13 ();
 sg13g2_fill_2 FILLER_31_24 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_87 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_106 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_1 FILLER_31_152 ();
 sg13g2_fill_2 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_169 ();
 sg13g2_fill_1 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_186 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_decap_8 FILLER_31_284 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_328 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_fill_1 FILLER_31_359 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_403 ();
 sg13g2_fill_2 FILLER_31_484 ();
 sg13g2_fill_2 FILLER_31_490 ();
 sg13g2_fill_1 FILLER_31_492 ();
 sg13g2_decap_8 FILLER_31_502 ();
 sg13g2_fill_1 FILLER_31_509 ();
 sg13g2_fill_2 FILLER_31_545 ();
 sg13g2_fill_1 FILLER_31_547 ();
 sg13g2_fill_1 FILLER_31_557 ();
 sg13g2_fill_1 FILLER_31_588 ();
 sg13g2_decap_4 FILLER_31_620 ();
 sg13g2_fill_2 FILLER_31_628 ();
 sg13g2_fill_2 FILLER_31_656 ();
 sg13g2_fill_1 FILLER_31_663 ();
 sg13g2_fill_2 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_697 ();
 sg13g2_fill_1 FILLER_31_711 ();
 sg13g2_fill_2 FILLER_31_716 ();
 sg13g2_fill_2 FILLER_31_722 ();
 sg13g2_fill_1 FILLER_31_724 ();
 sg13g2_fill_1 FILLER_31_729 ();
 sg13g2_fill_2 FILLER_31_734 ();
 sg13g2_fill_1 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_746 ();
 sg13g2_decap_8 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_760 ();
 sg13g2_fill_1 FILLER_31_791 ();
 sg13g2_fill_1 FILLER_31_797 ();
 sg13g2_fill_2 FILLER_31_803 ();
 sg13g2_decap_4 FILLER_31_899 ();
 sg13g2_decap_4 FILLER_31_907 ();
 sg13g2_decap_4 FILLER_31_915 ();
 sg13g2_decap_8 FILLER_31_923 ();
 sg13g2_fill_1 FILLER_31_930 ();
 sg13g2_fill_1 FILLER_31_985 ();
 sg13g2_fill_2 FILLER_31_990 ();
 sg13g2_fill_2 FILLER_31_1015 ();
 sg13g2_fill_2 FILLER_31_1040 ();
 sg13g2_fill_1 FILLER_31_1074 ();
 sg13g2_fill_2 FILLER_31_1112 ();
 sg13g2_fill_2 FILLER_31_1156 ();
 sg13g2_fill_2 FILLER_31_1196 ();
 sg13g2_decap_4 FILLER_31_1202 ();
 sg13g2_decap_8 FILLER_31_1214 ();
 sg13g2_fill_2 FILLER_31_1221 ();
 sg13g2_fill_1 FILLER_31_1223 ();
 sg13g2_fill_1 FILLER_31_1242 ();
 sg13g2_fill_1 FILLER_31_1247 ();
 sg13g2_fill_2 FILLER_31_1283 ();
 sg13g2_fill_2 FILLER_31_1289 ();
 sg13g2_fill_1 FILLER_31_1291 ();
 sg13g2_fill_1 FILLER_31_1296 ();
 sg13g2_fill_2 FILLER_31_1302 ();
 sg13g2_fill_2 FILLER_31_1308 ();
 sg13g2_fill_2 FILLER_31_1314 ();
 sg13g2_fill_2 FILLER_31_1320 ();
 sg13g2_fill_2 FILLER_31_1326 ();
 sg13g2_fill_1 FILLER_31_1328 ();
 sg13g2_fill_1 FILLER_31_1334 ();
 sg13g2_fill_2 FILLER_31_1339 ();
 sg13g2_fill_1 FILLER_31_1341 ();
 sg13g2_decap_8 FILLER_31_1368 ();
 sg13g2_fill_1 FILLER_31_1403 ();
 sg13g2_fill_1 FILLER_31_1415 ();
 sg13g2_fill_2 FILLER_31_1433 ();
 sg13g2_fill_2 FILLER_31_1440 ();
 sg13g2_fill_1 FILLER_31_1442 ();
 sg13g2_fill_1 FILLER_31_1447 ();
 sg13g2_fill_2 FILLER_31_1461 ();
 sg13g2_decap_4 FILLER_31_1470 ();
 sg13g2_decap_8 FILLER_31_1507 ();
 sg13g2_fill_2 FILLER_31_1514 ();
 sg13g2_fill_2 FILLER_31_1536 ();
 sg13g2_fill_2 FILLER_31_1550 ();
 sg13g2_decap_4 FILLER_31_1556 ();
 sg13g2_fill_2 FILLER_31_1560 ();
 sg13g2_decap_8 FILLER_31_1567 ();
 sg13g2_fill_1 FILLER_31_1574 ();
 sg13g2_fill_1 FILLER_31_1597 ();
 sg13g2_fill_2 FILLER_31_1608 ();
 sg13g2_fill_1 FILLER_31_1610 ();
 sg13g2_decap_8 FILLER_31_1648 ();
 sg13g2_fill_2 FILLER_31_1660 ();
 sg13g2_fill_1 FILLER_31_1662 ();
 sg13g2_fill_2 FILLER_31_1675 ();
 sg13g2_fill_1 FILLER_31_1677 ();
 sg13g2_fill_1 FILLER_31_1686 ();
 sg13g2_fill_2 FILLER_31_1692 ();
 sg13g2_fill_1 FILLER_31_1694 ();
 sg13g2_fill_2 FILLER_31_1708 ();
 sg13g2_decap_4 FILLER_31_1714 ();
 sg13g2_fill_1 FILLER_31_1745 ();
 sg13g2_fill_2 FILLER_31_1751 ();
 sg13g2_fill_1 FILLER_31_1758 ();
 sg13g2_fill_1 FILLER_31_1764 ();
 sg13g2_decap_4 FILLER_31_1770 ();
 sg13g2_fill_1 FILLER_32_41 ();
 sg13g2_fill_1 FILLER_32_47 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_114 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_314 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_382 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_427 ();
 sg13g2_fill_2 FILLER_32_431 ();
 sg13g2_decap_4 FILLER_32_443 ();
 sg13g2_fill_2 FILLER_32_447 ();
 sg13g2_fill_1 FILLER_32_480 ();
 sg13g2_fill_1 FILLER_32_485 ();
 sg13g2_fill_2 FILLER_32_491 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_2 FILLER_32_503 ();
 sg13g2_fill_1 FILLER_32_535 ();
 sg13g2_fill_2 FILLER_32_541 ();
 sg13g2_fill_1 FILLER_32_548 ();
 sg13g2_fill_2 FILLER_32_554 ();
 sg13g2_fill_2 FILLER_32_582 ();
 sg13g2_fill_1 FILLER_32_584 ();
 sg13g2_fill_1 FILLER_32_589 ();
 sg13g2_fill_1 FILLER_32_595 ();
 sg13g2_fill_2 FILLER_32_604 ();
 sg13g2_fill_2 FILLER_32_610 ();
 sg13g2_fill_1 FILLER_32_616 ();
 sg13g2_fill_1 FILLER_32_635 ();
 sg13g2_decap_4 FILLER_32_663 ();
 sg13g2_fill_2 FILLER_32_690 ();
 sg13g2_fill_1 FILLER_32_701 ();
 sg13g2_fill_2 FILLER_32_779 ();
 sg13g2_fill_2 FILLER_32_791 ();
 sg13g2_fill_2 FILLER_32_808 ();
 sg13g2_fill_1 FILLER_32_836 ();
 sg13g2_fill_2 FILLER_32_845 ();
 sg13g2_fill_1 FILLER_32_873 ();
 sg13g2_fill_1 FILLER_32_879 ();
 sg13g2_fill_1 FILLER_32_906 ();
 sg13g2_fill_2 FILLER_32_911 ();
 sg13g2_fill_1 FILLER_32_927 ();
 sg13g2_fill_1 FILLER_32_932 ();
 sg13g2_fill_2 FILLER_32_971 ();
 sg13g2_fill_2 FILLER_32_1032 ();
 sg13g2_fill_2 FILLER_32_1053 ();
 sg13g2_fill_1 FILLER_32_1085 ();
 sg13g2_fill_1 FILLER_32_1116 ();
 sg13g2_fill_1 FILLER_32_1139 ();
 sg13g2_fill_2 FILLER_32_1180 ();
 sg13g2_fill_1 FILLER_32_1196 ();
 sg13g2_fill_2 FILLER_32_1223 ();
 sg13g2_fill_2 FILLER_32_1264 ();
 sg13g2_fill_1 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1340 ();
 sg13g2_fill_1 FILLER_32_1347 ();
 sg13g2_fill_2 FILLER_32_1360 ();
 sg13g2_fill_1 FILLER_32_1362 ();
 sg13g2_decap_4 FILLER_32_1367 ();
 sg13g2_fill_2 FILLER_32_1371 ();
 sg13g2_fill_1 FILLER_32_1381 ();
 sg13g2_fill_2 FILLER_32_1398 ();
 sg13g2_fill_1 FILLER_32_1400 ();
 sg13g2_fill_1 FILLER_32_1406 ();
 sg13g2_fill_1 FILLER_32_1415 ();
 sg13g2_fill_1 FILLER_32_1424 ();
 sg13g2_fill_1 FILLER_32_1438 ();
 sg13g2_fill_1 FILLER_32_1446 ();
 sg13g2_fill_1 FILLER_32_1453 ();
 sg13g2_fill_2 FILLER_32_1462 ();
 sg13g2_fill_2 FILLER_32_1469 ();
 sg13g2_fill_2 FILLER_32_1476 ();
 sg13g2_fill_1 FILLER_32_1478 ();
 sg13g2_decap_8 FILLER_32_1487 ();
 sg13g2_fill_2 FILLER_32_1494 ();
 sg13g2_fill_1 FILLER_32_1496 ();
 sg13g2_fill_1 FILLER_32_1502 ();
 sg13g2_decap_8 FILLER_32_1507 ();
 sg13g2_decap_8 FILLER_32_1514 ();
 sg13g2_fill_2 FILLER_32_1529 ();
 sg13g2_fill_1 FILLER_32_1535 ();
 sg13g2_decap_4 FILLER_32_1570 ();
 sg13g2_fill_1 FILLER_32_1587 ();
 sg13g2_decap_4 FILLER_32_1601 ();
 sg13g2_fill_1 FILLER_32_1605 ();
 sg13g2_decap_4 FILLER_32_1610 ();
 sg13g2_fill_2 FILLER_32_1614 ();
 sg13g2_fill_2 FILLER_32_1653 ();
 sg13g2_fill_1 FILLER_32_1655 ();
 sg13g2_fill_1 FILLER_32_1661 ();
 sg13g2_fill_2 FILLER_32_1670 ();
 sg13g2_fill_1 FILLER_32_1741 ();
 sg13g2_fill_1 FILLER_32_1747 ();
 sg13g2_fill_1 FILLER_32_1753 ();
 sg13g2_fill_2 FILLER_32_1758 ();
 sg13g2_decap_8 FILLER_32_1764 ();
 sg13g2_fill_2 FILLER_32_1771 ();
 sg13g2_fill_1 FILLER_32_1773 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_150 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_254 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_decap_4 FILLER_33_368 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_2 FILLER_33_432 ();
 sg13g2_fill_1 FILLER_33_434 ();
 sg13g2_fill_2 FILLER_33_438 ();
 sg13g2_fill_1 FILLER_33_445 ();
 sg13g2_fill_2 FILLER_33_450 ();
 sg13g2_fill_2 FILLER_33_457 ();
 sg13g2_fill_2 FILLER_33_463 ();
 sg13g2_fill_1 FILLER_33_465 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_fill_1 FILLER_33_520 ();
 sg13g2_fill_2 FILLER_33_547 ();
 sg13g2_fill_2 FILLER_33_558 ();
 sg13g2_fill_2 FILLER_33_565 ();
 sg13g2_fill_1 FILLER_33_567 ();
 sg13g2_fill_2 FILLER_33_577 ();
 sg13g2_fill_2 FILLER_33_583 ();
 sg13g2_fill_1 FILLER_33_630 ();
 sg13g2_fill_1 FILLER_33_639 ();
 sg13g2_fill_1 FILLER_33_645 ();
 sg13g2_fill_1 FILLER_33_650 ();
 sg13g2_fill_1 FILLER_33_656 ();
 sg13g2_fill_1 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_678 ();
 sg13g2_fill_1 FILLER_33_690 ();
 sg13g2_fill_1 FILLER_33_701 ();
 sg13g2_decap_4 FILLER_33_708 ();
 sg13g2_fill_1 FILLER_33_712 ();
 sg13g2_fill_1 FILLER_33_717 ();
 sg13g2_fill_2 FILLER_33_726 ();
 sg13g2_fill_2 FILLER_33_744 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_fill_1 FILLER_33_761 ();
 sg13g2_fill_1 FILLER_33_766 ();
 sg13g2_fill_1 FILLER_33_771 ();
 sg13g2_fill_1 FILLER_33_777 ();
 sg13g2_fill_1 FILLER_33_785 ();
 sg13g2_fill_1 FILLER_33_803 ();
 sg13g2_fill_1 FILLER_33_809 ();
 sg13g2_fill_1 FILLER_33_827 ();
 sg13g2_fill_1 FILLER_33_866 ();
 sg13g2_fill_1 FILLER_33_875 ();
 sg13g2_decap_4 FILLER_33_886 ();
 sg13g2_fill_2 FILLER_33_890 ();
 sg13g2_fill_1 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_933 ();
 sg13g2_fill_2 FILLER_33_940 ();
 sg13g2_fill_1 FILLER_33_942 ();
 sg13g2_fill_1 FILLER_33_947 ();
 sg13g2_fill_1 FILLER_33_953 ();
 sg13g2_fill_1 FILLER_33_959 ();
 sg13g2_fill_2 FILLER_33_985 ();
 sg13g2_fill_1 FILLER_33_987 ();
 sg13g2_fill_1 FILLER_33_1005 ();
 sg13g2_fill_2 FILLER_33_1036 ();
 sg13g2_fill_1 FILLER_33_1042 ();
 sg13g2_fill_2 FILLER_33_1048 ();
 sg13g2_fill_1 FILLER_33_1054 ();
 sg13g2_fill_1 FILLER_33_1059 ();
 sg13g2_fill_2 FILLER_33_1069 ();
 sg13g2_fill_1 FILLER_33_1071 ();
 sg13g2_fill_2 FILLER_33_1084 ();
 sg13g2_fill_1 FILLER_33_1086 ();
 sg13g2_fill_1 FILLER_33_1101 ();
 sg13g2_fill_1 FILLER_33_1111 ();
 sg13g2_fill_2 FILLER_33_1117 ();
 sg13g2_fill_2 FILLER_33_1157 ();
 sg13g2_fill_2 FILLER_33_1198 ();
 sg13g2_fill_1 FILLER_33_1200 ();
 sg13g2_fill_1 FILLER_33_1272 ();
 sg13g2_fill_1 FILLER_33_1277 ();
 sg13g2_fill_1 FILLER_33_1283 ();
 sg13g2_fill_2 FILLER_33_1288 ();
 sg13g2_fill_2 FILLER_33_1303 ();
 sg13g2_fill_2 FILLER_33_1310 ();
 sg13g2_fill_1 FILLER_33_1312 ();
 sg13g2_fill_1 FILLER_33_1330 ();
 sg13g2_fill_1 FILLER_33_1363 ();
 sg13g2_fill_2 FILLER_33_1369 ();
 sg13g2_fill_1 FILLER_33_1371 ();
 sg13g2_decap_4 FILLER_33_1386 ();
 sg13g2_fill_1 FILLER_33_1390 ();
 sg13g2_decap_4 FILLER_33_1396 ();
 sg13g2_fill_1 FILLER_33_1400 ();
 sg13g2_fill_2 FILLER_33_1414 ();
 sg13g2_decap_8 FILLER_33_1436 ();
 sg13g2_decap_4 FILLER_33_1443 ();
 sg13g2_fill_2 FILLER_33_1447 ();
 sg13g2_decap_4 FILLER_33_1457 ();
 sg13g2_fill_1 FILLER_33_1461 ();
 sg13g2_fill_1 FILLER_33_1470 ();
 sg13g2_fill_2 FILLER_33_1513 ();
 sg13g2_fill_1 FILLER_33_1530 ();
 sg13g2_decap_4 FILLER_33_1560 ();
 sg13g2_fill_2 FILLER_33_1611 ();
 sg13g2_fill_1 FILLER_33_1626 ();
 sg13g2_fill_1 FILLER_33_1632 ();
 sg13g2_fill_2 FILLER_33_1638 ();
 sg13g2_fill_1 FILLER_33_1648 ();
 sg13g2_fill_1 FILLER_33_1659 ();
 sg13g2_fill_2 FILLER_33_1664 ();
 sg13g2_fill_1 FILLER_33_1666 ();
 sg13g2_fill_2 FILLER_33_1676 ();
 sg13g2_fill_1 FILLER_33_1678 ();
 sg13g2_fill_1 FILLER_33_1686 ();
 sg13g2_fill_2 FILLER_33_1692 ();
 sg13g2_fill_1 FILLER_33_1703 ();
 sg13g2_fill_1 FILLER_33_1714 ();
 sg13g2_fill_2 FILLER_33_1719 ();
 sg13g2_fill_1 FILLER_33_1726 ();
 sg13g2_fill_1 FILLER_33_1734 ();
 sg13g2_fill_2 FILLER_33_1740 ();
 sg13g2_fill_2 FILLER_33_1750 ();
 sg13g2_fill_2 FILLER_33_1756 ();
 sg13g2_fill_2 FILLER_33_1771 ();
 sg13g2_fill_1 FILLER_33_1773 ();
 sg13g2_fill_2 FILLER_34_26 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_113 ();
 sg13g2_fill_1 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_fill_2 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_decap_8 FILLER_34_268 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_decap_4 FILLER_34_482 ();
 sg13g2_fill_2 FILLER_34_486 ();
 sg13g2_fill_1 FILLER_34_497 ();
 sg13g2_fill_1 FILLER_34_524 ();
 sg13g2_fill_2 FILLER_34_533 ();
 sg13g2_fill_1 FILLER_34_569 ();
 sg13g2_fill_2 FILLER_34_579 ();
 sg13g2_fill_1 FILLER_34_597 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_decap_4 FILLER_34_607 ();
 sg13g2_fill_1 FILLER_34_611 ();
 sg13g2_fill_1 FILLER_34_626 ();
 sg13g2_fill_1 FILLER_34_632 ();
 sg13g2_fill_1 FILLER_34_651 ();
 sg13g2_fill_2 FILLER_34_672 ();
 sg13g2_fill_1 FILLER_34_679 ();
 sg13g2_fill_2 FILLER_34_685 ();
 sg13g2_fill_1 FILLER_34_701 ();
 sg13g2_fill_2 FILLER_34_723 ();
 sg13g2_fill_2 FILLER_34_764 ();
 sg13g2_fill_1 FILLER_34_766 ();
 sg13g2_fill_1 FILLER_34_783 ();
 sg13g2_decap_4 FILLER_34_788 ();
 sg13g2_fill_2 FILLER_34_792 ();
 sg13g2_decap_4 FILLER_34_809 ();
 sg13g2_fill_2 FILLER_34_813 ();
 sg13g2_fill_1 FILLER_34_858 ();
 sg13g2_fill_2 FILLER_34_889 ();
 sg13g2_decap_4 FILLER_34_895 ();
 sg13g2_fill_2 FILLER_34_899 ();
 sg13g2_fill_2 FILLER_34_951 ();
 sg13g2_fill_1 FILLER_34_953 ();
 sg13g2_fill_2 FILLER_34_977 ();
 sg13g2_fill_2 FILLER_34_999 ();
 sg13g2_fill_1 FILLER_34_1001 ();
 sg13g2_fill_1 FILLER_34_1006 ();
 sg13g2_fill_1 FILLER_34_1041 ();
 sg13g2_fill_1 FILLER_34_1046 ();
 sg13g2_fill_1 FILLER_34_1052 ();
 sg13g2_fill_1 FILLER_34_1058 ();
 sg13g2_fill_1 FILLER_34_1063 ();
 sg13g2_fill_1 FILLER_34_1072 ();
 sg13g2_decap_4 FILLER_34_1113 ();
 sg13g2_fill_1 FILLER_34_1134 ();
 sg13g2_fill_1 FILLER_34_1179 ();
 sg13g2_fill_2 FILLER_34_1191 ();
 sg13g2_fill_1 FILLER_34_1193 ();
 sg13g2_fill_2 FILLER_34_1265 ();
 sg13g2_fill_1 FILLER_34_1267 ();
 sg13g2_fill_2 FILLER_34_1347 ();
 sg13g2_fill_1 FILLER_34_1349 ();
 sg13g2_decap_8 FILLER_34_1380 ();
 sg13g2_decap_4 FILLER_34_1387 ();
 sg13g2_fill_2 FILLER_34_1391 ();
 sg13g2_fill_2 FILLER_34_1397 ();
 sg13g2_fill_2 FILLER_34_1408 ();
 sg13g2_fill_1 FILLER_34_1410 ();
 sg13g2_fill_2 FILLER_34_1437 ();
 sg13g2_fill_2 FILLER_34_1456 ();
 sg13g2_fill_1 FILLER_34_1458 ();
 sg13g2_fill_2 FILLER_34_1464 ();
 sg13g2_decap_4 FILLER_34_1470 ();
 sg13g2_fill_2 FILLER_34_1474 ();
 sg13g2_fill_1 FILLER_34_1487 ();
 sg13g2_decap_4 FILLER_34_1493 ();
 sg13g2_fill_1 FILLER_34_1513 ();
 sg13g2_fill_1 FILLER_34_1531 ();
 sg13g2_fill_2 FILLER_34_1548 ();
 sg13g2_fill_1 FILLER_34_1550 ();
 sg13g2_fill_2 FILLER_34_1573 ();
 sg13g2_fill_2 FILLER_34_1597 ();
 sg13g2_fill_1 FILLER_34_1608 ();
 sg13g2_fill_1 FILLER_34_1614 ();
 sg13g2_decap_4 FILLER_34_1647 ();
 sg13g2_fill_2 FILLER_34_1665 ();
 sg13g2_decap_8 FILLER_34_1672 ();
 sg13g2_fill_2 FILLER_34_1679 ();
 sg13g2_fill_1 FILLER_34_1681 ();
 sg13g2_fill_2 FILLER_34_1704 ();
 sg13g2_fill_2 FILLER_34_1711 ();
 sg13g2_fill_2 FILLER_34_1718 ();
 sg13g2_fill_2 FILLER_34_1724 ();
 sg13g2_fill_1 FILLER_34_1736 ();
 sg13g2_fill_1 FILLER_34_1742 ();
 sg13g2_fill_1 FILLER_34_1748 ();
 sg13g2_fill_2 FILLER_34_1753 ();
 sg13g2_fill_1 FILLER_34_1755 ();
 sg13g2_decap_8 FILLER_34_1763 ();
 sg13g2_decap_4 FILLER_34_1770 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_80 ();
 sg13g2_fill_1 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_154 ();
 sg13g2_fill_2 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_291 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_decap_4 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_fill_2 FILLER_35_354 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_2 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_420 ();
 sg13g2_fill_2 FILLER_35_427 ();
 sg13g2_fill_1 FILLER_35_442 ();
 sg13g2_fill_2 FILLER_35_455 ();
 sg13g2_fill_2 FILLER_35_542 ();
 sg13g2_fill_2 FILLER_35_552 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_566 ();
 sg13g2_fill_1 FILLER_35_588 ();
 sg13g2_fill_1 FILLER_35_602 ();
 sg13g2_fill_1 FILLER_35_629 ();
 sg13g2_fill_1 FILLER_35_682 ();
 sg13g2_fill_2 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_695 ();
 sg13g2_fill_2 FILLER_35_701 ();
 sg13g2_fill_2 FILLER_35_737 ();
 sg13g2_fill_1 FILLER_35_750 ();
 sg13g2_fill_1 FILLER_35_755 ();
 sg13g2_fill_2 FILLER_35_781 ();
 sg13g2_fill_2 FILLER_35_834 ();
 sg13g2_fill_2 FILLER_35_840 ();
 sg13g2_fill_1 FILLER_35_842 ();
 sg13g2_fill_1 FILLER_35_856 ();
 sg13g2_fill_1 FILLER_35_879 ();
 sg13g2_fill_1 FILLER_35_895 ();
 sg13g2_fill_1 FILLER_35_926 ();
 sg13g2_fill_2 FILLER_35_941 ();
 sg13g2_fill_1 FILLER_35_948 ();
 sg13g2_fill_1 FILLER_35_954 ();
 sg13g2_fill_1 FILLER_35_960 ();
 sg13g2_fill_2 FILLER_35_966 ();
 sg13g2_fill_2 FILLER_35_994 ();
 sg13g2_fill_2 FILLER_35_1000 ();
 sg13g2_fill_2 FILLER_35_1021 ();
 sg13g2_fill_2 FILLER_35_1032 ();
 sg13g2_fill_1 FILLER_35_1034 ();
 sg13g2_fill_1 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1055 ();
 sg13g2_fill_2 FILLER_35_1091 ();
 sg13g2_fill_1 FILLER_35_1093 ();
 sg13g2_fill_1 FILLER_35_1103 ();
 sg13g2_fill_1 FILLER_35_1109 ();
 sg13g2_fill_1 FILLER_35_1192 ();
 sg13g2_decap_4 FILLER_35_1235 ();
 sg13g2_fill_1 FILLER_35_1243 ();
 sg13g2_fill_1 FILLER_35_1252 ();
 sg13g2_fill_1 FILLER_35_1257 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_fill_2 FILLER_35_1319 ();
 sg13g2_decap_4 FILLER_35_1326 ();
 sg13g2_fill_1 FILLER_35_1330 ();
 sg13g2_fill_2 FILLER_35_1361 ();
 sg13g2_fill_1 FILLER_35_1363 ();
 sg13g2_fill_2 FILLER_35_1382 ();
 sg13g2_decap_8 FILLER_35_1389 ();
 sg13g2_decap_4 FILLER_35_1396 ();
 sg13g2_fill_2 FILLER_35_1400 ();
 sg13g2_decap_4 FILLER_35_1415 ();
 sg13g2_fill_1 FILLER_35_1424 ();
 sg13g2_fill_2 FILLER_35_1430 ();
 sg13g2_fill_2 FILLER_35_1437 ();
 sg13g2_fill_1 FILLER_35_1439 ();
 sg13g2_fill_2 FILLER_35_1444 ();
 sg13g2_fill_2 FILLER_35_1459 ();
 sg13g2_fill_1 FILLER_35_1465 ();
 sg13g2_fill_1 FILLER_35_1471 ();
 sg13g2_decap_8 FILLER_35_1492 ();
 sg13g2_fill_1 FILLER_35_1513 ();
 sg13g2_decap_4 FILLER_35_1523 ();
 sg13g2_fill_1 FILLER_35_1533 ();
 sg13g2_fill_1 FILLER_35_1551 ();
 sg13g2_fill_2 FILLER_35_1617 ();
 sg13g2_fill_1 FILLER_35_1643 ();
 sg13g2_fill_2 FILLER_35_1651 ();
 sg13g2_fill_1 FILLER_35_1653 ();
 sg13g2_fill_1 FILLER_35_1667 ();
 sg13g2_fill_1 FILLER_35_1685 ();
 sg13g2_fill_1 FILLER_35_1695 ();
 sg13g2_fill_1 FILLER_35_1700 ();
 sg13g2_fill_1 FILLER_35_1709 ();
 sg13g2_fill_2 FILLER_35_1745 ();
 sg13g2_fill_2 FILLER_35_1771 ();
 sg13g2_fill_1 FILLER_35_1773 ();
 sg13g2_fill_1 FILLER_36_112 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_fill_1 FILLER_36_137 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_244 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_decap_4 FILLER_36_360 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_378 ();
 sg13g2_fill_2 FILLER_36_389 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_fill_1 FILLER_36_464 ();
 sg13g2_fill_1 FILLER_36_470 ();
 sg13g2_fill_2 FILLER_36_485 ();
 sg13g2_fill_2 FILLER_36_493 ();
 sg13g2_fill_1 FILLER_36_543 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_2 FILLER_36_562 ();
 sg13g2_fill_1 FILLER_36_564 ();
 sg13g2_fill_2 FILLER_36_586 ();
 sg13g2_fill_2 FILLER_36_592 ();
 sg13g2_fill_1 FILLER_36_594 ();
 sg13g2_fill_1 FILLER_36_621 ();
 sg13g2_fill_1 FILLER_36_631 ();
 sg13g2_fill_1 FILLER_36_636 ();
 sg13g2_fill_1 FILLER_36_641 ();
 sg13g2_decap_4 FILLER_36_674 ();
 sg13g2_fill_2 FILLER_36_678 ();
 sg13g2_fill_2 FILLER_36_685 ();
 sg13g2_fill_1 FILLER_36_692 ();
 sg13g2_fill_1 FILLER_36_701 ();
 sg13g2_fill_2 FILLER_36_737 ();
 sg13g2_fill_1 FILLER_36_759 ();
 sg13g2_fill_1 FILLER_36_819 ();
 sg13g2_fill_2 FILLER_36_877 ();
 sg13g2_fill_2 FILLER_36_893 ();
 sg13g2_fill_2 FILLER_36_909 ();
 sg13g2_fill_1 FILLER_36_911 ();
 sg13g2_fill_2 FILLER_36_940 ();
 sg13g2_fill_1 FILLER_36_942 ();
 sg13g2_fill_1 FILLER_36_947 ();
 sg13g2_fill_1 FILLER_36_974 ();
 sg13g2_fill_2 FILLER_36_992 ();
 sg13g2_fill_2 FILLER_36_1003 ();
 sg13g2_fill_1 FILLER_36_1005 ();
 sg13g2_fill_1 FILLER_36_1049 ();
 sg13g2_fill_1 FILLER_36_1055 ();
 sg13g2_fill_1 FILLER_36_1061 ();
 sg13g2_fill_1 FILLER_36_1080 ();
 sg13g2_fill_2 FILLER_36_1111 ();
 sg13g2_fill_2 FILLER_36_1126 ();
 sg13g2_fill_1 FILLER_36_1132 ();
 sg13g2_fill_1 FILLER_36_1137 ();
 sg13g2_fill_1 FILLER_36_1170 ();
 sg13g2_fill_2 FILLER_36_1180 ();
 sg13g2_fill_1 FILLER_36_1199 ();
 sg13g2_fill_2 FILLER_36_1235 ();
 sg13g2_fill_1 FILLER_36_1237 ();
 sg13g2_fill_2 FILLER_36_1273 ();
 sg13g2_fill_1 FILLER_36_1279 ();
 sg13g2_fill_2 FILLER_36_1315 ();
 sg13g2_fill_1 FILLER_36_1386 ();
 sg13g2_fill_1 FILLER_36_1392 ();
 sg13g2_decap_4 FILLER_36_1409 ();
 sg13g2_fill_1 FILLER_36_1413 ();
 sg13g2_fill_2 FILLER_36_1444 ();
 sg13g2_fill_1 FILLER_36_1446 ();
 sg13g2_decap_4 FILLER_36_1455 ();
 sg13g2_fill_2 FILLER_36_1459 ();
 sg13g2_decap_4 FILLER_36_1476 ();
 sg13g2_fill_1 FILLER_36_1480 ();
 sg13g2_decap_8 FILLER_36_1511 ();
 sg13g2_decap_8 FILLER_36_1530 ();
 sg13g2_fill_2 FILLER_36_1537 ();
 sg13g2_fill_1 FILLER_36_1548 ();
 sg13g2_decap_4 FILLER_36_1554 ();
 sg13g2_fill_2 FILLER_36_1562 ();
 sg13g2_fill_1 FILLER_36_1587 ();
 sg13g2_decap_4 FILLER_36_1613 ();
 sg13g2_fill_2 FILLER_36_1634 ();
 sg13g2_fill_1 FILLER_36_1636 ();
 sg13g2_decap_8 FILLER_36_1651 ();
 sg13g2_fill_2 FILLER_36_1658 ();
 sg13g2_fill_1 FILLER_36_1660 ();
 sg13g2_decap_4 FILLER_36_1674 ();
 sg13g2_fill_1 FILLER_36_1678 ();
 sg13g2_fill_2 FILLER_36_1694 ();
 sg13g2_fill_1 FILLER_36_1696 ();
 sg13g2_fill_1 FILLER_36_1702 ();
 sg13g2_decap_4 FILLER_36_1707 ();
 sg13g2_fill_2 FILLER_36_1733 ();
 sg13g2_fill_1 FILLER_36_1756 ();
 sg13g2_fill_2 FILLER_36_1761 ();
 sg13g2_fill_1 FILLER_36_1763 ();
 sg13g2_decap_4 FILLER_36_1768 ();
 sg13g2_fill_2 FILLER_36_1772 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_17 ();
 sg13g2_fill_1 FILLER_37_95 ();
 sg13g2_fill_1 FILLER_37_100 ();
 sg13g2_fill_1 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_122 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_1 FILLER_37_161 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_2 FILLER_37_343 ();
 sg13g2_fill_2 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_425 ();
 sg13g2_fill_1 FILLER_37_427 ();
 sg13g2_fill_2 FILLER_37_432 ();
 sg13g2_fill_1 FILLER_37_434 ();
 sg13g2_fill_2 FILLER_37_444 ();
 sg13g2_fill_1 FILLER_37_456 ();
 sg13g2_fill_1 FILLER_37_464 ();
 sg13g2_decap_4 FILLER_37_469 ();
 sg13g2_fill_1 FILLER_37_473 ();
 sg13g2_fill_1 FILLER_37_500 ();
 sg13g2_decap_4 FILLER_37_515 ();
 sg13g2_fill_1 FILLER_37_519 ();
 sg13g2_fill_1 FILLER_37_524 ();
 sg13g2_fill_1 FILLER_37_530 ();
 sg13g2_fill_2 FILLER_37_543 ();
 sg13g2_fill_1 FILLER_37_545 ();
 sg13g2_fill_1 FILLER_37_580 ();
 sg13g2_fill_1 FILLER_37_595 ();
 sg13g2_fill_2 FILLER_37_600 ();
 sg13g2_fill_2 FILLER_37_609 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_fill_1 FILLER_37_623 ();
 sg13g2_fill_2 FILLER_37_652 ();
 sg13g2_fill_2 FILLER_37_691 ();
 sg13g2_fill_1 FILLER_37_698 ();
 sg13g2_fill_1 FILLER_37_716 ();
 sg13g2_fill_1 FILLER_37_722 ();
 sg13g2_fill_1 FILLER_37_727 ();
 sg13g2_fill_1 FILLER_37_733 ();
 sg13g2_fill_1 FILLER_37_739 ();
 sg13g2_decap_4 FILLER_37_761 ();
 sg13g2_fill_1 FILLER_37_765 ();
 sg13g2_fill_1 FILLER_37_780 ();
 sg13g2_fill_1 FILLER_37_786 ();
 sg13g2_fill_1 FILLER_37_792 ();
 sg13g2_fill_2 FILLER_37_802 ();
 sg13g2_fill_1 FILLER_37_804 ();
 sg13g2_fill_2 FILLER_37_809 ();
 sg13g2_fill_1 FILLER_37_811 ();
 sg13g2_fill_1 FILLER_37_830 ();
 sg13g2_fill_2 FILLER_37_835 ();
 sg13g2_fill_1 FILLER_37_841 ();
 sg13g2_fill_2 FILLER_37_850 ();
 sg13g2_fill_2 FILLER_37_857 ();
 sg13g2_decap_8 FILLER_37_863 ();
 sg13g2_decap_4 FILLER_37_893 ();
 sg13g2_fill_1 FILLER_37_897 ();
 sg13g2_fill_1 FILLER_37_903 ();
 sg13g2_fill_2 FILLER_37_939 ();
 sg13g2_fill_1 FILLER_37_941 ();
 sg13g2_fill_2 FILLER_37_947 ();
 sg13g2_fill_1 FILLER_37_975 ();
 sg13g2_fill_2 FILLER_37_1002 ();
 sg13g2_fill_1 FILLER_37_1004 ();
 sg13g2_fill_2 FILLER_37_1035 ();
 sg13g2_fill_1 FILLER_37_1041 ();
 sg13g2_decap_4 FILLER_37_1050 ();
 sg13g2_fill_2 FILLER_37_1097 ();
 sg13g2_fill_1 FILLER_37_1099 ();
 sg13g2_fill_1 FILLER_37_1104 ();
 sg13g2_fill_1 FILLER_37_1110 ();
 sg13g2_decap_4 FILLER_37_1115 ();
 sg13g2_fill_1 FILLER_37_1119 ();
 sg13g2_fill_1 FILLER_37_1129 ();
 sg13g2_fill_2 FILLER_37_1135 ();
 sg13g2_fill_1 FILLER_37_1137 ();
 sg13g2_fill_1 FILLER_37_1176 ();
 sg13g2_fill_2 FILLER_37_1182 ();
 sg13g2_fill_1 FILLER_37_1223 ();
 sg13g2_fill_2 FILLER_37_1246 ();
 sg13g2_fill_1 FILLER_37_1252 ();
 sg13g2_fill_2 FILLER_37_1257 ();
 sg13g2_fill_1 FILLER_37_1276 ();
 sg13g2_fill_1 FILLER_37_1282 ();
 sg13g2_fill_2 FILLER_37_1287 ();
 sg13g2_fill_2 FILLER_37_1293 ();
 sg13g2_fill_1 FILLER_37_1299 ();
 sg13g2_fill_1 FILLER_37_1304 ();
 sg13g2_fill_1 FILLER_37_1312 ();
 sg13g2_fill_1 FILLER_37_1317 ();
 sg13g2_fill_2 FILLER_37_1325 ();
 sg13g2_fill_1 FILLER_37_1327 ();
 sg13g2_fill_1 FILLER_37_1359 ();
 sg13g2_fill_1 FILLER_37_1364 ();
 sg13g2_fill_1 FILLER_37_1395 ();
 sg13g2_decap_4 FILLER_37_1401 ();
 sg13g2_fill_2 FILLER_37_1405 ();
 sg13g2_fill_2 FILLER_37_1436 ();
 sg13g2_fill_1 FILLER_37_1443 ();
 sg13g2_fill_2 FILLER_37_1460 ();
 sg13g2_fill_1 FILLER_37_1477 ();
 sg13g2_fill_1 FILLER_37_1488 ();
 sg13g2_fill_1 FILLER_37_1492 ();
 sg13g2_decap_8 FILLER_37_1509 ();
 sg13g2_decap_4 FILLER_37_1516 ();
 sg13g2_decap_8 FILLER_37_1545 ();
 sg13g2_fill_1 FILLER_37_1552 ();
 sg13g2_decap_8 FILLER_37_1571 ();
 sg13g2_decap_8 FILLER_37_1578 ();
 sg13g2_decap_8 FILLER_37_1585 ();
 sg13g2_fill_1 FILLER_37_1596 ();
 sg13g2_fill_1 FILLER_37_1638 ();
 sg13g2_fill_2 FILLER_37_1644 ();
 sg13g2_fill_1 FILLER_37_1650 ();
 sg13g2_fill_2 FILLER_37_1664 ();
 sg13g2_decap_8 FILLER_37_1670 ();
 sg13g2_decap_8 FILLER_37_1701 ();
 sg13g2_fill_1 FILLER_37_1708 ();
 sg13g2_fill_1 FILLER_37_1739 ();
 sg13g2_fill_1 FILLER_37_1748 ();
 sg13g2_fill_1 FILLER_37_1755 ();
 sg13g2_fill_1 FILLER_37_1766 ();
 sg13g2_fill_2 FILLER_37_1771 ();
 sg13g2_fill_1 FILLER_37_1773 ();
 sg13g2_fill_1 FILLER_38_3 ();
 sg13g2_fill_2 FILLER_38_47 ();
 sg13g2_fill_1 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_59 ();
 sg13g2_fill_2 FILLER_38_71 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_fill_1 FILLER_38_89 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_fill_2 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_378 ();
 sg13g2_fill_1 FILLER_38_409 ();
 sg13g2_fill_2 FILLER_38_414 ();
 sg13g2_fill_1 FILLER_38_416 ();
 sg13g2_fill_1 FILLER_38_459 ();
 sg13g2_fill_1 FILLER_38_478 ();
 sg13g2_decap_8 FILLER_38_494 ();
 sg13g2_fill_2 FILLER_38_501 ();
 sg13g2_fill_2 FILLER_38_524 ();
 sg13g2_decap_4 FILLER_38_530 ();
 sg13g2_fill_2 FILLER_38_534 ();
 sg13g2_fill_1 FILLER_38_540 ();
 sg13g2_fill_1 FILLER_38_545 ();
 sg13g2_fill_1 FILLER_38_554 ();
 sg13g2_fill_2 FILLER_38_590 ();
 sg13g2_fill_1 FILLER_38_597 ();
 sg13g2_decap_4 FILLER_38_613 ();
 sg13g2_fill_1 FILLER_38_617 ();
 sg13g2_fill_1 FILLER_38_651 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_fill_1 FILLER_38_672 ();
 sg13g2_fill_1 FILLER_38_677 ();
 sg13g2_fill_1 FILLER_38_683 ();
 sg13g2_fill_1 FILLER_38_687 ();
 sg13g2_fill_2 FILLER_38_703 ();
 sg13g2_decap_4 FILLER_38_710 ();
 sg13g2_decap_4 FILLER_38_718 ();
 sg13g2_fill_1 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_742 ();
 sg13g2_fill_1 FILLER_38_748 ();
 sg13g2_fill_1 FILLER_38_755 ();
 sg13g2_fill_1 FILLER_38_761 ();
 sg13g2_decap_4 FILLER_38_766 ();
 sg13g2_fill_1 FILLER_38_770 ();
 sg13g2_fill_1 FILLER_38_903 ();
 sg13g2_fill_2 FILLER_38_908 ();
 sg13g2_fill_1 FILLER_38_910 ();
 sg13g2_fill_2 FILLER_38_976 ();
 sg13g2_fill_2 FILLER_38_982 ();
 sg13g2_fill_2 FILLER_38_989 ();
 sg13g2_fill_1 FILLER_38_1004 ();
 sg13g2_fill_1 FILLER_38_1010 ();
 sg13g2_fill_1 FILLER_38_1015 ();
 sg13g2_fill_1 FILLER_38_1020 ();
 sg13g2_fill_1 FILLER_38_1030 ();
 sg13g2_fill_1 FILLER_38_1035 ();
 sg13g2_fill_2 FILLER_38_1040 ();
 sg13g2_fill_1 FILLER_38_1047 ();
 sg13g2_fill_2 FILLER_38_1065 ();
 sg13g2_fill_2 FILLER_38_1110 ();
 sg13g2_fill_1 FILLER_38_1112 ();
 sg13g2_fill_2 FILLER_38_1123 ();
 sg13g2_fill_2 FILLER_38_1142 ();
 sg13g2_fill_1 FILLER_38_1144 ();
 sg13g2_fill_2 FILLER_38_1149 ();
 sg13g2_fill_1 FILLER_38_1151 ();
 sg13g2_fill_2 FILLER_38_1173 ();
 sg13g2_fill_1 FILLER_38_1205 ();
 sg13g2_fill_1 FILLER_38_1210 ();
 sg13g2_fill_1 FILLER_38_1237 ();
 sg13g2_fill_1 FILLER_38_1264 ();
 sg13g2_fill_1 FILLER_38_1269 ();
 sg13g2_fill_1 FILLER_38_1275 ();
 sg13g2_fill_1 FILLER_38_1280 ();
 sg13g2_fill_1 FILLER_38_1285 ();
 sg13g2_fill_1 FILLER_38_1293 ();
 sg13g2_fill_2 FILLER_38_1298 ();
 sg13g2_fill_1 FILLER_38_1334 ();
 sg13g2_decap_4 FILLER_38_1370 ();
 sg13g2_fill_2 FILLER_38_1412 ();
 sg13g2_fill_2 FILLER_38_1423 ();
 sg13g2_fill_1 FILLER_38_1425 ();
 sg13g2_fill_2 FILLER_38_1441 ();
 sg13g2_fill_1 FILLER_38_1443 ();
 sg13g2_decap_8 FILLER_38_1456 ();
 sg13g2_fill_2 FILLER_38_1493 ();
 sg13g2_fill_2 FILLER_38_1523 ();
 sg13g2_fill_1 FILLER_38_1525 ();
 sg13g2_fill_2 FILLER_38_1539 ();
 sg13g2_fill_1 FILLER_38_1541 ();
 sg13g2_fill_1 FILLER_38_1546 ();
 sg13g2_decap_4 FILLER_38_1550 ();
 sg13g2_fill_1 FILLER_38_1554 ();
 sg13g2_decap_8 FILLER_38_1575 ();
 sg13g2_fill_2 FILLER_38_1582 ();
 sg13g2_decap_8 FILLER_38_1587 ();
 sg13g2_fill_1 FILLER_38_1594 ();
 sg13g2_fill_2 FILLER_38_1599 ();
 sg13g2_fill_1 FILLER_38_1620 ();
 sg13g2_fill_1 FILLER_38_1628 ();
 sg13g2_fill_1 FILLER_38_1633 ();
 sg13g2_fill_1 FILLER_38_1642 ();
 sg13g2_fill_1 FILLER_38_1651 ();
 sg13g2_fill_2 FILLER_38_1659 ();
 sg13g2_fill_2 FILLER_38_1682 ();
 sg13g2_decap_8 FILLER_38_1701 ();
 sg13g2_fill_2 FILLER_38_1708 ();
 sg13g2_decap_4 FILLER_38_1740 ();
 sg13g2_fill_1 FILLER_38_1744 ();
 sg13g2_fill_2 FILLER_38_1755 ();
 sg13g2_fill_1 FILLER_38_1757 ();
 sg13g2_decap_4 FILLER_38_1762 ();
 sg13g2_fill_1 FILLER_38_1766 ();
 sg13g2_fill_2 FILLER_38_1772 ();
 sg13g2_fill_2 FILLER_39_9 ();
 sg13g2_fill_1 FILLER_39_27 ();
 sg13g2_fill_1 FILLER_39_67 ();
 sg13g2_fill_2 FILLER_39_94 ();
 sg13g2_fill_1 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_152 ();
 sg13g2_fill_1 FILLER_39_158 ();
 sg13g2_fill_1 FILLER_39_164 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_decap_8 FILLER_39_184 ();
 sg13g2_fill_1 FILLER_39_191 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_fill_1 FILLER_39_215 ();
 sg13g2_decap_4 FILLER_39_242 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_312 ();
 sg13g2_fill_2 FILLER_39_358 ();
 sg13g2_fill_2 FILLER_39_391 ();
 sg13g2_fill_1 FILLER_39_393 ();
 sg13g2_decap_4 FILLER_39_402 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_fill_2 FILLER_39_429 ();
 sg13g2_fill_1 FILLER_39_482 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_fill_2 FILLER_39_506 ();
 sg13g2_decap_8 FILLER_39_563 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_fill_1 FILLER_39_581 ();
 sg13g2_fill_1 FILLER_39_587 ();
 sg13g2_fill_2 FILLER_39_592 ();
 sg13g2_fill_1 FILLER_39_594 ();
 sg13g2_fill_2 FILLER_39_604 ();
 sg13g2_fill_1 FILLER_39_606 ();
 sg13g2_fill_1 FILLER_39_624 ();
 sg13g2_fill_1 FILLER_39_629 ();
 sg13g2_fill_1 FILLER_39_665 ();
 sg13g2_decap_4 FILLER_39_682 ();
 sg13g2_fill_1 FILLER_39_686 ();
 sg13g2_fill_1 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_fill_2 FILLER_39_721 ();
 sg13g2_fill_1 FILLER_39_727 ();
 sg13g2_fill_1 FILLER_39_733 ();
 sg13g2_decap_4 FILLER_39_738 ();
 sg13g2_fill_2 FILLER_39_742 ();
 sg13g2_fill_2 FILLER_39_748 ();
 sg13g2_fill_1 FILLER_39_762 ();
 sg13g2_fill_1 FILLER_39_767 ();
 sg13g2_fill_2 FILLER_39_794 ();
 sg13g2_fill_1 FILLER_39_796 ();
 sg13g2_fill_2 FILLER_39_814 ();
 sg13g2_fill_1 FILLER_39_816 ();
 sg13g2_decap_4 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_843 ();
 sg13g2_fill_2 FILLER_39_867 ();
 sg13g2_fill_1 FILLER_39_869 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_fill_2 FILLER_39_934 ();
 sg13g2_fill_1 FILLER_39_936 ();
 sg13g2_fill_2 FILLER_39_947 ();
 sg13g2_fill_1 FILLER_39_949 ();
 sg13g2_fill_1 FILLER_39_994 ();
 sg13g2_fill_1 FILLER_39_1031 ();
 sg13g2_decap_4 FILLER_39_1042 ();
 sg13g2_fill_1 FILLER_39_1046 ();
 sg13g2_fill_2 FILLER_39_1060 ();
 sg13g2_fill_2 FILLER_39_1076 ();
 sg13g2_fill_1 FILLER_39_1087 ();
 sg13g2_fill_2 FILLER_39_1092 ();
 sg13g2_fill_1 FILLER_39_1099 ();
 sg13g2_fill_2 FILLER_39_1118 ();
 sg13g2_fill_2 FILLER_39_1129 ();
 sg13g2_fill_1 FILLER_39_1159 ();
 sg13g2_fill_2 FILLER_39_1195 ();
 sg13g2_fill_2 FILLER_39_1232 ();
 sg13g2_fill_1 FILLER_39_1234 ();
 sg13g2_decap_4 FILLER_39_1239 ();
 sg13g2_decap_8 FILLER_39_1256 ();
 sg13g2_decap_4 FILLER_39_1263 ();
 sg13g2_fill_2 FILLER_39_1267 ();
 sg13g2_fill_2 FILLER_39_1309 ();
 sg13g2_fill_1 FILLER_39_1315 ();
 sg13g2_fill_1 FILLER_39_1354 ();
 sg13g2_fill_1 FILLER_39_1368 ();
 sg13g2_fill_1 FILLER_39_1374 ();
 sg13g2_fill_1 FILLER_39_1380 ();
 sg13g2_fill_1 FILLER_39_1385 ();
 sg13g2_fill_2 FILLER_39_1390 ();
 sg13g2_fill_2 FILLER_39_1445 ();
 sg13g2_fill_1 FILLER_39_1447 ();
 sg13g2_fill_1 FILLER_39_1463 ();
 sg13g2_fill_2 FILLER_39_1469 ();
 sg13g2_decap_8 FILLER_39_1489 ();
 sg13g2_decap_4 FILLER_39_1496 ();
 sg13g2_decap_8 FILLER_39_1509 ();
 sg13g2_fill_2 FILLER_39_1516 ();
 sg13g2_fill_1 FILLER_39_1518 ();
 sg13g2_fill_1 FILLER_39_1527 ();
 sg13g2_fill_2 FILLER_39_1540 ();
 sg13g2_fill_1 FILLER_39_1598 ();
 sg13g2_fill_1 FILLER_39_1603 ();
 sg13g2_fill_1 FILLER_39_1608 ();
 sg13g2_fill_2 FILLER_39_1616 ();
 sg13g2_fill_2 FILLER_39_1624 ();
 sg13g2_fill_1 FILLER_39_1634 ();
 sg13g2_fill_2 FILLER_39_1657 ();
 sg13g2_fill_1 FILLER_39_1667 ();
 sg13g2_fill_1 FILLER_39_1673 ();
 sg13g2_decap_4 FILLER_39_1694 ();
 sg13g2_decap_8 FILLER_39_1702 ();
 sg13g2_decap_4 FILLER_39_1709 ();
 sg13g2_fill_1 FILLER_39_1729 ();
 sg13g2_decap_8 FILLER_39_1767 ();
 sg13g2_fill_2 FILLER_40_57 ();
 sg13g2_fill_2 FILLER_40_64 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_fill_2 FILLER_40_170 ();
 sg13g2_fill_1 FILLER_40_203 ();
 sg13g2_fill_2 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_211 ();
 sg13g2_fill_1 FILLER_40_252 ();
 sg13g2_fill_1 FILLER_40_258 ();
 sg13g2_fill_2 FILLER_40_263 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_decap_4 FILLER_40_341 ();
 sg13g2_fill_1 FILLER_40_345 ();
 sg13g2_fill_1 FILLER_40_354 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_fill_1 FILLER_40_390 ();
 sg13g2_fill_1 FILLER_40_421 ();
 sg13g2_fill_1 FILLER_40_448 ();
 sg13g2_fill_1 FILLER_40_453 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_fill_1 FILLER_40_467 ();
 sg13g2_decap_4 FILLER_40_472 ();
 sg13g2_fill_2 FILLER_40_476 ();
 sg13g2_fill_2 FILLER_40_485 ();
 sg13g2_fill_1 FILLER_40_487 ();
 sg13g2_fill_1 FILLER_40_518 ();
 sg13g2_fill_2 FILLER_40_527 ();
 sg13g2_fill_2 FILLER_40_555 ();
 sg13g2_fill_1 FILLER_40_557 ();
 sg13g2_fill_2 FILLER_40_567 ();
 sg13g2_fill_1 FILLER_40_569 ();
 sg13g2_fill_1 FILLER_40_605 ();
 sg13g2_fill_1 FILLER_40_624 ();
 sg13g2_fill_2 FILLER_40_658 ();
 sg13g2_fill_1 FILLER_40_690 ();
 sg13g2_decap_4 FILLER_40_699 ();
 sg13g2_fill_1 FILLER_40_703 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_decap_4 FILLER_40_766 ();
 sg13g2_fill_2 FILLER_40_770 ();
 sg13g2_fill_1 FILLER_40_780 ();
 sg13g2_decap_8 FILLER_40_825 ();
 sg13g2_fill_1 FILLER_40_858 ();
 sg13g2_fill_1 FILLER_40_867 ();
 sg13g2_fill_1 FILLER_40_872 ();
 sg13g2_fill_1 FILLER_40_877 ();
 sg13g2_fill_1 FILLER_40_883 ();
 sg13g2_fill_2 FILLER_40_889 ();
 sg13g2_fill_2 FILLER_40_895 ();
 sg13g2_fill_1 FILLER_40_897 ();
 sg13g2_fill_1 FILLER_40_947 ();
 sg13g2_fill_1 FILLER_40_979 ();
 sg13g2_decap_8 FILLER_40_985 ();
 sg13g2_fill_1 FILLER_40_992 ();
 sg13g2_fill_1 FILLER_40_1009 ();
 sg13g2_decap_8 FILLER_40_1018 ();
 sg13g2_decap_4 FILLER_40_1025 ();
 sg13g2_fill_1 FILLER_40_1029 ();
 sg13g2_fill_1 FILLER_40_1048 ();
 sg13g2_fill_1 FILLER_40_1079 ();
 sg13g2_decap_8 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1094 ();
 sg13g2_decap_4 FILLER_40_1121 ();
 sg13g2_decap_4 FILLER_40_1159 ();
 sg13g2_fill_1 FILLER_40_1163 ();
 sg13g2_fill_2 FILLER_40_1270 ();
 sg13g2_fill_1 FILLER_40_1281 ();
 sg13g2_fill_1 FILLER_40_1322 ();
 sg13g2_fill_2 FILLER_40_1328 ();
 sg13g2_decap_4 FILLER_40_1390 ();
 sg13g2_decap_8 FILLER_40_1399 ();
 sg13g2_fill_1 FILLER_40_1406 ();
 sg13g2_fill_2 FILLER_40_1411 ();
 sg13g2_fill_1 FILLER_40_1413 ();
 sg13g2_fill_2 FILLER_40_1424 ();
 sg13g2_fill_1 FILLER_40_1426 ();
 sg13g2_decap_8 FILLER_40_1431 ();
 sg13g2_decap_8 FILLER_40_1438 ();
 sg13g2_decap_8 FILLER_40_1445 ();
 sg13g2_decap_4 FILLER_40_1452 ();
 sg13g2_fill_2 FILLER_40_1456 ();
 sg13g2_fill_1 FILLER_40_1482 ();
 sg13g2_fill_2 FILLER_40_1487 ();
 sg13g2_fill_1 FILLER_40_1494 ();
 sg13g2_fill_2 FILLER_40_1505 ();
 sg13g2_fill_1 FILLER_40_1507 ();
 sg13g2_decap_4 FILLER_40_1516 ();
 sg13g2_fill_1 FILLER_40_1525 ();
 sg13g2_decap_8 FILLER_40_1538 ();
 sg13g2_fill_1 FILLER_40_1545 ();
 sg13g2_fill_1 FILLER_40_1551 ();
 sg13g2_fill_1 FILLER_40_1556 ();
 sg13g2_fill_1 FILLER_40_1562 ();
 sg13g2_fill_1 FILLER_40_1568 ();
 sg13g2_fill_1 FILLER_40_1584 ();
 sg13g2_fill_1 FILLER_40_1590 ();
 sg13g2_fill_1 FILLER_40_1601 ();
 sg13g2_fill_2 FILLER_40_1628 ();
 sg13g2_fill_1 FILLER_40_1630 ();
 sg13g2_fill_2 FILLER_40_1661 ();
 sg13g2_decap_8 FILLER_40_1688 ();
 sg13g2_fill_2 FILLER_40_1700 ();
 sg13g2_decap_8 FILLER_40_1710 ();
 sg13g2_fill_2 FILLER_40_1721 ();
 sg13g2_fill_1 FILLER_40_1723 ();
 sg13g2_decap_4 FILLER_40_1754 ();
 sg13g2_fill_2 FILLER_40_1771 ();
 sg13g2_fill_1 FILLER_40_1773 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_fill_2 FILLER_41_110 ();
 sg13g2_fill_1 FILLER_41_116 ();
 sg13g2_fill_1 FILLER_41_122 ();
 sg13g2_fill_1 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_fill_1 FILLER_41_228 ();
 sg13g2_fill_1 FILLER_41_233 ();
 sg13g2_fill_1 FILLER_41_260 ();
 sg13g2_fill_1 FILLER_41_266 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_1 FILLER_41_302 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_fill_2 FILLER_41_313 ();
 sg13g2_fill_2 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_372 ();
 sg13g2_decap_4 FILLER_41_379 ();
 sg13g2_fill_2 FILLER_41_401 ();
 sg13g2_decap_4 FILLER_41_419 ();
 sg13g2_fill_1 FILLER_41_437 ();
 sg13g2_decap_4 FILLER_41_468 ();
 sg13g2_fill_2 FILLER_41_472 ();
 sg13g2_decap_4 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_507 ();
 sg13g2_fill_2 FILLER_41_513 ();
 sg13g2_fill_1 FILLER_41_531 ();
 sg13g2_fill_1 FILLER_41_546 ();
 sg13g2_fill_1 FILLER_41_554 ();
 sg13g2_fill_1 FILLER_41_565 ();
 sg13g2_fill_2 FILLER_41_575 ();
 sg13g2_fill_2 FILLER_41_581 ();
 sg13g2_decap_4 FILLER_41_621 ();
 sg13g2_fill_2 FILLER_41_630 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_681 ();
 sg13g2_fill_2 FILLER_41_708 ();
 sg13g2_fill_2 FILLER_41_714 ();
 sg13g2_fill_2 FILLER_41_720 ();
 sg13g2_fill_1 FILLER_41_722 ();
 sg13g2_fill_2 FILLER_41_740 ();
 sg13g2_fill_2 FILLER_41_750 ();
 sg13g2_fill_1 FILLER_41_766 ();
 sg13g2_fill_1 FILLER_41_793 ();
 sg13g2_fill_2 FILLER_41_798 ();
 sg13g2_fill_2 FILLER_41_830 ();
 sg13g2_decap_8 FILLER_41_836 ();
 sg13g2_fill_1 FILLER_41_843 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_fill_1 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_867 ();
 sg13g2_fill_1 FILLER_41_874 ();
 sg13g2_fill_1 FILLER_41_884 ();
 sg13g2_fill_1 FILLER_41_921 ();
 sg13g2_decap_4 FILLER_41_949 ();
 sg13g2_decap_4 FILLER_41_967 ();
 sg13g2_fill_1 FILLER_41_1068 ();
 sg13g2_decap_4 FILLER_41_1077 ();
 sg13g2_fill_2 FILLER_41_1093 ();
 sg13g2_fill_2 FILLER_41_1107 ();
 sg13g2_fill_1 FILLER_41_1114 ();
 sg13g2_decap_4 FILLER_41_1123 ();
 sg13g2_fill_2 FILLER_41_1136 ();
 sg13g2_fill_1 FILLER_41_1138 ();
 sg13g2_fill_2 FILLER_41_1198 ();
 sg13g2_fill_1 FILLER_41_1200 ();
 sg13g2_decap_4 FILLER_41_1205 ();
 sg13g2_fill_1 FILLER_41_1213 ();
 sg13g2_decap_4 FILLER_41_1219 ();
 sg13g2_fill_1 FILLER_41_1223 ();
 sg13g2_fill_2 FILLER_41_1228 ();
 sg13g2_fill_1 FILLER_41_1242 ();
 sg13g2_fill_1 FILLER_41_1248 ();
 sg13g2_decap_4 FILLER_41_1253 ();
 sg13g2_decap_8 FILLER_41_1291 ();
 sg13g2_decap_4 FILLER_41_1298 ();
 sg13g2_fill_2 FILLER_41_1302 ();
 sg13g2_fill_2 FILLER_41_1308 ();
 sg13g2_decap_4 FILLER_41_1315 ();
 sg13g2_fill_1 FILLER_41_1323 ();
 sg13g2_fill_1 FILLER_41_1341 ();
 sg13g2_decap_8 FILLER_41_1346 ();
 sg13g2_decap_8 FILLER_41_1353 ();
 sg13g2_decap_8 FILLER_41_1360 ();
 sg13g2_fill_2 FILLER_41_1367 ();
 sg13g2_fill_1 FILLER_41_1409 ();
 sg13g2_fill_1 FILLER_41_1424 ();
 sg13g2_fill_1 FILLER_41_1451 ();
 sg13g2_decap_8 FILLER_41_1457 ();
 sg13g2_fill_1 FILLER_41_1464 ();
 sg13g2_fill_1 FILLER_41_1484 ();
 sg13g2_fill_1 FILLER_41_1490 ();
 sg13g2_fill_1 FILLER_41_1502 ();
 sg13g2_fill_2 FILLER_41_1508 ();
 sg13g2_fill_1 FILLER_41_1522 ();
 sg13g2_fill_2 FILLER_41_1528 ();
 sg13g2_fill_1 FILLER_41_1530 ();
 sg13g2_fill_1 FILLER_41_1540 ();
 sg13g2_fill_1 FILLER_41_1556 ();
 sg13g2_fill_1 FILLER_41_1562 ();
 sg13g2_fill_1 FILLER_41_1570 ();
 sg13g2_fill_1 FILLER_41_1577 ();
 sg13g2_fill_1 FILLER_41_1585 ();
 sg13g2_fill_1 FILLER_41_1593 ();
 sg13g2_fill_2 FILLER_41_1599 ();
 sg13g2_decap_8 FILLER_41_1606 ();
 sg13g2_fill_2 FILLER_41_1613 ();
 sg13g2_fill_2 FILLER_41_1619 ();
 sg13g2_fill_2 FILLER_41_1626 ();
 sg13g2_fill_1 FILLER_41_1628 ();
 sg13g2_decap_4 FILLER_41_1633 ();
 sg13g2_fill_2 FILLER_41_1637 ();
 sg13g2_fill_2 FILLER_41_1651 ();
 sg13g2_decap_4 FILLER_41_1657 ();
 sg13g2_fill_2 FILLER_41_1669 ();
 sg13g2_decap_4 FILLER_41_1686 ();
 sg13g2_fill_1 FILLER_41_1690 ();
 sg13g2_fill_2 FILLER_41_1712 ();
 sg13g2_fill_1 FILLER_41_1714 ();
 sg13g2_fill_2 FILLER_41_1731 ();
 sg13g2_fill_1 FILLER_41_1733 ();
 sg13g2_fill_2 FILLER_41_1739 ();
 sg13g2_fill_2 FILLER_41_1750 ();
 sg13g2_decap_4 FILLER_41_1756 ();
 sg13g2_decap_4 FILLER_41_1768 ();
 sg13g2_fill_2 FILLER_41_1772 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_27 ();
 sg13g2_fill_1 FILLER_42_33 ();
 sg13g2_fill_1 FILLER_42_42 ();
 sg13g2_fill_2 FILLER_42_51 ();
 sg13g2_fill_1 FILLER_42_88 ();
 sg13g2_fill_2 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_186 ();
 sg13g2_fill_1 FILLER_42_191 ();
 sg13g2_fill_1 FILLER_42_201 ();
 sg13g2_fill_1 FILLER_42_206 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_1 FILLER_42_216 ();
 sg13g2_fill_2 FILLER_42_221 ();
 sg13g2_fill_1 FILLER_42_254 ();
 sg13g2_fill_2 FILLER_42_260 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_283 ();
 sg13g2_decap_4 FILLER_42_290 ();
 sg13g2_decap_4 FILLER_42_333 ();
 sg13g2_decap_4 FILLER_42_349 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_decap_8 FILLER_42_373 ();
 sg13g2_decap_4 FILLER_42_380 ();
 sg13g2_fill_2 FILLER_42_384 ();
 sg13g2_fill_1 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_438 ();
 sg13g2_fill_2 FILLER_42_449 ();
 sg13g2_fill_1 FILLER_42_451 ();
 sg13g2_fill_1 FILLER_42_458 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_472 ();
 sg13g2_fill_1 FILLER_42_478 ();
 sg13g2_fill_2 FILLER_42_484 ();
 sg13g2_fill_1 FILLER_42_509 ();
 sg13g2_fill_1 FILLER_42_555 ();
 sg13g2_fill_2 FILLER_42_561 ();
 sg13g2_fill_1 FILLER_42_563 ();
 sg13g2_fill_2 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_601 ();
 sg13g2_decap_4 FILLER_42_608 ();
 sg13g2_fill_1 FILLER_42_612 ();
 sg13g2_decap_8 FILLER_42_622 ();
 sg13g2_fill_2 FILLER_42_629 ();
 sg13g2_decap_4 FILLER_42_636 ();
 sg13g2_fill_1 FILLER_42_640 ();
 sg13g2_fill_2 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_690 ();
 sg13g2_fill_2 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_759 ();
 sg13g2_decap_8 FILLER_42_766 ();
 sg13g2_fill_2 FILLER_42_773 ();
 sg13g2_fill_1 FILLER_42_779 ();
 sg13g2_fill_1 FILLER_42_814 ();
 sg13g2_fill_1 FILLER_42_825 ();
 sg13g2_fill_1 FILLER_42_852 ();
 sg13g2_fill_1 FILLER_42_863 ();
 sg13g2_decap_4 FILLER_42_869 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_fill_2 FILLER_42_885 ();
 sg13g2_fill_1 FILLER_42_887 ();
 sg13g2_fill_1 FILLER_42_892 ();
 sg13g2_decap_4 FILLER_42_902 ();
 sg13g2_fill_2 FILLER_42_936 ();
 sg13g2_fill_1 FILLER_42_979 ();
 sg13g2_decap_8 FILLER_42_989 ();
 sg13g2_fill_2 FILLER_42_996 ();
 sg13g2_decap_4 FILLER_42_1001 ();
 sg13g2_decap_4 FILLER_42_1028 ();
 sg13g2_fill_2 FILLER_42_1049 ();
 sg13g2_fill_1 FILLER_42_1051 ();
 sg13g2_fill_2 FILLER_42_1056 ();
 sg13g2_fill_1 FILLER_42_1058 ();
 sg13g2_fill_2 FILLER_42_1076 ();
 sg13g2_fill_1 FILLER_42_1078 ();
 sg13g2_fill_1 FILLER_42_1087 ();
 sg13g2_fill_1 FILLER_42_1093 ();
 sg13g2_fill_1 FILLER_42_1109 ();
 sg13g2_fill_2 FILLER_42_1119 ();
 sg13g2_fill_1 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1152 ();
 sg13g2_fill_2 FILLER_42_1159 ();
 sg13g2_fill_2 FILLER_42_1165 ();
 sg13g2_fill_1 FILLER_42_1171 ();
 sg13g2_decap_4 FILLER_42_1249 ();
 sg13g2_fill_2 FILLER_42_1253 ();
 sg13g2_fill_2 FILLER_42_1267 ();
 sg13g2_fill_1 FILLER_42_1269 ();
 sg13g2_fill_1 FILLER_42_1301 ();
 sg13g2_fill_1 FILLER_42_1306 ();
 sg13g2_decap_4 FILLER_42_1315 ();
 sg13g2_fill_1 FILLER_42_1319 ();
 sg13g2_fill_2 FILLER_42_1331 ();
 sg13g2_decap_8 FILLER_42_1376 ();
 sg13g2_fill_1 FILLER_42_1383 ();
 sg13g2_decap_4 FILLER_42_1392 ();
 sg13g2_fill_2 FILLER_42_1396 ();
 sg13g2_fill_2 FILLER_42_1427 ();
 sg13g2_decap_4 FILLER_42_1460 ();
 sg13g2_fill_1 FILLER_42_1464 ();
 sg13g2_decap_8 FILLER_42_1479 ();
 sg13g2_fill_2 FILLER_42_1520 ();
 sg13g2_fill_1 FILLER_42_1526 ();
 sg13g2_decap_8 FILLER_42_1549 ();
 sg13g2_decap_4 FILLER_42_1568 ();
 sg13g2_decap_8 FILLER_42_1576 ();
 sg13g2_fill_1 FILLER_42_1621 ();
 sg13g2_fill_2 FILLER_42_1635 ();
 sg13g2_fill_1 FILLER_42_1658 ();
 sg13g2_decap_8 FILLER_42_1667 ();
 sg13g2_decap_8 FILLER_42_1674 ();
 sg13g2_fill_1 FILLER_42_1681 ();
 sg13g2_fill_1 FILLER_42_1723 ();
 sg13g2_fill_1 FILLER_42_1729 ();
 sg13g2_fill_2 FILLER_42_1735 ();
 sg13g2_fill_2 FILLER_42_1742 ();
 sg13g2_fill_1 FILLER_42_1744 ();
 sg13g2_decap_8 FILLER_42_1757 ();
 sg13g2_decap_8 FILLER_42_1764 ();
 sg13g2_fill_2 FILLER_42_1771 ();
 sg13g2_fill_1 FILLER_42_1773 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_14 ();
 sg13g2_fill_1 FILLER_43_30 ();
 sg13g2_fill_1 FILLER_43_42 ();
 sg13g2_fill_2 FILLER_43_68 ();
 sg13g2_fill_1 FILLER_43_75 ();
 sg13g2_fill_1 FILLER_43_85 ();
 sg13g2_fill_1 FILLER_43_90 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_1 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_123 ();
 sg13g2_fill_2 FILLER_43_218 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_2 FILLER_43_292 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_decap_8 FILLER_43_317 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_decap_4 FILLER_43_377 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_fill_1 FILLER_43_392 ();
 sg13g2_fill_1 FILLER_43_402 ();
 sg13g2_fill_2 FILLER_43_411 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_424 ();
 sg13g2_fill_1 FILLER_43_426 ();
 sg13g2_fill_2 FILLER_43_432 ();
 sg13g2_fill_1 FILLER_43_434 ();
 sg13g2_fill_1 FILLER_43_465 ();
 sg13g2_fill_2 FILLER_43_469 ();
 sg13g2_fill_2 FILLER_43_500 ();
 sg13g2_fill_1 FILLER_43_502 ();
 sg13g2_fill_2 FILLER_43_511 ();
 sg13g2_fill_1 FILLER_43_513 ();
 sg13g2_fill_1 FILLER_43_523 ();
 sg13g2_decap_4 FILLER_43_528 ();
 sg13g2_fill_1 FILLER_43_532 ();
 sg13g2_fill_2 FILLER_43_537 ();
 sg13g2_decap_4 FILLER_43_544 ();
 sg13g2_fill_1 FILLER_43_552 ();
 sg13g2_fill_2 FILLER_43_557 ();
 sg13g2_fill_2 FILLER_43_567 ();
 sg13g2_fill_1 FILLER_43_569 ();
 sg13g2_fill_1 FILLER_43_579 ();
 sg13g2_fill_1 FILLER_43_584 ();
 sg13g2_decap_4 FILLER_43_590 ();
 sg13g2_fill_1 FILLER_43_594 ();
 sg13g2_decap_4 FILLER_43_676 ();
 sg13g2_fill_2 FILLER_43_703 ();
 sg13g2_fill_1 FILLER_43_705 ();
 sg13g2_decap_4 FILLER_43_750 ();
 sg13g2_fill_1 FILLER_43_754 ();
 sg13g2_fill_2 FILLER_43_780 ();
 sg13g2_fill_1 FILLER_43_789 ();
 sg13g2_fill_1 FILLER_43_794 ();
 sg13g2_fill_2 FILLER_43_799 ();
 sg13g2_fill_2 FILLER_43_811 ();
 sg13g2_fill_2 FILLER_43_818 ();
 sg13g2_fill_1 FILLER_43_825 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_decap_8 FILLER_43_849 ();
 sg13g2_fill_2 FILLER_43_856 ();
 sg13g2_fill_1 FILLER_43_895 ();
 sg13g2_fill_1 FILLER_43_908 ();
 sg13g2_fill_2 FILLER_43_922 ();
 sg13g2_fill_1 FILLER_43_924 ();
 sg13g2_fill_1 FILLER_43_930 ();
 sg13g2_fill_1 FILLER_43_935 ();
 sg13g2_fill_2 FILLER_43_941 ();
 sg13g2_fill_2 FILLER_43_947 ();
 sg13g2_fill_1 FILLER_43_949 ();
 sg13g2_fill_1 FILLER_43_954 ();
 sg13g2_fill_2 FILLER_43_959 ();
 sg13g2_fill_1 FILLER_43_966 ();
 sg13g2_fill_2 FILLER_43_971 ();
 sg13g2_fill_2 FILLER_43_981 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_fill_1 FILLER_43_1027 ();
 sg13g2_decap_4 FILLER_43_1069 ();
 sg13g2_fill_1 FILLER_43_1073 ();
 sg13g2_fill_2 FILLER_43_1094 ();
 sg13g2_decap_4 FILLER_43_1139 ();
 sg13g2_fill_1 FILLER_43_1151 ();
 sg13g2_fill_1 FILLER_43_1156 ();
 sg13g2_fill_1 FILLER_43_1168 ();
 sg13g2_fill_1 FILLER_43_1174 ();
 sg13g2_fill_1 FILLER_43_1180 ();
 sg13g2_fill_2 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1226 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_fill_2 FILLER_43_1272 ();
 sg13g2_fill_2 FILLER_43_1303 ();
 sg13g2_fill_1 FILLER_43_1305 ();
 sg13g2_decap_8 FILLER_43_1313 ();
 sg13g2_fill_1 FILLER_43_1338 ();
 sg13g2_fill_1 FILLER_43_1347 ();
 sg13g2_fill_1 FILLER_43_1352 ();
 sg13g2_fill_1 FILLER_43_1358 ();
 sg13g2_fill_1 FILLER_43_1366 ();
 sg13g2_fill_1 FILLER_43_1371 ();
 sg13g2_fill_1 FILLER_43_1408 ();
 sg13g2_fill_1 FILLER_43_1419 ();
 sg13g2_fill_1 FILLER_43_1424 ();
 sg13g2_fill_1 FILLER_43_1430 ();
 sg13g2_fill_2 FILLER_43_1440 ();
 sg13g2_fill_1 FILLER_43_1442 ();
 sg13g2_fill_2 FILLER_43_1447 ();
 sg13g2_fill_2 FILLER_43_1458 ();
 sg13g2_fill_1 FILLER_43_1460 ();
 sg13g2_decap_8 FILLER_43_1465 ();
 sg13g2_decap_8 FILLER_43_1472 ();
 sg13g2_decap_4 FILLER_43_1479 ();
 sg13g2_fill_1 FILLER_43_1483 ();
 sg13g2_fill_1 FILLER_43_1500 ();
 sg13g2_fill_2 FILLER_43_1515 ();
 sg13g2_decap_4 FILLER_43_1527 ();
 sg13g2_fill_1 FILLER_43_1540 ();
 sg13g2_fill_1 FILLER_43_1557 ();
 sg13g2_fill_1 FILLER_43_1587 ();
 sg13g2_decap_8 FILLER_43_1612 ();
 sg13g2_fill_1 FILLER_43_1619 ();
 sg13g2_fill_1 FILLER_43_1624 ();
 sg13g2_decap_8 FILLER_43_1630 ();
 sg13g2_fill_2 FILLER_43_1637 ();
 sg13g2_fill_1 FILLER_43_1644 ();
 sg13g2_fill_1 FILLER_43_1649 ();
 sg13g2_fill_1 FILLER_43_1653 ();
 sg13g2_fill_2 FILLER_43_1667 ();
 sg13g2_decap_4 FILLER_43_1674 ();
 sg13g2_fill_1 FILLER_43_1678 ();
 sg13g2_decap_8 FILLER_43_1689 ();
 sg13g2_decap_4 FILLER_43_1696 ();
 sg13g2_fill_2 FILLER_43_1700 ();
 sg13g2_fill_2 FILLER_43_1731 ();
 sg13g2_fill_1 FILLER_43_1741 ();
 sg13g2_decap_8 FILLER_43_1757 ();
 sg13g2_decap_8 FILLER_43_1764 ();
 sg13g2_fill_2 FILLER_43_1771 ();
 sg13g2_fill_1 FILLER_43_1773 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_60 ();
 sg13g2_fill_2 FILLER_44_118 ();
 sg13g2_fill_1 FILLER_44_172 ();
 sg13g2_fill_1 FILLER_44_177 ();
 sg13g2_fill_1 FILLER_44_182 ();
 sg13g2_fill_2 FILLER_44_188 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_fill_2 FILLER_44_221 ();
 sg13g2_fill_1 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_251 ();
 sg13g2_fill_1 FILLER_44_257 ();
 sg13g2_fill_2 FILLER_44_301 ();
 sg13g2_fill_1 FILLER_44_303 ();
 sg13g2_fill_1 FILLER_44_311 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_fill_1 FILLER_44_348 ();
 sg13g2_fill_2 FILLER_44_355 ();
 sg13g2_fill_2 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_373 ();
 sg13g2_decap_4 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_404 ();
 sg13g2_decap_4 FILLER_44_409 ();
 sg13g2_fill_1 FILLER_44_413 ();
 sg13g2_fill_2 FILLER_44_466 ();
 sg13g2_fill_1 FILLER_44_489 ();
 sg13g2_fill_2 FILLER_44_498 ();
 sg13g2_fill_1 FILLER_44_556 ();
 sg13g2_fill_1 FILLER_44_616 ();
 sg13g2_fill_2 FILLER_44_629 ();
 sg13g2_fill_1 FILLER_44_631 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_fill_1 FILLER_44_659 ();
 sg13g2_fill_2 FILLER_44_680 ();
 sg13g2_fill_1 FILLER_44_682 ();
 sg13g2_fill_2 FILLER_44_713 ();
 sg13g2_fill_2 FILLER_44_773 ();
 sg13g2_decap_4 FILLER_44_823 ();
 sg13g2_fill_2 FILLER_44_834 ();
 sg13g2_fill_1 FILLER_44_856 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_fill_2 FILLER_44_869 ();
 sg13g2_fill_1 FILLER_44_877 ();
 sg13g2_fill_2 FILLER_44_906 ();
 sg13g2_fill_1 FILLER_44_908 ();
 sg13g2_fill_2 FILLER_44_930 ();
 sg13g2_fill_1 FILLER_44_932 ();
 sg13g2_fill_2 FILLER_44_943 ();
 sg13g2_fill_1 FILLER_44_945 ();
 sg13g2_fill_2 FILLER_44_990 ();
 sg13g2_fill_1 FILLER_44_992 ();
 sg13g2_fill_2 FILLER_44_998 ();
 sg13g2_fill_1 FILLER_44_1000 ();
 sg13g2_fill_2 FILLER_44_1005 ();
 sg13g2_fill_1 FILLER_44_1007 ();
 sg13g2_fill_2 FILLER_44_1043 ();
 sg13g2_fill_2 FILLER_44_1054 ();
 sg13g2_fill_2 FILLER_44_1077 ();
 sg13g2_decap_8 FILLER_44_1083 ();
 sg13g2_fill_1 FILLER_44_1090 ();
 sg13g2_fill_1 FILLER_44_1117 ();
 sg13g2_fill_1 FILLER_44_1122 ();
 sg13g2_fill_1 FILLER_44_1149 ();
 sg13g2_fill_2 FILLER_44_1155 ();
 sg13g2_fill_1 FILLER_44_1195 ();
 sg13g2_fill_1 FILLER_44_1200 ();
 sg13g2_fill_1 FILLER_44_1214 ();
 sg13g2_fill_2 FILLER_44_1236 ();
 sg13g2_fill_1 FILLER_44_1238 ();
 sg13g2_fill_2 FILLER_44_1254 ();
 sg13g2_fill_1 FILLER_44_1256 ();
 sg13g2_fill_2 FILLER_44_1270 ();
 sg13g2_fill_2 FILLER_44_1280 ();
 sg13g2_fill_1 FILLER_44_1282 ();
 sg13g2_fill_1 FILLER_44_1295 ();
 sg13g2_fill_1 FILLER_44_1304 ();
 sg13g2_fill_2 FILLER_44_1331 ();
 sg13g2_fill_1 FILLER_44_1333 ();
 sg13g2_fill_2 FILLER_44_1351 ();
 sg13g2_fill_2 FILLER_44_1366 ();
 sg13g2_fill_1 FILLER_44_1368 ();
 sg13g2_fill_1 FILLER_44_1374 ();
 sg13g2_fill_2 FILLER_44_1387 ();
 sg13g2_fill_1 FILLER_44_1389 ();
 sg13g2_fill_2 FILLER_44_1411 ();
 sg13g2_fill_2 FILLER_44_1447 ();
 sg13g2_fill_1 FILLER_44_1449 ();
 sg13g2_fill_2 FILLER_44_1480 ();
 sg13g2_fill_1 FILLER_44_1482 ();
 sg13g2_decap_4 FILLER_44_1517 ();
 sg13g2_fill_1 FILLER_44_1521 ();
 sg13g2_fill_1 FILLER_44_1526 ();
 sg13g2_fill_1 FILLER_44_1531 ();
 sg13g2_fill_2 FILLER_44_1537 ();
 sg13g2_fill_1 FILLER_44_1539 ();
 sg13g2_decap_4 FILLER_44_1561 ();
 sg13g2_fill_1 FILLER_44_1565 ();
 sg13g2_fill_2 FILLER_44_1571 ();
 sg13g2_fill_1 FILLER_44_1573 ();
 sg13g2_fill_1 FILLER_44_1606 ();
 sg13g2_fill_2 FILLER_44_1615 ();
 sg13g2_fill_2 FILLER_44_1633 ();
 sg13g2_decap_8 FILLER_44_1658 ();
 sg13g2_fill_2 FILLER_44_1665 ();
 sg13g2_fill_1 FILLER_44_1667 ();
 sg13g2_fill_1 FILLER_44_1672 ();
 sg13g2_fill_1 FILLER_44_1678 ();
 sg13g2_fill_1 FILLER_44_1687 ();
 sg13g2_fill_1 FILLER_44_1697 ();
 sg13g2_fill_2 FILLER_44_1705 ();
 sg13g2_decap_4 FILLER_44_1717 ();
 sg13g2_fill_1 FILLER_44_1721 ();
 sg13g2_fill_2 FILLER_44_1725 ();
 sg13g2_decap_4 FILLER_44_1739 ();
 sg13g2_fill_1 FILLER_44_1743 ();
 sg13g2_decap_8 FILLER_44_1749 ();
 sg13g2_fill_1 FILLER_44_1756 ();
 sg13g2_fill_2 FILLER_44_1768 ();
 sg13g2_fill_1 FILLER_44_1773 ();
 sg13g2_fill_1 FILLER_45_15 ();
 sg13g2_fill_2 FILLER_45_20 ();
 sg13g2_fill_2 FILLER_45_27 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_fill_2 FILLER_45_43 ();
 sg13g2_fill_1 FILLER_45_49 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_1 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_80 ();
 sg13g2_fill_1 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_fill_2 FILLER_45_145 ();
 sg13g2_fill_2 FILLER_45_225 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_263 ();
 sg13g2_decap_4 FILLER_45_348 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_decap_8 FILLER_45_380 ();
 sg13g2_fill_2 FILLER_45_433 ();
 sg13g2_fill_1 FILLER_45_460 ();
 sg13g2_fill_1 FILLER_45_487 ();
 sg13g2_fill_1 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_501 ();
 sg13g2_fill_2 FILLER_45_510 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_523 ();
 sg13g2_fill_1 FILLER_45_530 ();
 sg13g2_fill_2 FILLER_45_535 ();
 sg13g2_fill_2 FILLER_45_551 ();
 sg13g2_fill_2 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_611 ();
 sg13g2_decap_4 FILLER_45_618 ();
 sg13g2_fill_2 FILLER_45_622 ();
 sg13g2_fill_1 FILLER_45_628 ();
 sg13g2_fill_1 FILLER_45_637 ();
 sg13g2_fill_2 FILLER_45_642 ();
 sg13g2_fill_1 FILLER_45_649 ();
 sg13g2_fill_2 FILLER_45_654 ();
 sg13g2_fill_2 FILLER_45_670 ();
 sg13g2_decap_8 FILLER_45_680 ();
 sg13g2_fill_2 FILLER_45_687 ();
 sg13g2_decap_4 FILLER_45_707 ();
 sg13g2_fill_2 FILLER_45_725 ();
 sg13g2_fill_1 FILLER_45_727 ();
 sg13g2_fill_1 FILLER_45_766 ();
 sg13g2_fill_2 FILLER_45_776 ();
 sg13g2_fill_1 FILLER_45_782 ();
 sg13g2_fill_2 FILLER_45_814 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_fill_2 FILLER_45_831 ();
 sg13g2_fill_1 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_863 ();
 sg13g2_decap_4 FILLER_45_870 ();
 sg13g2_fill_1 FILLER_45_879 ();
 sg13g2_fill_1 FILLER_45_906 ();
 sg13g2_fill_2 FILLER_45_912 ();
 sg13g2_fill_2 FILLER_45_990 ();
 sg13g2_fill_1 FILLER_45_1018 ();
 sg13g2_fill_1 FILLER_45_1034 ();
 sg13g2_fill_2 FILLER_45_1053 ();
 sg13g2_fill_2 FILLER_45_1065 ();
 sg13g2_fill_1 FILLER_45_1098 ();
 sg13g2_fill_1 FILLER_45_1122 ();
 sg13g2_fill_1 FILLER_45_1128 ();
 sg13g2_fill_1 FILLER_45_1137 ();
 sg13g2_fill_1 FILLER_45_1143 ();
 sg13g2_fill_2 FILLER_45_1149 ();
 sg13g2_fill_1 FILLER_45_1161 ();
 sg13g2_fill_2 FILLER_45_1168 ();
 sg13g2_fill_2 FILLER_45_1204 ();
 sg13g2_fill_2 FILLER_45_1247 ();
 sg13g2_fill_1 FILLER_45_1249 ();
 sg13g2_fill_1 FILLER_45_1266 ();
 sg13g2_fill_1 FILLER_45_1274 ();
 sg13g2_fill_2 FILLER_45_1288 ();
 sg13g2_fill_1 FILLER_45_1295 ();
 sg13g2_fill_1 FILLER_45_1341 ();
 sg13g2_fill_1 FILLER_45_1363 ();
 sg13g2_fill_1 FILLER_45_1390 ();
 sg13g2_fill_2 FILLER_45_1448 ();
 sg13g2_fill_1 FILLER_45_1450 ();
 sg13g2_decap_4 FILLER_45_1461 ();
 sg13g2_decap_8 FILLER_45_1469 ();
 sg13g2_decap_8 FILLER_45_1476 ();
 sg13g2_fill_2 FILLER_45_1494 ();
 sg13g2_fill_1 FILLER_45_1523 ();
 sg13g2_fill_2 FILLER_45_1545 ();
 sg13g2_fill_2 FILLER_45_1552 ();
 sg13g2_decap_8 FILLER_45_1558 ();
 sg13g2_fill_2 FILLER_45_1565 ();
 sg13g2_fill_1 FILLER_45_1567 ();
 sg13g2_fill_2 FILLER_45_1576 ();
 sg13g2_decap_8 FILLER_45_1599 ();
 sg13g2_decap_8 FILLER_45_1606 ();
 sg13g2_decap_4 FILLER_45_1613 ();
 sg13g2_fill_2 FILLER_45_1617 ();
 sg13g2_decap_4 FILLER_45_1632 ();
 sg13g2_fill_1 FILLER_45_1636 ();
 sg13g2_decap_8 FILLER_45_1651 ();
 sg13g2_fill_2 FILLER_45_1658 ();
 sg13g2_fill_1 FILLER_45_1660 ();
 sg13g2_fill_1 FILLER_45_1687 ();
 sg13g2_fill_1 FILLER_45_1696 ();
 sg13g2_fill_1 FILLER_45_1702 ();
 sg13g2_fill_1 FILLER_45_1708 ();
 sg13g2_decap_4 FILLER_45_1713 ();
 sg13g2_fill_2 FILLER_45_1717 ();
 sg13g2_decap_8 FILLER_45_1731 ();
 sg13g2_decap_8 FILLER_45_1738 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_27 ();
 sg13g2_fill_1 FILLER_46_36 ();
 sg13g2_fill_2 FILLER_46_48 ();
 sg13g2_fill_2 FILLER_46_75 ();
 sg13g2_fill_1 FILLER_46_103 ();
 sg13g2_fill_2 FILLER_46_161 ();
 sg13g2_fill_2 FILLER_46_229 ();
 sg13g2_fill_1 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_244 ();
 sg13g2_fill_2 FILLER_46_272 ();
 sg13g2_fill_1 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_353 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_fill_2 FILLER_46_377 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_decap_4 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_388 ();
 sg13g2_fill_2 FILLER_46_403 ();
 sg13g2_fill_1 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_46_411 ();
 sg13g2_fill_2 FILLER_46_432 ();
 sg13g2_fill_2 FILLER_46_453 ();
 sg13g2_fill_1 FILLER_46_473 ();
 sg13g2_fill_2 FILLER_46_484 ();
 sg13g2_fill_1 FILLER_46_486 ();
 sg13g2_decap_8 FILLER_46_502 ();
 sg13g2_decap_4 FILLER_46_509 ();
 sg13g2_decap_8 FILLER_46_524 ();
 sg13g2_fill_1 FILLER_46_557 ();
 sg13g2_fill_2 FILLER_46_585 ();
 sg13g2_fill_1 FILLER_46_617 ();
 sg13g2_fill_1 FILLER_46_649 ();
 sg13g2_fill_2 FILLER_46_682 ();
 sg13g2_fill_2 FILLER_46_688 ();
 sg13g2_fill_1 FILLER_46_703 ();
 sg13g2_fill_2 FILLER_46_753 ();
 sg13g2_fill_1 FILLER_46_766 ();
 sg13g2_fill_2 FILLER_46_793 ();
 sg13g2_fill_1 FILLER_46_799 ();
 sg13g2_fill_2 FILLER_46_816 ();
 sg13g2_fill_1 FILLER_46_818 ();
 sg13g2_fill_1 FILLER_46_824 ();
 sg13g2_fill_2 FILLER_46_832 ();
 sg13g2_fill_1 FILLER_46_842 ();
 sg13g2_fill_2 FILLER_46_855 ();
 sg13g2_fill_1 FILLER_46_857 ();
 sg13g2_fill_1 FILLER_46_862 ();
 sg13g2_fill_2 FILLER_46_892 ();
 sg13g2_fill_1 FILLER_46_898 ();
 sg13g2_fill_1 FILLER_46_903 ();
 sg13g2_fill_1 FILLER_46_908 ();
 sg13g2_fill_2 FILLER_46_913 ();
 sg13g2_fill_2 FILLER_46_919 ();
 sg13g2_fill_2 FILLER_46_925 ();
 sg13g2_fill_2 FILLER_46_948 ();
 sg13g2_fill_1 FILLER_46_950 ();
 sg13g2_fill_1 FILLER_46_960 ();
 sg13g2_fill_2 FILLER_46_970 ();
 sg13g2_fill_1 FILLER_46_982 ();
 sg13g2_fill_1 FILLER_46_1002 ();
 sg13g2_fill_1 FILLER_46_1011 ();
 sg13g2_fill_1 FILLER_46_1016 ();
 sg13g2_fill_2 FILLER_46_1043 ();
 sg13g2_fill_1 FILLER_46_1049 ();
 sg13g2_fill_2 FILLER_46_1058 ();
 sg13g2_fill_1 FILLER_46_1064 ();
 sg13g2_decap_8 FILLER_46_1075 ();
 sg13g2_decap_4 FILLER_46_1082 ();
 sg13g2_fill_2 FILLER_46_1086 ();
 sg13g2_fill_1 FILLER_46_1092 ();
 sg13g2_fill_2 FILLER_46_1101 ();
 sg13g2_fill_1 FILLER_46_1103 ();
 sg13g2_fill_1 FILLER_46_1107 ();
 sg13g2_fill_1 FILLER_46_1113 ();
 sg13g2_fill_1 FILLER_46_1122 ();
 sg13g2_fill_2 FILLER_46_1130 ();
 sg13g2_fill_1 FILLER_46_1201 ();
 sg13g2_fill_1 FILLER_46_1207 ();
 sg13g2_fill_1 FILLER_46_1215 ();
 sg13g2_fill_1 FILLER_46_1221 ();
 sg13g2_fill_1 FILLER_46_1227 ();
 sg13g2_fill_2 FILLER_46_1235 ();
 sg13g2_fill_1 FILLER_46_1253 ();
 sg13g2_fill_2 FILLER_46_1285 ();
 sg13g2_decap_8 FILLER_46_1294 ();
 sg13g2_decap_8 FILLER_46_1301 ();
 sg13g2_fill_1 FILLER_46_1313 ();
 sg13g2_fill_1 FILLER_46_1320 ();
 sg13g2_decap_4 FILLER_46_1357 ();
 sg13g2_decap_4 FILLER_46_1385 ();
 sg13g2_fill_2 FILLER_46_1389 ();
 sg13g2_decap_4 FILLER_46_1395 ();
 sg13g2_fill_2 FILLER_46_1399 ();
 sg13g2_fill_1 FILLER_46_1424 ();
 sg13g2_fill_1 FILLER_46_1457 ();
 sg13g2_decap_8 FILLER_46_1484 ();
 sg13g2_fill_2 FILLER_46_1491 ();
 sg13g2_fill_1 FILLER_46_1493 ();
 sg13g2_fill_1 FILLER_46_1505 ();
 sg13g2_decap_8 FILLER_46_1516 ();
 sg13g2_decap_8 FILLER_46_1523 ();
 sg13g2_fill_2 FILLER_46_1530 ();
 sg13g2_fill_1 FILLER_46_1532 ();
 sg13g2_decap_4 FILLER_46_1542 ();
 sg13g2_fill_1 FILLER_46_1546 ();
 sg13g2_decap_4 FILLER_46_1551 ();
 sg13g2_fill_1 FILLER_46_1555 ();
 sg13g2_decap_4 FILLER_46_1561 ();
 sg13g2_fill_2 FILLER_46_1565 ();
 sg13g2_decap_8 FILLER_46_1575 ();
 sg13g2_decap_8 FILLER_46_1582 ();
 sg13g2_decap_8 FILLER_46_1589 ();
 sg13g2_fill_1 FILLER_46_1600 ();
 sg13g2_fill_2 FILLER_46_1617 ();
 sg13g2_fill_2 FILLER_46_1635 ();
 sg13g2_fill_1 FILLER_46_1641 ();
 sg13g2_decap_8 FILLER_46_1650 ();
 sg13g2_fill_1 FILLER_46_1665 ();
 sg13g2_fill_1 FILLER_46_1670 ();
 sg13g2_fill_1 FILLER_46_1689 ();
 sg13g2_fill_1 FILLER_46_1694 ();
 sg13g2_fill_1 FILLER_46_1699 ();
 sg13g2_fill_1 FILLER_46_1705 ();
 sg13g2_decap_4 FILLER_46_1714 ();
 sg13g2_fill_2 FILLER_46_1718 ();
 sg13g2_fill_1 FILLER_46_1724 ();
 sg13g2_decap_8 FILLER_46_1748 ();
 sg13g2_fill_1 FILLER_46_1755 ();
 sg13g2_fill_1 FILLER_46_1765 ();
 sg13g2_fill_2 FILLER_46_1771 ();
 sg13g2_fill_1 FILLER_46_1773 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_46 ();
 sg13g2_fill_2 FILLER_47_62 ();
 sg13g2_fill_2 FILLER_47_81 ();
 sg13g2_fill_1 FILLER_47_92 ();
 sg13g2_fill_1 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_2 FILLER_47_291 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_331 ();
 sg13g2_fill_2 FILLER_47_336 ();
 sg13g2_fill_2 FILLER_47_368 ();
 sg13g2_fill_1 FILLER_47_405 ();
 sg13g2_fill_1 FILLER_47_432 ();
 sg13g2_fill_2 FILLER_47_497 ();
 sg13g2_fill_2 FILLER_47_507 ();
 sg13g2_fill_1 FILLER_47_509 ();
 sg13g2_fill_1 FILLER_47_518 ();
 sg13g2_fill_1 FILLER_47_523 ();
 sg13g2_fill_1 FILLER_47_554 ();
 sg13g2_fill_1 FILLER_47_559 ();
 sg13g2_fill_1 FILLER_47_586 ();
 sg13g2_fill_2 FILLER_47_605 ();
 sg13g2_fill_2 FILLER_47_616 ();
 sg13g2_fill_1 FILLER_47_618 ();
 sg13g2_fill_1 FILLER_47_623 ();
 sg13g2_fill_2 FILLER_47_659 ();
 sg13g2_fill_1 FILLER_47_666 ();
 sg13g2_fill_2 FILLER_47_703 ();
 sg13g2_fill_2 FILLER_47_713 ();
 sg13g2_fill_1 FILLER_47_735 ();
 sg13g2_fill_2 FILLER_47_752 ();
 sg13g2_fill_1 FILLER_47_761 ();
 sg13g2_fill_1 FILLER_47_774 ();
 sg13g2_fill_1 FILLER_47_815 ();
 sg13g2_decap_4 FILLER_47_824 ();
 sg13g2_fill_1 FILLER_47_828 ();
 sg13g2_decap_4 FILLER_47_833 ();
 sg13g2_decap_4 FILLER_47_868 ();
 sg13g2_fill_1 FILLER_47_872 ();
 sg13g2_fill_2 FILLER_47_881 ();
 sg13g2_fill_1 FILLER_47_907 ();
 sg13g2_fill_1 FILLER_47_912 ();
 sg13g2_fill_1 FILLER_47_918 ();
 sg13g2_fill_2 FILLER_47_927 ();
 sg13g2_fill_1 FILLER_47_929 ();
 sg13g2_decap_4 FILLER_47_934 ();
 sg13g2_fill_1 FILLER_47_947 ();
 sg13g2_fill_1 FILLER_47_954 ();
 sg13g2_fill_1 FILLER_47_967 ();
 sg13g2_fill_1 FILLER_47_1003 ();
 sg13g2_fill_1 FILLER_47_1017 ();
 sg13g2_fill_2 FILLER_47_1024 ();
 sg13g2_fill_2 FILLER_47_1030 ();
 sg13g2_fill_2 FILLER_47_1037 ();
 sg13g2_fill_2 FILLER_47_1042 ();
 sg13g2_fill_1 FILLER_47_1044 ();
 sg13g2_decap_4 FILLER_47_1049 ();
 sg13g2_fill_2 FILLER_47_1053 ();
 sg13g2_fill_2 FILLER_47_1059 ();
 sg13g2_fill_1 FILLER_47_1061 ();
 sg13g2_fill_2 FILLER_47_1066 ();
 sg13g2_fill_2 FILLER_47_1127 ();
 sg13g2_fill_2 FILLER_47_1235 ();
 sg13g2_fill_2 FILLER_47_1275 ();
 sg13g2_fill_1 FILLER_47_1277 ();
 sg13g2_fill_2 FILLER_47_1292 ();
 sg13g2_decap_4 FILLER_47_1303 ();
 sg13g2_fill_2 FILLER_47_1307 ();
 sg13g2_fill_2 FILLER_47_1336 ();
 sg13g2_fill_1 FILLER_47_1343 ();
 sg13g2_fill_1 FILLER_47_1350 ();
 sg13g2_fill_1 FILLER_47_1358 ();
 sg13g2_fill_2 FILLER_47_1363 ();
 sg13g2_fill_1 FILLER_47_1368 ();
 sg13g2_fill_1 FILLER_47_1375 ();
 sg13g2_fill_2 FILLER_47_1423 ();
 sg13g2_fill_2 FILLER_47_1449 ();
 sg13g2_decap_4 FILLER_47_1487 ();
 sg13g2_fill_1 FILLER_47_1491 ();
 sg13g2_fill_2 FILLER_47_1515 ();
 sg13g2_decap_4 FILLER_47_1525 ();
 sg13g2_fill_1 FILLER_47_1529 ();
 sg13g2_fill_2 FILLER_47_1560 ();
 sg13g2_fill_2 FILLER_47_1591 ();
 sg13g2_fill_1 FILLER_47_1593 ();
 sg13g2_fill_1 FILLER_47_1598 ();
 sg13g2_fill_1 FILLER_47_1607 ();
 sg13g2_fill_1 FILLER_47_1624 ();
 sg13g2_fill_1 FILLER_47_1630 ();
 sg13g2_fill_2 FILLER_47_1636 ();
 sg13g2_fill_2 FILLER_47_1642 ();
 sg13g2_fill_2 FILLER_47_1649 ();
 sg13g2_fill_2 FILLER_47_1656 ();
 sg13g2_fill_1 FILLER_47_1658 ();
 sg13g2_fill_2 FILLER_47_1663 ();
 sg13g2_fill_1 FILLER_47_1665 ();
 sg13g2_fill_2 FILLER_47_1670 ();
 sg13g2_fill_2 FILLER_47_1681 ();
 sg13g2_decap_8 FILLER_47_1686 ();
 sg13g2_fill_2 FILLER_47_1693 ();
 sg13g2_fill_2 FILLER_47_1703 ();
 sg13g2_fill_2 FILLER_47_1713 ();
 sg13g2_fill_1 FILLER_47_1715 ();
 sg13g2_fill_2 FILLER_47_1762 ();
 sg13g2_fill_2 FILLER_47_1772 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_11 ();
 sg13g2_fill_1 FILLER_48_38 ();
 sg13g2_fill_1 FILLER_48_67 ();
 sg13g2_fill_2 FILLER_48_94 ();
 sg13g2_fill_1 FILLER_48_122 ();
 sg13g2_fill_2 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_150 ();
 sg13g2_fill_1 FILLER_48_156 ();
 sg13g2_fill_1 FILLER_48_161 ();
 sg13g2_fill_2 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_248 ();
 sg13g2_fill_2 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_271 ();
 sg13g2_fill_1 FILLER_48_276 ();
 sg13g2_fill_1 FILLER_48_324 ();
 sg13g2_fill_2 FILLER_48_355 ();
 sg13g2_fill_1 FILLER_48_357 ();
 sg13g2_fill_2 FILLER_48_370 ();
 sg13g2_fill_1 FILLER_48_372 ();
 sg13g2_decap_4 FILLER_48_377 ();
 sg13g2_fill_2 FILLER_48_381 ();
 sg13g2_fill_2 FILLER_48_399 ();
 sg13g2_fill_1 FILLER_48_401 ();
 sg13g2_fill_2 FILLER_48_410 ();
 sg13g2_fill_1 FILLER_48_412 ();
 sg13g2_fill_1 FILLER_48_440 ();
 sg13g2_fill_1 FILLER_48_451 ();
 sg13g2_fill_1 FILLER_48_460 ();
 sg13g2_fill_1 FILLER_48_465 ();
 sg13g2_fill_2 FILLER_48_470 ();
 sg13g2_fill_1 FILLER_48_480 ();
 sg13g2_fill_1 FILLER_48_491 ();
 sg13g2_fill_2 FILLER_48_523 ();
 sg13g2_decap_8 FILLER_48_530 ();
 sg13g2_decap_4 FILLER_48_537 ();
 sg13g2_fill_1 FILLER_48_541 ();
 sg13g2_fill_1 FILLER_48_546 ();
 sg13g2_fill_1 FILLER_48_551 ();
 sg13g2_fill_1 FILLER_48_557 ();
 sg13g2_fill_2 FILLER_48_568 ();
 sg13g2_fill_1 FILLER_48_570 ();
 sg13g2_decap_4 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_618 ();
 sg13g2_fill_1 FILLER_48_637 ();
 sg13g2_fill_1 FILLER_48_667 ();
 sg13g2_fill_1 FILLER_48_674 ();
 sg13g2_fill_2 FILLER_48_686 ();
 sg13g2_fill_1 FILLER_48_700 ();
 sg13g2_fill_2 FILLER_48_720 ();
 sg13g2_fill_1 FILLER_48_743 ();
 sg13g2_fill_1 FILLER_48_748 ();
 sg13g2_fill_1 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_773 ();
 sg13g2_fill_2 FILLER_48_786 ();
 sg13g2_fill_2 FILLER_48_799 ();
 sg13g2_fill_1 FILLER_48_801 ();
 sg13g2_fill_1 FILLER_48_810 ();
 sg13g2_fill_2 FILLER_48_821 ();
 sg13g2_fill_1 FILLER_48_823 ();
 sg13g2_fill_2 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_831 ();
 sg13g2_fill_2 FILLER_48_889 ();
 sg13g2_fill_2 FILLER_48_895 ();
 sg13g2_fill_1 FILLER_48_897 ();
 sg13g2_fill_2 FILLER_48_901 ();
 sg13g2_fill_2 FILLER_48_908 ();
 sg13g2_fill_1 FILLER_48_910 ();
 sg13g2_fill_2 FILLER_48_941 ();
 sg13g2_fill_2 FILLER_48_965 ();
 sg13g2_fill_2 FILLER_48_971 ();
 sg13g2_fill_1 FILLER_48_973 ();
 sg13g2_fill_2 FILLER_48_1014 ();
 sg13g2_fill_2 FILLER_48_1021 ();
 sg13g2_fill_2 FILLER_48_1026 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_fill_1 FILLER_48_1064 ();
 sg13g2_fill_1 FILLER_48_1081 ();
 sg13g2_fill_2 FILLER_48_1086 ();
 sg13g2_fill_1 FILLER_48_1093 ();
 sg13g2_fill_2 FILLER_48_1099 ();
 sg13g2_fill_1 FILLER_48_1110 ();
 sg13g2_fill_1 FILLER_48_1116 ();
 sg13g2_fill_1 FILLER_48_1123 ();
 sg13g2_fill_1 FILLER_48_1141 ();
 sg13g2_decap_4 FILLER_48_1147 ();
 sg13g2_fill_1 FILLER_48_1228 ();
 sg13g2_fill_1 FILLER_48_1263 ();
 sg13g2_fill_2 FILLER_48_1269 ();
 sg13g2_fill_1 FILLER_48_1371 ();
 sg13g2_fill_1 FILLER_48_1376 ();
 sg13g2_fill_2 FILLER_48_1395 ();
 sg13g2_fill_1 FILLER_48_1397 ();
 sg13g2_fill_2 FILLER_48_1428 ();
 sg13g2_fill_1 FILLER_48_1430 ();
 sg13g2_fill_2 FILLER_48_1465 ();
 sg13g2_fill_1 FILLER_48_1467 ();
 sg13g2_decap_8 FILLER_48_1472 ();
 sg13g2_fill_1 FILLER_48_1483 ();
 sg13g2_fill_1 FILLER_48_1492 ();
 sg13g2_decap_8 FILLER_48_1502 ();
 sg13g2_fill_1 FILLER_48_1513 ();
 sg13g2_fill_1 FILLER_48_1519 ();
 sg13g2_fill_1 FILLER_48_1528 ();
 sg13g2_fill_2 FILLER_48_1537 ();
 sg13g2_fill_2 FILLER_48_1543 ();
 sg13g2_fill_2 FILLER_48_1549 ();
 sg13g2_decap_8 FILLER_48_1563 ();
 sg13g2_fill_2 FILLER_48_1596 ();
 sg13g2_fill_1 FILLER_48_1606 ();
 sg13g2_decap_4 FILLER_48_1615 ();
 sg13g2_fill_1 FILLER_48_1619 ();
 sg13g2_fill_1 FILLER_48_1637 ();
 sg13g2_fill_1 FILLER_48_1646 ();
 sg13g2_fill_1 FILLER_48_1655 ();
 sg13g2_fill_2 FILLER_48_1673 ();
 sg13g2_fill_1 FILLER_48_1675 ();
 sg13g2_fill_1 FILLER_48_1700 ();
 sg13g2_decap_4 FILLER_48_1728 ();
 sg13g2_fill_2 FILLER_48_1732 ();
 sg13g2_fill_1 FILLER_49_30 ();
 sg13g2_fill_1 FILLER_49_74 ();
 sg13g2_fill_1 FILLER_49_79 ();
 sg13g2_fill_2 FILLER_49_87 ();
 sg13g2_fill_1 FILLER_49_190 ();
 sg13g2_fill_1 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_239 ();
 sg13g2_fill_1 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_decap_4 FILLER_49_392 ();
 sg13g2_fill_1 FILLER_49_452 ();
 sg13g2_fill_1 FILLER_49_464 ();
 sg13g2_fill_2 FILLER_49_470 ();
 sg13g2_fill_1 FILLER_49_476 ();
 sg13g2_fill_1 FILLER_49_481 ();
 sg13g2_fill_2 FILLER_49_497 ();
 sg13g2_fill_1 FILLER_49_509 ();
 sg13g2_fill_1 FILLER_49_518 ();
 sg13g2_fill_1 FILLER_49_545 ();
 sg13g2_fill_1 FILLER_49_598 ();
 sg13g2_fill_1 FILLER_49_625 ();
 sg13g2_decap_4 FILLER_49_636 ();
 sg13g2_fill_2 FILLER_49_655 ();
 sg13g2_fill_2 FILLER_49_677 ();
 sg13g2_fill_2 FILLER_49_698 ();
 sg13g2_fill_2 FILLER_49_778 ();
 sg13g2_fill_1 FILLER_49_788 ();
 sg13g2_fill_1 FILLER_49_834 ();
 sg13g2_fill_1 FILLER_49_841 ();
 sg13g2_fill_1 FILLER_49_847 ();
 sg13g2_fill_1 FILLER_49_852 ();
 sg13g2_fill_1 FILLER_49_858 ();
 sg13g2_decap_4 FILLER_49_957 ();
 sg13g2_fill_1 FILLER_49_961 ();
 sg13g2_fill_2 FILLER_49_967 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_fill_2 FILLER_49_1002 ();
 sg13g2_fill_1 FILLER_49_1060 ();
 sg13g2_fill_1 FILLER_49_1082 ();
 sg13g2_fill_2 FILLER_49_1089 ();
 sg13g2_fill_2 FILLER_49_1138 ();
 sg13g2_fill_1 FILLER_49_1170 ();
 sg13g2_fill_1 FILLER_49_1196 ();
 sg13g2_fill_1 FILLER_49_1215 ();
 sg13g2_fill_2 FILLER_49_1229 ();
 sg13g2_fill_1 FILLER_49_1231 ();
 sg13g2_fill_1 FILLER_49_1241 ();
 sg13g2_fill_2 FILLER_49_1263 ();
 sg13g2_fill_1 FILLER_49_1272 ();
 sg13g2_fill_2 FILLER_49_1312 ();
 sg13g2_fill_1 FILLER_49_1314 ();
 sg13g2_fill_2 FILLER_49_1325 ();
 sg13g2_fill_1 FILLER_49_1327 ();
 sg13g2_fill_1 FILLER_49_1333 ();
 sg13g2_fill_2 FILLER_49_1339 ();
 sg13g2_fill_2 FILLER_49_1346 ();
 sg13g2_fill_1 FILLER_49_1348 ();
 sg13g2_fill_2 FILLER_49_1354 ();
 sg13g2_fill_1 FILLER_49_1364 ();
 sg13g2_fill_1 FILLER_49_1370 ();
 sg13g2_fill_1 FILLER_49_1384 ();
 sg13g2_fill_2 FILLER_49_1393 ();
 sg13g2_fill_2 FILLER_49_1401 ();
 sg13g2_fill_2 FILLER_49_1411 ();
 sg13g2_fill_1 FILLER_49_1418 ();
 sg13g2_fill_1 FILLER_49_1445 ();
 sg13g2_fill_2 FILLER_49_1450 ();
 sg13g2_fill_2 FILLER_49_1457 ();
 sg13g2_decap_8 FILLER_49_1464 ();
 sg13g2_fill_2 FILLER_49_1471 ();
 sg13g2_fill_1 FILLER_49_1473 ();
 sg13g2_fill_2 FILLER_49_1478 ();
 sg13g2_fill_1 FILLER_49_1480 ();
 sg13g2_decap_8 FILLER_49_1517 ();
 sg13g2_decap_8 FILLER_49_1524 ();
 sg13g2_fill_2 FILLER_49_1557 ();
 sg13g2_fill_1 FILLER_49_1567 ();
 sg13g2_decap_4 FILLER_49_1580 ();
 sg13g2_decap_8 FILLER_49_1630 ();
 sg13g2_fill_2 FILLER_49_1637 ();
 sg13g2_fill_1 FILLER_49_1639 ();
 sg13g2_fill_2 FILLER_49_1688 ();
 sg13g2_fill_1 FILLER_49_1698 ();
 sg13g2_fill_1 FILLER_49_1707 ();
 sg13g2_fill_2 FILLER_49_1713 ();
 sg13g2_fill_1 FILLER_49_1744 ();
 sg13g2_decap_4 FILLER_49_1750 ();
 sg13g2_fill_1 FILLER_49_1757 ();
 sg13g2_decap_4 FILLER_49_1770 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_48 ();
 sg13g2_fill_1 FILLER_50_54 ();
 sg13g2_fill_2 FILLER_50_66 ();
 sg13g2_fill_1 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_1 FILLER_50_141 ();
 sg13g2_fill_1 FILLER_50_146 ();
 sg13g2_fill_1 FILLER_50_152 ();
 sg13g2_fill_1 FILLER_50_157 ();
 sg13g2_fill_1 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_172 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_324 ();
 sg13g2_fill_2 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_fill_2 FILLER_50_377 ();
 sg13g2_fill_1 FILLER_50_379 ();
 sg13g2_fill_2 FILLER_50_384 ();
 sg13g2_fill_1 FILLER_50_386 ();
 sg13g2_fill_1 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_397 ();
 sg13g2_fill_2 FILLER_50_441 ();
 sg13g2_fill_2 FILLER_50_472 ();
 sg13g2_fill_1 FILLER_50_478 ();
 sg13g2_fill_1 FILLER_50_526 ();
 sg13g2_fill_1 FILLER_50_531 ();
 sg13g2_fill_1 FILLER_50_538 ();
 sg13g2_fill_1 FILLER_50_544 ();
 sg13g2_fill_2 FILLER_50_548 ();
 sg13g2_fill_1 FILLER_50_554 ();
 sg13g2_fill_1 FILLER_50_560 ();
 sg13g2_fill_2 FILLER_50_565 ();
 sg13g2_fill_1 FILLER_50_567 ();
 sg13g2_decap_4 FILLER_50_573 ();
 sg13g2_fill_1 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_582 ();
 sg13g2_fill_2 FILLER_50_588 ();
 sg13g2_fill_1 FILLER_50_590 ();
 sg13g2_fill_2 FILLER_50_595 ();
 sg13g2_fill_1 FILLER_50_597 ();
 sg13g2_fill_1 FILLER_50_602 ();
 sg13g2_fill_2 FILLER_50_612 ();
 sg13g2_fill_2 FILLER_50_618 ();
 sg13g2_fill_2 FILLER_50_644 ();
 sg13g2_fill_2 FILLER_50_667 ();
 sg13g2_fill_2 FILLER_50_682 ();
 sg13g2_fill_1 FILLER_50_684 ();
 sg13g2_fill_2 FILLER_50_708 ();
 sg13g2_fill_2 FILLER_50_715 ();
 sg13g2_fill_2 FILLER_50_722 ();
 sg13g2_fill_2 FILLER_50_732 ();
 sg13g2_fill_1 FILLER_50_734 ();
 sg13g2_decap_8 FILLER_50_739 ();
 sg13g2_fill_1 FILLER_50_746 ();
 sg13g2_fill_2 FILLER_50_763 ();
 sg13g2_fill_1 FILLER_50_777 ();
 sg13g2_fill_1 FILLER_50_809 ();
 sg13g2_fill_2 FILLER_50_880 ();
 sg13g2_fill_2 FILLER_50_890 ();
 sg13g2_fill_1 FILLER_50_892 ();
 sg13g2_fill_1 FILLER_50_919 ();
 sg13g2_decap_8 FILLER_50_924 ();
 sg13g2_fill_2 FILLER_50_935 ();
 sg13g2_fill_2 FILLER_50_941 ();
 sg13g2_fill_1 FILLER_50_943 ();
 sg13g2_decap_4 FILLER_50_988 ();
 sg13g2_fill_1 FILLER_50_998 ();
 sg13g2_fill_2 FILLER_50_1009 ();
 sg13g2_fill_2 FILLER_50_1041 ();
 sg13g2_fill_1 FILLER_50_1043 ();
 sg13g2_fill_1 FILLER_50_1051 ();
 sg13g2_fill_2 FILLER_50_1057 ();
 sg13g2_fill_2 FILLER_50_1068 ();
 sg13g2_fill_1 FILLER_50_1070 ();
 sg13g2_fill_2 FILLER_50_1105 ();
 sg13g2_decap_4 FILLER_50_1112 ();
 sg13g2_fill_2 FILLER_50_1116 ();
 sg13g2_fill_2 FILLER_50_1144 ();
 sg13g2_fill_1 FILLER_50_1158 ();
 sg13g2_fill_2 FILLER_50_1164 ();
 sg13g2_fill_2 FILLER_50_1171 ();
 sg13g2_fill_2 FILLER_50_1178 ();
 sg13g2_fill_2 FILLER_50_1186 ();
 sg13g2_fill_1 FILLER_50_1231 ();
 sg13g2_fill_2 FILLER_50_1249 ();
 sg13g2_fill_1 FILLER_50_1251 ();
 sg13g2_fill_2 FILLER_50_1272 ();
 sg13g2_fill_1 FILLER_50_1295 ();
 sg13g2_fill_1 FILLER_50_1301 ();
 sg13g2_fill_1 FILLER_50_1327 ();
 sg13g2_fill_2 FILLER_50_1338 ();
 sg13g2_fill_2 FILLER_50_1345 ();
 sg13g2_decap_4 FILLER_50_1389 ();
 sg13g2_fill_1 FILLER_50_1438 ();
 sg13g2_fill_1 FILLER_50_1444 ();
 sg13g2_fill_2 FILLER_50_1449 ();
 sg13g2_fill_2 FILLER_50_1455 ();
 sg13g2_fill_2 FILLER_50_1461 ();
 sg13g2_fill_1 FILLER_50_1463 ();
 sg13g2_fill_1 FILLER_50_1498 ();
 sg13g2_fill_1 FILLER_50_1504 ();
 sg13g2_fill_1 FILLER_50_1513 ();
 sg13g2_fill_2 FILLER_50_1526 ();
 sg13g2_fill_1 FILLER_50_1559 ();
 sg13g2_fill_1 FILLER_50_1573 ();
 sg13g2_decap_8 FILLER_50_1587 ();
 sg13g2_decap_4 FILLER_50_1594 ();
 sg13g2_fill_1 FILLER_50_1635 ();
 sg13g2_decap_8 FILLER_50_1640 ();
 sg13g2_fill_2 FILLER_50_1647 ();
 sg13g2_fill_2 FILLER_50_1657 ();
 sg13g2_decap_4 FILLER_50_1667 ();
 sg13g2_fill_2 FILLER_50_1694 ();
 sg13g2_fill_2 FILLER_50_1704 ();
 sg13g2_fill_1 FILLER_50_1710 ();
 sg13g2_fill_2 FILLER_50_1715 ();
 sg13g2_fill_2 FILLER_50_1733 ();
 sg13g2_fill_1 FILLER_50_1735 ();
 sg13g2_decap_8 FILLER_50_1739 ();
 sg13g2_decap_4 FILLER_50_1746 ();
 sg13g2_fill_1 FILLER_50_1773 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_95 ();
 sg13g2_fill_2 FILLER_51_179 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_fill_1 FILLER_51_280 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_304 ();
 sg13g2_fill_2 FILLER_51_318 ();
 sg13g2_fill_1 FILLER_51_354 ();
 sg13g2_fill_2 FILLER_51_381 ();
 sg13g2_fill_2 FILLER_51_402 ();
 sg13g2_fill_2 FILLER_51_414 ();
 sg13g2_fill_2 FILLER_51_440 ();
 sg13g2_fill_1 FILLER_51_447 ();
 sg13g2_fill_2 FILLER_51_456 ();
 sg13g2_decap_8 FILLER_51_468 ();
 sg13g2_decap_4 FILLER_51_475 ();
 sg13g2_fill_2 FILLER_51_479 ();
 sg13g2_decap_4 FILLER_51_499 ();
 sg13g2_fill_1 FILLER_51_528 ();
 sg13g2_fill_2 FILLER_51_539 ();
 sg13g2_fill_2 FILLER_51_567 ();
 sg13g2_fill_1 FILLER_51_569 ();
 sg13g2_fill_1 FILLER_51_575 ();
 sg13g2_fill_2 FILLER_51_602 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_fill_2 FILLER_51_631 ();
 sg13g2_fill_1 FILLER_51_668 ();
 sg13g2_fill_1 FILLER_51_733 ();
 sg13g2_fill_1 FILLER_51_739 ();
 sg13g2_fill_1 FILLER_51_749 ();
 sg13g2_fill_1 FILLER_51_755 ();
 sg13g2_fill_1 FILLER_51_776 ();
 sg13g2_fill_2 FILLER_51_793 ();
 sg13g2_fill_1 FILLER_51_799 ();
 sg13g2_fill_2 FILLER_51_843 ();
 sg13g2_fill_1 FILLER_51_845 ();
 sg13g2_fill_2 FILLER_51_872 ();
 sg13g2_fill_2 FILLER_51_900 ();
 sg13g2_fill_2 FILLER_51_906 ();
 sg13g2_fill_1 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_913 ();
 sg13g2_fill_1 FILLER_51_918 ();
 sg13g2_fill_1 FILLER_51_950 ();
 sg13g2_fill_2 FILLER_51_955 ();
 sg13g2_fill_2 FILLER_51_961 ();
 sg13g2_decap_8 FILLER_51_967 ();
 sg13g2_fill_1 FILLER_51_979 ();
 sg13g2_fill_1 FILLER_51_984 ();
 sg13g2_fill_1 FILLER_51_991 ();
 sg13g2_fill_1 FILLER_51_1004 ();
 sg13g2_fill_1 FILLER_51_1010 ();
 sg13g2_fill_1 FILLER_51_1083 ();
 sg13g2_fill_2 FILLER_51_1094 ();
 sg13g2_fill_2 FILLER_51_1102 ();
 sg13g2_fill_2 FILLER_51_1122 ();
 sg13g2_fill_1 FILLER_51_1124 ();
 sg13g2_fill_2 FILLER_51_1129 ();
 sg13g2_fill_2 FILLER_51_1136 ();
 sg13g2_fill_1 FILLER_51_1141 ();
 sg13g2_fill_2 FILLER_51_1183 ();
 sg13g2_fill_1 FILLER_51_1204 ();
 sg13g2_fill_1 FILLER_51_1211 ();
 sg13g2_fill_1 FILLER_51_1219 ();
 sg13g2_fill_1 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1270 ();
 sg13g2_fill_2 FILLER_51_1277 ();
 sg13g2_fill_1 FILLER_51_1279 ();
 sg13g2_fill_1 FILLER_51_1317 ();
 sg13g2_fill_1 FILLER_51_1358 ();
 sg13g2_fill_2 FILLER_51_1389 ();
 sg13g2_fill_1 FILLER_51_1391 ();
 sg13g2_decap_8 FILLER_51_1426 ();
 sg13g2_fill_2 FILLER_51_1445 ();
 sg13g2_fill_1 FILLER_51_1457 ();
 sg13g2_fill_2 FILLER_51_1462 ();
 sg13g2_fill_2 FILLER_51_1473 ();
 sg13g2_fill_1 FILLER_51_1480 ();
 sg13g2_fill_1 FILLER_51_1486 ();
 sg13g2_fill_2 FILLER_51_1495 ();
 sg13g2_decap_8 FILLER_51_1505 ();
 sg13g2_decap_4 FILLER_51_1512 ();
 sg13g2_fill_1 FILLER_51_1516 ();
 sg13g2_decap_8 FILLER_51_1526 ();
 sg13g2_decap_4 FILLER_51_1533 ();
 sg13g2_fill_1 FILLER_51_1547 ();
 sg13g2_decap_8 FILLER_51_1557 ();
 sg13g2_fill_1 FILLER_51_1564 ();
 sg13g2_fill_1 FILLER_51_1581 ();
 sg13g2_fill_2 FILLER_51_1586 ();
 sg13g2_fill_1 FILLER_51_1588 ();
 sg13g2_fill_2 FILLER_51_1644 ();
 sg13g2_decap_4 FILLER_51_1650 ();
 sg13g2_fill_1 FILLER_51_1654 ();
 sg13g2_fill_1 FILLER_51_1670 ();
 sg13g2_fill_2 FILLER_51_1685 ();
 sg13g2_fill_2 FILLER_51_1696 ();
 sg13g2_fill_1 FILLER_51_1698 ();
 sg13g2_decap_4 FILLER_51_1704 ();
 sg13g2_fill_1 FILLER_51_1712 ();
 sg13g2_decap_4 FILLER_51_1740 ();
 sg13g2_fill_2 FILLER_51_1744 ();
 sg13g2_decap_8 FILLER_51_1764 ();
 sg13g2_fill_2 FILLER_51_1771 ();
 sg13g2_fill_1 FILLER_51_1773 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_46 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_74 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_201 ();
 sg13g2_fill_1 FILLER_52_267 ();
 sg13g2_fill_2 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_309 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_2 FILLER_52_367 ();
 sg13g2_fill_2 FILLER_52_382 ();
 sg13g2_fill_1 FILLER_52_384 ();
 sg13g2_fill_1 FILLER_52_392 ();
 sg13g2_fill_1 FILLER_52_401 ();
 sg13g2_fill_1 FILLER_52_406 ();
 sg13g2_fill_2 FILLER_52_418 ();
 sg13g2_fill_2 FILLER_52_493 ();
 sg13g2_fill_2 FILLER_52_504 ();
 sg13g2_fill_1 FILLER_52_506 ();
 sg13g2_fill_2 FILLER_52_515 ();
 sg13g2_fill_2 FILLER_52_550 ();
 sg13g2_fill_1 FILLER_52_552 ();
 sg13g2_fill_2 FILLER_52_594 ();
 sg13g2_fill_2 FILLER_52_600 ();
 sg13g2_fill_1 FILLER_52_602 ();
 sg13g2_fill_2 FILLER_52_652 ();
 sg13g2_fill_2 FILLER_52_672 ();
 sg13g2_fill_2 FILLER_52_689 ();
 sg13g2_fill_2 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_718 ();
 sg13g2_fill_1 FILLER_52_729 ();
 sg13g2_fill_2 FILLER_52_765 ();
 sg13g2_fill_2 FILLER_52_786 ();
 sg13g2_decap_4 FILLER_52_828 ();
 sg13g2_decap_4 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_840 ();
 sg13g2_fill_2 FILLER_52_845 ();
 sg13g2_fill_1 FILLER_52_852 ();
 sg13g2_decap_8 FILLER_52_857 ();
 sg13g2_decap_8 FILLER_52_864 ();
 sg13g2_fill_2 FILLER_52_871 ();
 sg13g2_fill_1 FILLER_52_873 ();
 sg13g2_decap_4 FILLER_52_878 ();
 sg13g2_fill_1 FILLER_52_909 ();
 sg13g2_fill_2 FILLER_52_924 ();
 sg13g2_fill_1 FILLER_52_930 ();
 sg13g2_fill_2 FILLER_52_935 ();
 sg13g2_fill_1 FILLER_52_941 ();
 sg13g2_fill_2 FILLER_52_947 ();
 sg13g2_fill_2 FILLER_52_953 ();
 sg13g2_fill_1 FILLER_52_955 ();
 sg13g2_fill_1 FILLER_52_982 ();
 sg13g2_fill_1 FILLER_52_987 ();
 sg13g2_fill_2 FILLER_52_999 ();
 sg13g2_decap_4 FILLER_52_1006 ();
 sg13g2_fill_2 FILLER_52_1030 ();
 sg13g2_fill_1 FILLER_52_1032 ();
 sg13g2_fill_2 FILLER_52_1040 ();
 sg13g2_fill_1 FILLER_52_1042 ();
 sg13g2_fill_1 FILLER_52_1049 ();
 sg13g2_fill_1 FILLER_52_1055 ();
 sg13g2_fill_1 FILLER_52_1065 ();
 sg13g2_fill_2 FILLER_52_1071 ();
 sg13g2_fill_1 FILLER_52_1077 ();
 sg13g2_fill_2 FILLER_52_1133 ();
 sg13g2_fill_2 FILLER_52_1139 ();
 sg13g2_fill_1 FILLER_52_1141 ();
 sg13g2_fill_2 FILLER_52_1155 ();
 sg13g2_fill_1 FILLER_52_1157 ();
 sg13g2_fill_1 FILLER_52_1228 ();
 sg13g2_fill_2 FILLER_52_1239 ();
 sg13g2_fill_2 FILLER_52_1248 ();
 sg13g2_fill_1 FILLER_52_1267 ();
 sg13g2_decap_8 FILLER_52_1272 ();
 sg13g2_decap_8 FILLER_52_1293 ();
 sg13g2_fill_2 FILLER_52_1300 ();
 sg13g2_fill_1 FILLER_52_1302 ();
 sg13g2_fill_1 FILLER_52_1312 ();
 sg13g2_fill_1 FILLER_52_1321 ();
 sg13g2_fill_1 FILLER_52_1348 ();
 sg13g2_fill_1 FILLER_52_1358 ();
 sg13g2_fill_2 FILLER_52_1363 ();
 sg13g2_decap_4 FILLER_52_1405 ();
 sg13g2_fill_2 FILLER_52_1409 ();
 sg13g2_fill_2 FILLER_52_1422 ();
 sg13g2_decap_4 FILLER_52_1429 ();
 sg13g2_fill_1 FILLER_52_1433 ();
 sg13g2_fill_1 FILLER_52_1438 ();
 sg13g2_fill_2 FILLER_52_1450 ();
 sg13g2_fill_2 FILLER_52_1457 ();
 sg13g2_fill_1 FILLER_52_1485 ();
 sg13g2_fill_1 FILLER_52_1491 ();
 sg13g2_decap_4 FILLER_52_1500 ();
 sg13g2_fill_2 FILLER_52_1504 ();
 sg13g2_decap_8 FILLER_52_1527 ();
 sg13g2_decap_4 FILLER_52_1554 ();
 sg13g2_fill_1 FILLER_52_1558 ();
 sg13g2_fill_1 FILLER_52_1635 ();
 sg13g2_fill_2 FILLER_52_1640 ();
 sg13g2_decap_4 FILLER_52_1651 ();
 sg13g2_decap_4 FILLER_52_1664 ();
 sg13g2_fill_1 FILLER_52_1730 ();
 sg13g2_decap_4 FILLER_52_1736 ();
 sg13g2_fill_2 FILLER_52_1744 ();
 sg13g2_fill_2 FILLER_52_1767 ();
 sg13g2_fill_1 FILLER_52_1769 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_27 ();
 sg13g2_fill_2 FILLER_53_33 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_fill_1 FILLER_53_116 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_129 ();
 sg13g2_fill_2 FILLER_53_135 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_2 FILLER_53_219 ();
 sg13g2_fill_1 FILLER_53_231 ();
 sg13g2_fill_1 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_fill_1 FILLER_53_312 ();
 sg13g2_fill_2 FILLER_53_339 ();
 sg13g2_fill_2 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_386 ();
 sg13g2_fill_1 FILLER_53_388 ();
 sg13g2_fill_2 FILLER_53_394 ();
 sg13g2_fill_2 FILLER_53_401 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_fill_1 FILLER_53_409 ();
 sg13g2_fill_2 FILLER_53_445 ();
 sg13g2_fill_2 FILLER_53_452 ();
 sg13g2_fill_2 FILLER_53_458 ();
 sg13g2_fill_1 FILLER_53_460 ();
 sg13g2_fill_2 FILLER_53_465 ();
 sg13g2_fill_1 FILLER_53_467 ();
 sg13g2_fill_2 FILLER_53_472 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_2 FILLER_53_480 ();
 sg13g2_fill_2 FILLER_53_486 ();
 sg13g2_fill_1 FILLER_53_488 ();
 sg13g2_fill_2 FILLER_53_497 ();
 sg13g2_fill_2 FILLER_53_515 ();
 sg13g2_fill_1 FILLER_53_517 ();
 sg13g2_fill_1 FILLER_53_547 ();
 sg13g2_fill_1 FILLER_53_552 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_fill_1 FILLER_53_622 ();
 sg13g2_fill_1 FILLER_53_649 ();
 sg13g2_fill_1 FILLER_53_654 ();
 sg13g2_fill_2 FILLER_53_681 ();
 sg13g2_fill_1 FILLER_53_713 ();
 sg13g2_fill_1 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_723 ();
 sg13g2_fill_2 FILLER_53_727 ();
 sg13g2_fill_1 FILLER_53_766 ();
 sg13g2_fill_2 FILLER_53_772 ();
 sg13g2_fill_2 FILLER_53_779 ();
 sg13g2_decap_8 FILLER_53_831 ();
 sg13g2_fill_2 FILLER_53_838 ();
 sg13g2_fill_1 FILLER_53_840 ();
 sg13g2_fill_1 FILLER_53_849 ();
 sg13g2_fill_1 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_859 ();
 sg13g2_decap_4 FILLER_53_868 ();
 sg13g2_fill_2 FILLER_53_932 ();
 sg13g2_fill_2 FILLER_53_938 ();
 sg13g2_fill_1 FILLER_53_940 ();
 sg13g2_fill_1 FILLER_53_967 ();
 sg13g2_fill_2 FILLER_53_972 ();
 sg13g2_fill_1 FILLER_53_974 ();
 sg13g2_fill_1 FILLER_53_979 ();
 sg13g2_fill_2 FILLER_53_989 ();
 sg13g2_fill_1 FILLER_53_998 ();
 sg13g2_fill_2 FILLER_53_1023 ();
 sg13g2_fill_1 FILLER_53_1025 ();
 sg13g2_fill_2 FILLER_53_1078 ();
 sg13g2_fill_2 FILLER_53_1084 ();
 sg13g2_fill_1 FILLER_53_1090 ();
 sg13g2_fill_1 FILLER_53_1117 ();
 sg13g2_fill_1 FILLER_53_1170 ();
 sg13g2_fill_2 FILLER_53_1175 ();
 sg13g2_fill_1 FILLER_53_1186 ();
 sg13g2_fill_1 FILLER_53_1191 ();
 sg13g2_fill_2 FILLER_53_1201 ();
 sg13g2_decap_8 FILLER_53_1342 ();
 sg13g2_decap_4 FILLER_53_1349 ();
 sg13g2_decap_4 FILLER_53_1383 ();
 sg13g2_fill_2 FILLER_53_1400 ();
 sg13g2_fill_1 FILLER_53_1402 ();
 sg13g2_fill_2 FILLER_53_1419 ();
 sg13g2_fill_1 FILLER_53_1421 ();
 sg13g2_fill_1 FILLER_53_1440 ();
 sg13g2_fill_1 FILLER_53_1459 ();
 sg13g2_fill_2 FILLER_53_1480 ();
 sg13g2_fill_2 FILLER_53_1486 ();
 sg13g2_decap_4 FILLER_53_1498 ();
 sg13g2_fill_1 FILLER_53_1502 ();
 sg13g2_decap_4 FILLER_53_1511 ();
 sg13g2_fill_2 FILLER_53_1515 ();
 sg13g2_fill_1 FILLER_53_1525 ();
 sg13g2_fill_2 FILLER_53_1534 ();
 sg13g2_fill_1 FILLER_53_1536 ();
 sg13g2_fill_1 FILLER_53_1558 ();
 sg13g2_fill_2 FILLER_53_1571 ();
 sg13g2_fill_1 FILLER_53_1573 ();
 sg13g2_decap_4 FILLER_53_1577 ();
 sg13g2_fill_1 FILLER_53_1585 ();
 sg13g2_fill_1 FILLER_53_1590 ();
 sg13g2_fill_1 FILLER_53_1596 ();
 sg13g2_fill_1 FILLER_53_1609 ();
 sg13g2_fill_2 FILLER_53_1629 ();
 sg13g2_fill_1 FILLER_53_1631 ();
 sg13g2_fill_2 FILLER_53_1636 ();
 sg13g2_fill_1 FILLER_53_1638 ();
 sg13g2_decap_8 FILLER_53_1668 ();
 sg13g2_decap_4 FILLER_53_1675 ();
 sg13g2_fill_1 FILLER_53_1679 ();
 sg13g2_decap_4 FILLER_53_1684 ();
 sg13g2_fill_1 FILLER_53_1692 ();
 sg13g2_fill_1 FILLER_53_1698 ();
 sg13g2_fill_1 FILLER_53_1715 ();
 sg13g2_fill_1 FILLER_53_1721 ();
 sg13g2_fill_2 FILLER_53_1746 ();
 sg13g2_fill_1 FILLER_53_1748 ();
 sg13g2_fill_1 FILLER_53_1773 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_11 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_2 FILLER_54_114 ();
 sg13g2_fill_1 FILLER_54_165 ();
 sg13g2_fill_1 FILLER_54_200 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_fill_2 FILLER_54_378 ();
 sg13g2_fill_1 FILLER_54_417 ();
 sg13g2_fill_1 FILLER_54_421 ();
 sg13g2_decap_4 FILLER_54_441 ();
 sg13g2_fill_2 FILLER_54_445 ();
 sg13g2_fill_2 FILLER_54_451 ();
 sg13g2_fill_1 FILLER_54_453 ();
 sg13g2_fill_2 FILLER_54_484 ();
 sg13g2_decap_4 FILLER_54_490 ();
 sg13g2_fill_1 FILLER_54_494 ();
 sg13g2_fill_2 FILLER_54_498 ();
 sg13g2_fill_1 FILLER_54_516 ();
 sg13g2_fill_1 FILLER_54_523 ();
 sg13g2_fill_2 FILLER_54_579 ();
 sg13g2_fill_1 FILLER_54_594 ();
 sg13g2_fill_1 FILLER_54_621 ();
 sg13g2_fill_2 FILLER_54_643 ();
 sg13g2_fill_1 FILLER_54_645 ();
 sg13g2_fill_1 FILLER_54_663 ();
 sg13g2_fill_1 FILLER_54_685 ();
 sg13g2_fill_2 FILLER_54_699 ();
 sg13g2_fill_1 FILLER_54_701 ();
 sg13g2_fill_2 FILLER_54_745 ();
 sg13g2_fill_1 FILLER_54_823 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_fill_1 FILLER_54_846 ();
 sg13g2_fill_1 FILLER_54_858 ();
 sg13g2_fill_1 FILLER_54_864 ();
 sg13g2_decap_4 FILLER_54_869 ();
 sg13g2_fill_1 FILLER_54_873 ();
 sg13g2_fill_1 FILLER_54_886 ();
 sg13g2_fill_1 FILLER_54_899 ();
 sg13g2_fill_1 FILLER_54_904 ();
 sg13g2_fill_1 FILLER_54_936 ();
 sg13g2_fill_1 FILLER_54_941 ();
 sg13g2_fill_1 FILLER_54_963 ();
 sg13g2_fill_1 FILLER_54_968 ();
 sg13g2_fill_1 FILLER_54_1007 ();
 sg13g2_fill_1 FILLER_54_1017 ();
 sg13g2_fill_1 FILLER_54_1022 ();
 sg13g2_fill_1 FILLER_54_1027 ();
 sg13g2_fill_1 FILLER_54_1058 ();
 sg13g2_decap_4 FILLER_54_1089 ();
 sg13g2_fill_1 FILLER_54_1093 ();
 sg13g2_fill_1 FILLER_54_1120 ();
 sg13g2_fill_1 FILLER_54_1130 ();
 sg13g2_fill_1 FILLER_54_1135 ();
 sg13g2_fill_1 FILLER_54_1141 ();
 sg13g2_fill_1 FILLER_54_1147 ();
 sg13g2_fill_1 FILLER_54_1153 ();
 sg13g2_fill_1 FILLER_54_1158 ();
 sg13g2_fill_1 FILLER_54_1178 ();
 sg13g2_fill_2 FILLER_54_1184 ();
 sg13g2_fill_2 FILLER_54_1220 ();
 sg13g2_fill_2 FILLER_54_1225 ();
 sg13g2_fill_2 FILLER_54_1235 ();
 sg13g2_fill_1 FILLER_54_1242 ();
 sg13g2_fill_2 FILLER_54_1262 ();
 sg13g2_fill_1 FILLER_54_1264 ();
 sg13g2_fill_2 FILLER_54_1269 ();
 sg13g2_decap_8 FILLER_54_1275 ();
 sg13g2_fill_1 FILLER_54_1282 ();
 sg13g2_fill_2 FILLER_54_1287 ();
 sg13g2_fill_1 FILLER_54_1289 ();
 sg13g2_decap_4 FILLER_54_1298 ();
 sg13g2_fill_1 FILLER_54_1302 ();
 sg13g2_decap_8 FILLER_54_1307 ();
 sg13g2_fill_1 FILLER_54_1314 ();
 sg13g2_fill_1 FILLER_54_1319 ();
 sg13g2_fill_1 FILLER_54_1324 ();
 sg13g2_decap_4 FILLER_54_1351 ();
 sg13g2_fill_2 FILLER_54_1355 ();
 sg13g2_fill_2 FILLER_54_1361 ();
 sg13g2_decap_4 FILLER_54_1372 ();
 sg13g2_decap_8 FILLER_54_1381 ();
 sg13g2_decap_8 FILLER_54_1388 ();
 sg13g2_decap_4 FILLER_54_1395 ();
 sg13g2_fill_1 FILLER_54_1406 ();
 sg13g2_fill_1 FILLER_54_1415 ();
 sg13g2_decap_4 FILLER_54_1424 ();
 sg13g2_fill_1 FILLER_54_1447 ();
 sg13g2_fill_1 FILLER_54_1457 ();
 sg13g2_fill_1 FILLER_54_1463 ();
 sg13g2_fill_1 FILLER_54_1482 ();
 sg13g2_fill_1 FILLER_54_1514 ();
 sg13g2_fill_1 FILLER_54_1547 ();
 sg13g2_fill_1 FILLER_54_1556 ();
 sg13g2_fill_1 FILLER_54_1562 ();
 sg13g2_fill_1 FILLER_54_1567 ();
 sg13g2_fill_1 FILLER_54_1572 ();
 sg13g2_fill_1 FILLER_54_1577 ();
 sg13g2_fill_2 FILLER_54_1615 ();
 sg13g2_fill_1 FILLER_54_1617 ();
 sg13g2_fill_2 FILLER_54_1630 ();
 sg13g2_fill_1 FILLER_54_1636 ();
 sg13g2_fill_2 FILLER_54_1645 ();
 sg13g2_fill_2 FILLER_54_1677 ();
 sg13g2_fill_1 FILLER_54_1692 ();
 sg13g2_fill_1 FILLER_54_1702 ();
 sg13g2_fill_1 FILLER_54_1708 ();
 sg13g2_fill_1 FILLER_54_1717 ();
 sg13g2_fill_1 FILLER_54_1733 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_fill_1 FILLER_54_1752 ();
 sg13g2_fill_1 FILLER_54_1761 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_7 ();
 sg13g2_fill_2 FILLER_55_78 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_fill_1 FILLER_55_156 ();
 sg13g2_fill_1 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_204 ();
 sg13g2_fill_1 FILLER_55_227 ();
 sg13g2_fill_2 FILLER_55_232 ();
 sg13g2_fill_2 FILLER_55_312 ();
 sg13g2_fill_1 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_385 ();
 sg13g2_fill_2 FILLER_55_389 ();
 sg13g2_fill_2 FILLER_55_395 ();
 sg13g2_fill_2 FILLER_55_456 ();
 sg13g2_fill_2 FILLER_55_505 ();
 sg13g2_fill_1 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_636 ();
 sg13g2_fill_2 FILLER_55_663 ();
 sg13g2_fill_2 FILLER_55_691 ();
 sg13g2_decap_8 FILLER_55_698 ();
 sg13g2_decap_8 FILLER_55_739 ();
 sg13g2_decap_4 FILLER_55_746 ();
 sg13g2_fill_1 FILLER_55_750 ();
 sg13g2_fill_2 FILLER_55_810 ();
 sg13g2_fill_1 FILLER_55_812 ();
 sg13g2_fill_2 FILLER_55_817 ();
 sg13g2_fill_1 FILLER_55_827 ();
 sg13g2_fill_2 FILLER_55_866 ();
 sg13g2_fill_1 FILLER_55_868 ();
 sg13g2_fill_1 FILLER_55_899 ();
 sg13g2_fill_2 FILLER_55_930 ();
 sg13g2_fill_1 FILLER_55_997 ();
 sg13g2_fill_2 FILLER_55_1024 ();
 sg13g2_fill_1 FILLER_55_1026 ();
 sg13g2_fill_1 FILLER_55_1057 ();
 sg13g2_fill_2 FILLER_55_1063 ();
 sg13g2_fill_1 FILLER_55_1073 ();
 sg13g2_fill_1 FILLER_55_1079 ();
 sg13g2_fill_1 FILLER_55_1084 ();
 sg13g2_fill_2 FILLER_55_1090 ();
 sg13g2_fill_1 FILLER_55_1100 ();
 sg13g2_fill_2 FILLER_55_1122 ();
 sg13g2_fill_1 FILLER_55_1128 ();
 sg13g2_decap_8 FILLER_55_1141 ();
 sg13g2_fill_1 FILLER_55_1148 ();
 sg13g2_fill_2 FILLER_55_1190 ();
 sg13g2_fill_1 FILLER_55_1196 ();
 sg13g2_fill_1 FILLER_55_1213 ();
 sg13g2_fill_1 FILLER_55_1218 ();
 sg13g2_decap_4 FILLER_55_1228 ();
 sg13g2_fill_2 FILLER_55_1232 ();
 sg13g2_fill_2 FILLER_55_1261 ();
 sg13g2_fill_1 FILLER_55_1263 ();
 sg13g2_fill_2 FILLER_55_1268 ();
 sg13g2_fill_1 FILLER_55_1270 ();
 sg13g2_decap_4 FILLER_55_1312 ();
 sg13g2_fill_1 FILLER_55_1316 ();
 sg13g2_decap_4 FILLER_55_1321 ();
 sg13g2_fill_1 FILLER_55_1325 ();
 sg13g2_fill_1 FILLER_55_1331 ();
 sg13g2_fill_1 FILLER_55_1340 ();
 sg13g2_decap_4 FILLER_55_1350 ();
 sg13g2_fill_2 FILLER_55_1354 ();
 sg13g2_fill_1 FILLER_55_1361 ();
 sg13g2_fill_1 FILLER_55_1374 ();
 sg13g2_fill_2 FILLER_55_1383 ();
 sg13g2_fill_2 FILLER_55_1406 ();
 sg13g2_decap_8 FILLER_55_1412 ();
 sg13g2_decap_4 FILLER_55_1419 ();
 sg13g2_fill_1 FILLER_55_1423 ();
 sg13g2_fill_2 FILLER_55_1467 ();
 sg13g2_fill_1 FILLER_55_1469 ();
 sg13g2_fill_2 FILLER_55_1490 ();
 sg13g2_fill_1 FILLER_55_1492 ();
 sg13g2_decap_4 FILLER_55_1517 ();
 sg13g2_fill_2 FILLER_55_1521 ();
 sg13g2_decap_8 FILLER_55_1543 ();
 sg13g2_fill_2 FILLER_55_1550 ();
 sg13g2_fill_2 FILLER_55_1564 ();
 sg13g2_fill_2 FILLER_55_1628 ();
 sg13g2_fill_2 FILLER_55_1638 ();
 sg13g2_fill_2 FILLER_55_1644 ();
 sg13g2_fill_2 FILLER_55_1663 ();
 sg13g2_fill_1 FILLER_55_1682 ();
 sg13g2_fill_2 FILLER_55_1688 ();
 sg13g2_fill_2 FILLER_55_1695 ();
 sg13g2_fill_1 FILLER_55_1697 ();
 sg13g2_fill_2 FILLER_55_1726 ();
 sg13g2_fill_1 FILLER_55_1728 ();
 sg13g2_fill_2 FILLER_55_1746 ();
 sg13g2_fill_1 FILLER_55_1753 ();
 sg13g2_fill_1 FILLER_55_1767 ();
 sg13g2_fill_2 FILLER_56_26 ();
 sg13g2_fill_1 FILLER_56_49 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_fill_1 FILLER_56_74 ();
 sg13g2_fill_1 FILLER_56_79 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_133 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_fill_1 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_185 ();
 sg13g2_fill_1 FILLER_56_213 ();
 sg13g2_fill_2 FILLER_56_238 ();
 sg13g2_fill_1 FILLER_56_308 ();
 sg13g2_fill_2 FILLER_56_313 ();
 sg13g2_fill_1 FILLER_56_319 ();
 sg13g2_fill_1 FILLER_56_324 ();
 sg13g2_fill_2 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_362 ();
 sg13g2_fill_1 FILLER_56_369 ();
 sg13g2_fill_1 FILLER_56_380 ();
 sg13g2_fill_1 FILLER_56_407 ();
 sg13g2_fill_1 FILLER_56_412 ();
 sg13g2_fill_2 FILLER_56_423 ();
 sg13g2_fill_2 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_516 ();
 sg13g2_fill_1 FILLER_56_572 ();
 sg13g2_fill_1 FILLER_56_586 ();
 sg13g2_fill_2 FILLER_56_615 ();
 sg13g2_fill_1 FILLER_56_655 ();
 sg13g2_fill_1 FILLER_56_660 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_fill_1 FILLER_56_690 ();
 sg13g2_fill_1 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_718 ();
 sg13g2_fill_2 FILLER_56_725 ();
 sg13g2_fill_2 FILLER_56_757 ();
 sg13g2_fill_1 FILLER_56_759 ();
 sg13g2_fill_2 FILLER_56_828 ();
 sg13g2_fill_1 FILLER_56_838 ();
 sg13g2_fill_2 FILLER_56_865 ();
 sg13g2_decap_4 FILLER_56_871 ();
 sg13g2_fill_2 FILLER_56_875 ();
 sg13g2_fill_2 FILLER_56_882 ();
 sg13g2_fill_1 FILLER_56_884 ();
 sg13g2_fill_2 FILLER_56_889 ();
 sg13g2_decap_8 FILLER_56_895 ();
 sg13g2_decap_8 FILLER_56_902 ();
 sg13g2_fill_1 FILLER_56_934 ();
 sg13g2_fill_1 FILLER_56_944 ();
 sg13g2_fill_1 FILLER_56_950 ();
 sg13g2_fill_1 FILLER_56_956 ();
 sg13g2_fill_2 FILLER_56_962 ();
 sg13g2_fill_2 FILLER_56_990 ();
 sg13g2_fill_1 FILLER_56_997 ();
 sg13g2_fill_2 FILLER_56_1032 ();
 sg13g2_fill_1 FILLER_56_1034 ();
 sg13g2_fill_1 FILLER_56_1056 ();
 sg13g2_fill_1 FILLER_56_1061 ();
 sg13g2_fill_1 FILLER_56_1091 ();
 sg13g2_fill_2 FILLER_56_1096 ();
 sg13g2_fill_1 FILLER_56_1102 ();
 sg13g2_fill_1 FILLER_56_1108 ();
 sg13g2_fill_2 FILLER_56_1117 ();
 sg13g2_decap_4 FILLER_56_1123 ();
 sg13g2_fill_1 FILLER_56_1127 ();
 sg13g2_fill_2 FILLER_56_1163 ();
 sg13g2_fill_1 FILLER_56_1165 ();
 sg13g2_fill_1 FILLER_56_1195 ();
 sg13g2_fill_2 FILLER_56_1201 ();
 sg13g2_fill_1 FILLER_56_1203 ();
 sg13g2_fill_2 FILLER_56_1207 ();
 sg13g2_fill_2 FILLER_56_1243 ();
 sg13g2_fill_1 FILLER_56_1250 ();
 sg13g2_fill_2 FILLER_56_1254 ();
 sg13g2_fill_2 FILLER_56_1275 ();
 sg13g2_fill_1 FILLER_56_1277 ();
 sg13g2_fill_1 FILLER_56_1287 ();
 sg13g2_decap_4 FILLER_56_1292 ();
 sg13g2_fill_1 FILLER_56_1296 ();
 sg13g2_fill_1 FILLER_56_1313 ();
 sg13g2_fill_2 FILLER_56_1357 ();
 sg13g2_fill_2 FILLER_56_1381 ();
 sg13g2_fill_1 FILLER_56_1383 ();
 sg13g2_decap_4 FILLER_56_1417 ();
 sg13g2_fill_2 FILLER_56_1421 ();
 sg13g2_decap_4 FILLER_56_1451 ();
 sg13g2_fill_1 FILLER_56_1455 ();
 sg13g2_fill_2 FILLER_56_1464 ();
 sg13g2_fill_1 FILLER_56_1466 ();
 sg13g2_fill_1 FILLER_56_1470 ();
 sg13g2_decap_4 FILLER_56_1490 ();
 sg13g2_decap_8 FILLER_56_1504 ();
 sg13g2_decap_8 FILLER_56_1511 ();
 sg13g2_decap_8 FILLER_56_1518 ();
 sg13g2_fill_1 FILLER_56_1525 ();
 sg13g2_fill_1 FILLER_56_1534 ();
 sg13g2_fill_2 FILLER_56_1543 ();
 sg13g2_fill_2 FILLER_56_1549 ();
 sg13g2_fill_2 FILLER_56_1564 ();
 sg13g2_decap_8 FILLER_56_1613 ();
 sg13g2_decap_8 FILLER_56_1620 ();
 sg13g2_decap_8 FILLER_56_1627 ();
 sg13g2_decap_8 FILLER_56_1634 ();
 sg13g2_decap_4 FILLER_56_1641 ();
 sg13g2_fill_2 FILLER_56_1645 ();
 sg13g2_fill_1 FILLER_56_1651 ();
 sg13g2_fill_1 FILLER_56_1662 ();
 sg13g2_decap_8 FILLER_56_1667 ();
 sg13g2_fill_2 FILLER_56_1679 ();
 sg13g2_fill_2 FILLER_56_1688 ();
 sg13g2_fill_1 FILLER_56_1690 ();
 sg13g2_fill_1 FILLER_56_1701 ();
 sg13g2_fill_2 FILLER_56_1706 ();
 sg13g2_fill_1 FILLER_56_1708 ();
 sg13g2_decap_4 FILLER_56_1723 ();
 sg13g2_fill_1 FILLER_56_1741 ();
 sg13g2_fill_1 FILLER_56_1753 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_5 ();
 sg13g2_fill_2 FILLER_57_17 ();
 sg13g2_fill_1 FILLER_57_23 ();
 sg13g2_fill_2 FILLER_57_50 ();
 sg13g2_fill_2 FILLER_57_78 ();
 sg13g2_fill_2 FILLER_57_84 ();
 sg13g2_fill_1 FILLER_57_96 ();
 sg13g2_fill_1 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_193 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_333 ();
 sg13g2_fill_1 FILLER_57_359 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_405 ();
 sg13g2_fill_2 FILLER_57_449 ();
 sg13g2_fill_2 FILLER_57_458 ();
 sg13g2_fill_2 FILLER_57_510 ();
 sg13g2_fill_1 FILLER_57_512 ();
 sg13g2_decap_8 FILLER_57_552 ();
 sg13g2_decap_4 FILLER_57_559 ();
 sg13g2_fill_1 FILLER_57_610 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_1 FILLER_57_630 ();
 sg13g2_fill_1 FILLER_57_636 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_fill_1 FILLER_57_722 ();
 sg13g2_fill_1 FILLER_57_734 ();
 sg13g2_fill_1 FILLER_57_743 ();
 sg13g2_fill_1 FILLER_57_768 ();
 sg13g2_fill_1 FILLER_57_774 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_fill_2 FILLER_57_801 ();
 sg13g2_fill_1 FILLER_57_803 ();
 sg13g2_fill_2 FILLER_57_807 ();
 sg13g2_fill_2 FILLER_57_813 ();
 sg13g2_fill_1 FILLER_57_815 ();
 sg13g2_fill_2 FILLER_57_923 ();
 sg13g2_fill_1 FILLER_57_925 ();
 sg13g2_fill_1 FILLER_57_947 ();
 sg13g2_fill_1 FILLER_57_974 ();
 sg13g2_fill_2 FILLER_57_980 ();
 sg13g2_fill_2 FILLER_57_1024 ();
 sg13g2_fill_2 FILLER_57_1033 ();
 sg13g2_fill_2 FILLER_57_1040 ();
 sg13g2_fill_1 FILLER_57_1042 ();
 sg13g2_fill_1 FILLER_57_1048 ();
 sg13g2_fill_2 FILLER_57_1053 ();
 sg13g2_fill_1 FILLER_57_1055 ();
 sg13g2_fill_2 FILLER_57_1060 ();
 sg13g2_fill_1 FILLER_57_1079 ();
 sg13g2_fill_1 FILLER_57_1087 ();
 sg13g2_fill_2 FILLER_57_1116 ();
 sg13g2_fill_1 FILLER_57_1146 ();
 sg13g2_fill_1 FILLER_57_1151 ();
 sg13g2_fill_1 FILLER_57_1156 ();
 sg13g2_fill_1 FILLER_57_1165 ();
 sg13g2_fill_1 FILLER_57_1171 ();
 sg13g2_fill_2 FILLER_57_1212 ();
 sg13g2_fill_1 FILLER_57_1214 ();
 sg13g2_fill_1 FILLER_57_1238 ();
 sg13g2_fill_2 FILLER_57_1289 ();
 sg13g2_fill_1 FILLER_57_1295 ();
 sg13g2_fill_1 FILLER_57_1304 ();
 sg13g2_fill_1 FILLER_57_1315 ();
 sg13g2_fill_1 FILLER_57_1320 ();
 sg13g2_fill_2 FILLER_57_1326 ();
 sg13g2_fill_2 FILLER_57_1332 ();
 sg13g2_fill_1 FILLER_57_1349 ();
 sg13g2_decap_4 FILLER_57_1366 ();
 sg13g2_decap_4 FILLER_57_1383 ();
 sg13g2_fill_2 FILLER_57_1408 ();
 sg13g2_fill_1 FILLER_57_1410 ();
 sg13g2_decap_4 FILLER_57_1415 ();
 sg13g2_decap_4 FILLER_57_1436 ();
 sg13g2_decap_8 FILLER_57_1444 ();
 sg13g2_fill_1 FILLER_57_1460 ();
 sg13g2_fill_1 FILLER_57_1466 ();
 sg13g2_fill_1 FILLER_57_1475 ();
 sg13g2_fill_2 FILLER_57_1481 ();
 sg13g2_fill_2 FILLER_57_1491 ();
 sg13g2_fill_1 FILLER_57_1501 ();
 sg13g2_fill_2 FILLER_57_1522 ();
 sg13g2_fill_2 FILLER_57_1545 ();
 sg13g2_fill_1 FILLER_57_1555 ();
 sg13g2_decap_4 FILLER_57_1568 ();
 sg13g2_decap_8 FILLER_57_1576 ();
 sg13g2_fill_1 FILLER_57_1588 ();
 sg13g2_fill_1 FILLER_57_1593 ();
 sg13g2_fill_1 FILLER_57_1599 ();
 sg13g2_fill_1 FILLER_57_1605 ();
 sg13g2_fill_2 FILLER_57_1611 ();
 sg13g2_fill_1 FILLER_57_1621 ();
 sg13g2_fill_2 FILLER_57_1652 ();
 sg13g2_fill_2 FILLER_57_1676 ();
 sg13g2_fill_1 FILLER_57_1678 ();
 sg13g2_fill_1 FILLER_57_1693 ();
 sg13g2_fill_1 FILLER_57_1699 ();
 sg13g2_fill_1 FILLER_57_1712 ();
 sg13g2_decap_8 FILLER_57_1725 ();
 sg13g2_fill_2 FILLER_57_1732 ();
 sg13g2_decap_4 FILLER_57_1738 ();
 sg13g2_fill_2 FILLER_57_1742 ();
 sg13g2_decap_4 FILLER_57_1768 ();
 sg13g2_fill_2 FILLER_57_1772 ();
 sg13g2_fill_1 FILLER_58_71 ();
 sg13g2_fill_2 FILLER_58_98 ();
 sg13g2_fill_1 FILLER_58_121 ();
 sg13g2_fill_1 FILLER_58_359 ();
 sg13g2_fill_2 FILLER_58_398 ();
 sg13g2_fill_1 FILLER_58_518 ();
 sg13g2_fill_1 FILLER_58_529 ();
 sg13g2_fill_1 FILLER_58_556 ();
 sg13g2_fill_1 FILLER_58_561 ();
 sg13g2_fill_1 FILLER_58_566 ();
 sg13g2_fill_2 FILLER_58_572 ();
 sg13g2_fill_1 FILLER_58_578 ();
 sg13g2_fill_2 FILLER_58_592 ();
 sg13g2_fill_2 FILLER_58_633 ();
 sg13g2_fill_1 FILLER_58_696 ();
 sg13g2_fill_1 FILLER_58_728 ();
 sg13g2_fill_2 FILLER_58_739 ();
 sg13g2_fill_1 FILLER_58_746 ();
 sg13g2_fill_2 FILLER_58_782 ();
 sg13g2_fill_1 FILLER_58_784 ();
 sg13g2_fill_2 FILLER_58_812 ();
 sg13g2_fill_2 FILLER_58_830 ();
 sg13g2_fill_2 FILLER_58_837 ();
 sg13g2_fill_1 FILLER_58_839 ();
 sg13g2_fill_1 FILLER_58_866 ();
 sg13g2_fill_1 FILLER_58_872 ();
 sg13g2_fill_1 FILLER_58_877 ();
 sg13g2_fill_2 FILLER_58_882 ();
 sg13g2_fill_2 FILLER_58_918 ();
 sg13g2_fill_1 FILLER_58_954 ();
 sg13g2_fill_2 FILLER_58_978 ();
 sg13g2_fill_2 FILLER_58_988 ();
 sg13g2_fill_2 FILLER_58_998 ();
 sg13g2_fill_2 FILLER_58_1020 ();
 sg13g2_fill_1 FILLER_58_1048 ();
 sg13g2_fill_2 FILLER_58_1053 ();
 sg13g2_fill_2 FILLER_58_1068 ();
 sg13g2_fill_1 FILLER_58_1093 ();
 sg13g2_fill_1 FILLER_58_1098 ();
 sg13g2_fill_1 FILLER_58_1120 ();
 sg13g2_fill_2 FILLER_58_1145 ();
 sg13g2_fill_2 FILLER_58_1155 ();
 sg13g2_fill_1 FILLER_58_1165 ();
 sg13g2_fill_1 FILLER_58_1170 ();
 sg13g2_fill_1 FILLER_58_1179 ();
 sg13g2_fill_1 FILLER_58_1185 ();
 sg13g2_fill_1 FILLER_58_1194 ();
 sg13g2_fill_1 FILLER_58_1199 ();
 sg13g2_fill_1 FILLER_58_1217 ();
 sg13g2_fill_1 FILLER_58_1223 ();
 sg13g2_decap_4 FILLER_58_1235 ();
 sg13g2_fill_1 FILLER_58_1273 ();
 sg13g2_fill_1 FILLER_58_1278 ();
 sg13g2_fill_1 FILLER_58_1283 ();
 sg13g2_fill_1 FILLER_58_1293 ();
 sg13g2_fill_1 FILLER_58_1300 ();
 sg13g2_fill_1 FILLER_58_1311 ();
 sg13g2_fill_2 FILLER_58_1317 ();
 sg13g2_fill_1 FILLER_58_1319 ();
 sg13g2_fill_2 FILLER_58_1336 ();
 sg13g2_fill_1 FILLER_58_1338 ();
 sg13g2_fill_1 FILLER_58_1376 ();
 sg13g2_fill_2 FILLER_58_1381 ();
 sg13g2_fill_2 FILLER_58_1387 ();
 sg13g2_fill_2 FILLER_58_1393 ();
 sg13g2_fill_1 FILLER_58_1395 ();
 sg13g2_fill_1 FILLER_58_1424 ();
 sg13g2_decap_4 FILLER_58_1433 ();
 sg13g2_fill_2 FILLER_58_1437 ();
 sg13g2_fill_2 FILLER_58_1447 ();
 sg13g2_fill_1 FILLER_58_1449 ();
 sg13g2_fill_1 FILLER_58_1480 ();
 sg13g2_fill_2 FILLER_58_1501 ();
 sg13g2_fill_2 FILLER_58_1507 ();
 sg13g2_fill_1 FILLER_58_1509 ();
 sg13g2_fill_2 FILLER_58_1523 ();
 sg13g2_fill_1 FILLER_58_1533 ();
 sg13g2_decap_8 FILLER_58_1547 ();
 sg13g2_fill_1 FILLER_58_1554 ();
 sg13g2_fill_2 FILLER_58_1606 ();
 sg13g2_fill_2 FILLER_58_1612 ();
 sg13g2_fill_2 FILLER_58_1664 ();
 sg13g2_fill_1 FILLER_58_1670 ();
 sg13g2_fill_1 FILLER_58_1691 ();
 sg13g2_fill_1 FILLER_58_1713 ();
 sg13g2_fill_2 FILLER_58_1735 ();
 sg13g2_fill_1 FILLER_58_1761 ();
 sg13g2_fill_2 FILLER_58_1772 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_11 ();
 sg13g2_fill_2 FILLER_59_23 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_106 ();
 sg13g2_fill_1 FILLER_59_117 ();
 sg13g2_fill_1 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_229 ();
 sg13g2_fill_2 FILLER_59_247 ();
 sg13g2_fill_2 FILLER_59_259 ();
 sg13g2_fill_1 FILLER_59_297 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_fill_2 FILLER_59_419 ();
 sg13g2_fill_1 FILLER_59_425 ();
 sg13g2_fill_2 FILLER_59_436 ();
 sg13g2_fill_1 FILLER_59_480 ();
 sg13g2_fill_1 FILLER_59_537 ();
 sg13g2_fill_2 FILLER_59_559 ();
 sg13g2_fill_2 FILLER_59_584 ();
 sg13g2_fill_2 FILLER_59_607 ();
 sg13g2_fill_1 FILLER_59_613 ();
 sg13g2_decap_4 FILLER_59_626 ();
 sg13g2_fill_2 FILLER_59_630 ();
 sg13g2_fill_1 FILLER_59_639 ();
 sg13g2_fill_1 FILLER_59_647 ();
 sg13g2_fill_1 FILLER_59_697 ();
 sg13g2_decap_4 FILLER_59_737 ();
 sg13g2_fill_2 FILLER_59_741 ();
 sg13g2_fill_2 FILLER_59_781 ();
 sg13g2_fill_1 FILLER_59_791 ();
 sg13g2_fill_2 FILLER_59_800 ();
 sg13g2_fill_1 FILLER_59_838 ();
 sg13g2_decap_4 FILLER_59_843 ();
 sg13g2_fill_2 FILLER_59_851 ();
 sg13g2_fill_1 FILLER_59_922 ();
 sg13g2_fill_1 FILLER_59_988 ();
 sg13g2_fill_2 FILLER_59_1002 ();
 sg13g2_fill_2 FILLER_59_1029 ();
 sg13g2_decap_8 FILLER_59_1041 ();
 sg13g2_fill_1 FILLER_59_1048 ();
 sg13g2_fill_1 FILLER_59_1073 ();
 sg13g2_fill_2 FILLER_59_1079 ();
 sg13g2_fill_1 FILLER_59_1081 ();
 sg13g2_fill_2 FILLER_59_1095 ();
 sg13g2_fill_1 FILLER_59_1097 ();
 sg13g2_fill_1 FILLER_59_1157 ();
 sg13g2_fill_2 FILLER_59_1162 ();
 sg13g2_fill_2 FILLER_59_1169 ();
 sg13g2_fill_2 FILLER_59_1175 ();
 sg13g2_fill_1 FILLER_59_1181 ();
 sg13g2_fill_2 FILLER_59_1190 ();
 sg13g2_decap_8 FILLER_59_1229 ();
 sg13g2_decap_4 FILLER_59_1244 ();
 sg13g2_decap_8 FILLER_59_1261 ();
 sg13g2_decap_4 FILLER_59_1268 ();
 sg13g2_fill_2 FILLER_59_1272 ();
 sg13g2_fill_2 FILLER_59_1295 ();
 sg13g2_fill_1 FILLER_59_1297 ();
 sg13g2_fill_2 FILLER_59_1337 ();
 sg13g2_fill_1 FILLER_59_1352 ();
 sg13g2_fill_2 FILLER_59_1381 ();
 sg13g2_fill_2 FILLER_59_1396 ();
 sg13g2_fill_2 FILLER_59_1403 ();
 sg13g2_fill_1 FILLER_59_1409 ();
 sg13g2_fill_1 FILLER_59_1418 ();
 sg13g2_fill_1 FILLER_59_1424 ();
 sg13g2_decap_4 FILLER_59_1451 ();
 sg13g2_fill_1 FILLER_59_1459 ();
 sg13g2_fill_1 FILLER_59_1468 ();
 sg13g2_fill_1 FILLER_59_1479 ();
 sg13g2_decap_4 FILLER_59_1492 ();
 sg13g2_fill_2 FILLER_59_1496 ();
 sg13g2_fill_1 FILLER_59_1521 ();
 sg13g2_decap_4 FILLER_59_1526 ();
 sg13g2_fill_2 FILLER_59_1530 ();
 sg13g2_decap_4 FILLER_59_1540 ();
 sg13g2_fill_2 FILLER_59_1544 ();
 sg13g2_fill_2 FILLER_59_1576 ();
 sg13g2_fill_1 FILLER_59_1591 ();
 sg13g2_decap_4 FILLER_59_1607 ();
 sg13g2_fill_1 FILLER_59_1649 ();
 sg13g2_fill_2 FILLER_59_1666 ();
 sg13g2_fill_2 FILLER_59_1676 ();
 sg13g2_fill_1 FILLER_59_1686 ();
 sg13g2_fill_1 FILLER_59_1692 ();
 sg13g2_fill_2 FILLER_59_1701 ();
 sg13g2_fill_2 FILLER_59_1707 ();
 sg13g2_decap_8 FILLER_59_1712 ();
 sg13g2_fill_2 FILLER_59_1719 ();
 sg13g2_fill_1 FILLER_59_1721 ();
 sg13g2_decap_8 FILLER_59_1735 ();
 sg13g2_fill_2 FILLER_59_1742 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_157 ();
 sg13g2_fill_1 FILLER_60_214 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_fill_2 FILLER_60_334 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_1 FILLER_60_373 ();
 sg13g2_fill_2 FILLER_60_380 ();
 sg13g2_fill_2 FILLER_60_387 ();
 sg13g2_fill_2 FILLER_60_393 ();
 sg13g2_fill_1 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_470 ();
 sg13g2_fill_1 FILLER_60_512 ();
 sg13g2_decap_4 FILLER_60_523 ();
 sg13g2_fill_2 FILLER_60_527 ();
 sg13g2_decap_8 FILLER_60_541 ();
 sg13g2_decap_8 FILLER_60_548 ();
 sg13g2_fill_2 FILLER_60_555 ();
 sg13g2_fill_1 FILLER_60_557 ();
 sg13g2_fill_1 FILLER_60_563 ();
 sg13g2_fill_1 FILLER_60_570 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_fill_2 FILLER_60_594 ();
 sg13g2_fill_2 FILLER_60_616 ();
 sg13g2_fill_1 FILLER_60_627 ();
 sg13g2_fill_1 FILLER_60_664 ();
 sg13g2_fill_1 FILLER_60_675 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_fill_2 FILLER_60_697 ();
 sg13g2_fill_1 FILLER_60_713 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_4 FILLER_60_759 ();
 sg13g2_fill_1 FILLER_60_763 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_fill_2 FILLER_60_782 ();
 sg13g2_fill_1 FILLER_60_784 ();
 sg13g2_fill_1 FILLER_60_799 ();
 sg13g2_decap_4 FILLER_60_810 ();
 sg13g2_fill_1 FILLER_60_814 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_fill_2 FILLER_60_834 ();
 sg13g2_fill_1 FILLER_60_836 ();
 sg13g2_decap_4 FILLER_60_840 ();
 sg13g2_fill_1 FILLER_60_844 ();
 sg13g2_fill_1 FILLER_60_849 ();
 sg13g2_fill_2 FILLER_60_872 ();
 sg13g2_fill_1 FILLER_60_882 ();
 sg13g2_fill_1 FILLER_60_891 ();
 sg13g2_fill_1 FILLER_60_897 ();
 sg13g2_fill_1 FILLER_60_955 ();
 sg13g2_fill_1 FILLER_60_960 ();
 sg13g2_fill_1 FILLER_60_965 ();
 sg13g2_fill_2 FILLER_60_971 ();
 sg13g2_fill_1 FILLER_60_982 ();
 sg13g2_fill_2 FILLER_60_1037 ();
 sg13g2_fill_1 FILLER_60_1039 ();
 sg13g2_fill_1 FILLER_60_1044 ();
 sg13g2_fill_2 FILLER_60_1062 ();
 sg13g2_fill_1 FILLER_60_1064 ();
 sg13g2_fill_1 FILLER_60_1069 ();
 sg13g2_fill_1 FILLER_60_1085 ();
 sg13g2_decap_4 FILLER_60_1102 ();
 sg13g2_fill_1 FILLER_60_1106 ();
 sg13g2_fill_1 FILLER_60_1119 ();
 sg13g2_fill_1 FILLER_60_1125 ();
 sg13g2_decap_4 FILLER_60_1130 ();
 sg13g2_fill_1 FILLER_60_1134 ();
 sg13g2_fill_2 FILLER_60_1176 ();
 sg13g2_fill_2 FILLER_60_1211 ();
 sg13g2_fill_1 FILLER_60_1223 ();
 sg13g2_fill_2 FILLER_60_1245 ();
 sg13g2_fill_1 FILLER_60_1255 ();
 sg13g2_fill_2 FILLER_60_1262 ();
 sg13g2_fill_1 FILLER_60_1264 ();
 sg13g2_fill_1 FILLER_60_1318 ();
 sg13g2_fill_1 FILLER_60_1323 ();
 sg13g2_fill_1 FILLER_60_1332 ();
 sg13g2_decap_8 FILLER_60_1341 ();
 sg13g2_decap_8 FILLER_60_1348 ();
 sg13g2_fill_2 FILLER_60_1360 ();
 sg13g2_fill_1 FILLER_60_1374 ();
 sg13g2_fill_1 FILLER_60_1422 ();
 sg13g2_fill_1 FILLER_60_1431 ();
 sg13g2_fill_1 FILLER_60_1437 ();
 sg13g2_decap_4 FILLER_60_1453 ();
 sg13g2_fill_1 FILLER_60_1457 ();
 sg13g2_decap_8 FILLER_60_1490 ();
 sg13g2_decap_4 FILLER_60_1497 ();
 sg13g2_fill_1 FILLER_60_1501 ();
 sg13g2_fill_2 FILLER_60_1518 ();
 sg13g2_fill_1 FILLER_60_1520 ();
 sg13g2_decap_8 FILLER_60_1533 ();
 sg13g2_fill_2 FILLER_60_1540 ();
 sg13g2_fill_1 FILLER_60_1547 ();
 sg13g2_fill_1 FILLER_60_1564 ();
 sg13g2_decap_8 FILLER_60_1570 ();
 sg13g2_fill_1 FILLER_60_1577 ();
 sg13g2_fill_2 FILLER_60_1587 ();
 sg13g2_fill_1 FILLER_60_1589 ();
 sg13g2_decap_4 FILLER_60_1602 ();
 sg13g2_fill_2 FILLER_60_1615 ();
 sg13g2_fill_1 FILLER_60_1617 ();
 sg13g2_decap_8 FILLER_60_1622 ();
 sg13g2_fill_2 FILLER_60_1629 ();
 sg13g2_fill_1 FILLER_60_1631 ();
 sg13g2_decap_8 FILLER_60_1648 ();
 sg13g2_fill_2 FILLER_60_1655 ();
 sg13g2_fill_1 FILLER_60_1657 ();
 sg13g2_decap_4 FILLER_60_1682 ();
 sg13g2_fill_2 FILLER_60_1686 ();
 sg13g2_fill_1 FILLER_60_1692 ();
 sg13g2_fill_1 FILLER_60_1698 ();
 sg13g2_fill_1 FILLER_60_1711 ();
 sg13g2_fill_1 FILLER_60_1720 ();
 sg13g2_fill_1 FILLER_60_1729 ();
 sg13g2_fill_1 FILLER_60_1734 ();
 sg13g2_fill_2 FILLER_60_1751 ();
 sg13g2_fill_1 FILLER_60_1753 ();
 sg13g2_fill_1 FILLER_60_1762 ();
 sg13g2_fill_2 FILLER_60_1772 ();
 sg13g2_fill_2 FILLER_61_153 ();
 sg13g2_fill_2 FILLER_61_168 ();
 sg13g2_fill_1 FILLER_61_218 ();
 sg13g2_fill_1 FILLER_61_225 ();
 sg13g2_fill_1 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_258 ();
 sg13g2_fill_1 FILLER_61_332 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_426 ();
 sg13g2_fill_1 FILLER_61_443 ();
 sg13g2_fill_1 FILLER_61_599 ();
 sg13g2_fill_1 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_618 ();
 sg13g2_fill_2 FILLER_61_666 ();
 sg13g2_fill_1 FILLER_61_700 ();
 sg13g2_fill_2 FILLER_61_714 ();
 sg13g2_decap_4 FILLER_61_762 ();
 sg13g2_fill_1 FILLER_61_766 ();
 sg13g2_fill_2 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_815 ();
 sg13g2_fill_2 FILLER_61_822 ();
 sg13g2_fill_1 FILLER_61_824 ();
 sg13g2_fill_2 FILLER_61_851 ();
 sg13g2_fill_2 FILLER_61_857 ();
 sg13g2_fill_1 FILLER_61_864 ();
 sg13g2_fill_1 FILLER_61_910 ();
 sg13g2_fill_2 FILLER_61_952 ();
 sg13g2_fill_1 FILLER_61_987 ();
 sg13g2_fill_1 FILLER_61_1005 ();
 sg13g2_fill_1 FILLER_61_1013 ();
 sg13g2_fill_1 FILLER_61_1019 ();
 sg13g2_fill_2 FILLER_61_1057 ();
 sg13g2_fill_1 FILLER_61_1059 ();
 sg13g2_decap_8 FILLER_61_1065 ();
 sg13g2_decap_4 FILLER_61_1072 ();
 sg13g2_fill_2 FILLER_61_1076 ();
 sg13g2_decap_4 FILLER_61_1088 ();
 sg13g2_fill_2 FILLER_61_1092 ();
 sg13g2_decap_8 FILLER_61_1107 ();
 sg13g2_decap_4 FILLER_61_1122 ();
 sg13g2_fill_2 FILLER_61_1134 ();
 sg13g2_decap_8 FILLER_61_1151 ();
 sg13g2_fill_2 FILLER_61_1158 ();
 sg13g2_fill_1 FILLER_61_1173 ();
 sg13g2_fill_2 FILLER_61_1191 ();
 sg13g2_fill_2 FILLER_61_1213 ();
 sg13g2_fill_1 FILLER_61_1223 ();
 sg13g2_fill_1 FILLER_61_1229 ();
 sg13g2_fill_1 FILLER_61_1246 ();
 sg13g2_fill_1 FILLER_61_1252 ();
 sg13g2_fill_1 FILLER_61_1260 ();
 sg13g2_decap_4 FILLER_61_1273 ();
 sg13g2_fill_1 FILLER_61_1277 ();
 sg13g2_decap_4 FILLER_61_1283 ();
 sg13g2_fill_1 FILLER_61_1287 ();
 sg13g2_fill_1 FILLER_61_1292 ();
 sg13g2_fill_2 FILLER_61_1313 ();
 sg13g2_fill_1 FILLER_61_1319 ();
 sg13g2_fill_2 FILLER_61_1326 ();
 sg13g2_fill_1 FILLER_61_1353 ();
 sg13g2_decap_4 FILLER_61_1361 ();
 sg13g2_fill_2 FILLER_61_1369 ();
 sg13g2_fill_2 FILLER_61_1393 ();
 sg13g2_fill_1 FILLER_61_1395 ();
 sg13g2_fill_1 FILLER_61_1420 ();
 sg13g2_decap_8 FILLER_61_1441 ();
 sg13g2_decap_8 FILLER_61_1448 ();
 sg13g2_fill_2 FILLER_61_1455 ();
 sg13g2_fill_1 FILLER_61_1461 ();
 sg13g2_fill_1 FILLER_61_1466 ();
 sg13g2_fill_1 FILLER_61_1488 ();
 sg13g2_decap_8 FILLER_61_1493 ();
 sg13g2_decap_4 FILLER_61_1500 ();
 sg13g2_fill_2 FILLER_61_1504 ();
 sg13g2_decap_8 FILLER_61_1510 ();
 sg13g2_fill_1 FILLER_61_1517 ();
 sg13g2_decap_4 FILLER_61_1538 ();
 sg13g2_fill_1 FILLER_61_1554 ();
 sg13g2_fill_1 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1575 ();
 sg13g2_fill_1 FILLER_61_1596 ();
 sg13g2_fill_2 FILLER_61_1601 ();
 sg13g2_fill_1 FILLER_61_1627 ();
 sg13g2_fill_1 FILLER_61_1645 ();
 sg13g2_fill_2 FILLER_61_1650 ();
 sg13g2_fill_2 FILLER_61_1660 ();
 sg13g2_decap_8 FILLER_61_1672 ();
 sg13g2_decap_8 FILLER_61_1703 ();
 sg13g2_decap_4 FILLER_61_1710 ();
 sg13g2_fill_1 FILLER_61_1721 ();
 sg13g2_fill_1 FILLER_61_1730 ();
 sg13g2_fill_2 FILLER_61_1747 ();
 sg13g2_fill_1 FILLER_61_1749 ();
 sg13g2_fill_2 FILLER_61_1766 ();
 sg13g2_fill_2 FILLER_61_1771 ();
 sg13g2_fill_1 FILLER_61_1773 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_154 ();
 sg13g2_fill_2 FILLER_62_181 ();
 sg13g2_fill_1 FILLER_62_187 ();
 sg13g2_fill_2 FILLER_62_214 ();
 sg13g2_fill_1 FILLER_62_226 ();
 sg13g2_fill_1 FILLER_62_231 ();
 sg13g2_fill_1 FILLER_62_242 ();
 sg13g2_fill_1 FILLER_62_269 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_1 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_fill_1 FILLER_62_433 ();
 sg13g2_fill_1 FILLER_62_482 ();
 sg13g2_fill_1 FILLER_62_600 ();
 sg13g2_fill_1 FILLER_62_611 ();
 sg13g2_fill_2 FILLER_62_673 ();
 sg13g2_fill_1 FILLER_62_680 ();
 sg13g2_fill_1 FILLER_62_690 ();
 sg13g2_fill_1 FILLER_62_696 ();
 sg13g2_fill_1 FILLER_62_718 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_fill_2 FILLER_62_732 ();
 sg13g2_fill_2 FILLER_62_742 ();
 sg13g2_fill_2 FILLER_62_749 ();
 sg13g2_fill_1 FILLER_62_751 ();
 sg13g2_fill_1 FILLER_62_843 ();
 sg13g2_fill_2 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_855 ();
 sg13g2_fill_2 FILLER_62_862 ();
 sg13g2_fill_1 FILLER_62_864 ();
 sg13g2_fill_2 FILLER_62_870 ();
 sg13g2_fill_1 FILLER_62_872 ();
 sg13g2_fill_2 FILLER_62_877 ();
 sg13g2_fill_1 FILLER_62_896 ();
 sg13g2_fill_2 FILLER_62_955 ();
 sg13g2_fill_2 FILLER_62_979 ();
 sg13g2_fill_1 FILLER_62_1019 ();
 sg13g2_decap_8 FILLER_62_1037 ();
 sg13g2_decap_4 FILLER_62_1044 ();
 sg13g2_fill_1 FILLER_62_1048 ();
 sg13g2_fill_2 FILLER_62_1062 ();
 sg13g2_fill_2 FILLER_62_1088 ();
 sg13g2_fill_2 FILLER_62_1124 ();
 sg13g2_fill_1 FILLER_62_1126 ();
 sg13g2_fill_1 FILLER_62_1139 ();
 sg13g2_fill_2 FILLER_62_1148 ();
 sg13g2_fill_2 FILLER_62_1168 ();
 sg13g2_fill_2 FILLER_62_1177 ();
 sg13g2_fill_1 FILLER_62_1179 ();
 sg13g2_fill_1 FILLER_62_1211 ();
 sg13g2_fill_1 FILLER_62_1226 ();
 sg13g2_fill_2 FILLER_62_1294 ();
 sg13g2_fill_1 FILLER_62_1296 ();
 sg13g2_fill_1 FILLER_62_1312 ();
 sg13g2_fill_1 FILLER_62_1341 ();
 sg13g2_fill_1 FILLER_62_1357 ();
 sg13g2_fill_2 FILLER_62_1363 ();
 sg13g2_fill_2 FILLER_62_1369 ();
 sg13g2_fill_2 FILLER_62_1384 ();
 sg13g2_fill_2 FILLER_62_1391 ();
 sg13g2_fill_1 FILLER_62_1406 ();
 sg13g2_fill_1 FILLER_62_1412 ();
 sg13g2_fill_1 FILLER_62_1421 ();
 sg13g2_decap_8 FILLER_62_1445 ();
 sg13g2_decap_8 FILLER_62_1452 ();
 sg13g2_fill_2 FILLER_62_1459 ();
 sg13g2_fill_2 FILLER_62_1496 ();
 sg13g2_fill_2 FILLER_62_1536 ();
 sg13g2_fill_1 FILLER_62_1538 ();
 sg13g2_fill_2 FILLER_62_1551 ();
 sg13g2_fill_1 FILLER_62_1553 ();
 sg13g2_fill_2 FILLER_62_1566 ();
 sg13g2_fill_1 FILLER_62_1610 ();
 sg13g2_fill_2 FILLER_62_1631 ();
 sg13g2_fill_1 FILLER_62_1649 ();
 sg13g2_fill_1 FILLER_62_1654 ();
 sg13g2_fill_2 FILLER_62_1690 ();
 sg13g2_fill_1 FILLER_62_1696 ();
 sg13g2_decap_4 FILLER_62_1705 ();
 sg13g2_fill_2 FILLER_62_1709 ();
 sg13g2_fill_2 FILLER_62_1745 ();
 sg13g2_fill_1 FILLER_62_1747 ();
 sg13g2_decap_4 FILLER_62_1769 ();
 sg13g2_fill_1 FILLER_62_1773 ();
 sg13g2_fill_2 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_97 ();
 sg13g2_fill_1 FILLER_63_158 ();
 sg13g2_fill_2 FILLER_63_176 ();
 sg13g2_fill_2 FILLER_63_191 ();
 sg13g2_fill_1 FILLER_63_197 ();
 sg13g2_fill_1 FILLER_63_219 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_256 ();
 sg13g2_fill_2 FILLER_63_267 ();
 sg13g2_fill_2 FILLER_63_298 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_1 FILLER_63_393 ();
 sg13g2_fill_2 FILLER_63_418 ();
 sg13g2_fill_1 FILLER_63_577 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_640 ();
 sg13g2_fill_1 FILLER_63_671 ();
 sg13g2_fill_1 FILLER_63_677 ();
 sg13g2_fill_1 FILLER_63_704 ();
 sg13g2_fill_1 FILLER_63_709 ();
 sg13g2_fill_1 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_760 ();
 sg13g2_fill_1 FILLER_63_807 ();
 sg13g2_decap_4 FILLER_63_836 ();
 sg13g2_fill_2 FILLER_63_840 ();
 sg13g2_fill_2 FILLER_63_861 ();
 sg13g2_fill_1 FILLER_63_863 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_decap_8 FILLER_63_875 ();
 sg13g2_fill_1 FILLER_63_882 ();
 sg13g2_decap_4 FILLER_63_899 ();
 sg13g2_decap_4 FILLER_63_916 ();
 sg13g2_fill_1 FILLER_63_920 ();
 sg13g2_fill_2 FILLER_63_951 ();
 sg13g2_fill_2 FILLER_63_1013 ();
 sg13g2_fill_1 FILLER_63_1015 ();
 sg13g2_fill_1 FILLER_63_1073 ();
 sg13g2_fill_1 FILLER_63_1078 ();
 sg13g2_fill_2 FILLER_63_1086 ();
 sg13g2_fill_1 FILLER_63_1088 ();
 sg13g2_decap_8 FILLER_63_1097 ();
 sg13g2_fill_1 FILLER_63_1149 ();
 sg13g2_fill_1 FILLER_63_1164 ();
 sg13g2_decap_4 FILLER_63_1179 ();
 sg13g2_fill_1 FILLER_63_1189 ();
 sg13g2_decap_8 FILLER_63_1200 ();
 sg13g2_fill_2 FILLER_63_1207 ();
 sg13g2_fill_1 FILLER_63_1221 ();
 sg13g2_fill_1 FILLER_63_1230 ();
 sg13g2_fill_1 FILLER_63_1260 ();
 sg13g2_fill_1 FILLER_63_1266 ();
 sg13g2_fill_1 FILLER_63_1272 ();
 sg13g2_fill_1 FILLER_63_1278 ();
 sg13g2_fill_2 FILLER_63_1303 ();
 sg13g2_decap_8 FILLER_63_1309 ();
 sg13g2_fill_1 FILLER_63_1316 ();
 sg13g2_fill_1 FILLER_63_1322 ();
 sg13g2_fill_1 FILLER_63_1333 ();
 sg13g2_fill_2 FILLER_63_1340 ();
 sg13g2_fill_1 FILLER_63_1346 ();
 sg13g2_fill_2 FILLER_63_1355 ();
 sg13g2_fill_2 FILLER_63_1361 ();
 sg13g2_fill_1 FILLER_63_1363 ();
 sg13g2_decap_4 FILLER_63_1369 ();
 sg13g2_decap_4 FILLER_63_1381 ();
 sg13g2_fill_1 FILLER_63_1385 ();
 sg13g2_fill_1 FILLER_63_1390 ();
 sg13g2_fill_1 FILLER_63_1399 ();
 sg13g2_fill_1 FILLER_63_1409 ();
 sg13g2_fill_1 FILLER_63_1418 ();
 sg13g2_decap_4 FILLER_63_1432 ();
 sg13g2_fill_2 FILLER_63_1473 ();
 sg13g2_fill_1 FILLER_63_1475 ();
 sg13g2_fill_1 FILLER_63_1536 ();
 sg13g2_fill_2 FILLER_63_1571 ();
 sg13g2_fill_1 FILLER_63_1573 ();
 sg13g2_decap_8 FILLER_63_1578 ();
 sg13g2_fill_2 FILLER_63_1585 ();
 sg13g2_fill_1 FILLER_63_1595 ();
 sg13g2_decap_8 FILLER_63_1605 ();
 sg13g2_decap_4 FILLER_63_1612 ();
 sg13g2_fill_2 FILLER_63_1628 ();
 sg13g2_decap_8 FILLER_63_1680 ();
 sg13g2_fill_1 FILLER_63_1691 ();
 sg13g2_fill_2 FILLER_63_1737 ();
 sg13g2_fill_1 FILLER_63_1739 ();
 sg13g2_fill_2 FILLER_63_1758 ();
 sg13g2_fill_1 FILLER_63_1773 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_98 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_fill_2 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_fill_1 FILLER_64_144 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_fill_1 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_224 ();
 sg13g2_fill_1 FILLER_64_287 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_389 ();
 sg13g2_fill_2 FILLER_64_451 ();
 sg13g2_fill_1 FILLER_64_463 ();
 sg13g2_fill_1 FILLER_64_490 ();
 sg13g2_fill_1 FILLER_64_517 ();
 sg13g2_fill_2 FILLER_64_544 ();
 sg13g2_fill_2 FILLER_64_567 ();
 sg13g2_fill_2 FILLER_64_658 ();
 sg13g2_fill_1 FILLER_64_724 ();
 sg13g2_fill_1 FILLER_64_765 ();
 sg13g2_fill_1 FILLER_64_792 ();
 sg13g2_fill_2 FILLER_64_824 ();
 sg13g2_fill_1 FILLER_64_826 ();
 sg13g2_fill_1 FILLER_64_840 ();
 sg13g2_fill_1 FILLER_64_890 ();
 sg13g2_fill_2 FILLER_64_906 ();
 sg13g2_fill_1 FILLER_64_908 ();
 sg13g2_fill_1 FILLER_64_918 ();
 sg13g2_fill_2 FILLER_64_923 ();
 sg13g2_fill_2 FILLER_64_929 ();
 sg13g2_fill_2 FILLER_64_935 ();
 sg13g2_fill_1 FILLER_64_954 ();
 sg13g2_fill_2 FILLER_64_964 ();
 sg13g2_decap_4 FILLER_64_974 ();
 sg13g2_fill_1 FILLER_64_1008 ();
 sg13g2_decap_4 FILLER_64_1013 ();
 sg13g2_decap_4 FILLER_64_1021 ();
 sg13g2_fill_1 FILLER_64_1037 ();
 sg13g2_decap_8 FILLER_64_1042 ();
 sg13g2_fill_2 FILLER_64_1049 ();
 sg13g2_fill_2 FILLER_64_1062 ();
 sg13g2_fill_2 FILLER_64_1125 ();
 sg13g2_fill_1 FILLER_64_1137 ();
 sg13g2_fill_1 FILLER_64_1160 ();
 sg13g2_fill_1 FILLER_64_1165 ();
 sg13g2_fill_1 FILLER_64_1171 ();
 sg13g2_fill_2 FILLER_64_1176 ();
 sg13g2_decap_8 FILLER_64_1203 ();
 sg13g2_fill_2 FILLER_64_1210 ();
 sg13g2_fill_2 FILLER_64_1216 ();
 sg13g2_fill_1 FILLER_64_1218 ();
 sg13g2_fill_1 FILLER_64_1238 ();
 sg13g2_fill_1 FILLER_64_1253 ();
 sg13g2_fill_2 FILLER_64_1259 ();
 sg13g2_fill_1 FILLER_64_1265 ();
 sg13g2_fill_1 FILLER_64_1271 ();
 sg13g2_fill_2 FILLER_64_1304 ();
 sg13g2_fill_1 FILLER_64_1318 ();
 sg13g2_fill_1 FILLER_64_1331 ();
 sg13g2_fill_1 FILLER_64_1342 ();
 sg13g2_fill_1 FILLER_64_1386 ();
 sg13g2_fill_1 FILLER_64_1392 ();
 sg13g2_fill_1 FILLER_64_1401 ();
 sg13g2_fill_2 FILLER_64_1436 ();
 sg13g2_decap_8 FILLER_64_1466 ();
 sg13g2_decap_8 FILLER_64_1473 ();
 sg13g2_fill_2 FILLER_64_1480 ();
 sg13g2_decap_8 FILLER_64_1495 ();
 sg13g2_decap_8 FILLER_64_1502 ();
 sg13g2_decap_8 FILLER_64_1509 ();
 sg13g2_fill_2 FILLER_64_1529 ();
 sg13g2_fill_2 FILLER_64_1543 ();
 sg13g2_fill_2 FILLER_64_1553 ();
 sg13g2_decap_4 FILLER_64_1575 ();
 sg13g2_fill_1 FILLER_64_1603 ();
 sg13g2_fill_1 FILLER_64_1608 ();
 sg13g2_decap_8 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1633 ();
 sg13g2_fill_1 FILLER_64_1640 ();
 sg13g2_fill_2 FILLER_64_1649 ();
 sg13g2_fill_1 FILLER_64_1651 ();
 sg13g2_fill_1 FILLER_64_1693 ();
 sg13g2_fill_2 FILLER_64_1731 ();
 sg13g2_decap_4 FILLER_64_1741 ();
 sg13g2_decap_8 FILLER_64_1755 ();
 sg13g2_decap_4 FILLER_64_1770 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_1 FILLER_65_27 ();
 sg13g2_fill_1 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_133 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_fill_2 FILLER_65_222 ();
 sg13g2_fill_2 FILLER_65_241 ();
 sg13g2_fill_1 FILLER_65_283 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_407 ();
 sg13g2_fill_1 FILLER_65_413 ();
 sg13g2_fill_1 FILLER_65_458 ();
 sg13g2_fill_1 FILLER_65_471 ();
 sg13g2_fill_2 FILLER_65_476 ();
 sg13g2_fill_2 FILLER_65_488 ();
 sg13g2_fill_2 FILLER_65_494 ();
 sg13g2_fill_1 FILLER_65_501 ();
 sg13g2_fill_1 FILLER_65_509 ();
 sg13g2_fill_1 FILLER_65_634 ();
 sg13g2_fill_1 FILLER_65_670 ();
 sg13g2_fill_2 FILLER_65_676 ();
 sg13g2_fill_2 FILLER_65_697 ();
 sg13g2_fill_1 FILLER_65_768 ();
 sg13g2_fill_2 FILLER_65_830 ();
 sg13g2_fill_1 FILLER_65_832 ();
 sg13g2_fill_2 FILLER_65_850 ();
 sg13g2_fill_2 FILLER_65_867 ();
 sg13g2_fill_1 FILLER_65_873 ();
 sg13g2_fill_2 FILLER_65_878 ();
 sg13g2_fill_1 FILLER_65_923 ();
 sg13g2_fill_2 FILLER_65_929 ();
 sg13g2_fill_1 FILLER_65_965 ();
 sg13g2_fill_2 FILLER_65_971 ();
 sg13g2_fill_2 FILLER_65_977 ();
 sg13g2_fill_2 FILLER_65_983 ();
 sg13g2_fill_2 FILLER_65_1019 ();
 sg13g2_decap_4 FILLER_65_1070 ();
 sg13g2_decap_8 FILLER_65_1107 ();
 sg13g2_fill_1 FILLER_65_1114 ();
 sg13g2_decap_4 FILLER_65_1120 ();
 sg13g2_fill_1 FILLER_65_1124 ();
 sg13g2_fill_1 FILLER_65_1130 ();
 sg13g2_fill_1 FILLER_65_1135 ();
 sg13g2_fill_1 FILLER_65_1145 ();
 sg13g2_decap_4 FILLER_65_1154 ();
 sg13g2_fill_1 FILLER_65_1158 ();
 sg13g2_fill_2 FILLER_65_1188 ();
 sg13g2_fill_1 FILLER_65_1232 ();
 sg13g2_fill_1 FILLER_65_1291 ();
 sg13g2_fill_1 FILLER_65_1297 ();
 sg13g2_fill_1 FILLER_65_1302 ();
 sg13g2_fill_1 FILLER_65_1308 ();
 sg13g2_fill_2 FILLER_65_1336 ();
 sg13g2_fill_1 FILLER_65_1386 ();
 sg13g2_fill_1 FILLER_65_1430 ();
 sg13g2_fill_1 FILLER_65_1435 ();
 sg13g2_fill_1 FILLER_65_1441 ();
 sg13g2_fill_1 FILLER_65_1446 ();
 sg13g2_fill_2 FILLER_65_1471 ();
 sg13g2_fill_1 FILLER_65_1473 ();
 sg13g2_fill_2 FILLER_65_1490 ();
 sg13g2_fill_1 FILLER_65_1492 ();
 sg13g2_fill_1 FILLER_65_1518 ();
 sg13g2_fill_1 FILLER_65_1537 ();
 sg13g2_fill_1 FILLER_65_1542 ();
 sg13g2_fill_1 FILLER_65_1548 ();
 sg13g2_decap_4 FILLER_65_1553 ();
 sg13g2_fill_2 FILLER_65_1557 ();
 sg13g2_fill_1 FILLER_65_1594 ();
 sg13g2_fill_1 FILLER_65_1600 ();
 sg13g2_fill_1 FILLER_65_1628 ();
 sg13g2_decap_4 FILLER_65_1637 ();
 sg13g2_fill_2 FILLER_65_1658 ();
 sg13g2_fill_2 FILLER_65_1665 ();
 sg13g2_fill_1 FILLER_65_1667 ();
 sg13g2_fill_2 FILLER_65_1701 ();
 sg13g2_decap_8 FILLER_65_1713 ();
 sg13g2_decap_8 FILLER_65_1720 ();
 sg13g2_decap_4 FILLER_65_1732 ();
 sg13g2_fill_2 FILLER_65_1736 ();
 sg13g2_decap_4 FILLER_65_1755 ();
 sg13g2_fill_1 FILLER_65_1759 ();
 sg13g2_fill_2 FILLER_65_1764 ();
 sg13g2_fill_2 FILLER_66_66 ();
 sg13g2_fill_1 FILLER_66_89 ();
 sg13g2_fill_1 FILLER_66_133 ();
 sg13g2_fill_2 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_290 ();
 sg13g2_fill_2 FILLER_66_317 ();
 sg13g2_fill_2 FILLER_66_329 ();
 sg13g2_fill_2 FILLER_66_335 ();
 sg13g2_fill_2 FILLER_66_341 ();
 sg13g2_fill_1 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_384 ();
 sg13g2_fill_1 FILLER_66_395 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_2 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_464 ();
 sg13g2_fill_1 FILLER_66_597 ();
 sg13g2_fill_1 FILLER_66_606 ();
 sg13g2_fill_1 FILLER_66_617 ();
 sg13g2_fill_1 FILLER_66_633 ();
 sg13g2_fill_1 FILLER_66_660 ();
 sg13g2_fill_2 FILLER_66_718 ();
 sg13g2_fill_1 FILLER_66_728 ();
 sg13g2_fill_1 FILLER_66_743 ();
 sg13g2_fill_2 FILLER_66_754 ();
 sg13g2_fill_2 FILLER_66_806 ();
 sg13g2_fill_2 FILLER_66_989 ();
 sg13g2_fill_1 FILLER_66_991 ();
 sg13g2_fill_1 FILLER_66_1018 ();
 sg13g2_fill_1 FILLER_66_1023 ();
 sg13g2_decap_4 FILLER_66_1050 ();
 sg13g2_fill_2 FILLER_66_1078 ();
 sg13g2_decap_4 FILLER_66_1088 ();
 sg13g2_fill_1 FILLER_66_1092 ();
 sg13g2_fill_1 FILLER_66_1114 ();
 sg13g2_fill_1 FILLER_66_1127 ();
 sg13g2_fill_1 FILLER_66_1180 ();
 sg13g2_decap_4 FILLER_66_1195 ();
 sg13g2_fill_2 FILLER_66_1211 ();
 sg13g2_fill_1 FILLER_66_1213 ();
 sg13g2_fill_2 FILLER_66_1222 ();
 sg13g2_fill_1 FILLER_66_1224 ();
 sg13g2_fill_2 FILLER_66_1234 ();
 sg13g2_fill_2 FILLER_66_1247 ();
 sg13g2_decap_4 FILLER_66_1297 ();
 sg13g2_fill_1 FILLER_66_1301 ();
 sg13g2_fill_1 FILLER_66_1307 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_fill_2 FILLER_66_1352 ();
 sg13g2_fill_1 FILLER_66_1354 ();
 sg13g2_fill_2 FILLER_66_1391 ();
 sg13g2_fill_2 FILLER_66_1402 ();
 sg13g2_fill_2 FILLER_66_1409 ();
 sg13g2_fill_1 FILLER_66_1411 ();
 sg13g2_fill_1 FILLER_66_1417 ();
 sg13g2_fill_1 FILLER_66_1423 ();
 sg13g2_fill_1 FILLER_66_1432 ();
 sg13g2_fill_1 FILLER_66_1440 ();
 sg13g2_fill_2 FILLER_66_1446 ();
 sg13g2_fill_2 FILLER_66_1456 ();
 sg13g2_decap_8 FILLER_66_1461 ();
 sg13g2_decap_4 FILLER_66_1468 ();
 sg13g2_fill_2 FILLER_66_1472 ();
 sg13g2_decap_8 FILLER_66_1482 ();
 sg13g2_decap_4 FILLER_66_1489 ();
 sg13g2_fill_1 FILLER_66_1498 ();
 sg13g2_fill_1 FILLER_66_1520 ();
 sg13g2_fill_2 FILLER_66_1551 ();
 sg13g2_decap_4 FILLER_66_1561 ();
 sg13g2_fill_2 FILLER_66_1585 ();
 sg13g2_fill_2 FILLER_66_1591 ();
 sg13g2_fill_1 FILLER_66_1593 ();
 sg13g2_fill_1 FILLER_66_1602 ();
 sg13g2_fill_1 FILLER_66_1611 ();
 sg13g2_fill_1 FILLER_66_1620 ();
 sg13g2_fill_1 FILLER_66_1625 ();
 sg13g2_fill_1 FILLER_66_1630 ();
 sg13g2_fill_1 FILLER_66_1636 ();
 sg13g2_fill_1 FILLER_66_1641 ();
 sg13g2_fill_1 FILLER_66_1666 ();
 sg13g2_fill_2 FILLER_66_1686 ();
 sg13g2_decap_8 FILLER_66_1692 ();
 sg13g2_fill_1 FILLER_66_1720 ();
 sg13g2_decap_8 FILLER_66_1734 ();
 sg13g2_decap_4 FILLER_66_1749 ();
 sg13g2_fill_2 FILLER_66_1753 ();
 sg13g2_fill_2 FILLER_66_1764 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_120 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_1 FILLER_67_169 ();
 sg13g2_fill_1 FILLER_67_301 ();
 sg13g2_fill_2 FILLER_67_362 ();
 sg13g2_fill_2 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_67_442 ();
 sg13g2_fill_2 FILLER_67_523 ();
 sg13g2_fill_2 FILLER_67_545 ();
 sg13g2_fill_1 FILLER_67_574 ();
 sg13g2_fill_1 FILLER_67_594 ();
 sg13g2_fill_1 FILLER_67_621 ();
 sg13g2_fill_1 FILLER_67_647 ();
 sg13g2_fill_1 FILLER_67_652 ();
 sg13g2_fill_2 FILLER_67_663 ();
 sg13g2_fill_2 FILLER_67_686 ();
 sg13g2_fill_2 FILLER_67_765 ();
 sg13g2_fill_1 FILLER_67_793 ();
 sg13g2_decap_4 FILLER_67_807 ();
 sg13g2_fill_2 FILLER_67_824 ();
 sg13g2_fill_1 FILLER_67_826 ();
 sg13g2_fill_2 FILLER_67_879 ();
 sg13g2_fill_1 FILLER_67_933 ();
 sg13g2_fill_1 FILLER_67_938 ();
 sg13g2_fill_1 FILLER_67_943 ();
 sg13g2_fill_1 FILLER_67_948 ();
 sg13g2_fill_2 FILLER_67_961 ();
 sg13g2_fill_1 FILLER_67_963 ();
 sg13g2_fill_2 FILLER_67_1017 ();
 sg13g2_fill_1 FILLER_67_1052 ();
 sg13g2_fill_1 FILLER_67_1061 ();
 sg13g2_fill_2 FILLER_67_1066 ();
 sg13g2_fill_1 FILLER_67_1080 ();
 sg13g2_fill_1 FILLER_67_1097 ();
 sg13g2_fill_1 FILLER_67_1103 ();
 sg13g2_fill_2 FILLER_67_1112 ();
 sg13g2_fill_2 FILLER_67_1118 ();
 sg13g2_fill_1 FILLER_67_1120 ();
 sg13g2_fill_1 FILLER_67_1142 ();
 sg13g2_fill_2 FILLER_67_1151 ();
 sg13g2_decap_4 FILLER_67_1165 ();
 sg13g2_fill_2 FILLER_67_1169 ();
 sg13g2_fill_1 FILLER_67_1204 ();
 sg13g2_fill_2 FILLER_67_1245 ();
 sg13g2_fill_1 FILLER_67_1247 ();
 sg13g2_fill_1 FILLER_67_1257 ();
 sg13g2_fill_1 FILLER_67_1264 ();
 sg13g2_fill_2 FILLER_67_1270 ();
 sg13g2_fill_1 FILLER_67_1272 ();
 sg13g2_fill_1 FILLER_67_1295 ();
 sg13g2_fill_1 FILLER_67_1306 ();
 sg13g2_fill_2 FILLER_67_1340 ();
 sg13g2_fill_1 FILLER_67_1347 ();
 sg13g2_fill_1 FILLER_67_1357 ();
 sg13g2_decap_8 FILLER_67_1366 ();
 sg13g2_decap_8 FILLER_67_1383 ();
 sg13g2_decap_4 FILLER_67_1390 ();
 sg13g2_fill_2 FILLER_67_1394 ();
 sg13g2_decap_8 FILLER_67_1421 ();
 sg13g2_decap_4 FILLER_67_1428 ();
 sg13g2_fill_1 FILLER_67_1432 ();
 sg13g2_fill_2 FILLER_67_1449 ();
 sg13g2_fill_2 FILLER_67_1473 ();
 sg13g2_fill_1 FILLER_67_1500 ();
 sg13g2_decap_8 FILLER_67_1524 ();
 sg13g2_decap_4 FILLER_67_1531 ();
 sg13g2_decap_4 FILLER_67_1539 ();
 sg13g2_decap_8 FILLER_67_1547 ();
 sg13g2_fill_1 FILLER_67_1554 ();
 sg13g2_decap_8 FILLER_67_1559 ();
 sg13g2_fill_2 FILLER_67_1566 ();
 sg13g2_fill_1 FILLER_67_1613 ();
 sg13g2_fill_1 FILLER_67_1622 ();
 sg13g2_fill_2 FILLER_67_1654 ();
 sg13g2_fill_1 FILLER_67_1656 ();
 sg13g2_fill_2 FILLER_67_1669 ();
 sg13g2_fill_2 FILLER_67_1679 ();
 sg13g2_fill_2 FILLER_67_1689 ();
 sg13g2_fill_1 FILLER_67_1707 ();
 sg13g2_fill_1 FILLER_67_1732 ();
 sg13g2_fill_2 FILLER_67_1741 ();
 sg13g2_fill_2 FILLER_67_1751 ();
 sg13g2_fill_2 FILLER_67_1761 ();
 sg13g2_fill_2 FILLER_67_1771 ();
 sg13g2_fill_1 FILLER_67_1773 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_20 ();
 sg13g2_fill_1 FILLER_68_74 ();
 sg13g2_fill_2 FILLER_68_105 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_fill_1 FILLER_68_278 ();
 sg13g2_fill_1 FILLER_68_369 ();
 sg13g2_fill_1 FILLER_68_400 ();
 sg13g2_fill_1 FILLER_68_406 ();
 sg13g2_fill_2 FILLER_68_421 ();
 sg13g2_fill_1 FILLER_68_462 ();
 sg13g2_fill_1 FILLER_68_489 ();
 sg13g2_fill_1 FILLER_68_500 ();
 sg13g2_fill_1 FILLER_68_511 ();
 sg13g2_fill_1 FILLER_68_533 ();
 sg13g2_fill_2 FILLER_68_560 ();
 sg13g2_fill_1 FILLER_68_628 ();
 sg13g2_fill_1 FILLER_68_668 ();
 sg13g2_fill_2 FILLER_68_676 ();
 sg13g2_fill_1 FILLER_68_764 ();
 sg13g2_fill_2 FILLER_68_770 ();
 sg13g2_decap_4 FILLER_68_813 ();
 sg13g2_decap_4 FILLER_68_846 ();
 sg13g2_fill_2 FILLER_68_857 ();
 sg13g2_fill_1 FILLER_68_893 ();
 sg13g2_fill_2 FILLER_68_933 ();
 sg13g2_fill_2 FILLER_68_1038 ();
 sg13g2_fill_2 FILLER_68_1048 ();
 sg13g2_fill_2 FILLER_68_1058 ();
 sg13g2_fill_2 FILLER_68_1064 ();
 sg13g2_fill_1 FILLER_68_1074 ();
 sg13g2_decap_4 FILLER_68_1088 ();
 sg13g2_fill_2 FILLER_68_1092 ();
 sg13g2_fill_1 FILLER_68_1102 ();
 sg13g2_fill_1 FILLER_68_1107 ();
 sg13g2_fill_1 FILLER_68_1112 ();
 sg13g2_fill_1 FILLER_68_1121 ();
 sg13g2_fill_2 FILLER_68_1126 ();
 sg13g2_fill_2 FILLER_68_1153 ();
 sg13g2_fill_2 FILLER_68_1174 ();
 sg13g2_fill_1 FILLER_68_1185 ();
 sg13g2_fill_1 FILLER_68_1200 ();
 sg13g2_fill_1 FILLER_68_1213 ();
 sg13g2_fill_1 FILLER_68_1219 ();
 sg13g2_fill_2 FILLER_68_1245 ();
 sg13g2_fill_1 FILLER_68_1247 ();
 sg13g2_fill_1 FILLER_68_1261 ();
 sg13g2_fill_2 FILLER_68_1269 ();
 sg13g2_fill_2 FILLER_68_1296 ();
 sg13g2_fill_1 FILLER_68_1298 ();
 sg13g2_fill_2 FILLER_68_1311 ();
 sg13g2_fill_1 FILLER_68_1313 ();
 sg13g2_fill_2 FILLER_68_1319 ();
 sg13g2_fill_1 FILLER_68_1346 ();
 sg13g2_fill_1 FILLER_68_1367 ();
 sg13g2_fill_2 FILLER_68_1388 ();
 sg13g2_fill_2 FILLER_68_1395 ();
 sg13g2_fill_1 FILLER_68_1402 ();
 sg13g2_fill_2 FILLER_68_1419 ();
 sg13g2_decap_4 FILLER_68_1425 ();
 sg13g2_fill_2 FILLER_68_1429 ();
 sg13g2_fill_2 FILLER_68_1499 ();
 sg13g2_fill_1 FILLER_68_1501 ();
 sg13g2_fill_2 FILLER_68_1515 ();
 sg13g2_decap_8 FILLER_68_1525 ();
 sg13g2_decap_4 FILLER_68_1532 ();
 sg13g2_fill_1 FILLER_68_1536 ();
 sg13g2_fill_1 FILLER_68_1549 ();
 sg13g2_decap_4 FILLER_68_1559 ();
 sg13g2_fill_1 FILLER_68_1591 ();
 sg13g2_fill_1 FILLER_68_1603 ();
 sg13g2_fill_2 FILLER_68_1608 ();
 sg13g2_fill_2 FILLER_68_1614 ();
 sg13g2_fill_2 FILLER_68_1624 ();
 sg13g2_fill_1 FILLER_68_1626 ();
 sg13g2_fill_1 FILLER_68_1635 ();
 sg13g2_fill_2 FILLER_68_1648 ();
 sg13g2_fill_1 FILLER_68_1650 ();
 sg13g2_fill_2 FILLER_68_1674 ();
 sg13g2_fill_1 FILLER_68_1676 ();
 sg13g2_fill_1 FILLER_68_1681 ();
 sg13g2_fill_1 FILLER_68_1691 ();
 sg13g2_decap_8 FILLER_68_1697 ();
 sg13g2_fill_2 FILLER_68_1704 ();
 sg13g2_fill_1 FILLER_68_1706 ();
 sg13g2_decap_8 FILLER_68_1715 ();
 sg13g2_fill_1 FILLER_68_1722 ();
 sg13g2_decap_4 FILLER_68_1733 ();
 sg13g2_fill_2 FILLER_68_1737 ();
 sg13g2_fill_1 FILLER_69_190 ();
 sg13g2_fill_1 FILLER_69_196 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_1 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_285 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_1 FILLER_69_305 ();
 sg13g2_fill_2 FILLER_69_332 ();
 sg13g2_fill_1 FILLER_69_348 ();
 sg13g2_fill_1 FILLER_69_389 ();
 sg13g2_fill_1 FILLER_69_397 ();
 sg13g2_fill_1 FILLER_69_464 ();
 sg13g2_fill_1 FILLER_69_469 ();
 sg13g2_fill_1 FILLER_69_474 ();
 sg13g2_fill_1 FILLER_69_501 ();
 sg13g2_fill_1 FILLER_69_528 ();
 sg13g2_fill_2 FILLER_69_592 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_fill_1 FILLER_69_707 ();
 sg13g2_fill_1 FILLER_69_718 ();
 sg13g2_fill_1 FILLER_69_723 ();
 sg13g2_fill_1 FILLER_69_749 ();
 sg13g2_fill_1 FILLER_69_755 ();
 sg13g2_fill_1 FILLER_69_792 ();
 sg13g2_fill_1 FILLER_69_829 ();
 sg13g2_fill_1 FILLER_69_894 ();
 sg13g2_decap_4 FILLER_69_940 ();
 sg13g2_fill_1 FILLER_69_944 ();
 sg13g2_decap_4 FILLER_69_949 ();
 sg13g2_fill_1 FILLER_69_953 ();
 sg13g2_decap_4 FILLER_69_957 ();
 sg13g2_fill_1 FILLER_69_961 ();
 sg13g2_fill_2 FILLER_69_966 ();
 sg13g2_fill_1 FILLER_69_968 ();
 sg13g2_decap_4 FILLER_69_989 ();
 sg13g2_fill_1 FILLER_69_993 ();
 sg13g2_fill_1 FILLER_69_1002 ();
 sg13g2_fill_1 FILLER_69_1011 ();
 sg13g2_fill_1 FILLER_69_1028 ();
 sg13g2_decap_8 FILLER_69_1040 ();
 sg13g2_fill_2 FILLER_69_1047 ();
 sg13g2_fill_1 FILLER_69_1053 ();
 sg13g2_fill_1 FILLER_69_1059 ();
 sg13g2_fill_1 FILLER_69_1068 ();
 sg13g2_fill_2 FILLER_69_1074 ();
 sg13g2_fill_2 FILLER_69_1080 ();
 sg13g2_fill_2 FILLER_69_1090 ();
 sg13g2_fill_1 FILLER_69_1096 ();
 sg13g2_fill_1 FILLER_69_1128 ();
 sg13g2_fill_2 FILLER_69_1174 ();
 sg13g2_fill_1 FILLER_69_1204 ();
 sg13g2_fill_2 FILLER_69_1209 ();
 sg13g2_fill_1 FILLER_69_1211 ();
 sg13g2_fill_1 FILLER_69_1221 ();
 sg13g2_fill_1 FILLER_69_1238 ();
 sg13g2_fill_2 FILLER_69_1243 ();
 sg13g2_fill_1 FILLER_69_1245 ();
 sg13g2_fill_1 FILLER_69_1271 ();
 sg13g2_fill_1 FILLER_69_1282 ();
 sg13g2_fill_1 FILLER_69_1295 ();
 sg13g2_fill_1 FILLER_69_1304 ();
 sg13g2_fill_2 FILLER_69_1312 ();
 sg13g2_fill_1 FILLER_69_1347 ();
 sg13g2_fill_1 FILLER_69_1356 ();
 sg13g2_fill_1 FILLER_69_1361 ();
 sg13g2_fill_2 FILLER_69_1366 ();
 sg13g2_fill_1 FILLER_69_1372 ();
 sg13g2_fill_1 FILLER_69_1381 ();
 sg13g2_fill_1 FILLER_69_1390 ();
 sg13g2_fill_1 FILLER_69_1396 ();
 sg13g2_fill_1 FILLER_69_1401 ();
 sg13g2_fill_1 FILLER_69_1410 ();
 sg13g2_fill_2 FILLER_69_1416 ();
 sg13g2_fill_2 FILLER_69_1422 ();
 sg13g2_fill_1 FILLER_69_1481 ();
 sg13g2_fill_1 FILLER_69_1500 ();
 sg13g2_fill_2 FILLER_69_1505 ();
 sg13g2_fill_2 FILLER_69_1511 ();
 sg13g2_fill_2 FILLER_69_1517 ();
 sg13g2_decap_4 FILLER_69_1523 ();
 sg13g2_fill_1 FILLER_69_1531 ();
 sg13g2_fill_2 FILLER_69_1548 ();
 sg13g2_fill_1 FILLER_69_1563 ();
 sg13g2_fill_1 FILLER_69_1569 ();
 sg13g2_fill_1 FILLER_69_1578 ();
 sg13g2_fill_2 FILLER_69_1583 ();
 sg13g2_decap_8 FILLER_69_1589 ();
 sg13g2_fill_1 FILLER_69_1596 ();
 sg13g2_fill_2 FILLER_69_1601 ();
 sg13g2_fill_1 FILLER_69_1603 ();
 sg13g2_decap_4 FILLER_69_1609 ();
 sg13g2_fill_2 FILLER_69_1613 ();
 sg13g2_fill_2 FILLER_69_1624 ();
 sg13g2_fill_1 FILLER_69_1634 ();
 sg13g2_fill_2 FILLER_69_1639 ();
 sg13g2_fill_1 FILLER_69_1649 ();
 sg13g2_fill_2 FILLER_69_1654 ();
 sg13g2_fill_2 FILLER_69_1676 ();
 sg13g2_fill_1 FILLER_69_1678 ();
 sg13g2_decap_4 FILLER_69_1683 ();
 sg13g2_fill_1 FILLER_69_1687 ();
 sg13g2_fill_1 FILLER_69_1703 ();
 sg13g2_fill_1 FILLER_69_1712 ();
 sg13g2_fill_2 FILLER_69_1717 ();
 sg13g2_fill_2 FILLER_69_1726 ();
 sg13g2_fill_2 FILLER_69_1736 ();
 sg13g2_fill_1 FILLER_69_1738 ();
 sg13g2_decap_8 FILLER_69_1767 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_29 ();
 sg13g2_fill_1 FILLER_70_40 ();
 sg13g2_fill_2 FILLER_70_67 ();
 sg13g2_fill_2 FILLER_70_93 ();
 sg13g2_fill_2 FILLER_70_149 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_1 FILLER_70_289 ();
 sg13g2_fill_2 FILLER_70_331 ();
 sg13g2_fill_2 FILLER_70_359 ();
 sg13g2_fill_2 FILLER_70_453 ();
 sg13g2_fill_1 FILLER_70_485 ();
 sg13g2_fill_2 FILLER_70_496 ();
 sg13g2_fill_2 FILLER_70_502 ();
 sg13g2_fill_2 FILLER_70_541 ();
 sg13g2_fill_1 FILLER_70_573 ();
 sg13g2_fill_1 FILLER_70_646 ();
 sg13g2_fill_1 FILLER_70_668 ();
 sg13g2_fill_1 FILLER_70_712 ();
 sg13g2_fill_1 FILLER_70_772 ();
 sg13g2_fill_1 FILLER_70_806 ();
 sg13g2_fill_1 FILLER_70_819 ();
 sg13g2_fill_2 FILLER_70_823 ();
 sg13g2_fill_1 FILLER_70_833 ();
 sg13g2_fill_2 FILLER_70_883 ();
 sg13g2_decap_8 FILLER_70_939 ();
 sg13g2_fill_2 FILLER_70_946 ();
 sg13g2_fill_1 FILLER_70_948 ();
 sg13g2_fill_1 FILLER_70_1014 ();
 sg13g2_decap_8 FILLER_70_1059 ();
 sg13g2_fill_1 FILLER_70_1079 ();
 sg13g2_fill_1 FILLER_70_1088 ();
 sg13g2_fill_1 FILLER_70_1098 ();
 sg13g2_fill_1 FILLER_70_1107 ();
 sg13g2_fill_1 FILLER_70_1120 ();
 sg13g2_decap_8 FILLER_70_1126 ();
 sg13g2_fill_1 FILLER_70_1145 ();
 sg13g2_fill_1 FILLER_70_1155 ();
 sg13g2_fill_1 FILLER_70_1161 ();
 sg13g2_fill_1 FILLER_70_1166 ();
 sg13g2_fill_1 FILLER_70_1171 ();
 sg13g2_fill_1 FILLER_70_1178 ();
 sg13g2_fill_1 FILLER_70_1187 ();
 sg13g2_fill_1 FILLER_70_1198 ();
 sg13g2_fill_2 FILLER_70_1225 ();
 sg13g2_fill_1 FILLER_70_1237 ();
 sg13g2_decap_4 FILLER_70_1251 ();
 sg13g2_fill_2 FILLER_70_1255 ();
 sg13g2_fill_1 FILLER_70_1261 ();
 sg13g2_fill_1 FILLER_70_1279 ();
 sg13g2_fill_1 FILLER_70_1289 ();
 sg13g2_fill_1 FILLER_70_1294 ();
 sg13g2_fill_1 FILLER_70_1316 ();
 sg13g2_fill_1 FILLER_70_1339 ();
 sg13g2_fill_1 FILLER_70_1358 ();
 sg13g2_fill_1 FILLER_70_1363 ();
 sg13g2_fill_2 FILLER_70_1373 ();
 sg13g2_fill_1 FILLER_70_1375 ();
 sg13g2_fill_2 FILLER_70_1380 ();
 sg13g2_fill_1 FILLER_70_1382 ();
 sg13g2_fill_2 FILLER_70_1391 ();
 sg13g2_fill_1 FILLER_70_1393 ();
 sg13g2_decap_4 FILLER_70_1414 ();
 sg13g2_fill_2 FILLER_70_1446 ();
 sg13g2_fill_2 FILLER_70_1513 ();
 sg13g2_fill_2 FILLER_70_1527 ();
 sg13g2_fill_1 FILLER_70_1541 ();
 sg13g2_fill_1 FILLER_70_1547 ();
 sg13g2_fill_1 FILLER_70_1560 ();
 sg13g2_fill_1 FILLER_70_1565 ();
 sg13g2_fill_1 FILLER_70_1578 ();
 sg13g2_fill_1 FILLER_70_1584 ();
 sg13g2_fill_1 FILLER_70_1589 ();
 sg13g2_fill_1 FILLER_70_1598 ();
 sg13g2_fill_2 FILLER_70_1604 ();
 sg13g2_fill_2 FILLER_70_1619 ();
 sg13g2_fill_1 FILLER_70_1643 ();
 sg13g2_decap_8 FILLER_70_1658 ();
 sg13g2_fill_1 FILLER_70_1669 ();
 sg13g2_decap_4 FILLER_70_1674 ();
 sg13g2_fill_2 FILLER_70_1678 ();
 sg13g2_fill_2 FILLER_70_1688 ();
 sg13g2_fill_1 FILLER_70_1698 ();
 sg13g2_fill_2 FILLER_70_1707 ();
 sg13g2_fill_2 FILLER_70_1713 ();
 sg13g2_fill_2 FILLER_70_1723 ();
 sg13g2_fill_2 FILLER_70_1729 ();
 sg13g2_fill_2 FILLER_70_1739 ();
 sg13g2_fill_2 FILLER_70_1747 ();
 sg13g2_fill_2 FILLER_70_1763 ();
 sg13g2_fill_1 FILLER_70_1765 ();
 sg13g2_fill_1 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_74 ();
 sg13g2_fill_2 FILLER_71_193 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_fill_2 FILLER_71_233 ();
 sg13g2_fill_1 FILLER_71_295 ();
 sg13g2_fill_2 FILLER_71_344 ();
 sg13g2_fill_2 FILLER_71_446 ();
 sg13g2_fill_1 FILLER_71_467 ();
 sg13g2_fill_2 FILLER_71_574 ();
 sg13g2_fill_2 FILLER_71_626 ();
 sg13g2_fill_2 FILLER_71_686 ();
 sg13g2_fill_1 FILLER_71_688 ();
 sg13g2_fill_1 FILLER_71_699 ();
 sg13g2_fill_2 FILLER_71_805 ();
 sg13g2_fill_1 FILLER_71_820 ();
 sg13g2_fill_2 FILLER_71_873 ();
 sg13g2_fill_1 FILLER_71_875 ();
 sg13g2_fill_1 FILLER_71_889 ();
 sg13g2_fill_1 FILLER_71_920 ();
 sg13g2_fill_1 FILLER_71_942 ();
 sg13g2_fill_2 FILLER_71_953 ();
 sg13g2_fill_2 FILLER_71_959 ();
 sg13g2_fill_1 FILLER_71_1032 ();
 sg13g2_fill_1 FILLER_71_1037 ();
 sg13g2_fill_1 FILLER_71_1047 ();
 sg13g2_fill_2 FILLER_71_1066 ();
 sg13g2_fill_2 FILLER_71_1076 ();
 sg13g2_fill_1 FILLER_71_1078 ();
 sg13g2_decap_8 FILLER_71_1095 ();
 sg13g2_decap_4 FILLER_71_1110 ();
 sg13g2_fill_2 FILLER_71_1135 ();
 sg13g2_fill_2 FILLER_71_1158 ();
 sg13g2_fill_1 FILLER_71_1160 ();
 sg13g2_fill_1 FILLER_71_1169 ();
 sg13g2_fill_1 FILLER_71_1183 ();
 sg13g2_decap_4 FILLER_71_1195 ();
 sg13g2_decap_8 FILLER_71_1216 ();
 sg13g2_fill_1 FILLER_71_1227 ();
 sg13g2_fill_1 FILLER_71_1232 ();
 sg13g2_fill_2 FILLER_71_1241 ();
 sg13g2_fill_1 FILLER_71_1248 ();
 sg13g2_fill_2 FILLER_71_1274 ();
 sg13g2_fill_1 FILLER_71_1292 ();
 sg13g2_fill_2 FILLER_71_1298 ();
 sg13g2_fill_1 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1309 ();
 sg13g2_fill_2 FILLER_71_1320 ();
 sg13g2_decap_4 FILLER_71_1335 ();
 sg13g2_fill_2 FILLER_71_1339 ();
 sg13g2_fill_2 FILLER_71_1354 ();
 sg13g2_fill_1 FILLER_71_1356 ();
 sg13g2_fill_2 FILLER_71_1369 ();
 sg13g2_fill_2 FILLER_71_1392 ();
 sg13g2_fill_1 FILLER_71_1402 ();
 sg13g2_fill_1 FILLER_71_1407 ();
 sg13g2_decap_4 FILLER_71_1421 ();
 sg13g2_decap_8 FILLER_71_1437 ();
 sg13g2_fill_1 FILLER_71_1444 ();
 sg13g2_fill_2 FILLER_71_1460 ();
 sg13g2_fill_1 FILLER_71_1480 ();
 sg13g2_fill_1 FILLER_71_1485 ();
 sg13g2_fill_1 FILLER_71_1493 ();
 sg13g2_fill_1 FILLER_71_1502 ();
 sg13g2_fill_1 FILLER_71_1511 ();
 sg13g2_fill_1 FILLER_71_1517 ();
 sg13g2_decap_8 FILLER_71_1522 ();
 sg13g2_fill_2 FILLER_71_1529 ();
 sg13g2_fill_1 FILLER_71_1531 ();
 sg13g2_fill_2 FILLER_71_1548 ();
 sg13g2_fill_1 FILLER_71_1555 ();
 sg13g2_decap_4 FILLER_71_1560 ();
 sg13g2_fill_2 FILLER_71_1576 ();
 sg13g2_decap_4 FILLER_71_1586 ();
 sg13g2_fill_1 FILLER_71_1590 ();
 sg13g2_fill_1 FILLER_71_1615 ();
 sg13g2_decap_4 FILLER_71_1621 ();
 sg13g2_fill_2 FILLER_71_1625 ();
 sg13g2_fill_1 FILLER_71_1631 ();
 sg13g2_fill_2 FILLER_71_1648 ();
 sg13g2_fill_1 FILLER_71_1672 ();
 sg13g2_fill_1 FILLER_71_1681 ();
 sg13g2_fill_2 FILLER_71_1686 ();
 sg13g2_fill_1 FILLER_71_1688 ();
 sg13g2_fill_2 FILLER_71_1727 ();
 sg13g2_fill_1 FILLER_71_1733 ();
 sg13g2_decap_8 FILLER_71_1739 ();
 sg13g2_fill_2 FILLER_71_1746 ();
 sg13g2_fill_1 FILLER_71_1748 ();
 sg13g2_fill_1 FILLER_71_1765 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_118 ();
 sg13g2_fill_1 FILLER_72_123 ();
 sg13g2_fill_1 FILLER_72_150 ();
 sg13g2_fill_2 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_223 ();
 sg13g2_fill_1 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_434 ();
 sg13g2_fill_1 FILLER_72_583 ();
 sg13g2_fill_2 FILLER_72_614 ();
 sg13g2_fill_2 FILLER_72_621 ();
 sg13g2_fill_2 FILLER_72_631 ();
 sg13g2_fill_1 FILLER_72_690 ();
 sg13g2_fill_1 FILLER_72_695 ();
 sg13g2_fill_1 FILLER_72_722 ();
 sg13g2_fill_2 FILLER_72_727 ();
 sg13g2_fill_1 FILLER_72_765 ();
 sg13g2_fill_1 FILLER_72_776 ();
 sg13g2_fill_1 FILLER_72_813 ();
 sg13g2_fill_1 FILLER_72_837 ();
 sg13g2_fill_2 FILLER_72_898 ();
 sg13g2_decap_8 FILLER_72_929 ();
 sg13g2_decap_8 FILLER_72_936 ();
 sg13g2_fill_1 FILLER_72_943 ();
 sg13g2_fill_1 FILLER_72_984 ();
 sg13g2_decap_4 FILLER_72_1046 ();
 sg13g2_fill_2 FILLER_72_1050 ();
 sg13g2_fill_2 FILLER_72_1057 ();
 sg13g2_decap_4 FILLER_72_1079 ();
 sg13g2_fill_2 FILLER_72_1083 ();
 sg13g2_fill_1 FILLER_72_1143 ();
 sg13g2_decap_8 FILLER_72_1154 ();
 sg13g2_fill_1 FILLER_72_1177 ();
 sg13g2_fill_1 FILLER_72_1183 ();
 sg13g2_fill_1 FILLER_72_1189 ();
 sg13g2_fill_1 FILLER_72_1194 ();
 sg13g2_fill_2 FILLER_72_1211 ();
 sg13g2_fill_2 FILLER_72_1217 ();
 sg13g2_fill_2 FILLER_72_1235 ();
 sg13g2_fill_2 FILLER_72_1245 ();
 sg13g2_decap_8 FILLER_72_1252 ();
 sg13g2_fill_1 FILLER_72_1267 ();
 sg13g2_fill_1 FILLER_72_1273 ();
 sg13g2_fill_1 FILLER_72_1278 ();
 sg13g2_fill_1 FILLER_72_1284 ();
 sg13g2_fill_1 FILLER_72_1290 ();
 sg13g2_fill_1 FILLER_72_1344 ();
 sg13g2_fill_1 FILLER_72_1350 ();
 sg13g2_fill_1 FILLER_72_1363 ();
 sg13g2_fill_1 FILLER_72_1380 ();
 sg13g2_fill_1 FILLER_72_1389 ();
 sg13g2_fill_1 FILLER_72_1411 ();
 sg13g2_fill_2 FILLER_72_1420 ();
 sg13g2_fill_2 FILLER_72_1447 ();
 sg13g2_fill_1 FILLER_72_1461 ();
 sg13g2_fill_1 FILLER_72_1483 ();
 sg13g2_fill_1 FILLER_72_1489 ();
 sg13g2_fill_2 FILLER_72_1505 ();
 sg13g2_fill_1 FILLER_72_1507 ();
 sg13g2_fill_1 FILLER_72_1520 ();
 sg13g2_fill_2 FILLER_72_1547 ();
 sg13g2_fill_1 FILLER_72_1575 ();
 sg13g2_fill_1 FILLER_72_1584 ();
 sg13g2_fill_1 FILLER_72_1596 ();
 sg13g2_decap_4 FILLER_72_1613 ();
 sg13g2_fill_1 FILLER_72_1621 ();
 sg13g2_fill_1 FILLER_72_1634 ();
 sg13g2_fill_2 FILLER_72_1658 ();
 sg13g2_fill_1 FILLER_72_1669 ();
 sg13g2_fill_2 FILLER_72_1687 ();
 sg13g2_fill_2 FILLER_72_1701 ();
 sg13g2_fill_2 FILLER_72_1707 ();
 sg13g2_decap_8 FILLER_72_1713 ();
 sg13g2_fill_2 FILLER_72_1720 ();
 sg13g2_decap_8 FILLER_72_1766 ();
 sg13g2_fill_1 FILLER_72_1773 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_34 ();
 sg13g2_fill_2 FILLER_73_92 ();
 sg13g2_fill_1 FILLER_73_151 ();
 sg13g2_fill_1 FILLER_73_185 ();
 sg13g2_fill_1 FILLER_73_220 ();
 sg13g2_fill_2 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_2 FILLER_73_305 ();
 sg13g2_fill_1 FILLER_73_363 ();
 sg13g2_fill_1 FILLER_73_390 ();
 sg13g2_fill_1 FILLER_73_424 ();
 sg13g2_fill_1 FILLER_73_465 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_fill_2 FILLER_73_620 ();
 sg13g2_fill_2 FILLER_73_626 ();
 sg13g2_fill_1 FILLER_73_703 ();
 sg13g2_fill_1 FILLER_73_712 ();
 sg13g2_fill_2 FILLER_73_751 ();
 sg13g2_fill_2 FILLER_73_773 ();
 sg13g2_fill_2 FILLER_73_814 ();
 sg13g2_fill_2 FILLER_73_845 ();
 sg13g2_fill_2 FILLER_73_930 ();
 sg13g2_decap_4 FILLER_73_936 ();
 sg13g2_fill_2 FILLER_73_940 ();
 sg13g2_fill_1 FILLER_73_952 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_fill_2 FILLER_73_998 ();
 sg13g2_decap_8 FILLER_73_1036 ();
 sg13g2_decap_8 FILLER_73_1043 ();
 sg13g2_decap_4 FILLER_73_1050 ();
 sg13g2_fill_2 FILLER_73_1054 ();
 sg13g2_fill_1 FILLER_73_1060 ();
 sg13g2_fill_2 FILLER_73_1081 ();
 sg13g2_fill_2 FILLER_73_1088 ();
 sg13g2_decap_4 FILLER_73_1117 ();
 sg13g2_decap_4 FILLER_73_1137 ();
 sg13g2_decap_4 FILLER_73_1174 ();
 sg13g2_fill_2 FILLER_73_1190 ();
 sg13g2_fill_2 FILLER_73_1208 ();
 sg13g2_fill_2 FILLER_73_1218 ();
 sg13g2_fill_1 FILLER_73_1220 ();
 sg13g2_fill_1 FILLER_73_1229 ();
 sg13g2_fill_1 FILLER_73_1234 ();
 sg13g2_fill_2 FILLER_73_1249 ();
 sg13g2_fill_1 FILLER_73_1251 ();
 sg13g2_fill_2 FILLER_73_1260 ();
 sg13g2_fill_1 FILLER_73_1262 ();
 sg13g2_fill_2 FILLER_73_1279 ();
 sg13g2_fill_1 FILLER_73_1281 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_fill_2 FILLER_73_1333 ();
 sg13g2_decap_8 FILLER_73_1368 ();
 sg13g2_fill_2 FILLER_73_1375 ();
 sg13g2_fill_1 FILLER_73_1377 ();
 sg13g2_fill_2 FILLER_73_1382 ();
 sg13g2_decap_4 FILLER_73_1392 ();
 sg13g2_decap_4 FILLER_73_1404 ();
 sg13g2_fill_1 FILLER_73_1408 ();
 sg13g2_decap_8 FILLER_73_1424 ();
 sg13g2_decap_4 FILLER_73_1431 ();
 sg13g2_fill_1 FILLER_73_1460 ();
 sg13g2_fill_1 FILLER_73_1510 ();
 sg13g2_fill_1 FILLER_73_1544 ();
 sg13g2_fill_2 FILLER_73_1549 ();
 sg13g2_decap_8 FILLER_73_1555 ();
 sg13g2_decap_8 FILLER_73_1562 ();
 sg13g2_decap_4 FILLER_73_1581 ();
 sg13g2_decap_4 FILLER_73_1628 ();
 sg13g2_fill_1 FILLER_73_1632 ();
 sg13g2_fill_1 FILLER_73_1650 ();
 sg13g2_fill_2 FILLER_73_1659 ();
 sg13g2_fill_1 FILLER_73_1670 ();
 sg13g2_fill_2 FILLER_73_1675 ();
 sg13g2_fill_1 FILLER_73_1681 ();
 sg13g2_fill_2 FILLER_73_1687 ();
 sg13g2_fill_1 FILLER_73_1694 ();
 sg13g2_fill_1 FILLER_73_1703 ();
 sg13g2_fill_1 FILLER_73_1708 ();
 sg13g2_fill_1 FILLER_73_1714 ();
 sg13g2_fill_1 FILLER_73_1724 ();
 sg13g2_fill_1 FILLER_73_1739 ();
 sg13g2_fill_2 FILLER_73_1745 ();
 sg13g2_fill_1 FILLER_73_1747 ();
 sg13g2_decap_8 FILLER_73_1767 ();
 sg13g2_fill_1 FILLER_74_50 ();
 sg13g2_fill_2 FILLER_74_144 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_fill_2 FILLER_74_307 ();
 sg13g2_fill_1 FILLER_74_326 ();
 sg13g2_fill_2 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_393 ();
 sg13g2_fill_2 FILLER_74_448 ();
 sg13g2_fill_1 FILLER_74_465 ();
 sg13g2_fill_2 FILLER_74_477 ();
 sg13g2_fill_1 FILLER_74_483 ();
 sg13g2_fill_2 FILLER_74_491 ();
 sg13g2_fill_2 FILLER_74_534 ();
 sg13g2_fill_1 FILLER_74_581 ();
 sg13g2_fill_1 FILLER_74_590 ();
 sg13g2_fill_1 FILLER_74_617 ();
 sg13g2_fill_1 FILLER_74_639 ();
 sg13g2_fill_1 FILLER_74_666 ();
 sg13g2_fill_1 FILLER_74_677 ();
 sg13g2_fill_1 FILLER_74_734 ();
 sg13g2_fill_1 FILLER_74_812 ();
 sg13g2_fill_1 FILLER_74_823 ();
 sg13g2_fill_1 FILLER_74_828 ();
 sg13g2_fill_2 FILLER_74_855 ();
 sg13g2_fill_2 FILLER_74_865 ();
 sg13g2_fill_2 FILLER_74_871 ();
 sg13g2_fill_2 FILLER_74_912 ();
 sg13g2_fill_1 FILLER_74_965 ();
 sg13g2_fill_2 FILLER_74_1020 ();
 sg13g2_fill_2 FILLER_74_1047 ();
 sg13g2_fill_2 FILLER_74_1053 ();
 sg13g2_fill_1 FILLER_74_1055 ();
 sg13g2_decap_8 FILLER_74_1059 ();
 sg13g2_decap_4 FILLER_74_1066 ();
 sg13g2_decap_8 FILLER_74_1096 ();
 sg13g2_decap_8 FILLER_74_1103 ();
 sg13g2_fill_2 FILLER_74_1110 ();
 sg13g2_fill_1 FILLER_74_1112 ();
 sg13g2_decap_4 FILLER_74_1133 ();
 sg13g2_fill_2 FILLER_74_1163 ();
 sg13g2_fill_2 FILLER_74_1213 ();
 sg13g2_decap_8 FILLER_74_1227 ();
 sg13g2_decap_8 FILLER_74_1234 ();
 sg13g2_decap_8 FILLER_74_1241 ();
 sg13g2_fill_1 FILLER_74_1248 ();
 sg13g2_fill_1 FILLER_74_1257 ();
 sg13g2_fill_1 FILLER_74_1263 ();
 sg13g2_fill_1 FILLER_74_1272 ();
 sg13g2_fill_1 FILLER_74_1277 ();
 sg13g2_fill_1 FILLER_74_1283 ();
 sg13g2_fill_1 FILLER_74_1296 ();
 sg13g2_decap_4 FILLER_74_1337 ();
 sg13g2_fill_1 FILLER_74_1341 ();
 sg13g2_fill_2 FILLER_74_1357 ();
 sg13g2_fill_1 FILLER_74_1371 ();
 sg13g2_fill_1 FILLER_74_1380 ();
 sg13g2_fill_1 FILLER_74_1389 ();
 sg13g2_fill_1 FILLER_74_1394 ();
 sg13g2_fill_2 FILLER_74_1403 ();
 sg13g2_fill_2 FILLER_74_1409 ();
 sg13g2_fill_2 FILLER_74_1424 ();
 sg13g2_fill_1 FILLER_74_1426 ();
 sg13g2_fill_2 FILLER_74_1431 ();
 sg13g2_fill_2 FILLER_74_1491 ();
 sg13g2_fill_1 FILLER_74_1493 ();
 sg13g2_fill_1 FILLER_74_1499 ();
 sg13g2_fill_1 FILLER_74_1504 ();
 sg13g2_fill_1 FILLER_74_1509 ();
 sg13g2_fill_1 FILLER_74_1532 ();
 sg13g2_fill_2 FILLER_74_1553 ();
 sg13g2_fill_1 FILLER_74_1555 ();
 sg13g2_fill_2 FILLER_74_1593 ();
 sg13g2_fill_2 FILLER_74_1613 ();
 sg13g2_fill_2 FILLER_74_1624 ();
 sg13g2_fill_1 FILLER_74_1626 ();
 sg13g2_fill_1 FILLER_74_1646 ();
 sg13g2_fill_1 FILLER_74_1651 ();
 sg13g2_decap_4 FILLER_74_1665 ();
 sg13g2_fill_1 FILLER_74_1669 ();
 sg13g2_fill_1 FILLER_74_1682 ();
 sg13g2_decap_4 FILLER_74_1688 ();
 sg13g2_fill_1 FILLER_74_1692 ();
 sg13g2_decap_8 FILLER_74_1728 ();
 sg13g2_fill_2 FILLER_74_1735 ();
 sg13g2_fill_2 FILLER_74_1750 ();
 sg13g2_fill_1 FILLER_74_1765 ();
 sg13g2_fill_2 FILLER_74_1771 ();
 sg13g2_fill_1 FILLER_74_1773 ();
 sg13g2_fill_1 FILLER_75_80 ();
 sg13g2_fill_1 FILLER_75_119 ();
 sg13g2_fill_1 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_2 FILLER_75_190 ();
 sg13g2_fill_2 FILLER_75_249 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_370 ();
 sg13g2_fill_2 FILLER_75_375 ();
 sg13g2_fill_2 FILLER_75_381 ();
 sg13g2_fill_2 FILLER_75_393 ();
 sg13g2_fill_2 FILLER_75_409 ();
 sg13g2_fill_1 FILLER_75_451 ();
 sg13g2_fill_1 FILLER_75_502 ();
 sg13g2_fill_1 FILLER_75_508 ();
 sg13g2_fill_1 FILLER_75_514 ();
 sg13g2_fill_1 FILLER_75_519 ();
 sg13g2_fill_1 FILLER_75_524 ();
 sg13g2_fill_1 FILLER_75_587 ();
 sg13g2_fill_1 FILLER_75_598 ();
 sg13g2_fill_1 FILLER_75_625 ();
 sg13g2_fill_1 FILLER_75_658 ();
 sg13g2_fill_1 FILLER_75_664 ();
 sg13g2_fill_1 FILLER_75_671 ();
 sg13g2_fill_2 FILLER_75_682 ();
 sg13g2_fill_1 FILLER_75_694 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_767 ();
 sg13g2_fill_1 FILLER_75_832 ();
 sg13g2_fill_1 FILLER_75_837 ();
 sg13g2_fill_2 FILLER_75_848 ();
 sg13g2_fill_1 FILLER_75_889 ();
 sg13g2_fill_1 FILLER_75_894 ();
 sg13g2_fill_1 FILLER_75_899 ();
 sg13g2_fill_1 FILLER_75_921 ();
 sg13g2_fill_1 FILLER_75_927 ();
 sg13g2_fill_2 FILLER_75_941 ();
 sg13g2_fill_1 FILLER_75_993 ();
 sg13g2_fill_2 FILLER_75_1030 ();
 sg13g2_decap_4 FILLER_75_1076 ();
 sg13g2_fill_1 FILLER_75_1080 ();
 sg13g2_fill_1 FILLER_75_1098 ();
 sg13g2_decap_8 FILLER_75_1107 ();
 sg13g2_decap_4 FILLER_75_1126 ();
 sg13g2_fill_1 FILLER_75_1138 ();
 sg13g2_fill_1 FILLER_75_1152 ();
 sg13g2_fill_1 FILLER_75_1158 ();
 sg13g2_fill_1 FILLER_75_1163 ();
 sg13g2_fill_2 FILLER_75_1172 ();
 sg13g2_fill_1 FILLER_75_1179 ();
 sg13g2_fill_2 FILLER_75_1184 ();
 sg13g2_fill_1 FILLER_75_1194 ();
 sg13g2_fill_1 FILLER_75_1199 ();
 sg13g2_fill_1 FILLER_75_1208 ();
 sg13g2_fill_2 FILLER_75_1213 ();
 sg13g2_decap_4 FILLER_75_1219 ();
 sg13g2_fill_2 FILLER_75_1265 ();
 sg13g2_decap_8 FILLER_75_1284 ();
 sg13g2_fill_2 FILLER_75_1291 ();
 sg13g2_fill_1 FILLER_75_1349 ();
 sg13g2_fill_2 FILLER_75_1355 ();
 sg13g2_fill_1 FILLER_75_1370 ();
 sg13g2_fill_1 FILLER_75_1379 ();
 sg13g2_fill_1 FILLER_75_1384 ();
 sg13g2_fill_1 FILLER_75_1390 ();
 sg13g2_fill_1 FILLER_75_1401 ();
 sg13g2_fill_2 FILLER_75_1406 ();
 sg13g2_fill_1 FILLER_75_1412 ();
 sg13g2_fill_2 FILLER_75_1421 ();
 sg13g2_fill_2 FILLER_75_1427 ();
 sg13g2_fill_1 FILLER_75_1429 ();
 sg13g2_fill_2 FILLER_75_1434 ();
 sg13g2_fill_1 FILLER_75_1436 ();
 sg13g2_decap_8 FILLER_75_1441 ();
 sg13g2_fill_1 FILLER_75_1448 ();
 sg13g2_fill_1 FILLER_75_1474 ();
 sg13g2_fill_1 FILLER_75_1500 ();
 sg13g2_fill_1 FILLER_75_1518 ();
 sg13g2_decap_4 FILLER_75_1523 ();
 sg13g2_fill_1 FILLER_75_1527 ();
 sg13g2_fill_2 FILLER_75_1533 ();
 sg13g2_fill_1 FILLER_75_1535 ();
 sg13g2_fill_1 FILLER_75_1550 ();
 sg13g2_decap_4 FILLER_75_1563 ();
 sg13g2_fill_1 FILLER_75_1572 ();
 sg13g2_fill_1 FILLER_75_1577 ();
 sg13g2_fill_1 FILLER_75_1582 ();
 sg13g2_fill_2 FILLER_75_1601 ();
 sg13g2_fill_1 FILLER_75_1603 ();
 sg13g2_decap_4 FILLER_75_1623 ();
 sg13g2_fill_1 FILLER_75_1627 ();
 sg13g2_fill_1 FILLER_75_1648 ();
 sg13g2_fill_1 FILLER_75_1653 ();
 sg13g2_fill_1 FILLER_75_1659 ();
 sg13g2_fill_2 FILLER_75_1665 ();
 sg13g2_fill_1 FILLER_75_1671 ();
 sg13g2_fill_1 FILLER_75_1713 ();
 sg13g2_fill_2 FILLER_75_1718 ();
 sg13g2_fill_2 FILLER_75_1724 ();
 sg13g2_fill_1 FILLER_75_1726 ();
 sg13g2_fill_1 FILLER_75_1748 ();
 sg13g2_fill_2 FILLER_75_1761 ();
 sg13g2_decap_8 FILLER_75_1767 ();
 sg13g2_fill_2 FILLER_76_65 ();
 sg13g2_fill_1 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_190 ();
 sg13g2_fill_1 FILLER_76_202 ();
 sg13g2_fill_1 FILLER_76_277 ();
 sg13g2_fill_1 FILLER_76_389 ();
 sg13g2_fill_1 FILLER_76_400 ();
 sg13g2_fill_1 FILLER_76_437 ();
 sg13g2_fill_2 FILLER_76_477 ();
 sg13g2_fill_1 FILLER_76_544 ();
 sg13g2_fill_2 FILLER_76_579 ();
 sg13g2_fill_2 FILLER_76_670 ();
 sg13g2_fill_1 FILLER_76_680 ();
 sg13g2_fill_2 FILLER_76_719 ();
 sg13g2_fill_2 FILLER_76_757 ();
 sg13g2_fill_1 FILLER_76_799 ();
 sg13g2_fill_1 FILLER_76_808 ();
 sg13g2_fill_1 FILLER_76_814 ();
 sg13g2_fill_1 FILLER_76_841 ();
 sg13g2_fill_1 FILLER_76_852 ();
 sg13g2_fill_2 FILLER_76_953 ();
 sg13g2_fill_2 FILLER_76_981 ();
 sg13g2_fill_1 FILLER_76_1009 ();
 sg13g2_fill_1 FILLER_76_1058 ();
 sg13g2_fill_1 FILLER_76_1069 ();
 sg13g2_decap_4 FILLER_76_1084 ();
 sg13g2_fill_2 FILLER_76_1088 ();
 sg13g2_decap_4 FILLER_76_1107 ();
 sg13g2_decap_8 FILLER_76_1129 ();
 sg13g2_decap_4 FILLER_76_1136 ();
 sg13g2_fill_1 FILLER_76_1176 ();
 sg13g2_fill_2 FILLER_76_1205 ();
 sg13g2_fill_1 FILLER_76_1232 ();
 sg13g2_decap_4 FILLER_76_1245 ();
 sg13g2_fill_1 FILLER_76_1249 ();
 sg13g2_decap_4 FILLER_76_1285 ();
 sg13g2_fill_2 FILLER_76_1289 ();
 sg13g2_fill_1 FILLER_76_1299 ();
 sg13g2_decap_4 FILLER_76_1317 ();
 sg13g2_fill_2 FILLER_76_1346 ();
 sg13g2_fill_2 FILLER_76_1361 ();
 sg13g2_fill_1 FILLER_76_1363 ();
 sg13g2_fill_2 FILLER_76_1372 ();
 sg13g2_decap_8 FILLER_76_1386 ();
 sg13g2_decap_4 FILLER_76_1393 ();
 sg13g2_fill_2 FILLER_76_1397 ();
 sg13g2_fill_1 FILLER_76_1411 ();
 sg13g2_fill_2 FILLER_76_1417 ();
 sg13g2_fill_1 FILLER_76_1423 ();
 sg13g2_fill_1 FILLER_76_1437 ();
 sg13g2_fill_1 FILLER_76_1442 ();
 sg13g2_fill_1 FILLER_76_1447 ();
 sg13g2_fill_2 FILLER_76_1453 ();
 sg13g2_fill_1 FILLER_76_1473 ();
 sg13g2_fill_2 FILLER_76_1493 ();
 sg13g2_fill_1 FILLER_76_1495 ();
 sg13g2_fill_2 FILLER_76_1545 ();
 sg13g2_decap_4 FILLER_76_1559 ();
 sg13g2_fill_2 FILLER_76_1563 ();
 sg13g2_decap_8 FILLER_76_1586 ();
 sg13g2_fill_1 FILLER_76_1593 ();
 sg13g2_fill_2 FILLER_76_1603 ();
 sg13g2_fill_1 FILLER_76_1613 ();
 sg13g2_fill_1 FILLER_76_1623 ();
 sg13g2_fill_1 FILLER_76_1642 ();
 sg13g2_fill_1 FILLER_76_1651 ();
 sg13g2_fill_2 FILLER_76_1660 ();
 sg13g2_decap_8 FILLER_76_1670 ();
 sg13g2_decap_8 FILLER_76_1689 ();
 sg13g2_fill_2 FILLER_76_1704 ();
 sg13g2_fill_1 FILLER_76_1733 ();
 sg13g2_fill_1 FILLER_76_1738 ();
 sg13g2_fill_2 FILLER_76_1743 ();
 sg13g2_fill_2 FILLER_76_1753 ();
 sg13g2_fill_2 FILLER_76_1764 ();
 sg13g2_decap_4 FILLER_76_1770 ();
 sg13g2_fill_1 FILLER_77_22 ();
 sg13g2_fill_1 FILLER_77_98 ();
 sg13g2_fill_1 FILLER_77_149 ();
 sg13g2_fill_2 FILLER_77_167 ();
 sg13g2_fill_1 FILLER_77_320 ();
 sg13g2_fill_2 FILLER_77_370 ();
 sg13g2_fill_2 FILLER_77_398 ();
 sg13g2_fill_1 FILLER_77_436 ();
 sg13g2_fill_2 FILLER_77_445 ();
 sg13g2_fill_2 FILLER_77_480 ();
 sg13g2_fill_1 FILLER_77_529 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_fill_1 FILLER_77_593 ();
 sg13g2_fill_1 FILLER_77_655 ();
 sg13g2_fill_2 FILLER_77_661 ();
 sg13g2_fill_1 FILLER_77_667 ();
 sg13g2_fill_2 FILLER_77_672 ();
 sg13g2_fill_1 FILLER_77_769 ();
 sg13g2_fill_1 FILLER_77_796 ();
 sg13g2_fill_2 FILLER_77_811 ();
 sg13g2_fill_2 FILLER_77_823 ();
 sg13g2_fill_1 FILLER_77_846 ();
 sg13g2_fill_2 FILLER_77_855 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_1 FILLER_77_956 ();
 sg13g2_fill_1 FILLER_77_967 ();
 sg13g2_fill_1 FILLER_77_1052 ();
 sg13g2_decap_8 FILLER_77_1089 ();
 sg13g2_fill_2 FILLER_77_1103 ();
 sg13g2_decap_8 FILLER_77_1117 ();
 sg13g2_decap_8 FILLER_77_1124 ();
 sg13g2_decap_4 FILLER_77_1131 ();
 sg13g2_decap_8 FILLER_77_1155 ();
 sg13g2_decap_8 FILLER_77_1162 ();
 sg13g2_fill_2 FILLER_77_1169 ();
 sg13g2_fill_1 FILLER_77_1171 ();
 sg13g2_decap_4 FILLER_77_1185 ();
 sg13g2_decap_8 FILLER_77_1194 ();
 sg13g2_decap_4 FILLER_77_1201 ();
 sg13g2_fill_2 FILLER_77_1218 ();
 sg13g2_fill_1 FILLER_77_1220 ();
 sg13g2_decap_4 FILLER_77_1243 ();
 sg13g2_fill_2 FILLER_77_1247 ();
 sg13g2_fill_2 FILLER_77_1265 ();
 sg13g2_fill_1 FILLER_77_1267 ();
 sg13g2_decap_4 FILLER_77_1284 ();
 sg13g2_fill_1 FILLER_77_1296 ();
 sg13g2_fill_2 FILLER_77_1314 ();
 sg13g2_fill_1 FILLER_77_1316 ();
 sg13g2_fill_2 FILLER_77_1364 ();
 sg13g2_decap_4 FILLER_77_1390 ();
 sg13g2_fill_1 FILLER_77_1394 ();
 sg13g2_fill_1 FILLER_77_1412 ();
 sg13g2_decap_4 FILLER_77_1416 ();
 sg13g2_fill_2 FILLER_77_1425 ();
 sg13g2_fill_2 FILLER_77_1456 ();
 sg13g2_decap_8 FILLER_77_1470 ();
 sg13g2_decap_4 FILLER_77_1477 ();
 sg13g2_fill_1 FILLER_77_1481 ();
 sg13g2_fill_2 FILLER_77_1510 ();
 sg13g2_fill_1 FILLER_77_1520 ();
 sg13g2_fill_2 FILLER_77_1525 ();
 sg13g2_fill_1 FILLER_77_1527 ();
 sg13g2_fill_2 FILLER_77_1532 ();
 sg13g2_fill_1 FILLER_77_1538 ();
 sg13g2_decap_4 FILLER_77_1559 ();
 sg13g2_fill_1 FILLER_77_1563 ();
 sg13g2_decap_4 FILLER_77_1568 ();
 sg13g2_fill_1 FILLER_77_1596 ();
 sg13g2_decap_4 FILLER_77_1602 ();
 sg13g2_fill_1 FILLER_77_1627 ();
 sg13g2_fill_2 FILLER_77_1652 ();
 sg13g2_fill_1 FILLER_77_1671 ();
 sg13g2_fill_1 FILLER_77_1676 ();
 sg13g2_fill_1 FILLER_77_1682 ();
 sg13g2_fill_1 FILLER_77_1688 ();
 sg13g2_fill_1 FILLER_77_1708 ();
 sg13g2_fill_2 FILLER_77_1718 ();
 sg13g2_fill_2 FILLER_77_1733 ();
 sg13g2_fill_1 FILLER_77_1735 ();
 sg13g2_fill_1 FILLER_77_1768 ();
 sg13g2_fill_1 FILLER_77_1773 ();
 sg13g2_fill_1 FILLER_78_0 ();
 sg13g2_fill_2 FILLER_78_74 ();
 sg13g2_fill_1 FILLER_78_183 ();
 sg13g2_fill_2 FILLER_78_224 ();
 sg13g2_fill_1 FILLER_78_294 ();
 sg13g2_fill_1 FILLER_78_387 ();
 sg13g2_fill_2 FILLER_78_405 ();
 sg13g2_fill_2 FILLER_78_486 ();
 sg13g2_fill_1 FILLER_78_522 ();
 sg13g2_fill_1 FILLER_78_562 ();
 sg13g2_fill_2 FILLER_78_607 ();
 sg13g2_fill_2 FILLER_78_623 ();
 sg13g2_fill_1 FILLER_78_711 ();
 sg13g2_fill_2 FILLER_78_748 ();
 sg13g2_fill_1 FILLER_78_754 ();
 sg13g2_fill_1 FILLER_78_804 ();
 sg13g2_fill_2 FILLER_78_817 ();
 sg13g2_fill_1 FILLER_78_845 ();
 sg13g2_fill_1 FILLER_78_850 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_fill_1 FILLER_78_955 ();
 sg13g2_fill_2 FILLER_78_960 ();
 sg13g2_fill_1 FILLER_78_1006 ();
 sg13g2_fill_1 FILLER_78_1111 ();
 sg13g2_fill_2 FILLER_78_1128 ();
 sg13g2_fill_2 FILLER_78_1147 ();
 sg13g2_fill_1 FILLER_78_1149 ();
 sg13g2_fill_2 FILLER_78_1158 ();
 sg13g2_fill_2 FILLER_78_1164 ();
 sg13g2_decap_4 FILLER_78_1190 ();
 sg13g2_fill_1 FILLER_78_1194 ();
 sg13g2_fill_1 FILLER_78_1223 ();
 sg13g2_decap_8 FILLER_78_1232 ();
 sg13g2_decap_4 FILLER_78_1239 ();
 sg13g2_fill_1 FILLER_78_1243 ();
 sg13g2_fill_2 FILLER_78_1257 ();
 sg13g2_fill_1 FILLER_78_1259 ();
 sg13g2_fill_2 FILLER_78_1264 ();
 sg13g2_fill_1 FILLER_78_1279 ();
 sg13g2_fill_1 FILLER_78_1285 ();
 sg13g2_fill_1 FILLER_78_1294 ();
 sg13g2_fill_1 FILLER_78_1303 ();
 sg13g2_fill_1 FILLER_78_1309 ();
 sg13g2_fill_1 FILLER_78_1314 ();
 sg13g2_fill_2 FILLER_78_1319 ();
 sg13g2_fill_1 FILLER_78_1325 ();
 sg13g2_fill_1 FILLER_78_1334 ();
 sg13g2_fill_1 FILLER_78_1342 ();
 sg13g2_fill_1 FILLER_78_1347 ();
 sg13g2_decap_4 FILLER_78_1369 ();
 sg13g2_fill_1 FILLER_78_1373 ();
 sg13g2_decap_8 FILLER_78_1415 ();
 sg13g2_decap_4 FILLER_78_1422 ();
 sg13g2_fill_1 FILLER_78_1426 ();
 sg13g2_fill_1 FILLER_78_1440 ();
 sg13g2_fill_1 FILLER_78_1450 ();
 sg13g2_fill_1 FILLER_78_1459 ();
 sg13g2_decap_4 FILLER_78_1485 ();
 sg13g2_fill_2 FILLER_78_1489 ();
 sg13g2_fill_2 FILLER_78_1507 ();
 sg13g2_decap_8 FILLER_78_1531 ();
 sg13g2_fill_2 FILLER_78_1538 ();
 sg13g2_fill_1 FILLER_78_1544 ();
 sg13g2_decap_4 FILLER_78_1559 ();
 sg13g2_fill_2 FILLER_78_1584 ();
 sg13g2_fill_1 FILLER_78_1594 ();
 sg13g2_fill_2 FILLER_78_1602 ();
 sg13g2_fill_2 FILLER_78_1609 ();
 sg13g2_fill_1 FILLER_78_1611 ();
 sg13g2_decap_8 FILLER_78_1628 ();
 sg13g2_fill_1 FILLER_78_1635 ();
 sg13g2_decap_8 FILLER_78_1656 ();
 sg13g2_fill_1 FILLER_78_1663 ();
 sg13g2_fill_1 FILLER_78_1686 ();
 sg13g2_fill_2 FILLER_78_1695 ();
 sg13g2_decap_4 FILLER_78_1713 ();
 sg13g2_decap_4 FILLER_78_1721 ();
 sg13g2_fill_1 FILLER_78_1725 ();
 sg13g2_decap_8 FILLER_78_1735 ();
 sg13g2_decap_4 FILLER_78_1742 ();
 sg13g2_fill_2 FILLER_78_1746 ();
 sg13g2_fill_1 FILLER_78_1756 ();
 sg13g2_decap_8 FILLER_78_1766 ();
 sg13g2_fill_1 FILLER_78_1773 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_171 ();
 sg13g2_fill_2 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_232 ();
 sg13g2_fill_1 FILLER_79_329 ();
 sg13g2_fill_1 FILLER_79_344 ();
 sg13g2_fill_1 FILLER_79_431 ();
 sg13g2_fill_2 FILLER_79_458 ();
 sg13g2_fill_1 FILLER_79_490 ();
 sg13g2_fill_1 FILLER_79_585 ();
 sg13g2_fill_1 FILLER_79_612 ();
 sg13g2_fill_1 FILLER_79_649 ();
 sg13g2_fill_1 FILLER_79_686 ();
 sg13g2_fill_2 FILLER_79_691 ();
 sg13g2_fill_2 FILLER_79_697 ();
 sg13g2_fill_2 FILLER_79_709 ();
 sg13g2_fill_1 FILLER_79_761 ();
 sg13g2_fill_1 FILLER_79_881 ();
 sg13g2_fill_1 FILLER_79_886 ();
 sg13g2_fill_1 FILLER_79_908 ();
 sg13g2_fill_2 FILLER_79_913 ();
 sg13g2_fill_2 FILLER_79_975 ();
 sg13g2_fill_1 FILLER_79_977 ();
 sg13g2_fill_2 FILLER_79_1047 ();
 sg13g2_fill_1 FILLER_79_1068 ();
 sg13g2_fill_1 FILLER_79_1108 ();
 sg13g2_fill_2 FILLER_79_1114 ();
 sg13g2_fill_1 FILLER_79_1151 ();
 sg13g2_fill_2 FILLER_79_1155 ();
 sg13g2_fill_2 FILLER_79_1174 ();
 sg13g2_decap_8 FILLER_79_1184 ();
 sg13g2_decap_8 FILLER_79_1191 ();
 sg13g2_decap_8 FILLER_79_1198 ();
 sg13g2_decap_4 FILLER_79_1205 ();
 sg13g2_fill_2 FILLER_79_1218 ();
 sg13g2_fill_1 FILLER_79_1220 ();
 sg13g2_decap_8 FILLER_79_1230 ();
 sg13g2_decap_4 FILLER_79_1237 ();
 sg13g2_fill_2 FILLER_79_1241 ();
 sg13g2_fill_1 FILLER_79_1251 ();
 sg13g2_fill_2 FILLER_79_1256 ();
 sg13g2_fill_2 FILLER_79_1263 ();
 sg13g2_fill_1 FILLER_79_1269 ();
 sg13g2_fill_1 FILLER_79_1278 ();
 sg13g2_fill_1 FILLER_79_1284 ();
 sg13g2_fill_2 FILLER_79_1293 ();
 sg13g2_fill_1 FILLER_79_1328 ();
 sg13g2_fill_1 FILLER_79_1334 ();
 sg13g2_fill_2 FILLER_79_1340 ();
 sg13g2_fill_1 FILLER_79_1342 ();
 sg13g2_fill_1 FILLER_79_1347 ();
 sg13g2_fill_2 FILLER_79_1360 ();
 sg13g2_fill_2 FILLER_79_1369 ();
 sg13g2_fill_2 FILLER_79_1404 ();
 sg13g2_fill_2 FILLER_79_1410 ();
 sg13g2_fill_1 FILLER_79_1412 ();
 sg13g2_decap_4 FILLER_79_1426 ();
 sg13g2_fill_1 FILLER_79_1430 ();
 sg13g2_fill_1 FILLER_79_1460 ();
 sg13g2_fill_1 FILLER_79_1469 ();
 sg13g2_fill_1 FILLER_79_1474 ();
 sg13g2_fill_1 FILLER_79_1479 ();
 sg13g2_fill_2 FILLER_79_1488 ();
 sg13g2_fill_1 FILLER_79_1516 ();
 sg13g2_decap_8 FILLER_79_1525 ();
 sg13g2_decap_8 FILLER_79_1532 ();
 sg13g2_fill_1 FILLER_79_1539 ();
 sg13g2_fill_1 FILLER_79_1546 ();
 sg13g2_fill_1 FILLER_79_1551 ();
 sg13g2_fill_1 FILLER_79_1556 ();
 sg13g2_decap_4 FILLER_79_1562 ();
 sg13g2_fill_1 FILLER_79_1652 ();
 sg13g2_fill_2 FILLER_79_1658 ();
 sg13g2_fill_2 FILLER_79_1668 ();
 sg13g2_decap_8 FILLER_79_1678 ();
 sg13g2_fill_2 FILLER_79_1689 ();
 sg13g2_fill_1 FILLER_79_1691 ();
 sg13g2_fill_2 FILLER_79_1696 ();
 sg13g2_fill_1 FILLER_79_1719 ();
 sg13g2_fill_2 FILLER_79_1732 ();
 sg13g2_fill_1 FILLER_79_1734 ();
 sg13g2_decap_8 FILLER_79_1740 ();
 sg13g2_decap_8 FILLER_79_1747 ();
 sg13g2_fill_2 FILLER_79_1754 ();
 sg13g2_decap_8 FILLER_79_1760 ();
 sg13g2_decap_8 FILLER_79_1767 ();
 sg13g2_fill_1 FILLER_80_35 ();
 sg13g2_fill_1 FILLER_80_130 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_fill_2 FILLER_80_270 ();
 sg13g2_fill_2 FILLER_80_294 ();
 sg13g2_fill_1 FILLER_80_326 ();
 sg13g2_fill_1 FILLER_80_358 ();
 sg13g2_fill_2 FILLER_80_368 ();
 sg13g2_fill_2 FILLER_80_391 ();
 sg13g2_fill_2 FILLER_80_468 ();
 sg13g2_fill_2 FILLER_80_510 ();
 sg13g2_fill_2 FILLER_80_516 ();
 sg13g2_fill_1 FILLER_80_525 ();
 sg13g2_fill_1 FILLER_80_530 ();
 sg13g2_fill_1 FILLER_80_557 ();
 sg13g2_fill_1 FILLER_80_575 ();
 sg13g2_fill_2 FILLER_80_676 ();
 sg13g2_fill_1 FILLER_80_736 ();
 sg13g2_fill_1 FILLER_80_795 ();
 sg13g2_fill_1 FILLER_80_806 ();
 sg13g2_fill_2 FILLER_80_817 ();
 sg13g2_fill_2 FILLER_80_906 ();
 sg13g2_fill_1 FILLER_80_918 ();
 sg13g2_fill_1 FILLER_80_923 ();
 sg13g2_decap_4 FILLER_80_954 ();
 sg13g2_fill_1 FILLER_80_958 ();
 sg13g2_fill_1 FILLER_80_998 ();
 sg13g2_fill_1 FILLER_80_1011 ();
 sg13g2_fill_1 FILLER_80_1042 ();
 sg13g2_fill_2 FILLER_80_1107 ();
 sg13g2_fill_1 FILLER_80_1114 ();
 sg13g2_fill_1 FILLER_80_1119 ();
 sg13g2_decap_4 FILLER_80_1147 ();
 sg13g2_fill_1 FILLER_80_1151 ();
 sg13g2_fill_2 FILLER_80_1157 ();
 sg13g2_fill_1 FILLER_80_1166 ();
 sg13g2_fill_2 FILLER_80_1183 ();
 sg13g2_decap_8 FILLER_80_1232 ();
 sg13g2_decap_4 FILLER_80_1239 ();
 sg13g2_fill_1 FILLER_80_1263 ();
 sg13g2_fill_2 FILLER_80_1268 ();
 sg13g2_fill_2 FILLER_80_1282 ();
 sg13g2_fill_1 FILLER_80_1284 ();
 sg13g2_decap_8 FILLER_80_1289 ();
 sg13g2_fill_2 FILLER_80_1296 ();
 sg13g2_fill_2 FILLER_80_1306 ();
 sg13g2_decap_8 FILLER_80_1312 ();
 sg13g2_fill_2 FILLER_80_1319 ();
 sg13g2_fill_1 FILLER_80_1321 ();
 sg13g2_decap_4 FILLER_80_1326 ();
 sg13g2_fill_1 FILLER_80_1330 ();
 sg13g2_decap_8 FILLER_80_1360 ();
 sg13g2_decap_4 FILLER_80_1367 ();
 sg13g2_fill_2 FILLER_80_1371 ();
 sg13g2_decap_4 FILLER_80_1377 ();
 sg13g2_decap_8 FILLER_80_1384 ();
 sg13g2_decap_4 FILLER_80_1391 ();
 sg13g2_fill_1 FILLER_80_1395 ();
 sg13g2_fill_2 FILLER_80_1408 ();
 sg13g2_fill_2 FILLER_80_1426 ();
 sg13g2_decap_4 FILLER_80_1446 ();
 sg13g2_fill_2 FILLER_80_1450 ();
 sg13g2_decap_8 FILLER_80_1460 ();
 sg13g2_decap_4 FILLER_80_1467 ();
 sg13g2_fill_1 FILLER_80_1471 ();
 sg13g2_decap_8 FILLER_80_1484 ();
 sg13g2_decap_8 FILLER_80_1491 ();
 sg13g2_decap_8 FILLER_80_1514 ();
 sg13g2_decap_8 FILLER_80_1521 ();
 sg13g2_decap_8 FILLER_80_1528 ();
 sg13g2_decap_8 FILLER_80_1535 ();
 sg13g2_fill_2 FILLER_80_1542 ();
 sg13g2_fill_1 FILLER_80_1561 ();
 sg13g2_fill_1 FILLER_80_1570 ();
 sg13g2_decap_8 FILLER_80_1595 ();
 sg13g2_decap_8 FILLER_80_1602 ();
 sg13g2_decap_8 FILLER_80_1609 ();
 sg13g2_fill_2 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1638 ();
 sg13g2_decap_8 FILLER_80_1645 ();
 sg13g2_fill_2 FILLER_80_1652 ();
 sg13g2_decap_4 FILLER_80_1662 ();
 sg13g2_fill_2 FILLER_80_1679 ();
 sg13g2_fill_1 FILLER_80_1681 ();
 sg13g2_decap_4 FILLER_80_1695 ();
 sg13g2_fill_1 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1708 ();
 sg13g2_decap_4 FILLER_80_1715 ();
 sg13g2_fill_1 FILLER_80_1719 ();
 sg13g2_fill_1 FILLER_80_1732 ();
 sg13g2_decap_8 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1749 ();
 sg13g2_decap_8 FILLER_80_1756 ();
 sg13g2_decap_8 FILLER_80_1763 ();
 sg13g2_decap_4 FILLER_80_1770 ();
endmodule
