module tt_um_jamesrosssharp_1bitam (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire COMP_OUT;
 wire PWM_OUT;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire clknet_leaf_0_clk;
 wire net390;
 wire \am_sdr0.I_out[0] ;
 wire \am_sdr0.I_out[1] ;
 wire \am_sdr0.I_out[2] ;
 wire \am_sdr0.I_out[3] ;
 wire \am_sdr0.I_out[4] ;
 wire \am_sdr0.I_out[5] ;
 wire \am_sdr0.I_out[6] ;
 wire \am_sdr0.I_out[7] ;
 wire \am_sdr0.Q_out[0] ;
 wire \am_sdr0.Q_out[1] ;
 wire \am_sdr0.Q_out[2] ;
 wire \am_sdr0.Q_out[3] ;
 wire \am_sdr0.Q_out[4] ;
 wire \am_sdr0.Q_out[5] ;
 wire \am_sdr0.Q_out[6] ;
 wire \am_sdr0.Q_out[7] ;
 wire \am_sdr0.am0.I_in[0] ;
 wire \am_sdr0.am0.I_in[1] ;
 wire \am_sdr0.am0.I_in[2] ;
 wire \am_sdr0.am0.I_in[3] ;
 wire \am_sdr0.am0.I_in[4] ;
 wire \am_sdr0.am0.I_in[5] ;
 wire \am_sdr0.am0.I_in[6] ;
 wire \am_sdr0.am0.I_in[7] ;
 wire \am_sdr0.am0.Q_in[0] ;
 wire \am_sdr0.am0.Q_in[1] ;
 wire \am_sdr0.am0.Q_in[2] ;
 wire \am_sdr0.am0.Q_in[3] ;
 wire \am_sdr0.am0.Q_in[4] ;
 wire \am_sdr0.am0.Q_in[5] ;
 wire \am_sdr0.am0.Q_in[6] ;
 wire \am_sdr0.am0.Q_in[7] ;
 wire \am_sdr0.am0.a[0] ;
 wire \am_sdr0.am0.a[10] ;
 wire \am_sdr0.am0.a[11] ;
 wire \am_sdr0.am0.a[12] ;
 wire \am_sdr0.am0.a[13] ;
 wire \am_sdr0.am0.a[14] ;
 wire \am_sdr0.am0.a[15] ;
 wire \am_sdr0.am0.a[1] ;
 wire \am_sdr0.am0.a[2] ;
 wire \am_sdr0.am0.a[3] ;
 wire \am_sdr0.am0.a[4] ;
 wire \am_sdr0.am0.a[5] ;
 wire \am_sdr0.am0.a[6] ;
 wire \am_sdr0.am0.a[7] ;
 wire \am_sdr0.am0.a[8] ;
 wire \am_sdr0.am0.a[9] ;
 wire \am_sdr0.am0.count2[0] ;
 wire \am_sdr0.am0.count2[1] ;
 wire \am_sdr0.am0.count2[2] ;
 wire \am_sdr0.am0.count2[3] ;
 wire \am_sdr0.am0.count[0] ;
 wire \am_sdr0.am0.count[1] ;
 wire \am_sdr0.am0.demod_out[10] ;
 wire \am_sdr0.am0.demod_out[11] ;
 wire \am_sdr0.am0.demod_out[12] ;
 wire \am_sdr0.am0.demod_out[13] ;
 wire \am_sdr0.am0.demod_out[14] ;
 wire \am_sdr0.am0.demod_out[15] ;
 wire \am_sdr0.am0.demod_out[8] ;
 wire \am_sdr0.am0.demod_out[9] ;
 wire \am_sdr0.am0.left[0] ;
 wire \am_sdr0.am0.left[1] ;
 wire \am_sdr0.am0.left[2] ;
 wire \am_sdr0.am0.left[3] ;
 wire \am_sdr0.am0.left[4] ;
 wire \am_sdr0.am0.left[5] ;
 wire \am_sdr0.am0.left[6] ;
 wire \am_sdr0.am0.left[7] ;
 wire \am_sdr0.am0.left[8] ;
 wire \am_sdr0.am0.left[9] ;
 wire \am_sdr0.am0.load_tick ;
 wire \am_sdr0.am0.m_count[0] ;
 wire \am_sdr0.am0.m_count[1] ;
 wire \am_sdr0.am0.m_count[2] ;
 wire \am_sdr0.am0.m_count[3] ;
 wire \am_sdr0.am0.multA[0] ;
 wire \am_sdr0.am0.multA[10] ;
 wire \am_sdr0.am0.multA[11] ;
 wire \am_sdr0.am0.multA[12] ;
 wire \am_sdr0.am0.multA[13] ;
 wire \am_sdr0.am0.multA[14] ;
 wire \am_sdr0.am0.multA[15] ;
 wire \am_sdr0.am0.multA[16] ;
 wire \am_sdr0.am0.multA[1] ;
 wire \am_sdr0.am0.multA[2] ;
 wire \am_sdr0.am0.multA[3] ;
 wire \am_sdr0.am0.multA[4] ;
 wire \am_sdr0.am0.multA[5] ;
 wire \am_sdr0.am0.multA[6] ;
 wire \am_sdr0.am0.multA[7] ;
 wire \am_sdr0.am0.multA[8] ;
 wire \am_sdr0.am0.multA[9] ;
 wire \am_sdr0.am0.multB[0] ;
 wire \am_sdr0.am0.multB[1] ;
 wire \am_sdr0.am0.multB[2] ;
 wire \am_sdr0.am0.multB[3] ;
 wire \am_sdr0.am0.multB[4] ;
 wire \am_sdr0.am0.multB[5] ;
 wire \am_sdr0.am0.multB[6] ;
 wire \am_sdr0.am0.multB[7] ;
 wire \am_sdr0.am0.q[0] ;
 wire \am_sdr0.am0.q[1] ;
 wire \am_sdr0.am0.q[2] ;
 wire \am_sdr0.am0.q[3] ;
 wire \am_sdr0.am0.q[4] ;
 wire \am_sdr0.am0.q[5] ;
 wire \am_sdr0.am0.q[6] ;
 wire \am_sdr0.am0.q[7] ;
 wire \am_sdr0.am0.r[0] ;
 wire \am_sdr0.am0.r[1] ;
 wire \am_sdr0.am0.r[2] ;
 wire \am_sdr0.am0.r[3] ;
 wire \am_sdr0.am0.r[4] ;
 wire \am_sdr0.am0.r[5] ;
 wire \am_sdr0.am0.r[6] ;
 wire \am_sdr0.am0.r[7] ;
 wire \am_sdr0.am0.r[9] ;
 wire \am_sdr0.am0.right[0] ;
 wire \am_sdr0.am0.right[1] ;
 wire \am_sdr0.am0.right[2] ;
 wire \am_sdr0.am0.right[3] ;
 wire \am_sdr0.am0.right[4] ;
 wire \am_sdr0.am0.right[5] ;
 wire \am_sdr0.am0.right[6] ;
 wire \am_sdr0.am0.right[7] ;
 wire \am_sdr0.am0.right[8] ;
 wire \am_sdr0.am0.right[9] ;
 wire \am_sdr0.am0.sqrt_done ;
 wire \am_sdr0.am0.sqrt_state[0] ;
 wire \am_sdr0.am0.sqrt_state[1] ;
 wire \am_sdr0.am0.state[0] ;
 wire \am_sdr0.am0.state[1] ;
 wire \am_sdr0.am0.state[2] ;
 wire \am_sdr0.am0.state[3] ;
 wire \am_sdr0.am0.state[4] ;
 wire \am_sdr0.am0.state[5] ;
 wire \am_sdr0.am0.state[6] ;
 wire \am_sdr0.am0.sum[0] ;
 wire \am_sdr0.am0.sum[10] ;
 wire \am_sdr0.am0.sum[11] ;
 wire \am_sdr0.am0.sum[12] ;
 wire \am_sdr0.am0.sum[13] ;
 wire \am_sdr0.am0.sum[14] ;
 wire \am_sdr0.am0.sum[15] ;
 wire \am_sdr0.am0.sum[16] ;
 wire \am_sdr0.am0.sum[1] ;
 wire \am_sdr0.am0.sum[2] ;
 wire \am_sdr0.am0.sum[3] ;
 wire \am_sdr0.am0.sum[4] ;
 wire \am_sdr0.am0.sum[5] ;
 wire \am_sdr0.am0.sum[6] ;
 wire \am_sdr0.am0.sum[7] ;
 wire \am_sdr0.am0.sum[8] ;
 wire \am_sdr0.am0.sum[9] ;
 wire \am_sdr0.cic0.comb1[0] ;
 wire \am_sdr0.cic0.comb1[10] ;
 wire \am_sdr0.cic0.comb1[11] ;
 wire \am_sdr0.cic0.comb1[12] ;
 wire \am_sdr0.cic0.comb1[13] ;
 wire \am_sdr0.cic0.comb1[14] ;
 wire \am_sdr0.cic0.comb1[15] ;
 wire \am_sdr0.cic0.comb1[16] ;
 wire \am_sdr0.cic0.comb1[17] ;
 wire \am_sdr0.cic0.comb1[18] ;
 wire \am_sdr0.cic0.comb1[19] ;
 wire \am_sdr0.cic0.comb1[1] ;
 wire \am_sdr0.cic0.comb1[2] ;
 wire \am_sdr0.cic0.comb1[3] ;
 wire \am_sdr0.cic0.comb1[4] ;
 wire \am_sdr0.cic0.comb1[5] ;
 wire \am_sdr0.cic0.comb1[6] ;
 wire \am_sdr0.cic0.comb1[7] ;
 wire \am_sdr0.cic0.comb1[8] ;
 wire \am_sdr0.cic0.comb1[9] ;
 wire \am_sdr0.cic0.comb1_in_del[0] ;
 wire \am_sdr0.cic0.comb1_in_del[10] ;
 wire \am_sdr0.cic0.comb1_in_del[11] ;
 wire \am_sdr0.cic0.comb1_in_del[12] ;
 wire \am_sdr0.cic0.comb1_in_del[13] ;
 wire \am_sdr0.cic0.comb1_in_del[14] ;
 wire \am_sdr0.cic0.comb1_in_del[15] ;
 wire \am_sdr0.cic0.comb1_in_del[16] ;
 wire \am_sdr0.cic0.comb1_in_del[17] ;
 wire \am_sdr0.cic0.comb1_in_del[18] ;
 wire \am_sdr0.cic0.comb1_in_del[19] ;
 wire \am_sdr0.cic0.comb1_in_del[1] ;
 wire \am_sdr0.cic0.comb1_in_del[2] ;
 wire \am_sdr0.cic0.comb1_in_del[3] ;
 wire \am_sdr0.cic0.comb1_in_del[4] ;
 wire \am_sdr0.cic0.comb1_in_del[5] ;
 wire \am_sdr0.cic0.comb1_in_del[6] ;
 wire \am_sdr0.cic0.comb1_in_del[7] ;
 wire \am_sdr0.cic0.comb1_in_del[8] ;
 wire \am_sdr0.cic0.comb1_in_del[9] ;
 wire \am_sdr0.cic0.comb2[0] ;
 wire \am_sdr0.cic0.comb2[10] ;
 wire \am_sdr0.cic0.comb2[11] ;
 wire \am_sdr0.cic0.comb2[12] ;
 wire \am_sdr0.cic0.comb2[13] ;
 wire \am_sdr0.cic0.comb2[14] ;
 wire \am_sdr0.cic0.comb2[15] ;
 wire \am_sdr0.cic0.comb2[16] ;
 wire \am_sdr0.cic0.comb2[17] ;
 wire \am_sdr0.cic0.comb2[18] ;
 wire \am_sdr0.cic0.comb2[19] ;
 wire \am_sdr0.cic0.comb2[1] ;
 wire \am_sdr0.cic0.comb2[2] ;
 wire \am_sdr0.cic0.comb2[3] ;
 wire \am_sdr0.cic0.comb2[4] ;
 wire \am_sdr0.cic0.comb2[5] ;
 wire \am_sdr0.cic0.comb2[6] ;
 wire \am_sdr0.cic0.comb2[7] ;
 wire \am_sdr0.cic0.comb2[8] ;
 wire \am_sdr0.cic0.comb2[9] ;
 wire \am_sdr0.cic0.comb2_in_del[0] ;
 wire \am_sdr0.cic0.comb2_in_del[10] ;
 wire \am_sdr0.cic0.comb2_in_del[11] ;
 wire \am_sdr0.cic0.comb2_in_del[12] ;
 wire \am_sdr0.cic0.comb2_in_del[13] ;
 wire \am_sdr0.cic0.comb2_in_del[14] ;
 wire \am_sdr0.cic0.comb2_in_del[15] ;
 wire \am_sdr0.cic0.comb2_in_del[16] ;
 wire \am_sdr0.cic0.comb2_in_del[17] ;
 wire \am_sdr0.cic0.comb2_in_del[18] ;
 wire \am_sdr0.cic0.comb2_in_del[19] ;
 wire \am_sdr0.cic0.comb2_in_del[1] ;
 wire \am_sdr0.cic0.comb2_in_del[2] ;
 wire \am_sdr0.cic0.comb2_in_del[3] ;
 wire \am_sdr0.cic0.comb2_in_del[4] ;
 wire \am_sdr0.cic0.comb2_in_del[5] ;
 wire \am_sdr0.cic0.comb2_in_del[6] ;
 wire \am_sdr0.cic0.comb2_in_del[7] ;
 wire \am_sdr0.cic0.comb2_in_del[8] ;
 wire \am_sdr0.cic0.comb2_in_del[9] ;
 wire \am_sdr0.cic0.comb3[12] ;
 wire \am_sdr0.cic0.comb3[13] ;
 wire \am_sdr0.cic0.comb3[14] ;
 wire \am_sdr0.cic0.comb3[15] ;
 wire \am_sdr0.cic0.comb3[16] ;
 wire \am_sdr0.cic0.comb3[17] ;
 wire \am_sdr0.cic0.comb3[18] ;
 wire \am_sdr0.cic0.comb3[19] ;
 wire \am_sdr0.cic0.comb3_in_del[0] ;
 wire \am_sdr0.cic0.comb3_in_del[10] ;
 wire \am_sdr0.cic0.comb3_in_del[11] ;
 wire \am_sdr0.cic0.comb3_in_del[12] ;
 wire \am_sdr0.cic0.comb3_in_del[13] ;
 wire \am_sdr0.cic0.comb3_in_del[14] ;
 wire \am_sdr0.cic0.comb3_in_del[15] ;
 wire \am_sdr0.cic0.comb3_in_del[16] ;
 wire \am_sdr0.cic0.comb3_in_del[17] ;
 wire \am_sdr0.cic0.comb3_in_del[18] ;
 wire \am_sdr0.cic0.comb3_in_del[19] ;
 wire \am_sdr0.cic0.comb3_in_del[1] ;
 wire \am_sdr0.cic0.comb3_in_del[2] ;
 wire \am_sdr0.cic0.comb3_in_del[3] ;
 wire \am_sdr0.cic0.comb3_in_del[4] ;
 wire \am_sdr0.cic0.comb3_in_del[5] ;
 wire \am_sdr0.cic0.comb3_in_del[6] ;
 wire \am_sdr0.cic0.comb3_in_del[7] ;
 wire \am_sdr0.cic0.comb3_in_del[8] ;
 wire \am_sdr0.cic0.comb3_in_del[9] ;
 wire \am_sdr0.cic0.count[0] ;
 wire \am_sdr0.cic0.count[1] ;
 wire \am_sdr0.cic0.count[2] ;
 wire \am_sdr0.cic0.count[3] ;
 wire \am_sdr0.cic0.count[4] ;
 wire \am_sdr0.cic0.count[5] ;
 wire \am_sdr0.cic0.count[6] ;
 wire \am_sdr0.cic0.count[7] ;
 wire \am_sdr0.cic0.integ1[0] ;
 wire \am_sdr0.cic0.integ1[10] ;
 wire \am_sdr0.cic0.integ1[11] ;
 wire \am_sdr0.cic0.integ1[12] ;
 wire \am_sdr0.cic0.integ1[13] ;
 wire \am_sdr0.cic0.integ1[14] ;
 wire \am_sdr0.cic0.integ1[15] ;
 wire \am_sdr0.cic0.integ1[16] ;
 wire \am_sdr0.cic0.integ1[17] ;
 wire \am_sdr0.cic0.integ1[18] ;
 wire \am_sdr0.cic0.integ1[19] ;
 wire \am_sdr0.cic0.integ1[1] ;
 wire \am_sdr0.cic0.integ1[20] ;
 wire \am_sdr0.cic0.integ1[21] ;
 wire \am_sdr0.cic0.integ1[22] ;
 wire \am_sdr0.cic0.integ1[23] ;
 wire \am_sdr0.cic0.integ1[24] ;
 wire \am_sdr0.cic0.integ1[25] ;
 wire \am_sdr0.cic0.integ1[2] ;
 wire \am_sdr0.cic0.integ1[3] ;
 wire \am_sdr0.cic0.integ1[4] ;
 wire \am_sdr0.cic0.integ1[5] ;
 wire \am_sdr0.cic0.integ1[6] ;
 wire \am_sdr0.cic0.integ1[7] ;
 wire \am_sdr0.cic0.integ1[8] ;
 wire \am_sdr0.cic0.integ1[9] ;
 wire \am_sdr0.cic0.integ2[0] ;
 wire \am_sdr0.cic0.integ2[10] ;
 wire \am_sdr0.cic0.integ2[11] ;
 wire \am_sdr0.cic0.integ2[12] ;
 wire \am_sdr0.cic0.integ2[13] ;
 wire \am_sdr0.cic0.integ2[14] ;
 wire \am_sdr0.cic0.integ2[15] ;
 wire \am_sdr0.cic0.integ2[16] ;
 wire \am_sdr0.cic0.integ2[17] ;
 wire \am_sdr0.cic0.integ2[18] ;
 wire \am_sdr0.cic0.integ2[19] ;
 wire \am_sdr0.cic0.integ2[1] ;
 wire \am_sdr0.cic0.integ2[20] ;
 wire \am_sdr0.cic0.integ2[21] ;
 wire \am_sdr0.cic0.integ2[22] ;
 wire \am_sdr0.cic0.integ2[2] ;
 wire \am_sdr0.cic0.integ2[3] ;
 wire \am_sdr0.cic0.integ2[4] ;
 wire \am_sdr0.cic0.integ2[5] ;
 wire \am_sdr0.cic0.integ2[6] ;
 wire \am_sdr0.cic0.integ2[7] ;
 wire \am_sdr0.cic0.integ2[8] ;
 wire \am_sdr0.cic0.integ2[9] ;
 wire \am_sdr0.cic0.integ3[0] ;
 wire \am_sdr0.cic0.integ3[10] ;
 wire \am_sdr0.cic0.integ3[11] ;
 wire \am_sdr0.cic0.integ3[12] ;
 wire \am_sdr0.cic0.integ3[13] ;
 wire \am_sdr0.cic0.integ3[14] ;
 wire \am_sdr0.cic0.integ3[15] ;
 wire \am_sdr0.cic0.integ3[16] ;
 wire \am_sdr0.cic0.integ3[17] ;
 wire \am_sdr0.cic0.integ3[18] ;
 wire \am_sdr0.cic0.integ3[19] ;
 wire \am_sdr0.cic0.integ3[1] ;
 wire \am_sdr0.cic0.integ3[2] ;
 wire \am_sdr0.cic0.integ3[3] ;
 wire \am_sdr0.cic0.integ3[4] ;
 wire \am_sdr0.cic0.integ3[5] ;
 wire \am_sdr0.cic0.integ3[6] ;
 wire \am_sdr0.cic0.integ3[7] ;
 wire \am_sdr0.cic0.integ3[8] ;
 wire \am_sdr0.cic0.integ3[9] ;
 wire \am_sdr0.cic0.integ_sample[0] ;
 wire \am_sdr0.cic0.integ_sample[10] ;
 wire \am_sdr0.cic0.integ_sample[11] ;
 wire \am_sdr0.cic0.integ_sample[12] ;
 wire \am_sdr0.cic0.integ_sample[13] ;
 wire \am_sdr0.cic0.integ_sample[14] ;
 wire \am_sdr0.cic0.integ_sample[15] ;
 wire \am_sdr0.cic0.integ_sample[16] ;
 wire \am_sdr0.cic0.integ_sample[17] ;
 wire \am_sdr0.cic0.integ_sample[18] ;
 wire \am_sdr0.cic0.integ_sample[19] ;
 wire \am_sdr0.cic0.integ_sample[1] ;
 wire \am_sdr0.cic0.integ_sample[2] ;
 wire \am_sdr0.cic0.integ_sample[3] ;
 wire \am_sdr0.cic0.integ_sample[4] ;
 wire \am_sdr0.cic0.integ_sample[5] ;
 wire \am_sdr0.cic0.integ_sample[6] ;
 wire \am_sdr0.cic0.integ_sample[7] ;
 wire \am_sdr0.cic0.integ_sample[8] ;
 wire \am_sdr0.cic0.integ_sample[9] ;
 wire \am_sdr0.cic0.out_tick ;
 wire \am_sdr0.cic0.sample ;
 wire \am_sdr0.cic0.x_out[10] ;
 wire \am_sdr0.cic0.x_out[11] ;
 wire \am_sdr0.cic0.x_out[12] ;
 wire \am_sdr0.cic0.x_out[13] ;
 wire \am_sdr0.cic0.x_out[14] ;
 wire \am_sdr0.cic0.x_out[15] ;
 wire \am_sdr0.cic0.x_out[8] ;
 wire \am_sdr0.cic0.x_out[9] ;
 wire \am_sdr0.cic1.comb1[0] ;
 wire \am_sdr0.cic1.comb1[10] ;
 wire \am_sdr0.cic1.comb1[11] ;
 wire \am_sdr0.cic1.comb1[12] ;
 wire \am_sdr0.cic1.comb1[13] ;
 wire \am_sdr0.cic1.comb1[14] ;
 wire \am_sdr0.cic1.comb1[15] ;
 wire \am_sdr0.cic1.comb1[16] ;
 wire \am_sdr0.cic1.comb1[17] ;
 wire \am_sdr0.cic1.comb1[18] ;
 wire \am_sdr0.cic1.comb1[19] ;
 wire \am_sdr0.cic1.comb1[1] ;
 wire \am_sdr0.cic1.comb1[2] ;
 wire \am_sdr0.cic1.comb1[3] ;
 wire \am_sdr0.cic1.comb1[4] ;
 wire \am_sdr0.cic1.comb1[5] ;
 wire \am_sdr0.cic1.comb1[6] ;
 wire \am_sdr0.cic1.comb1[7] ;
 wire \am_sdr0.cic1.comb1[8] ;
 wire \am_sdr0.cic1.comb1[9] ;
 wire \am_sdr0.cic1.comb1_in_del[0] ;
 wire \am_sdr0.cic1.comb1_in_del[10] ;
 wire \am_sdr0.cic1.comb1_in_del[11] ;
 wire \am_sdr0.cic1.comb1_in_del[12] ;
 wire \am_sdr0.cic1.comb1_in_del[13] ;
 wire \am_sdr0.cic1.comb1_in_del[14] ;
 wire \am_sdr0.cic1.comb1_in_del[15] ;
 wire \am_sdr0.cic1.comb1_in_del[16] ;
 wire \am_sdr0.cic1.comb1_in_del[17] ;
 wire \am_sdr0.cic1.comb1_in_del[18] ;
 wire \am_sdr0.cic1.comb1_in_del[19] ;
 wire \am_sdr0.cic1.comb1_in_del[1] ;
 wire \am_sdr0.cic1.comb1_in_del[2] ;
 wire \am_sdr0.cic1.comb1_in_del[3] ;
 wire \am_sdr0.cic1.comb1_in_del[4] ;
 wire \am_sdr0.cic1.comb1_in_del[5] ;
 wire \am_sdr0.cic1.comb1_in_del[6] ;
 wire \am_sdr0.cic1.comb1_in_del[7] ;
 wire \am_sdr0.cic1.comb1_in_del[8] ;
 wire \am_sdr0.cic1.comb1_in_del[9] ;
 wire \am_sdr0.cic1.comb2[0] ;
 wire \am_sdr0.cic1.comb2[10] ;
 wire \am_sdr0.cic1.comb2[11] ;
 wire \am_sdr0.cic1.comb2[12] ;
 wire \am_sdr0.cic1.comb2[13] ;
 wire \am_sdr0.cic1.comb2[14] ;
 wire \am_sdr0.cic1.comb2[15] ;
 wire \am_sdr0.cic1.comb2[16] ;
 wire \am_sdr0.cic1.comb2[17] ;
 wire \am_sdr0.cic1.comb2[18] ;
 wire \am_sdr0.cic1.comb2[19] ;
 wire \am_sdr0.cic1.comb2[1] ;
 wire \am_sdr0.cic1.comb2[2] ;
 wire \am_sdr0.cic1.comb2[3] ;
 wire \am_sdr0.cic1.comb2[4] ;
 wire \am_sdr0.cic1.comb2[5] ;
 wire \am_sdr0.cic1.comb2[6] ;
 wire \am_sdr0.cic1.comb2[7] ;
 wire \am_sdr0.cic1.comb2[8] ;
 wire \am_sdr0.cic1.comb2[9] ;
 wire \am_sdr0.cic1.comb2_in_del[0] ;
 wire \am_sdr0.cic1.comb2_in_del[10] ;
 wire \am_sdr0.cic1.comb2_in_del[11] ;
 wire \am_sdr0.cic1.comb2_in_del[12] ;
 wire \am_sdr0.cic1.comb2_in_del[13] ;
 wire \am_sdr0.cic1.comb2_in_del[14] ;
 wire \am_sdr0.cic1.comb2_in_del[15] ;
 wire \am_sdr0.cic1.comb2_in_del[16] ;
 wire \am_sdr0.cic1.comb2_in_del[17] ;
 wire \am_sdr0.cic1.comb2_in_del[18] ;
 wire \am_sdr0.cic1.comb2_in_del[19] ;
 wire \am_sdr0.cic1.comb2_in_del[1] ;
 wire \am_sdr0.cic1.comb2_in_del[2] ;
 wire \am_sdr0.cic1.comb2_in_del[3] ;
 wire \am_sdr0.cic1.comb2_in_del[4] ;
 wire \am_sdr0.cic1.comb2_in_del[5] ;
 wire \am_sdr0.cic1.comb2_in_del[6] ;
 wire \am_sdr0.cic1.comb2_in_del[7] ;
 wire \am_sdr0.cic1.comb2_in_del[8] ;
 wire \am_sdr0.cic1.comb2_in_del[9] ;
 wire \am_sdr0.cic1.comb3[12] ;
 wire \am_sdr0.cic1.comb3[13] ;
 wire \am_sdr0.cic1.comb3[14] ;
 wire \am_sdr0.cic1.comb3[15] ;
 wire \am_sdr0.cic1.comb3[16] ;
 wire \am_sdr0.cic1.comb3[17] ;
 wire \am_sdr0.cic1.comb3[18] ;
 wire \am_sdr0.cic1.comb3[19] ;
 wire \am_sdr0.cic1.comb3_in_del[0] ;
 wire \am_sdr0.cic1.comb3_in_del[10] ;
 wire \am_sdr0.cic1.comb3_in_del[11] ;
 wire \am_sdr0.cic1.comb3_in_del[12] ;
 wire \am_sdr0.cic1.comb3_in_del[13] ;
 wire \am_sdr0.cic1.comb3_in_del[14] ;
 wire \am_sdr0.cic1.comb3_in_del[15] ;
 wire \am_sdr0.cic1.comb3_in_del[16] ;
 wire \am_sdr0.cic1.comb3_in_del[17] ;
 wire \am_sdr0.cic1.comb3_in_del[18] ;
 wire \am_sdr0.cic1.comb3_in_del[19] ;
 wire \am_sdr0.cic1.comb3_in_del[1] ;
 wire \am_sdr0.cic1.comb3_in_del[2] ;
 wire \am_sdr0.cic1.comb3_in_del[3] ;
 wire \am_sdr0.cic1.comb3_in_del[4] ;
 wire \am_sdr0.cic1.comb3_in_del[5] ;
 wire \am_sdr0.cic1.comb3_in_del[6] ;
 wire \am_sdr0.cic1.comb3_in_del[7] ;
 wire \am_sdr0.cic1.comb3_in_del[8] ;
 wire \am_sdr0.cic1.comb3_in_del[9] ;
 wire \am_sdr0.cic1.count[0] ;
 wire \am_sdr0.cic1.count[1] ;
 wire \am_sdr0.cic1.count[2] ;
 wire \am_sdr0.cic1.count[3] ;
 wire \am_sdr0.cic1.count[4] ;
 wire \am_sdr0.cic1.count[5] ;
 wire \am_sdr0.cic1.count[6] ;
 wire \am_sdr0.cic1.count[7] ;
 wire \am_sdr0.cic1.integ1[0] ;
 wire \am_sdr0.cic1.integ1[10] ;
 wire \am_sdr0.cic1.integ1[11] ;
 wire \am_sdr0.cic1.integ1[12] ;
 wire \am_sdr0.cic1.integ1[13] ;
 wire \am_sdr0.cic1.integ1[14] ;
 wire \am_sdr0.cic1.integ1[15] ;
 wire \am_sdr0.cic1.integ1[16] ;
 wire \am_sdr0.cic1.integ1[17] ;
 wire \am_sdr0.cic1.integ1[18] ;
 wire \am_sdr0.cic1.integ1[19] ;
 wire \am_sdr0.cic1.integ1[1] ;
 wire \am_sdr0.cic1.integ1[20] ;
 wire \am_sdr0.cic1.integ1[21] ;
 wire \am_sdr0.cic1.integ1[22] ;
 wire \am_sdr0.cic1.integ1[23] ;
 wire \am_sdr0.cic1.integ1[24] ;
 wire \am_sdr0.cic1.integ1[25] ;
 wire \am_sdr0.cic1.integ1[2] ;
 wire \am_sdr0.cic1.integ1[3] ;
 wire \am_sdr0.cic1.integ1[4] ;
 wire \am_sdr0.cic1.integ1[5] ;
 wire \am_sdr0.cic1.integ1[6] ;
 wire \am_sdr0.cic1.integ1[7] ;
 wire \am_sdr0.cic1.integ1[8] ;
 wire \am_sdr0.cic1.integ1[9] ;
 wire \am_sdr0.cic1.integ2[0] ;
 wire \am_sdr0.cic1.integ2[10] ;
 wire \am_sdr0.cic1.integ2[11] ;
 wire \am_sdr0.cic1.integ2[12] ;
 wire \am_sdr0.cic1.integ2[13] ;
 wire \am_sdr0.cic1.integ2[14] ;
 wire \am_sdr0.cic1.integ2[15] ;
 wire \am_sdr0.cic1.integ2[16] ;
 wire \am_sdr0.cic1.integ2[17] ;
 wire \am_sdr0.cic1.integ2[18] ;
 wire \am_sdr0.cic1.integ2[19] ;
 wire \am_sdr0.cic1.integ2[1] ;
 wire \am_sdr0.cic1.integ2[20] ;
 wire \am_sdr0.cic1.integ2[21] ;
 wire \am_sdr0.cic1.integ2[22] ;
 wire \am_sdr0.cic1.integ2[2] ;
 wire \am_sdr0.cic1.integ2[3] ;
 wire \am_sdr0.cic1.integ2[4] ;
 wire \am_sdr0.cic1.integ2[5] ;
 wire \am_sdr0.cic1.integ2[6] ;
 wire \am_sdr0.cic1.integ2[7] ;
 wire \am_sdr0.cic1.integ2[8] ;
 wire \am_sdr0.cic1.integ2[9] ;
 wire \am_sdr0.cic1.integ3[0] ;
 wire \am_sdr0.cic1.integ3[10] ;
 wire \am_sdr0.cic1.integ3[11] ;
 wire \am_sdr0.cic1.integ3[12] ;
 wire \am_sdr0.cic1.integ3[13] ;
 wire \am_sdr0.cic1.integ3[14] ;
 wire \am_sdr0.cic1.integ3[15] ;
 wire \am_sdr0.cic1.integ3[16] ;
 wire \am_sdr0.cic1.integ3[17] ;
 wire \am_sdr0.cic1.integ3[18] ;
 wire \am_sdr0.cic1.integ3[19] ;
 wire \am_sdr0.cic1.integ3[1] ;
 wire \am_sdr0.cic1.integ3[2] ;
 wire \am_sdr0.cic1.integ3[3] ;
 wire \am_sdr0.cic1.integ3[4] ;
 wire \am_sdr0.cic1.integ3[5] ;
 wire \am_sdr0.cic1.integ3[6] ;
 wire \am_sdr0.cic1.integ3[7] ;
 wire \am_sdr0.cic1.integ3[8] ;
 wire \am_sdr0.cic1.integ3[9] ;
 wire \am_sdr0.cic1.integ_sample[0] ;
 wire \am_sdr0.cic1.integ_sample[10] ;
 wire \am_sdr0.cic1.integ_sample[11] ;
 wire \am_sdr0.cic1.integ_sample[12] ;
 wire \am_sdr0.cic1.integ_sample[13] ;
 wire \am_sdr0.cic1.integ_sample[14] ;
 wire \am_sdr0.cic1.integ_sample[15] ;
 wire \am_sdr0.cic1.integ_sample[16] ;
 wire \am_sdr0.cic1.integ_sample[17] ;
 wire \am_sdr0.cic1.integ_sample[18] ;
 wire \am_sdr0.cic1.integ_sample[19] ;
 wire \am_sdr0.cic1.integ_sample[1] ;
 wire \am_sdr0.cic1.integ_sample[2] ;
 wire \am_sdr0.cic1.integ_sample[3] ;
 wire \am_sdr0.cic1.integ_sample[4] ;
 wire \am_sdr0.cic1.integ_sample[5] ;
 wire \am_sdr0.cic1.integ_sample[6] ;
 wire \am_sdr0.cic1.integ_sample[7] ;
 wire \am_sdr0.cic1.integ_sample[8] ;
 wire \am_sdr0.cic1.integ_sample[9] ;
 wire \am_sdr0.cic1.out_tick ;
 wire \am_sdr0.cic1.sample ;
 wire \am_sdr0.cic1.x_out[10] ;
 wire \am_sdr0.cic1.x_out[11] ;
 wire \am_sdr0.cic1.x_out[12] ;
 wire \am_sdr0.cic1.x_out[13] ;
 wire \am_sdr0.cic1.x_out[14] ;
 wire \am_sdr0.cic1.x_out[15] ;
 wire \am_sdr0.cic1.x_out[8] ;
 wire \am_sdr0.cic1.x_out[9] ;
 wire \am_sdr0.cic2.comb1[0] ;
 wire \am_sdr0.cic2.comb1[10] ;
 wire \am_sdr0.cic2.comb1[11] ;
 wire \am_sdr0.cic2.comb1[12] ;
 wire \am_sdr0.cic2.comb1[13] ;
 wire \am_sdr0.cic2.comb1[14] ;
 wire \am_sdr0.cic2.comb1[15] ;
 wire \am_sdr0.cic2.comb1[16] ;
 wire \am_sdr0.cic2.comb1[17] ;
 wire \am_sdr0.cic2.comb1[18] ;
 wire \am_sdr0.cic2.comb1[19] ;
 wire \am_sdr0.cic2.comb1[1] ;
 wire \am_sdr0.cic2.comb1[2] ;
 wire \am_sdr0.cic2.comb1[3] ;
 wire \am_sdr0.cic2.comb1[4] ;
 wire \am_sdr0.cic2.comb1[5] ;
 wire \am_sdr0.cic2.comb1[6] ;
 wire \am_sdr0.cic2.comb1[7] ;
 wire \am_sdr0.cic2.comb1[8] ;
 wire \am_sdr0.cic2.comb1[9] ;
 wire \am_sdr0.cic2.comb1_in_del[0] ;
 wire \am_sdr0.cic2.comb1_in_del[10] ;
 wire \am_sdr0.cic2.comb1_in_del[11] ;
 wire \am_sdr0.cic2.comb1_in_del[12] ;
 wire \am_sdr0.cic2.comb1_in_del[13] ;
 wire \am_sdr0.cic2.comb1_in_del[14] ;
 wire \am_sdr0.cic2.comb1_in_del[15] ;
 wire \am_sdr0.cic2.comb1_in_del[16] ;
 wire \am_sdr0.cic2.comb1_in_del[17] ;
 wire \am_sdr0.cic2.comb1_in_del[18] ;
 wire \am_sdr0.cic2.comb1_in_del[19] ;
 wire \am_sdr0.cic2.comb1_in_del[1] ;
 wire \am_sdr0.cic2.comb1_in_del[2] ;
 wire \am_sdr0.cic2.comb1_in_del[3] ;
 wire \am_sdr0.cic2.comb1_in_del[4] ;
 wire \am_sdr0.cic2.comb1_in_del[5] ;
 wire \am_sdr0.cic2.comb1_in_del[6] ;
 wire \am_sdr0.cic2.comb1_in_del[7] ;
 wire \am_sdr0.cic2.comb1_in_del[8] ;
 wire \am_sdr0.cic2.comb1_in_del[9] ;
 wire \am_sdr0.cic2.comb2[0] ;
 wire \am_sdr0.cic2.comb2[10] ;
 wire \am_sdr0.cic2.comb2[11] ;
 wire \am_sdr0.cic2.comb2[12] ;
 wire \am_sdr0.cic2.comb2[13] ;
 wire \am_sdr0.cic2.comb2[14] ;
 wire \am_sdr0.cic2.comb2[15] ;
 wire \am_sdr0.cic2.comb2[16] ;
 wire \am_sdr0.cic2.comb2[17] ;
 wire \am_sdr0.cic2.comb2[18] ;
 wire \am_sdr0.cic2.comb2[19] ;
 wire \am_sdr0.cic2.comb2[1] ;
 wire \am_sdr0.cic2.comb2[2] ;
 wire \am_sdr0.cic2.comb2[3] ;
 wire \am_sdr0.cic2.comb2[4] ;
 wire \am_sdr0.cic2.comb2[5] ;
 wire \am_sdr0.cic2.comb2[6] ;
 wire \am_sdr0.cic2.comb2[7] ;
 wire \am_sdr0.cic2.comb2[8] ;
 wire \am_sdr0.cic2.comb2[9] ;
 wire \am_sdr0.cic2.comb2_in_del[0] ;
 wire \am_sdr0.cic2.comb2_in_del[10] ;
 wire \am_sdr0.cic2.comb2_in_del[11] ;
 wire \am_sdr0.cic2.comb2_in_del[12] ;
 wire \am_sdr0.cic2.comb2_in_del[13] ;
 wire \am_sdr0.cic2.comb2_in_del[14] ;
 wire \am_sdr0.cic2.comb2_in_del[15] ;
 wire \am_sdr0.cic2.comb2_in_del[16] ;
 wire \am_sdr0.cic2.comb2_in_del[17] ;
 wire \am_sdr0.cic2.comb2_in_del[18] ;
 wire \am_sdr0.cic2.comb2_in_del[19] ;
 wire \am_sdr0.cic2.comb2_in_del[1] ;
 wire \am_sdr0.cic2.comb2_in_del[2] ;
 wire \am_sdr0.cic2.comb2_in_del[3] ;
 wire \am_sdr0.cic2.comb2_in_del[4] ;
 wire \am_sdr0.cic2.comb2_in_del[5] ;
 wire \am_sdr0.cic2.comb2_in_del[6] ;
 wire \am_sdr0.cic2.comb2_in_del[7] ;
 wire \am_sdr0.cic2.comb2_in_del[8] ;
 wire \am_sdr0.cic2.comb2_in_del[9] ;
 wire \am_sdr0.cic2.comb3[12] ;
 wire \am_sdr0.cic2.comb3[13] ;
 wire \am_sdr0.cic2.comb3[14] ;
 wire \am_sdr0.cic2.comb3[15] ;
 wire \am_sdr0.cic2.comb3[16] ;
 wire \am_sdr0.cic2.comb3[17] ;
 wire \am_sdr0.cic2.comb3[18] ;
 wire \am_sdr0.cic2.comb3[19] ;
 wire \am_sdr0.cic2.comb3_in_del[0] ;
 wire \am_sdr0.cic2.comb3_in_del[10] ;
 wire \am_sdr0.cic2.comb3_in_del[11] ;
 wire \am_sdr0.cic2.comb3_in_del[12] ;
 wire \am_sdr0.cic2.comb3_in_del[13] ;
 wire \am_sdr0.cic2.comb3_in_del[14] ;
 wire \am_sdr0.cic2.comb3_in_del[15] ;
 wire \am_sdr0.cic2.comb3_in_del[16] ;
 wire \am_sdr0.cic2.comb3_in_del[17] ;
 wire \am_sdr0.cic2.comb3_in_del[18] ;
 wire \am_sdr0.cic2.comb3_in_del[19] ;
 wire \am_sdr0.cic2.comb3_in_del[1] ;
 wire \am_sdr0.cic2.comb3_in_del[2] ;
 wire \am_sdr0.cic2.comb3_in_del[3] ;
 wire \am_sdr0.cic2.comb3_in_del[4] ;
 wire \am_sdr0.cic2.comb3_in_del[5] ;
 wire \am_sdr0.cic2.comb3_in_del[6] ;
 wire \am_sdr0.cic2.comb3_in_del[7] ;
 wire \am_sdr0.cic2.comb3_in_del[8] ;
 wire \am_sdr0.cic2.comb3_in_del[9] ;
 wire \am_sdr0.cic2.count[0] ;
 wire \am_sdr0.cic2.count[1] ;
 wire \am_sdr0.cic2.count[2] ;
 wire \am_sdr0.cic2.count[3] ;
 wire \am_sdr0.cic2.count[4] ;
 wire \am_sdr0.cic2.count[5] ;
 wire \am_sdr0.cic2.count[6] ;
 wire \am_sdr0.cic2.count[7] ;
 wire \am_sdr0.cic2.integ1[0] ;
 wire \am_sdr0.cic2.integ1[10] ;
 wire \am_sdr0.cic2.integ1[11] ;
 wire \am_sdr0.cic2.integ1[12] ;
 wire \am_sdr0.cic2.integ1[13] ;
 wire \am_sdr0.cic2.integ1[14] ;
 wire \am_sdr0.cic2.integ1[15] ;
 wire \am_sdr0.cic2.integ1[16] ;
 wire \am_sdr0.cic2.integ1[17] ;
 wire \am_sdr0.cic2.integ1[18] ;
 wire \am_sdr0.cic2.integ1[19] ;
 wire \am_sdr0.cic2.integ1[1] ;
 wire \am_sdr0.cic2.integ1[20] ;
 wire \am_sdr0.cic2.integ1[21] ;
 wire \am_sdr0.cic2.integ1[22] ;
 wire \am_sdr0.cic2.integ1[23] ;
 wire \am_sdr0.cic2.integ1[24] ;
 wire \am_sdr0.cic2.integ1[25] ;
 wire \am_sdr0.cic2.integ1[2] ;
 wire \am_sdr0.cic2.integ1[3] ;
 wire \am_sdr0.cic2.integ1[4] ;
 wire \am_sdr0.cic2.integ1[5] ;
 wire \am_sdr0.cic2.integ1[6] ;
 wire \am_sdr0.cic2.integ1[7] ;
 wire \am_sdr0.cic2.integ1[8] ;
 wire \am_sdr0.cic2.integ1[9] ;
 wire \am_sdr0.cic2.integ2[0] ;
 wire \am_sdr0.cic2.integ2[10] ;
 wire \am_sdr0.cic2.integ2[11] ;
 wire \am_sdr0.cic2.integ2[12] ;
 wire \am_sdr0.cic2.integ2[13] ;
 wire \am_sdr0.cic2.integ2[14] ;
 wire \am_sdr0.cic2.integ2[15] ;
 wire \am_sdr0.cic2.integ2[16] ;
 wire \am_sdr0.cic2.integ2[17] ;
 wire \am_sdr0.cic2.integ2[18] ;
 wire \am_sdr0.cic2.integ2[19] ;
 wire \am_sdr0.cic2.integ2[1] ;
 wire \am_sdr0.cic2.integ2[20] ;
 wire \am_sdr0.cic2.integ2[21] ;
 wire \am_sdr0.cic2.integ2[22] ;
 wire \am_sdr0.cic2.integ2[2] ;
 wire \am_sdr0.cic2.integ2[3] ;
 wire \am_sdr0.cic2.integ2[4] ;
 wire \am_sdr0.cic2.integ2[5] ;
 wire \am_sdr0.cic2.integ2[6] ;
 wire \am_sdr0.cic2.integ2[7] ;
 wire \am_sdr0.cic2.integ2[8] ;
 wire \am_sdr0.cic2.integ2[9] ;
 wire \am_sdr0.cic2.integ3[0] ;
 wire \am_sdr0.cic2.integ3[10] ;
 wire \am_sdr0.cic2.integ3[11] ;
 wire \am_sdr0.cic2.integ3[12] ;
 wire \am_sdr0.cic2.integ3[13] ;
 wire \am_sdr0.cic2.integ3[14] ;
 wire \am_sdr0.cic2.integ3[15] ;
 wire \am_sdr0.cic2.integ3[16] ;
 wire \am_sdr0.cic2.integ3[17] ;
 wire \am_sdr0.cic2.integ3[18] ;
 wire \am_sdr0.cic2.integ3[19] ;
 wire \am_sdr0.cic2.integ3[1] ;
 wire \am_sdr0.cic2.integ3[2] ;
 wire \am_sdr0.cic2.integ3[3] ;
 wire \am_sdr0.cic2.integ3[4] ;
 wire \am_sdr0.cic2.integ3[5] ;
 wire \am_sdr0.cic2.integ3[6] ;
 wire \am_sdr0.cic2.integ3[7] ;
 wire \am_sdr0.cic2.integ3[8] ;
 wire \am_sdr0.cic2.integ3[9] ;
 wire \am_sdr0.cic2.integ_sample[0] ;
 wire \am_sdr0.cic2.integ_sample[10] ;
 wire \am_sdr0.cic2.integ_sample[11] ;
 wire \am_sdr0.cic2.integ_sample[12] ;
 wire \am_sdr0.cic2.integ_sample[13] ;
 wire \am_sdr0.cic2.integ_sample[14] ;
 wire \am_sdr0.cic2.integ_sample[15] ;
 wire \am_sdr0.cic2.integ_sample[16] ;
 wire \am_sdr0.cic2.integ_sample[17] ;
 wire \am_sdr0.cic2.integ_sample[18] ;
 wire \am_sdr0.cic2.integ_sample[19] ;
 wire \am_sdr0.cic2.integ_sample[1] ;
 wire \am_sdr0.cic2.integ_sample[2] ;
 wire \am_sdr0.cic2.integ_sample[3] ;
 wire \am_sdr0.cic2.integ_sample[4] ;
 wire \am_sdr0.cic2.integ_sample[5] ;
 wire \am_sdr0.cic2.integ_sample[6] ;
 wire \am_sdr0.cic2.integ_sample[7] ;
 wire \am_sdr0.cic2.integ_sample[8] ;
 wire \am_sdr0.cic2.integ_sample[9] ;
 wire \am_sdr0.cic2.sample ;
 wire \am_sdr0.cic3.comb1[0] ;
 wire \am_sdr0.cic3.comb1[10] ;
 wire \am_sdr0.cic3.comb1[11] ;
 wire \am_sdr0.cic3.comb1[12] ;
 wire \am_sdr0.cic3.comb1[13] ;
 wire \am_sdr0.cic3.comb1[14] ;
 wire \am_sdr0.cic3.comb1[15] ;
 wire \am_sdr0.cic3.comb1[16] ;
 wire \am_sdr0.cic3.comb1[17] ;
 wire \am_sdr0.cic3.comb1[18] ;
 wire \am_sdr0.cic3.comb1[19] ;
 wire \am_sdr0.cic3.comb1[1] ;
 wire \am_sdr0.cic3.comb1[2] ;
 wire \am_sdr0.cic3.comb1[3] ;
 wire \am_sdr0.cic3.comb1[4] ;
 wire \am_sdr0.cic3.comb1[5] ;
 wire \am_sdr0.cic3.comb1[6] ;
 wire \am_sdr0.cic3.comb1[7] ;
 wire \am_sdr0.cic3.comb1[8] ;
 wire \am_sdr0.cic3.comb1[9] ;
 wire \am_sdr0.cic3.comb1_in_del[0] ;
 wire \am_sdr0.cic3.comb1_in_del[10] ;
 wire \am_sdr0.cic3.comb1_in_del[11] ;
 wire \am_sdr0.cic3.comb1_in_del[12] ;
 wire \am_sdr0.cic3.comb1_in_del[13] ;
 wire \am_sdr0.cic3.comb1_in_del[14] ;
 wire \am_sdr0.cic3.comb1_in_del[15] ;
 wire \am_sdr0.cic3.comb1_in_del[16] ;
 wire \am_sdr0.cic3.comb1_in_del[17] ;
 wire \am_sdr0.cic3.comb1_in_del[18] ;
 wire \am_sdr0.cic3.comb1_in_del[19] ;
 wire \am_sdr0.cic3.comb1_in_del[1] ;
 wire \am_sdr0.cic3.comb1_in_del[2] ;
 wire \am_sdr0.cic3.comb1_in_del[3] ;
 wire \am_sdr0.cic3.comb1_in_del[4] ;
 wire \am_sdr0.cic3.comb1_in_del[5] ;
 wire \am_sdr0.cic3.comb1_in_del[6] ;
 wire \am_sdr0.cic3.comb1_in_del[7] ;
 wire \am_sdr0.cic3.comb1_in_del[8] ;
 wire \am_sdr0.cic3.comb1_in_del[9] ;
 wire \am_sdr0.cic3.comb2[0] ;
 wire \am_sdr0.cic3.comb2[10] ;
 wire \am_sdr0.cic3.comb2[11] ;
 wire \am_sdr0.cic3.comb2[12] ;
 wire \am_sdr0.cic3.comb2[13] ;
 wire \am_sdr0.cic3.comb2[14] ;
 wire \am_sdr0.cic3.comb2[15] ;
 wire \am_sdr0.cic3.comb2[16] ;
 wire \am_sdr0.cic3.comb2[17] ;
 wire \am_sdr0.cic3.comb2[18] ;
 wire \am_sdr0.cic3.comb2[19] ;
 wire \am_sdr0.cic3.comb2[1] ;
 wire \am_sdr0.cic3.comb2[2] ;
 wire \am_sdr0.cic3.comb2[3] ;
 wire \am_sdr0.cic3.comb2[4] ;
 wire \am_sdr0.cic3.comb2[5] ;
 wire \am_sdr0.cic3.comb2[6] ;
 wire \am_sdr0.cic3.comb2[7] ;
 wire \am_sdr0.cic3.comb2[8] ;
 wire \am_sdr0.cic3.comb2[9] ;
 wire \am_sdr0.cic3.comb2_in_del[0] ;
 wire \am_sdr0.cic3.comb2_in_del[10] ;
 wire \am_sdr0.cic3.comb2_in_del[11] ;
 wire \am_sdr0.cic3.comb2_in_del[12] ;
 wire \am_sdr0.cic3.comb2_in_del[13] ;
 wire \am_sdr0.cic3.comb2_in_del[14] ;
 wire \am_sdr0.cic3.comb2_in_del[15] ;
 wire \am_sdr0.cic3.comb2_in_del[16] ;
 wire \am_sdr0.cic3.comb2_in_del[17] ;
 wire \am_sdr0.cic3.comb2_in_del[18] ;
 wire \am_sdr0.cic3.comb2_in_del[19] ;
 wire \am_sdr0.cic3.comb2_in_del[1] ;
 wire \am_sdr0.cic3.comb2_in_del[2] ;
 wire \am_sdr0.cic3.comb2_in_del[3] ;
 wire \am_sdr0.cic3.comb2_in_del[4] ;
 wire \am_sdr0.cic3.comb2_in_del[5] ;
 wire \am_sdr0.cic3.comb2_in_del[6] ;
 wire \am_sdr0.cic3.comb2_in_del[7] ;
 wire \am_sdr0.cic3.comb2_in_del[8] ;
 wire \am_sdr0.cic3.comb2_in_del[9] ;
 wire \am_sdr0.cic3.comb3[12] ;
 wire \am_sdr0.cic3.comb3[13] ;
 wire \am_sdr0.cic3.comb3[14] ;
 wire \am_sdr0.cic3.comb3[15] ;
 wire \am_sdr0.cic3.comb3[16] ;
 wire \am_sdr0.cic3.comb3[17] ;
 wire \am_sdr0.cic3.comb3[18] ;
 wire \am_sdr0.cic3.comb3[19] ;
 wire \am_sdr0.cic3.comb3_in_del[0] ;
 wire \am_sdr0.cic3.comb3_in_del[10] ;
 wire \am_sdr0.cic3.comb3_in_del[11] ;
 wire \am_sdr0.cic3.comb3_in_del[12] ;
 wire \am_sdr0.cic3.comb3_in_del[13] ;
 wire \am_sdr0.cic3.comb3_in_del[14] ;
 wire \am_sdr0.cic3.comb3_in_del[15] ;
 wire \am_sdr0.cic3.comb3_in_del[16] ;
 wire \am_sdr0.cic3.comb3_in_del[17] ;
 wire \am_sdr0.cic3.comb3_in_del[18] ;
 wire \am_sdr0.cic3.comb3_in_del[19] ;
 wire \am_sdr0.cic3.comb3_in_del[1] ;
 wire \am_sdr0.cic3.comb3_in_del[2] ;
 wire \am_sdr0.cic3.comb3_in_del[3] ;
 wire \am_sdr0.cic3.comb3_in_del[4] ;
 wire \am_sdr0.cic3.comb3_in_del[5] ;
 wire \am_sdr0.cic3.comb3_in_del[6] ;
 wire \am_sdr0.cic3.comb3_in_del[7] ;
 wire \am_sdr0.cic3.comb3_in_del[8] ;
 wire \am_sdr0.cic3.comb3_in_del[9] ;
 wire \am_sdr0.cic3.count[0] ;
 wire \am_sdr0.cic3.count[1] ;
 wire \am_sdr0.cic3.count[2] ;
 wire \am_sdr0.cic3.count[3] ;
 wire \am_sdr0.cic3.count[4] ;
 wire \am_sdr0.cic3.count[5] ;
 wire \am_sdr0.cic3.count[6] ;
 wire \am_sdr0.cic3.count[7] ;
 wire \am_sdr0.cic3.integ1[0] ;
 wire \am_sdr0.cic3.integ1[10] ;
 wire \am_sdr0.cic3.integ1[11] ;
 wire \am_sdr0.cic3.integ1[12] ;
 wire \am_sdr0.cic3.integ1[13] ;
 wire \am_sdr0.cic3.integ1[14] ;
 wire \am_sdr0.cic3.integ1[15] ;
 wire \am_sdr0.cic3.integ1[16] ;
 wire \am_sdr0.cic3.integ1[17] ;
 wire \am_sdr0.cic3.integ1[18] ;
 wire \am_sdr0.cic3.integ1[19] ;
 wire \am_sdr0.cic3.integ1[1] ;
 wire \am_sdr0.cic3.integ1[20] ;
 wire \am_sdr0.cic3.integ1[21] ;
 wire \am_sdr0.cic3.integ1[22] ;
 wire \am_sdr0.cic3.integ1[23] ;
 wire \am_sdr0.cic3.integ1[24] ;
 wire \am_sdr0.cic3.integ1[25] ;
 wire \am_sdr0.cic3.integ1[2] ;
 wire \am_sdr0.cic3.integ1[3] ;
 wire \am_sdr0.cic3.integ1[4] ;
 wire \am_sdr0.cic3.integ1[5] ;
 wire \am_sdr0.cic3.integ1[6] ;
 wire \am_sdr0.cic3.integ1[7] ;
 wire \am_sdr0.cic3.integ1[8] ;
 wire \am_sdr0.cic3.integ1[9] ;
 wire \am_sdr0.cic3.integ2[0] ;
 wire \am_sdr0.cic3.integ2[10] ;
 wire \am_sdr0.cic3.integ2[11] ;
 wire \am_sdr0.cic3.integ2[12] ;
 wire \am_sdr0.cic3.integ2[13] ;
 wire \am_sdr0.cic3.integ2[14] ;
 wire \am_sdr0.cic3.integ2[15] ;
 wire \am_sdr0.cic3.integ2[16] ;
 wire \am_sdr0.cic3.integ2[17] ;
 wire \am_sdr0.cic3.integ2[18] ;
 wire \am_sdr0.cic3.integ2[19] ;
 wire \am_sdr0.cic3.integ2[1] ;
 wire \am_sdr0.cic3.integ2[20] ;
 wire \am_sdr0.cic3.integ2[21] ;
 wire \am_sdr0.cic3.integ2[22] ;
 wire \am_sdr0.cic3.integ2[2] ;
 wire \am_sdr0.cic3.integ2[3] ;
 wire \am_sdr0.cic3.integ2[4] ;
 wire \am_sdr0.cic3.integ2[5] ;
 wire \am_sdr0.cic3.integ2[6] ;
 wire \am_sdr0.cic3.integ2[7] ;
 wire \am_sdr0.cic3.integ2[8] ;
 wire \am_sdr0.cic3.integ2[9] ;
 wire \am_sdr0.cic3.integ3[0] ;
 wire \am_sdr0.cic3.integ3[10] ;
 wire \am_sdr0.cic3.integ3[11] ;
 wire \am_sdr0.cic3.integ3[12] ;
 wire \am_sdr0.cic3.integ3[13] ;
 wire \am_sdr0.cic3.integ3[14] ;
 wire \am_sdr0.cic3.integ3[15] ;
 wire \am_sdr0.cic3.integ3[16] ;
 wire \am_sdr0.cic3.integ3[17] ;
 wire \am_sdr0.cic3.integ3[18] ;
 wire \am_sdr0.cic3.integ3[19] ;
 wire \am_sdr0.cic3.integ3[1] ;
 wire \am_sdr0.cic3.integ3[2] ;
 wire \am_sdr0.cic3.integ3[3] ;
 wire \am_sdr0.cic3.integ3[4] ;
 wire \am_sdr0.cic3.integ3[5] ;
 wire \am_sdr0.cic3.integ3[6] ;
 wire \am_sdr0.cic3.integ3[7] ;
 wire \am_sdr0.cic3.integ3[8] ;
 wire \am_sdr0.cic3.integ3[9] ;
 wire \am_sdr0.cic3.integ_sample[0] ;
 wire \am_sdr0.cic3.integ_sample[10] ;
 wire \am_sdr0.cic3.integ_sample[11] ;
 wire \am_sdr0.cic3.integ_sample[12] ;
 wire \am_sdr0.cic3.integ_sample[13] ;
 wire \am_sdr0.cic3.integ_sample[14] ;
 wire \am_sdr0.cic3.integ_sample[15] ;
 wire \am_sdr0.cic3.integ_sample[16] ;
 wire \am_sdr0.cic3.integ_sample[17] ;
 wire \am_sdr0.cic3.integ_sample[18] ;
 wire \am_sdr0.cic3.integ_sample[19] ;
 wire \am_sdr0.cic3.integ_sample[1] ;
 wire \am_sdr0.cic3.integ_sample[2] ;
 wire \am_sdr0.cic3.integ_sample[3] ;
 wire \am_sdr0.cic3.integ_sample[4] ;
 wire \am_sdr0.cic3.integ_sample[5] ;
 wire \am_sdr0.cic3.integ_sample[6] ;
 wire \am_sdr0.cic3.integ_sample[7] ;
 wire \am_sdr0.cic3.integ_sample[8] ;
 wire \am_sdr0.cic3.integ_sample[9] ;
 wire \am_sdr0.cic3.sample ;
 wire \am_sdr0.cos[0] ;
 wire \am_sdr0.cos[1] ;
 wire \am_sdr0.cos[2] ;
 wire \am_sdr0.cos[3] ;
 wire \am_sdr0.cos[4] ;
 wire \am_sdr0.cos[5] ;
 wire \am_sdr0.cos[6] ;
 wire \am_sdr0.cos[7] ;
 wire \am_sdr0.count[0] ;
 wire \am_sdr0.count[1] ;
 wire \am_sdr0.count[2] ;
 wire \am_sdr0.count[3] ;
 wire \am_sdr0.count[4] ;
 wire \am_sdr0.count[5] ;
 wire \am_sdr0.count[6] ;
 wire \am_sdr0.count[7] ;
 wire \am_sdr0.gain_spi[0] ;
 wire \am_sdr0.gain_spi[1] ;
 wire \am_sdr0.gain_spi[2] ;
 wire \am_sdr0.mix0.RF_in_q ;
 wire \am_sdr0.mix0.RF_in_qq ;
 wire \am_sdr0.mix0.cos_q[0] ;
 wire \am_sdr0.mix0.cos_q[1] ;
 wire \am_sdr0.mix0.cos_q[2] ;
 wire \am_sdr0.mix0.cos_q[3] ;
 wire \am_sdr0.mix0.cos_q[4] ;
 wire \am_sdr0.mix0.cos_q[5] ;
 wire \am_sdr0.mix0.cos_q[6] ;
 wire \am_sdr0.mix0.cos_q[7] ;
 wire \am_sdr0.mix0.sin_in[0] ;
 wire \am_sdr0.mix0.sin_in[1] ;
 wire \am_sdr0.mix0.sin_in[2] ;
 wire \am_sdr0.mix0.sin_in[3] ;
 wire \am_sdr0.mix0.sin_in[4] ;
 wire \am_sdr0.mix0.sin_in[5] ;
 wire \am_sdr0.mix0.sin_in[6] ;
 wire \am_sdr0.mix0.sin_in[7] ;
 wire \am_sdr0.mix0.sin_q[0] ;
 wire \am_sdr0.mix0.sin_q[1] ;
 wire \am_sdr0.mix0.sin_q[2] ;
 wire \am_sdr0.mix0.sin_q[3] ;
 wire \am_sdr0.mix0.sin_q[4] ;
 wire \am_sdr0.mix0.sin_q[5] ;
 wire \am_sdr0.mix0.sin_q[6] ;
 wire \am_sdr0.mix0.sin_q[7] ;
 wire \am_sdr0.nco0.phase[0] ;
 wire \am_sdr0.nco0.phase[10] ;
 wire \am_sdr0.nco0.phase[11] ;
 wire \am_sdr0.nco0.phase[12] ;
 wire \am_sdr0.nco0.phase[13] ;
 wire \am_sdr0.nco0.phase[14] ;
 wire \am_sdr0.nco0.phase[15] ;
 wire \am_sdr0.nco0.phase[16] ;
 wire \am_sdr0.nco0.phase[17] ;
 wire \am_sdr0.nco0.phase[18] ;
 wire \am_sdr0.nco0.phase[19] ;
 wire \am_sdr0.nco0.phase[1] ;
 wire \am_sdr0.nco0.phase[20] ;
 wire \am_sdr0.nco0.phase[21] ;
 wire \am_sdr0.nco0.phase[22] ;
 wire \am_sdr0.nco0.phase[23] ;
 wire \am_sdr0.nco0.phase[24] ;
 wire \am_sdr0.nco0.phase[25] ;
 wire \am_sdr0.nco0.phase[2] ;
 wire \am_sdr0.nco0.phase[3] ;
 wire \am_sdr0.nco0.phase[4] ;
 wire \am_sdr0.nco0.phase[5] ;
 wire \am_sdr0.nco0.phase[6] ;
 wire \am_sdr0.nco0.phase[7] ;
 wire \am_sdr0.nco0.phase[8] ;
 wire \am_sdr0.nco0.phase[9] ;
 wire \am_sdr0.nco0.phase_inc[0] ;
 wire \am_sdr0.nco0.phase_inc[10] ;
 wire \am_sdr0.nco0.phase_inc[11] ;
 wire \am_sdr0.nco0.phase_inc[12] ;
 wire \am_sdr0.nco0.phase_inc[13] ;
 wire \am_sdr0.nco0.phase_inc[14] ;
 wire \am_sdr0.nco0.phase_inc[15] ;
 wire \am_sdr0.nco0.phase_inc[16] ;
 wire \am_sdr0.nco0.phase_inc[17] ;
 wire \am_sdr0.nco0.phase_inc[18] ;
 wire \am_sdr0.nco0.phase_inc[19] ;
 wire \am_sdr0.nco0.phase_inc[1] ;
 wire \am_sdr0.nco0.phase_inc[20] ;
 wire \am_sdr0.nco0.phase_inc[21] ;
 wire \am_sdr0.nco0.phase_inc[22] ;
 wire \am_sdr0.nco0.phase_inc[23] ;
 wire \am_sdr0.nco0.phase_inc[24] ;
 wire \am_sdr0.nco0.phase_inc[25] ;
 wire \am_sdr0.nco0.phase_inc[2] ;
 wire \am_sdr0.nco0.phase_inc[3] ;
 wire \am_sdr0.nco0.phase_inc[4] ;
 wire \am_sdr0.nco0.phase_inc[5] ;
 wire \am_sdr0.nco0.phase_inc[6] ;
 wire \am_sdr0.nco0.phase_inc[7] ;
 wire \am_sdr0.nco0.phase_inc[8] ;
 wire \am_sdr0.nco0.phase_inc[9] ;
 wire \am_sdr0.spi0.CS_q ;
 wire \am_sdr0.spi0.CS_qq ;
 wire \am_sdr0.spi0.CS_qqq ;
 wire \am_sdr0.spi0.MOSI_q ;
 wire \am_sdr0.spi0.MOSI_qq ;
 wire \am_sdr0.spi0.SCK_q ;
 wire \am_sdr0.spi0.SCK_qq ;
 wire \am_sdr0.spi0.SCK_qqq ;
 wire \am_sdr0.spi0.shift_reg[0] ;
 wire \am_sdr0.spi0.shift_reg[10] ;
 wire \am_sdr0.spi0.shift_reg[11] ;
 wire \am_sdr0.spi0.shift_reg[12] ;
 wire \am_sdr0.spi0.shift_reg[13] ;
 wire \am_sdr0.spi0.shift_reg[14] ;
 wire \am_sdr0.spi0.shift_reg[15] ;
 wire \am_sdr0.spi0.shift_reg[16] ;
 wire \am_sdr0.spi0.shift_reg[17] ;
 wire \am_sdr0.spi0.shift_reg[18] ;
 wire \am_sdr0.spi0.shift_reg[19] ;
 wire \am_sdr0.spi0.shift_reg[1] ;
 wire \am_sdr0.spi0.shift_reg[20] ;
 wire \am_sdr0.spi0.shift_reg[21] ;
 wire \am_sdr0.spi0.shift_reg[22] ;
 wire \am_sdr0.spi0.shift_reg[23] ;
 wire \am_sdr0.spi0.shift_reg[24] ;
 wire \am_sdr0.spi0.shift_reg[25] ;
 wire \am_sdr0.spi0.shift_reg[26] ;
 wire \am_sdr0.spi0.shift_reg[27] ;
 wire \am_sdr0.spi0.shift_reg[28] ;
 wire \am_sdr0.spi0.shift_reg[2] ;
 wire \am_sdr0.spi0.shift_reg[3] ;
 wire \am_sdr0.spi0.shift_reg[4] ;
 wire \am_sdr0.spi0.shift_reg[5] ;
 wire \am_sdr0.spi0.shift_reg[6] ;
 wire \am_sdr0.spi0.shift_reg[7] ;
 wire \am_sdr0.spi0.shift_reg[8] ;
 wire \am_sdr0.spi0.shift_reg[9] ;
 wire \am_sdr0.spi0.state[0] ;
 wire \am_sdr0.spi0.state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _09161_ (.A(rst_n),
    .X(_01442_));
 sg13g2_inv_1 _09162_ (.Y(_01443_),
    .A(_01442_));
 sg13g2_buf_1 _09163_ (.A(_01443_),
    .X(_01444_));
 sg13g2_buf_1 _09164_ (.A(net310),
    .X(_01445_));
 sg13g2_buf_1 _09165_ (.A(net259),
    .X(_01446_));
 sg13g2_buf_1 _09166_ (.A(net191),
    .X(_01447_));
 sg13g2_buf_1 _09167_ (.A(\am_sdr0.am0.state[2] ),
    .X(_01448_));
 sg13g2_buf_2 _09168_ (.A(\am_sdr0.am0.m_count[3] ),
    .X(_01449_));
 sg13g2_inv_1 _09169_ (.Y(_01450_),
    .A(_01449_));
 sg13g2_buf_1 _09170_ (.A(\am_sdr0.am0.m_count[1] ),
    .X(_01451_));
 sg13g2_buf_2 _09171_ (.A(\am_sdr0.am0.m_count[0] ),
    .X(_01452_));
 sg13g2_buf_1 _09172_ (.A(\am_sdr0.am0.m_count[2] ),
    .X(_01453_));
 sg13g2_and3_1 _09173_ (.X(_01454_),
    .A(_01451_),
    .B(_01452_),
    .C(_01453_));
 sg13g2_nand2_1 _09174_ (.Y(_01455_),
    .A(_01450_),
    .B(_01454_));
 sg13g2_buf_8 _09175_ (.A(_01455_),
    .X(_01456_));
 sg13g2_a21oi_1 _09176_ (.A1(_01448_),
    .A2(net190),
    .Y(_01457_),
    .B1(\am_sdr0.am0.state[4] ));
 sg13g2_nor2_1 _09177_ (.A(net139),
    .B(_01457_),
    .Y(_00020_));
 sg13g2_buf_1 _09178_ (.A(\am_sdr0.am0.sqrt_done ),
    .X(_01458_));
 sg13g2_inv_1 _09179_ (.Y(_01459_),
    .A(_01458_));
 sg13g2_a21oi_1 _09180_ (.A1(_01459_),
    .A2(\am_sdr0.am0.state[6] ),
    .Y(_01460_),
    .B1(\am_sdr0.am0.state[3] ));
 sg13g2_nor2_1 _09181_ (.A(_01447_),
    .B(_01460_),
    .Y(_00021_));
 sg13g2_buf_1 _09182_ (.A(\am_sdr0.am0.state[1] ),
    .X(_01461_));
 sg13g2_buf_1 _09183_ (.A(\am_sdr0.am0.state[5] ),
    .X(_01462_));
 sg13g2_buf_1 _09184_ (.A(net367),
    .X(_01463_));
 sg13g2_a21oi_1 _09185_ (.A1(_01461_),
    .A2(net190),
    .Y(_01464_),
    .B1(_01463_));
 sg13g2_nor2_1 _09186_ (.A(_01447_),
    .B(_01464_),
    .Y(_00019_));
 sg13g2_inv_1 _09187_ (.Y(_01465_),
    .A(\am_sdr0.am0.state[0] ));
 sg13g2_o21ai_1 _09188_ (.B1(_01442_),
    .Y(_01466_),
    .A1(_01465_),
    .A2(\am_sdr0.am0.load_tick ));
 sg13g2_buf_1 _09189_ (.A(_01466_),
    .X(_01467_));
 sg13g2_a21o_1 _09190_ (.A2(\am_sdr0.am0.state[6] ),
    .A1(_01458_),
    .B1(_01467_),
    .X(_00018_));
 sg13g2_buf_1 _09191_ (.A(\am_sdr0.mix0.RF_in_qq ),
    .X(_01468_));
 sg13g2_buf_1 _09192_ (.A(_01468_),
    .X(_01469_));
 sg13g2_inv_1 _09193_ (.Y(_01470_),
    .A(net308));
 sg13g2_nand2_1 _09194_ (.Y(_01471_),
    .A(\am_sdr0.mix0.sin_q[0] ),
    .B(_01470_));
 sg13g2_xnor2_1 _09195_ (.Y(_00030_),
    .A(\am_sdr0.mix0.sin_q[1] ),
    .B(_01471_));
 sg13g2_o21ai_1 _09196_ (.B1(_01470_),
    .Y(_01472_),
    .A1(\am_sdr0.mix0.sin_q[0] ),
    .A2(\am_sdr0.mix0.sin_q[1] ));
 sg13g2_xnor2_1 _09197_ (.Y(_00031_),
    .A(\am_sdr0.mix0.sin_q[2] ),
    .B(_01472_));
 sg13g2_nor3_1 _09198_ (.A(\am_sdr0.mix0.sin_q[0] ),
    .B(\am_sdr0.mix0.sin_q[1] ),
    .C(\am_sdr0.mix0.sin_q[2] ),
    .Y(_01473_));
 sg13g2_nor2_1 _09199_ (.A(_01469_),
    .B(_01473_),
    .Y(_01474_));
 sg13g2_xor2_1 _09200_ (.B(_01474_),
    .A(\am_sdr0.mix0.sin_q[3] ),
    .X(_00032_));
 sg13g2_inv_1 _09201_ (.Y(_01475_),
    .A(\am_sdr0.mix0.sin_q[4] ));
 sg13g2_nor2b_1 _09202_ (.A(\am_sdr0.mix0.sin_q[3] ),
    .B_N(_01473_),
    .Y(_01476_));
 sg13g2_nor2_1 _09203_ (.A(net308),
    .B(_01476_),
    .Y(_01477_));
 sg13g2_xnor2_1 _09204_ (.Y(_00033_),
    .A(_01475_),
    .B(_01477_));
 sg13g2_a21oi_1 _09205_ (.A1(_01475_),
    .A2(_01476_),
    .Y(_01478_),
    .B1(_01468_));
 sg13g2_xor2_1 _09206_ (.B(_01478_),
    .A(\am_sdr0.mix0.sin_q[5] ),
    .X(_00034_));
 sg13g2_inv_1 _09207_ (.Y(_01479_),
    .A(\am_sdr0.mix0.sin_q[6] ));
 sg13g2_nor2_1 _09208_ (.A(\am_sdr0.mix0.sin_q[5] ),
    .B(_01478_),
    .Y(_01480_));
 sg13g2_nor2_1 _09209_ (.A(net308),
    .B(_01480_),
    .Y(_01481_));
 sg13g2_xnor2_1 _09210_ (.Y(_00035_),
    .A(_01479_),
    .B(_01481_));
 sg13g2_a21oi_1 _09211_ (.A1(_01479_),
    .A2(_01480_),
    .Y(_01482_),
    .B1(net308));
 sg13g2_xor2_1 _09212_ (.B(_01482_),
    .A(\am_sdr0.mix0.sin_q[7] ),
    .X(_00036_));
 sg13g2_nand2_1 _09213_ (.Y(_01483_),
    .A(_01470_),
    .B(\am_sdr0.mix0.cos_q[0] ));
 sg13g2_xnor2_1 _09214_ (.Y(_00023_),
    .A(\am_sdr0.mix0.cos_q[1] ),
    .B(_01483_));
 sg13g2_o21ai_1 _09215_ (.B1(_01470_),
    .Y(_01484_),
    .A1(\am_sdr0.mix0.cos_q[0] ),
    .A2(\am_sdr0.mix0.cos_q[1] ));
 sg13g2_xnor2_1 _09216_ (.Y(_00024_),
    .A(\am_sdr0.mix0.cos_q[2] ),
    .B(_01484_));
 sg13g2_nor3_1 _09217_ (.A(\am_sdr0.mix0.cos_q[0] ),
    .B(\am_sdr0.mix0.cos_q[1] ),
    .C(\am_sdr0.mix0.cos_q[2] ),
    .Y(_01485_));
 sg13g2_nor2_1 _09218_ (.A(net308),
    .B(_01485_),
    .Y(_01486_));
 sg13g2_xor2_1 _09219_ (.B(_01486_),
    .A(\am_sdr0.mix0.cos_q[3] ),
    .X(_00025_));
 sg13g2_inv_1 _09220_ (.Y(_01487_),
    .A(\am_sdr0.mix0.cos_q[4] ));
 sg13g2_nor2b_1 _09221_ (.A(\am_sdr0.mix0.cos_q[3] ),
    .B_N(_01485_),
    .Y(_01488_));
 sg13g2_nor2_1 _09222_ (.A(net308),
    .B(_01488_),
    .Y(_01489_));
 sg13g2_xnor2_1 _09223_ (.Y(_00026_),
    .A(_01487_),
    .B(_01489_));
 sg13g2_a21oi_1 _09224_ (.A1(_01487_),
    .A2(_01488_),
    .Y(_01490_),
    .B1(_01468_));
 sg13g2_xor2_1 _09225_ (.B(_01490_),
    .A(\am_sdr0.mix0.cos_q[5] ),
    .X(_00027_));
 sg13g2_inv_1 _09226_ (.Y(_01491_),
    .A(\am_sdr0.mix0.cos_q[6] ));
 sg13g2_nor2_1 _09227_ (.A(\am_sdr0.mix0.cos_q[5] ),
    .B(_01490_),
    .Y(_01492_));
 sg13g2_nor2_1 _09228_ (.A(net308),
    .B(_01492_),
    .Y(_01493_));
 sg13g2_xnor2_1 _09229_ (.Y(_00028_),
    .A(_01491_),
    .B(_01493_));
 sg13g2_a21oi_1 _09230_ (.A1(_01491_),
    .A2(_01492_),
    .Y(_01494_),
    .B1(net308));
 sg13g2_xor2_1 _09231_ (.B(_01494_),
    .A(\am_sdr0.mix0.cos_q[7] ),
    .X(_00029_));
 sg13g2_buf_1 _09232_ (.A(\am_sdr0.nco0.phase[25] ),
    .X(_01495_));
 sg13g2_buf_1 _09233_ (.A(net366),
    .X(_01496_));
 sg13g2_nor2_1 _09234_ (.A(_00037_),
    .B(net307),
    .Y(_01497_));
 sg13g2_buf_1 _09235_ (.A(\am_sdr0.nco0.phase[24] ),
    .X(_01498_));
 sg13g2_buf_1 _09236_ (.A(_01498_),
    .X(_01499_));
 sg13g2_buf_1 _09237_ (.A(net306),
    .X(_01500_));
 sg13g2_buf_2 _09238_ (.A(\am_sdr0.nco0.phase[23] ),
    .X(_01501_));
 sg13g2_buf_1 _09239_ (.A(\am_sdr0.nco0.phase[22] ),
    .X(_01502_));
 sg13g2_nand2_1 _09240_ (.Y(_01503_),
    .A(_01501_),
    .B(net365));
 sg13g2_buf_1 _09241_ (.A(_00038_),
    .X(_01504_));
 sg13g2_nand2_1 _09242_ (.Y(_01505_),
    .A(_01504_),
    .B(net258));
 sg13g2_o21ai_1 _09243_ (.B1(_01505_),
    .Y(_01506_),
    .A1(net258),
    .A2(_01503_));
 sg13g2_nor2_1 _09244_ (.A(_01497_),
    .B(_01506_),
    .Y(_00000_));
 sg13g2_inv_2 _09245_ (.Y(_01507_),
    .A(_01501_));
 sg13g2_buf_1 _09246_ (.A(_00039_),
    .X(_01508_));
 sg13g2_nand2_1 _09247_ (.Y(_01509_),
    .A(net366),
    .B(_01508_));
 sg13g2_or2_1 _09248_ (.X(_01510_),
    .B(net366),
    .A(net306));
 sg13g2_inv_2 _09249_ (.Y(_01511_),
    .A(_01502_));
 sg13g2_mux2_1 _09250_ (.A0(_01509_),
    .A1(_01510_),
    .S(_01511_),
    .X(_01512_));
 sg13g2_buf_1 _09251_ (.A(net365),
    .X(_01513_));
 sg13g2_inv_2 _09252_ (.Y(_01514_),
    .A(net366));
 sg13g2_nand2_2 _09253_ (.Y(_01515_),
    .A(_01498_),
    .B(_01514_));
 sg13g2_o21ai_1 _09254_ (.B1(_01515_),
    .Y(_01516_),
    .A1(net305),
    .A2(_01509_));
 sg13g2_nor2_1 _09255_ (.A(_01507_),
    .B(_01516_),
    .Y(_01517_));
 sg13g2_a21oi_1 _09256_ (.A1(_01507_),
    .A2(_01512_),
    .Y(_00001_),
    .B1(_01517_));
 sg13g2_nor2_1 _09257_ (.A(_01499_),
    .B(_01495_),
    .Y(_01518_));
 sg13g2_nand2b_1 _09258_ (.Y(_01519_),
    .B(net366),
    .A_N(_01498_));
 sg13g2_buf_1 _09259_ (.A(_01519_),
    .X(_01520_));
 sg13g2_a21oi_1 _09260_ (.A1(_01515_),
    .A2(_01520_),
    .Y(_01521_),
    .B1(net365));
 sg13g2_nand3_1 _09261_ (.B(net306),
    .C(net366),
    .A(net365),
    .Y(_01522_));
 sg13g2_nand2b_1 _09262_ (.Y(_01523_),
    .B(_01522_),
    .A_N(_01521_));
 sg13g2_buf_1 _09263_ (.A(_01501_),
    .X(_01524_));
 sg13g2_a22oi_1 _09264_ (.Y(_01525_),
    .B1(_01523_),
    .B2(net304),
    .A2(_01518_),
    .A1(_01504_));
 sg13g2_inv_1 _09265_ (.Y(_00002_),
    .A(_01525_));
 sg13g2_nand2_1 _09266_ (.Y(_01526_),
    .A(_01501_),
    .B(net306));
 sg13g2_xnor2_1 _09267_ (.Y(_01527_),
    .A(net305),
    .B(_01496_));
 sg13g2_nand2_1 _09268_ (.Y(_01528_),
    .A(_01507_),
    .B(net366));
 sg13g2_nor2_1 _09269_ (.A(net365),
    .B(_01514_),
    .Y(_01529_));
 sg13g2_a21oi_1 _09270_ (.A1(net305),
    .A2(_01528_),
    .Y(_01530_),
    .B1(_01529_));
 sg13g2_nand2b_1 _09271_ (.Y(_01531_),
    .B(_01530_),
    .A_N(net258));
 sg13g2_o21ai_1 _09272_ (.B1(_01531_),
    .Y(_00003_),
    .A1(_01526_),
    .A2(_01527_));
 sg13g2_nor2_1 _09273_ (.A(net305),
    .B(net258),
    .Y(_01532_));
 sg13g2_nand2_1 _09274_ (.Y(_01533_),
    .A(net304),
    .B(net307));
 sg13g2_nor2_1 _09275_ (.A(net304),
    .B(_01511_),
    .Y(_01534_));
 sg13g2_a22oi_1 _09276_ (.Y(_01535_),
    .B1(_01520_),
    .B2(_01534_),
    .A2(_01508_),
    .A1(_01514_));
 sg13g2_o21ai_1 _09277_ (.B1(_01535_),
    .Y(_00004_),
    .A1(_01532_),
    .A2(_01533_));
 sg13g2_nand3_1 _09278_ (.B(_01515_),
    .C(_01520_),
    .A(net305),
    .Y(_01536_));
 sg13g2_o21ai_1 _09279_ (.B1(_01536_),
    .Y(_01537_),
    .A1(net304),
    .A2(_01510_));
 sg13g2_a21o_1 _09280_ (.A2(_01521_),
    .A1(net304),
    .B1(_01537_),
    .X(_00005_));
 sg13g2_nor2_1 _09281_ (.A(_01504_),
    .B(net307),
    .Y(_01538_));
 sg13g2_or2_1 _09282_ (.X(_01539_),
    .B(_01508_),
    .A(net366));
 sg13g2_a21oi_1 _09283_ (.A1(_01520_),
    .A2(_01539_),
    .Y(_01540_),
    .B1(net305));
 sg13g2_a221oi_1 _09284_ (.B2(net305),
    .C1(_01540_),
    .B1(_01538_),
    .A1(_01507_),
    .Y(_00006_),
    .A2(net307));
 sg13g2_nor2_1 _09285_ (.A(_01501_),
    .B(net365),
    .Y(_01541_));
 sg13g2_o21ai_1 _09286_ (.B1(_01509_),
    .Y(_00007_),
    .A1(_01515_),
    .A2(_01541_));
 sg13g2_nor2_1 _09287_ (.A(_01504_),
    .B(_01500_),
    .Y(_01542_));
 sg13g2_a21oi_1 _09288_ (.A1(_01500_),
    .A2(_01503_),
    .Y(_01543_),
    .B1(_01542_));
 sg13g2_nor2_1 _09289_ (.A(_01497_),
    .B(_01543_),
    .Y(_00008_));
 sg13g2_nand2_1 _09290_ (.Y(_01544_),
    .A(net365),
    .B(net306));
 sg13g2_xnor2_1 _09291_ (.Y(_01545_),
    .A(net304),
    .B(_01544_));
 sg13g2_nor2b_1 _09292_ (.A(_01539_),
    .B_N(_01541_),
    .Y(_01546_));
 sg13g2_a21o_1 _09293_ (.A2(_01545_),
    .A1(net307),
    .B1(_01546_),
    .X(_00009_));
 sg13g2_a21oi_1 _09294_ (.A1(net305),
    .A2(_01518_),
    .Y(_01547_),
    .B1(_01529_));
 sg13g2_nand3_1 _09295_ (.B(net258),
    .C(_01514_),
    .A(_01504_),
    .Y(_01548_));
 sg13g2_o21ai_1 _09296_ (.B1(_01548_),
    .Y(_00010_),
    .A1(_01507_),
    .A2(_01547_));
 sg13g2_nor2_1 _09297_ (.A(net304),
    .B(net258),
    .Y(_01549_));
 sg13g2_a21oi_1 _09298_ (.A1(net307),
    .A2(_01526_),
    .Y(_01550_),
    .B1(_01511_));
 sg13g2_nor3_1 _09299_ (.A(_01529_),
    .B(_01549_),
    .C(_01550_),
    .Y(_00011_));
 sg13g2_o21ai_1 _09300_ (.B1(_01513_),
    .Y(_01551_),
    .A1(_01507_),
    .A2(net258));
 sg13g2_a22oi_1 _09301_ (.Y(_01552_),
    .B1(_01508_),
    .B2(_01511_),
    .A2(net307),
    .A1(net258));
 sg13g2_nor2_1 _09302_ (.A(net304),
    .B(_01552_),
    .Y(_01553_));
 sg13g2_a21oi_1 _09303_ (.A1(net307),
    .A2(_01551_),
    .Y(_00012_),
    .B1(_01553_));
 sg13g2_nand2_1 _09304_ (.Y(_01554_),
    .A(_01507_),
    .B(net306));
 sg13g2_a21oi_1 _09305_ (.A1(_01511_),
    .A2(_01554_),
    .Y(_01555_),
    .B1(_01496_));
 sg13g2_a21o_1 _09306_ (.A2(_01529_),
    .A1(_01524_),
    .B1(_01555_),
    .X(_00013_));
 sg13g2_o21ai_1 _09307_ (.B1(_01520_),
    .Y(_01556_),
    .A1(_01511_),
    .A2(_01515_));
 sg13g2_a21oi_1 _09308_ (.A1(_01513_),
    .A2(_01554_),
    .Y(_01557_),
    .B1(_01514_));
 sg13g2_a221oi_1 _09309_ (.B2(_01524_),
    .C1(_01557_),
    .B1(_01556_),
    .A1(_01504_),
    .Y(_00014_),
    .A2(_01518_));
 sg13g2_buf_1 _09310_ (.A(_01442_),
    .X(_01558_));
 sg13g2_buf_1 _09311_ (.A(_01558_),
    .X(_01559_));
 sg13g2_buf_1 _09312_ (.A(net303),
    .X(_01560_));
 sg13g2_nand3_1 _09313_ (.B(_01452_),
    .C(_01453_),
    .A(_01451_),
    .Y(_01561_));
 sg13g2_buf_1 _09314_ (.A(_01561_),
    .X(_01562_));
 sg13g2_nor2_1 _09315_ (.A(_01449_),
    .B(_01562_),
    .Y(_01563_));
 sg13g2_buf_1 _09316_ (.A(_01563_),
    .X(_01564_));
 sg13g2_buf_1 _09317_ (.A(net138),
    .X(_01565_));
 sg13g2_buf_1 _09318_ (.A(net42),
    .X(_01566_));
 sg13g2_and3_1 _09319_ (.X(_00015_),
    .A(_01461_),
    .B(net257),
    .C(net33));
 sg13g2_and3_1 _09320_ (.X(_00016_),
    .A(net257),
    .B(\am_sdr0.am0.state[0] ),
    .C(\am_sdr0.am0.load_tick ));
 sg13g2_and3_1 _09321_ (.X(_00017_),
    .A(_01448_),
    .B(_01560_),
    .C(net33));
 sg13g2_buf_1 _09322_ (.A(\am_sdr0.am0.sum[1] ),
    .X(_01567_));
 sg13g2_buf_1 _09323_ (.A(\am_sdr0.am0.sqrt_state[0] ),
    .X(_01568_));
 sg13g2_inv_1 _09324_ (.Y(_01569_),
    .A(_01568_));
 sg13g2_buf_2 _09325_ (.A(\am_sdr0.am0.sqrt_state[1] ),
    .X(_01570_));
 sg13g2_nor3_1 _09326_ (.A(net310),
    .B(_01569_),
    .C(_01570_),
    .Y(_01571_));
 sg13g2_nand2_1 _09327_ (.Y(_01572_),
    .A(_01569_),
    .B(_01570_));
 sg13g2_buf_1 _09328_ (.A(_01572_),
    .X(_01573_));
 sg13g2_buf_1 _09329_ (.A(_01568_),
    .X(_01574_));
 sg13g2_nand2b_1 _09330_ (.Y(_01575_),
    .B(_01574_),
    .A_N(_01570_));
 sg13g2_a21oi_1 _09331_ (.A1(_01573_),
    .A2(_01575_),
    .Y(_01576_),
    .B1(net310));
 sg13g2_buf_1 _09332_ (.A(_01576_),
    .X(_00173_));
 sg13g2_buf_1 _09333_ (.A(\am_sdr0.am0.count[1] ),
    .X(_01577_));
 sg13g2_buf_1 _09334_ (.A(\am_sdr0.am0.count[0] ),
    .X(_01578_));
 sg13g2_nor2b_1 _09335_ (.A(_01568_),
    .B_N(_01570_),
    .Y(_01579_));
 sg13g2_buf_2 _09336_ (.A(_01579_),
    .X(_01580_));
 sg13g2_o21ai_1 _09337_ (.B1(_01580_),
    .Y(_01581_),
    .A1(_01577_),
    .A2(_01578_));
 sg13g2_nand2_1 _09338_ (.Y(_01582_),
    .A(net41),
    .B(_01581_));
 sg13g2_buf_1 _09339_ (.A(_01582_),
    .X(_01583_));
 sg13g2_a22oi_1 _09340_ (.Y(_01584_),
    .B1(_01583_),
    .B2(\am_sdr0.am0.a[0] ),
    .A2(_01571_),
    .A1(_01567_));
 sg13g2_inv_1 _09341_ (.Y(_00075_),
    .A(_01584_));
 sg13g2_and2_1 _09342_ (.A(net41),
    .B(_01581_),
    .X(_01585_));
 sg13g2_buf_1 _09343_ (.A(_01585_),
    .X(_01586_));
 sg13g2_buf_1 _09344_ (.A(_01586_),
    .X(_01587_));
 sg13g2_buf_1 _09345_ (.A(_01587_),
    .X(_01588_));
 sg13g2_buf_1 _09346_ (.A(_01580_),
    .X(_01589_));
 sg13g2_buf_1 _09347_ (.A(\am_sdr0.am0.sum[11] ),
    .X(_01590_));
 sg13g2_inv_1 _09348_ (.Y(_01591_),
    .A(_01590_));
 sg13g2_buf_1 _09349_ (.A(_01580_),
    .X(_01592_));
 sg13g2_nor2_1 _09350_ (.A(_01591_),
    .B(net188),
    .Y(_01593_));
 sg13g2_a21oi_1 _09351_ (.A1(\am_sdr0.am0.a[8] ),
    .A2(net189),
    .Y(_01594_),
    .B1(_01593_));
 sg13g2_buf_1 _09352_ (.A(_01586_),
    .X(_01595_));
 sg13g2_nor2_1 _09353_ (.A(\am_sdr0.am0.a[10] ),
    .B(net15),
    .Y(_01596_));
 sg13g2_a21oi_1 _09354_ (.A1(_01588_),
    .A2(_01594_),
    .Y(_00076_),
    .B1(_01596_));
 sg13g2_buf_1 _09355_ (.A(\am_sdr0.am0.sum[12] ),
    .X(_01597_));
 sg13g2_buf_1 _09356_ (.A(_01573_),
    .X(_01598_));
 sg13g2_buf_1 _09357_ (.A(_01580_),
    .X(_01599_));
 sg13g2_and2_1 _09358_ (.A(\am_sdr0.am0.a[9] ),
    .B(net187),
    .X(_01600_));
 sg13g2_a21oi_1 _09359_ (.A1(_01597_),
    .A2(net137),
    .Y(_01601_),
    .B1(_01600_));
 sg13g2_nor2_1 _09360_ (.A(\am_sdr0.am0.a[11] ),
    .B(net15),
    .Y(_01602_));
 sg13g2_a21oi_1 _09361_ (.A1(net9),
    .A2(_01601_),
    .Y(_00077_),
    .B1(_01602_));
 sg13g2_buf_1 _09362_ (.A(\am_sdr0.am0.sum[13] ),
    .X(_01603_));
 sg13g2_and2_1 _09363_ (.A(\am_sdr0.am0.a[10] ),
    .B(net187),
    .X(_01604_));
 sg13g2_a21oi_1 _09364_ (.A1(_01603_),
    .A2(net137),
    .Y(_01605_),
    .B1(_01604_));
 sg13g2_nor2_1 _09365_ (.A(\am_sdr0.am0.a[12] ),
    .B(net15),
    .Y(_01606_));
 sg13g2_a21oi_1 _09366_ (.A1(net9),
    .A2(_01605_),
    .Y(_00078_),
    .B1(_01606_));
 sg13g2_inv_1 _09367_ (.Y(_01607_),
    .A(\am_sdr0.am0.sum[14] ));
 sg13g2_nor2_1 _09368_ (.A(_01607_),
    .B(net188),
    .Y(_01608_));
 sg13g2_a21oi_1 _09369_ (.A1(\am_sdr0.am0.a[11] ),
    .A2(net189),
    .Y(_01609_),
    .B1(_01608_));
 sg13g2_nor2_1 _09370_ (.A(\am_sdr0.am0.a[13] ),
    .B(net15),
    .Y(_01610_));
 sg13g2_a21oi_1 _09371_ (.A1(net9),
    .A2(_01609_),
    .Y(_00079_),
    .B1(_01610_));
 sg13g2_buf_1 _09372_ (.A(\am_sdr0.am0.sum[15] ),
    .X(_01611_));
 sg13g2_and2_1 _09373_ (.A(\am_sdr0.am0.a[12] ),
    .B(net187),
    .X(_01612_));
 sg13g2_a21oi_1 _09374_ (.A1(_01611_),
    .A2(net137),
    .Y(_01613_),
    .B1(_01612_));
 sg13g2_nor2_1 _09375_ (.A(\am_sdr0.am0.a[14] ),
    .B(net15),
    .Y(_01614_));
 sg13g2_a21oi_1 _09376_ (.A1(net9),
    .A2(_01613_),
    .Y(_00080_),
    .B1(_01614_));
 sg13g2_and2_1 _09377_ (.A(\am_sdr0.am0.a[13] ),
    .B(net187),
    .X(_01615_));
 sg13g2_a21oi_1 _09378_ (.A1(\am_sdr0.am0.sum[16] ),
    .A2(net137),
    .Y(_01616_),
    .B1(_01615_));
 sg13g2_nor2_1 _09379_ (.A(\am_sdr0.am0.a[15] ),
    .B(net15),
    .Y(_01617_));
 sg13g2_a21oi_1 _09380_ (.A1(net9),
    .A2(_01616_),
    .Y(_00081_),
    .B1(_01617_));
 sg13g2_buf_1 _09381_ (.A(\am_sdr0.am0.sum[2] ),
    .X(_01618_));
 sg13g2_a22oi_1 _09382_ (.Y(_01619_),
    .B1(_01583_),
    .B2(\am_sdr0.am0.a[1] ),
    .A2(_01571_),
    .A1(_01618_));
 sg13g2_inv_1 _09383_ (.Y(_00082_),
    .A(_01619_));
 sg13g2_buf_1 _09384_ (.A(\am_sdr0.am0.sum[3] ),
    .X(_01620_));
 sg13g2_inv_1 _09385_ (.Y(_01621_),
    .A(_01620_));
 sg13g2_nor2_1 _09386_ (.A(_01621_),
    .B(net188),
    .Y(_01622_));
 sg13g2_a21oi_1 _09387_ (.A1(\am_sdr0.am0.a[0] ),
    .A2(net189),
    .Y(_01623_),
    .B1(_01622_));
 sg13g2_nor2_1 _09388_ (.A(\am_sdr0.am0.a[2] ),
    .B(net15),
    .Y(_01624_));
 sg13g2_a21oi_1 _09389_ (.A1(net9),
    .A2(_01623_),
    .Y(_00083_),
    .B1(_01624_));
 sg13g2_buf_2 _09390_ (.A(\am_sdr0.am0.sum[4] ),
    .X(_01625_));
 sg13g2_and2_1 _09391_ (.A(\am_sdr0.am0.a[1] ),
    .B(net187),
    .X(_01626_));
 sg13g2_a21oi_1 _09392_ (.A1(_01625_),
    .A2(net137),
    .Y(_01627_),
    .B1(_01626_));
 sg13g2_nor2_1 _09393_ (.A(\am_sdr0.am0.a[3] ),
    .B(net15),
    .Y(_01628_));
 sg13g2_a21oi_1 _09394_ (.A1(_01588_),
    .A2(_01627_),
    .Y(_00084_),
    .B1(_01628_));
 sg13g2_buf_2 _09395_ (.A(\am_sdr0.am0.sum[5] ),
    .X(_01629_));
 sg13g2_and2_1 _09396_ (.A(\am_sdr0.am0.a[2] ),
    .B(_01599_),
    .X(_01630_));
 sg13g2_a21oi_1 _09397_ (.A1(_01629_),
    .A2(net137),
    .Y(_01631_),
    .B1(_01630_));
 sg13g2_nor2_1 _09398_ (.A(\am_sdr0.am0.a[4] ),
    .B(_01595_),
    .Y(_01632_));
 sg13g2_a21oi_1 _09399_ (.A1(net9),
    .A2(_01631_),
    .Y(_00085_),
    .B1(_01632_));
 sg13g2_buf_1 _09400_ (.A(\am_sdr0.am0.sum[6] ),
    .X(_01633_));
 sg13g2_and2_1 _09401_ (.A(\am_sdr0.am0.a[3] ),
    .B(net187),
    .X(_01634_));
 sg13g2_a21oi_1 _09402_ (.A1(_01633_),
    .A2(_01598_),
    .Y(_01635_),
    .B1(_01634_));
 sg13g2_nor2_1 _09403_ (.A(\am_sdr0.am0.a[5] ),
    .B(_01595_),
    .Y(_01636_));
 sg13g2_a21oi_1 _09404_ (.A1(net9),
    .A2(_01635_),
    .Y(_00086_),
    .B1(_01636_));
 sg13g2_buf_1 _09405_ (.A(net16),
    .X(_01637_));
 sg13g2_inv_1 _09406_ (.Y(_01638_),
    .A(\am_sdr0.am0.sum[7] ));
 sg13g2_nor2_1 _09407_ (.A(_01638_),
    .B(_01592_),
    .Y(_01639_));
 sg13g2_a21oi_1 _09408_ (.A1(\am_sdr0.am0.a[4] ),
    .A2(net189),
    .Y(_01640_),
    .B1(_01639_));
 sg13g2_buf_1 _09409_ (.A(_01586_),
    .X(_01641_));
 sg13g2_nor2_1 _09410_ (.A(\am_sdr0.am0.a[6] ),
    .B(net14),
    .Y(_01642_));
 sg13g2_a21oi_1 _09411_ (.A1(_01637_),
    .A2(_01640_),
    .Y(_00087_),
    .B1(_01642_));
 sg13g2_buf_1 _09412_ (.A(\am_sdr0.am0.sum[8] ),
    .X(_01643_));
 sg13g2_inv_1 _09413_ (.Y(_01644_),
    .A(_01643_));
 sg13g2_nor2_1 _09414_ (.A(_01644_),
    .B(_01592_),
    .Y(_01645_));
 sg13g2_a21oi_1 _09415_ (.A1(\am_sdr0.am0.a[5] ),
    .A2(_01589_),
    .Y(_01646_),
    .B1(_01645_));
 sg13g2_nor2_1 _09416_ (.A(\am_sdr0.am0.a[7] ),
    .B(net14),
    .Y(_01647_));
 sg13g2_a21oi_1 _09417_ (.A1(net8),
    .A2(_01646_),
    .Y(_00088_),
    .B1(_01647_));
 sg13g2_buf_2 _09418_ (.A(\am_sdr0.am0.sum[9] ),
    .X(_01648_));
 sg13g2_and2_1 _09419_ (.A(\am_sdr0.am0.a[6] ),
    .B(net187),
    .X(_01649_));
 sg13g2_a21oi_1 _09420_ (.A1(_01648_),
    .A2(_01598_),
    .Y(_01650_),
    .B1(_01649_));
 sg13g2_nor2_1 _09421_ (.A(\am_sdr0.am0.a[8] ),
    .B(_01641_),
    .Y(_01651_));
 sg13g2_a21oi_1 _09422_ (.A1(net8),
    .A2(_01650_),
    .Y(_00089_),
    .B1(_01651_));
 sg13g2_buf_1 _09423_ (.A(\am_sdr0.am0.sum[10] ),
    .X(_01652_));
 sg13g2_inv_1 _09424_ (.Y(_01653_),
    .A(_01652_));
 sg13g2_nor2_1 _09425_ (.A(_01653_),
    .B(net187),
    .Y(_01654_));
 sg13g2_a21oi_1 _09426_ (.A1(\am_sdr0.am0.a[7] ),
    .A2(_01589_),
    .Y(_01655_),
    .B1(_01654_));
 sg13g2_nor2_1 _09427_ (.A(\am_sdr0.am0.a[9] ),
    .B(_01641_),
    .Y(_01656_));
 sg13g2_a21oi_1 _09428_ (.A1(net8),
    .A2(_01655_),
    .Y(_00090_),
    .B1(_01656_));
 sg13g2_buf_1 _09429_ (.A(\am_sdr0.am0.count2[0] ),
    .X(_01657_));
 sg13g2_inv_1 _09430_ (.Y(_01658_),
    .A(_01577_));
 sg13g2_nor2_1 _09431_ (.A(_01658_),
    .B(_01578_),
    .Y(_01659_));
 sg13g2_o21ai_1 _09432_ (.B1(net41),
    .Y(_01660_),
    .A1(_01573_),
    .A2(_01659_));
 sg13g2_buf_1 _09433_ (.A(_01660_),
    .X(_01661_));
 sg13g2_buf_1 _09434_ (.A(_01661_),
    .X(_01662_));
 sg13g2_nand2_1 _09435_ (.Y(_01663_),
    .A(net364),
    .B(_01569_));
 sg13g2_nand2_1 _09436_ (.Y(_01664_),
    .A(_01570_),
    .B(_01659_));
 sg13g2_nor2_2 _09437_ (.A(_01663_),
    .B(_01664_),
    .Y(_01665_));
 sg13g2_a22oi_1 _09438_ (.Y(_01666_),
    .B1(_01665_),
    .B2(_00070_),
    .A2(net13),
    .A1(_01657_));
 sg13g2_inv_1 _09439_ (.Y(_00091_),
    .A(_01666_));
 sg13g2_buf_1 _09440_ (.A(_01661_),
    .X(_01667_));
 sg13g2_buf_1 _09441_ (.A(\am_sdr0.am0.count2[1] ),
    .X(_01668_));
 sg13g2_nand3b_1 _09442_ (.B(_01657_),
    .C(net188),
    .Y(_01669_),
    .A_N(_01668_));
 sg13g2_nor2_1 _09443_ (.A(_01657_),
    .B(net137),
    .Y(_01670_));
 sg13g2_o21ai_1 _09444_ (.B1(_01668_),
    .Y(_01671_),
    .A1(net13),
    .A2(_01670_));
 sg13g2_o21ai_1 _09445_ (.B1(_01671_),
    .Y(_00092_),
    .A1(net12),
    .A2(_01669_));
 sg13g2_nand3_1 _09446_ (.B(_01657_),
    .C(_01665_),
    .A(_01668_),
    .Y(_01672_));
 sg13g2_a21oi_1 _09447_ (.A1(_01668_),
    .A2(_01657_),
    .Y(_01673_),
    .B1(net137));
 sg13g2_o21ai_1 _09448_ (.B1(\am_sdr0.am0.count2[2] ),
    .Y(_01674_),
    .A1(net13),
    .A2(_01673_));
 sg13g2_o21ai_1 _09449_ (.B1(_01674_),
    .Y(_00093_),
    .A1(\am_sdr0.am0.count2[2] ),
    .A2(_01672_));
 sg13g2_inv_1 _09450_ (.Y(_01675_),
    .A(\am_sdr0.am0.count2[3] ));
 sg13g2_nand3_1 _09451_ (.B(_01657_),
    .C(\am_sdr0.am0.count2[2] ),
    .A(_01668_),
    .Y(_01676_));
 sg13g2_a21oi_1 _09452_ (.A1(_01665_),
    .A2(_01676_),
    .Y(_01677_),
    .B1(net13));
 sg13g2_nand2b_1 _09453_ (.Y(_01678_),
    .B(_01675_),
    .A_N(_01676_));
 sg13g2_or3_1 _09454_ (.A(_01663_),
    .B(_01664_),
    .C(_01678_),
    .X(_01679_));
 sg13g2_o21ai_1 _09455_ (.B1(_01679_),
    .Y(_00094_),
    .A1(_01675_),
    .A2(_01677_));
 sg13g2_inv_1 _09456_ (.Y(_01680_),
    .A(_01578_));
 sg13g2_nor2_1 _09457_ (.A(_01577_),
    .B(_01573_),
    .Y(_01681_));
 sg13g2_nand3_1 _09458_ (.B(net41),
    .C(_01681_),
    .A(_00069_),
    .Y(_01682_));
 sg13g2_o21ai_1 _09459_ (.B1(_01682_),
    .Y(_00095_),
    .A1(_01680_),
    .A2(net41));
 sg13g2_nand3_1 _09460_ (.B(net41),
    .C(_01681_),
    .A(_01578_),
    .Y(_01683_));
 sg13g2_buf_1 _09461_ (.A(_01683_),
    .X(_01684_));
 sg13g2_o21ai_1 _09462_ (.B1(net24),
    .Y(_00096_),
    .A1(_01658_),
    .A2(net41));
 sg13g2_buf_1 _09463_ (.A(\am_sdr0.am0.left[0] ),
    .X(_01685_));
 sg13g2_inv_1 _09464_ (.Y(_01686_),
    .A(_01685_));
 sg13g2_buf_1 _09465_ (.A(_01599_),
    .X(_01687_));
 sg13g2_nand3_1 _09466_ (.B(net136),
    .C(net14),
    .A(\am_sdr0.am0.a[14] ),
    .Y(_01688_));
 sg13g2_o21ai_1 _09467_ (.B1(_01688_),
    .Y(_00105_),
    .A1(_01686_),
    .A2(net8));
 sg13g2_buf_1 _09468_ (.A(\am_sdr0.am0.left[1] ),
    .X(_01689_));
 sg13g2_inv_1 _09469_ (.Y(_01690_),
    .A(_01689_));
 sg13g2_nand3_1 _09470_ (.B(net136),
    .C(net14),
    .A(\am_sdr0.am0.a[15] ),
    .Y(_01691_));
 sg13g2_o21ai_1 _09471_ (.B1(_01691_),
    .Y(_00106_),
    .A1(_01690_),
    .A2(net8));
 sg13g2_inv_1 _09472_ (.Y(_01692_),
    .A(\am_sdr0.am0.left[2] ));
 sg13g2_nand3_1 _09473_ (.B(net136),
    .C(net14),
    .A(\am_sdr0.am0.r[0] ),
    .Y(_01693_));
 sg13g2_o21ai_1 _09474_ (.B1(_01693_),
    .Y(_00107_),
    .A1(_01692_),
    .A2(net8));
 sg13g2_inv_1 _09475_ (.Y(_01694_),
    .A(\am_sdr0.am0.left[3] ));
 sg13g2_nand3_1 _09476_ (.B(net136),
    .C(net14),
    .A(\am_sdr0.am0.r[1] ),
    .Y(_01695_));
 sg13g2_o21ai_1 _09477_ (.B1(_01695_),
    .Y(_00108_),
    .A1(_01694_),
    .A2(net8));
 sg13g2_inv_1 _09478_ (.Y(_01696_),
    .A(\am_sdr0.am0.left[4] ));
 sg13g2_nand3_1 _09479_ (.B(net136),
    .C(net14),
    .A(\am_sdr0.am0.r[2] ),
    .Y(_01697_));
 sg13g2_o21ai_1 _09480_ (.B1(_01697_),
    .Y(_00109_),
    .A1(_01696_),
    .A2(net8));
 sg13g2_inv_1 _09481_ (.Y(_01698_),
    .A(\am_sdr0.am0.left[5] ));
 sg13g2_nand3_1 _09482_ (.B(net136),
    .C(_01587_),
    .A(\am_sdr0.am0.r[3] ),
    .Y(_01699_));
 sg13g2_o21ai_1 _09483_ (.B1(_01699_),
    .Y(_00110_),
    .A1(_01698_),
    .A2(_01637_));
 sg13g2_inv_1 _09484_ (.Y(_01700_),
    .A(\am_sdr0.am0.left[6] ));
 sg13g2_buf_1 _09485_ (.A(net16),
    .X(_01701_));
 sg13g2_nand3_1 _09486_ (.B(_01687_),
    .C(net16),
    .A(\am_sdr0.am0.r[4] ),
    .Y(_01702_));
 sg13g2_o21ai_1 _09487_ (.B1(_01702_),
    .Y(_00111_),
    .A1(_01700_),
    .A2(_01701_));
 sg13g2_inv_1 _09488_ (.Y(_01703_),
    .A(\am_sdr0.am0.left[7] ));
 sg13g2_nand3_1 _09489_ (.B(net136),
    .C(net16),
    .A(\am_sdr0.am0.r[5] ),
    .Y(_01704_));
 sg13g2_o21ai_1 _09490_ (.B1(_01704_),
    .Y(_00112_),
    .A1(_01703_),
    .A2(net7));
 sg13g2_inv_1 _09491_ (.Y(_01705_),
    .A(\am_sdr0.am0.left[8] ));
 sg13g2_nand3_1 _09492_ (.B(net189),
    .C(net16),
    .A(\am_sdr0.am0.r[6] ),
    .Y(_01706_));
 sg13g2_o21ai_1 _09493_ (.B1(_01706_),
    .Y(_00113_),
    .A1(_01705_),
    .A2(_01701_));
 sg13g2_inv_1 _09494_ (.Y(_01707_),
    .A(\am_sdr0.am0.left[9] ));
 sg13g2_nand3_1 _09495_ (.B(net189),
    .C(net16),
    .A(\am_sdr0.am0.r[7] ),
    .Y(_01708_));
 sg13g2_o21ai_1 _09496_ (.B1(_01708_),
    .Y(_00114_),
    .A1(_01707_),
    .A2(net7));
 sg13g2_or2_1 _09497_ (.X(_01709_),
    .B(_01461_),
    .A(_01448_));
 sg13g2_buf_1 _09498_ (.A(_01709_),
    .X(_01710_));
 sg13g2_or2_1 _09499_ (.X(_01711_),
    .B(net367),
    .A(\am_sdr0.am0.state[4] ));
 sg13g2_o21ai_1 _09500_ (.B1(_01442_),
    .Y(_01712_),
    .A1(net256),
    .A2(_01711_));
 sg13g2_buf_1 _09501_ (.A(_01712_),
    .X(_01713_));
 sg13g2_buf_1 _09502_ (.A(_01713_),
    .X(_01714_));
 sg13g2_nand2_1 _09503_ (.Y(_01715_),
    .A(_01452_),
    .B(net40));
 sg13g2_buf_1 _09504_ (.A(net256),
    .X(_01716_));
 sg13g2_nand3_1 _09505_ (.B(_00071_),
    .C(net186),
    .A(_01560_),
    .Y(_01717_));
 sg13g2_nand2_1 _09506_ (.Y(_00115_),
    .A(_01715_),
    .B(_01717_));
 sg13g2_buf_1 _09507_ (.A(net364),
    .X(_01718_));
 sg13g2_buf_1 _09508_ (.A(net256),
    .X(_01719_));
 sg13g2_nand3_1 _09509_ (.B(_01452_),
    .C(net185),
    .A(net301),
    .Y(_01720_));
 sg13g2_buf_1 _09510_ (.A(_01713_),
    .X(_01721_));
 sg13g2_nor2_1 _09511_ (.A(_01448_),
    .B(_01461_),
    .Y(_01722_));
 sg13g2_buf_1 _09512_ (.A(_01722_),
    .X(_01723_));
 sg13g2_nor2_1 _09513_ (.A(_01452_),
    .B(net255),
    .Y(_01724_));
 sg13g2_o21ai_1 _09514_ (.B1(_01451_),
    .Y(_01725_),
    .A1(_01721_),
    .A2(_01724_));
 sg13g2_o21ai_1 _09515_ (.B1(_01725_),
    .Y(_00116_),
    .A1(_01451_),
    .A2(_01720_));
 sg13g2_nand4_1 _09516_ (.B(_01451_),
    .C(_01452_),
    .A(_01718_),
    .Y(_01726_),
    .D(net256));
 sg13g2_a21oi_1 _09517_ (.A1(_01451_),
    .A2(_01452_),
    .Y(_01727_),
    .B1(net255));
 sg13g2_o21ai_1 _09518_ (.B1(_01453_),
    .Y(_01728_),
    .A1(net39),
    .A2(_01727_));
 sg13g2_o21ai_1 _09519_ (.B1(_01728_),
    .Y(_00117_),
    .A1(_01453_),
    .A2(_01726_));
 sg13g2_buf_1 _09520_ (.A(_01713_),
    .X(_01729_));
 sg13g2_nand2_1 _09521_ (.Y(_01730_),
    .A(_01449_),
    .B(_01562_));
 sg13g2_o21ai_1 _09522_ (.B1(_01730_),
    .Y(_01731_),
    .A1(net190),
    .A2(_01713_));
 sg13g2_a22oi_1 _09523_ (.Y(_01732_),
    .B1(_01731_),
    .B2(_01716_),
    .A2(net38),
    .A1(_01449_));
 sg13g2_inv_1 _09524_ (.Y(_00118_),
    .A(_01732_));
 sg13g2_buf_1 _09525_ (.A(_01713_),
    .X(_01733_));
 sg13g2_nor2b_1 _09526_ (.A(net367),
    .B_N(\am_sdr0.am0.I_in[0] ),
    .Y(_01734_));
 sg13g2_a22oi_1 _09527_ (.Y(_01735_),
    .B1(net255),
    .B2(_01734_),
    .A2(\am_sdr0.am0.Q_in[0] ),
    .A1(net309));
 sg13g2_buf_8 _09528_ (.A(\am_sdr0.am0.multA[0] ),
    .X(_01736_));
 sg13g2_nand2_1 _09529_ (.Y(_01737_),
    .A(_01736_),
    .B(net40));
 sg13g2_o21ai_1 _09530_ (.B1(_01737_),
    .Y(_00119_),
    .A1(net37),
    .A2(_01735_));
 sg13g2_nor2b_1 _09531_ (.A(net367),
    .B_N(\am_sdr0.am0.I_in[7] ),
    .Y(_01738_));
 sg13g2_a22oi_1 _09532_ (.Y(_01739_),
    .B1(_01722_),
    .B2(_01738_),
    .A2(\am_sdr0.am0.Q_in[7] ),
    .A1(net367));
 sg13g2_or2_1 _09533_ (.X(_01740_),
    .B(_01739_),
    .A(_01713_));
 sg13g2_buf_1 _09534_ (.A(_01740_),
    .X(_01741_));
 sg13g2_buf_1 _09535_ (.A(_01741_),
    .X(_01742_));
 sg13g2_buf_1 _09536_ (.A(net303),
    .X(_01743_));
 sg13g2_buf_1 _09537_ (.A(\am_sdr0.am0.multA[9] ),
    .X(_01744_));
 sg13g2_nand3_1 _09538_ (.B(_01744_),
    .C(net186),
    .A(net254),
    .Y(_01745_));
 sg13g2_buf_1 _09539_ (.A(\am_sdr0.am0.multA[10] ),
    .X(_01746_));
 sg13g2_nand2_1 _09540_ (.Y(_01747_),
    .A(_01746_),
    .B(net38));
 sg13g2_nand3_1 _09541_ (.B(_01745_),
    .C(_01747_),
    .A(net23),
    .Y(_00120_));
 sg13g2_nand3_1 _09542_ (.B(_01746_),
    .C(net186),
    .A(net254),
    .Y(_01748_));
 sg13g2_buf_1 _09543_ (.A(\am_sdr0.am0.multA[11] ),
    .X(_01749_));
 sg13g2_nand2_1 _09544_ (.Y(_01750_),
    .A(_01749_),
    .B(net38));
 sg13g2_nand3_1 _09545_ (.B(_01748_),
    .C(_01750_),
    .A(net23),
    .Y(_00121_));
 sg13g2_nand3_1 _09546_ (.B(_01749_),
    .C(net186),
    .A(net254),
    .Y(_01751_));
 sg13g2_buf_1 _09547_ (.A(\am_sdr0.am0.multA[12] ),
    .X(_01752_));
 sg13g2_nand2_1 _09548_ (.Y(_01753_),
    .A(_01752_),
    .B(net39));
 sg13g2_nand3_1 _09549_ (.B(_01751_),
    .C(_01753_),
    .A(_01742_),
    .Y(_00122_));
 sg13g2_nand3_1 _09550_ (.B(_01752_),
    .C(net186),
    .A(net254),
    .Y(_01754_));
 sg13g2_buf_1 _09551_ (.A(\am_sdr0.am0.multA[13] ),
    .X(_01755_));
 sg13g2_nand2_1 _09552_ (.Y(_01756_),
    .A(_01755_),
    .B(net39));
 sg13g2_nand3_1 _09553_ (.B(_01754_),
    .C(_01756_),
    .A(net23),
    .Y(_00123_));
 sg13g2_nand3_1 _09554_ (.B(_01755_),
    .C(net186),
    .A(net254),
    .Y(_01757_));
 sg13g2_buf_1 _09555_ (.A(\am_sdr0.am0.multA[14] ),
    .X(_01758_));
 sg13g2_nand2_1 _09556_ (.Y(_01759_),
    .A(_01758_),
    .B(net39));
 sg13g2_nand3_1 _09557_ (.B(_01757_),
    .C(_01759_),
    .A(net23),
    .Y(_00124_));
 sg13g2_buf_1 _09558_ (.A(net303),
    .X(_01760_));
 sg13g2_nand3_1 _09559_ (.B(_01758_),
    .C(net186),
    .A(net253),
    .Y(_01761_));
 sg13g2_buf_1 _09560_ (.A(\am_sdr0.am0.multA[15] ),
    .X(_01762_));
 sg13g2_nand2_1 _09561_ (.Y(_01763_),
    .A(_01762_),
    .B(net39));
 sg13g2_nand3_1 _09562_ (.B(_01761_),
    .C(_01763_),
    .A(net23),
    .Y(_00125_));
 sg13g2_nand3_1 _09563_ (.B(_01762_),
    .C(net185),
    .A(net253),
    .Y(_01764_));
 sg13g2_nand2_1 _09564_ (.Y(_01765_),
    .A(\am_sdr0.am0.multA[16] ),
    .B(net39));
 sg13g2_nand3_1 _09565_ (.B(_01764_),
    .C(_01765_),
    .A(net23),
    .Y(_00126_));
 sg13g2_nand2_1 _09566_ (.Y(_01766_),
    .A(\am_sdr0.am0.I_in[1] ),
    .B(net255));
 sg13g2_nand2_1 _09567_ (.Y(_01767_),
    .A(net309),
    .B(\am_sdr0.am0.Q_in[1] ));
 sg13g2_o21ai_1 _09568_ (.B1(_01767_),
    .Y(_01768_),
    .A1(net309),
    .A2(_01766_));
 sg13g2_a21oi_1 _09569_ (.A1(net363),
    .A2(net185),
    .Y(_01769_),
    .B1(_01768_));
 sg13g2_buf_8 _09570_ (.A(\am_sdr0.am0.multA[1] ),
    .X(_01770_));
 sg13g2_nand2_1 _09571_ (.Y(_01771_),
    .A(_01770_),
    .B(net40));
 sg13g2_o21ai_1 _09572_ (.B1(_01771_),
    .Y(_00127_),
    .A1(net37),
    .A2(_01769_));
 sg13g2_nand2_1 _09573_ (.Y(_01772_),
    .A(\am_sdr0.am0.I_in[2] ),
    .B(net255));
 sg13g2_nand2_1 _09574_ (.Y(_01773_),
    .A(net367),
    .B(\am_sdr0.am0.Q_in[2] ));
 sg13g2_o21ai_1 _09575_ (.B1(_01773_),
    .Y(_01774_),
    .A1(net309),
    .A2(_01772_));
 sg13g2_a21oi_1 _09576_ (.A1(_01770_),
    .A2(net185),
    .Y(_01775_),
    .B1(_01774_));
 sg13g2_buf_8 _09577_ (.A(\am_sdr0.am0.multA[2] ),
    .X(_01776_));
 sg13g2_nand2_1 _09578_ (.Y(_01777_),
    .A(_01776_),
    .B(net40));
 sg13g2_o21ai_1 _09579_ (.B1(_01777_),
    .Y(_00128_),
    .A1(net37),
    .A2(_01775_));
 sg13g2_nand2_1 _09580_ (.Y(_01778_),
    .A(\am_sdr0.am0.I_in[3] ),
    .B(net255));
 sg13g2_nand2_1 _09581_ (.Y(_01779_),
    .A(net367),
    .B(\am_sdr0.am0.Q_in[3] ));
 sg13g2_o21ai_1 _09582_ (.B1(_01779_),
    .Y(_01780_),
    .A1(net309),
    .A2(_01778_));
 sg13g2_a21oi_1 _09583_ (.A1(_01776_),
    .A2(net185),
    .Y(_01781_),
    .B1(_01780_));
 sg13g2_buf_2 _09584_ (.A(\am_sdr0.am0.multA[3] ),
    .X(_01782_));
 sg13g2_nand2_1 _09585_ (.Y(_01783_),
    .A(_01782_),
    .B(net40));
 sg13g2_o21ai_1 _09586_ (.B1(_01783_),
    .Y(_00129_),
    .A1(net37),
    .A2(_01781_));
 sg13g2_nand2_1 _09587_ (.Y(_01784_),
    .A(\am_sdr0.am0.I_in[4] ),
    .B(_01723_));
 sg13g2_nand2_1 _09588_ (.Y(_01785_),
    .A(net367),
    .B(\am_sdr0.am0.Q_in[4] ));
 sg13g2_o21ai_1 _09589_ (.B1(_01785_),
    .Y(_01786_),
    .A1(net309),
    .A2(_01784_));
 sg13g2_a21oi_1 _09590_ (.A1(_01782_),
    .A2(_01719_),
    .Y(_01787_),
    .B1(_01786_));
 sg13g2_buf_2 _09591_ (.A(\am_sdr0.am0.multA[4] ),
    .X(_01788_));
 sg13g2_nand2_1 _09592_ (.Y(_01789_),
    .A(_01788_),
    .B(net38));
 sg13g2_o21ai_1 _09593_ (.B1(_01789_),
    .Y(_00130_),
    .A1(net37),
    .A2(_01787_));
 sg13g2_inv_1 _09594_ (.Y(_01790_),
    .A(\am_sdr0.am0.multA[5] ));
 sg13g2_nor2b_1 _09595_ (.A(net309),
    .B_N(\am_sdr0.am0.I_in[5] ),
    .Y(_01791_));
 sg13g2_a221oi_1 _09596_ (.B2(_01791_),
    .C1(_01713_),
    .B1(net255),
    .A1(_01463_),
    .Y(_01792_),
    .A2(\am_sdr0.am0.Q_in[5] ));
 sg13g2_nand2_1 _09597_ (.Y(_01793_),
    .A(_01788_),
    .B(_01716_));
 sg13g2_a22oi_1 _09598_ (.Y(_00131_),
    .B1(_01792_),
    .B2(_01793_),
    .A2(net37),
    .A1(_01790_));
 sg13g2_nand2_1 _09599_ (.Y(_01794_),
    .A(\am_sdr0.am0.I_in[6] ),
    .B(_01723_));
 sg13g2_nand2_1 _09600_ (.Y(_01795_),
    .A(_01462_),
    .B(\am_sdr0.am0.Q_in[6] ));
 sg13g2_o21ai_1 _09601_ (.B1(_01795_),
    .Y(_01796_),
    .A1(net309),
    .A2(_01794_));
 sg13g2_a21oi_1 _09602_ (.A1(\am_sdr0.am0.multA[5] ),
    .A2(_01719_),
    .Y(_01797_),
    .B1(_01796_));
 sg13g2_buf_2 _09603_ (.A(\am_sdr0.am0.multA[6] ),
    .X(_01798_));
 sg13g2_nand2_1 _09604_ (.Y(_01799_),
    .A(_01798_),
    .B(net38));
 sg13g2_o21ai_1 _09605_ (.B1(_01799_),
    .Y(_00132_),
    .A1(net37),
    .A2(_01797_));
 sg13g2_nand3_1 _09606_ (.B(_01798_),
    .C(net185),
    .A(net253),
    .Y(_01800_));
 sg13g2_buf_1 _09607_ (.A(\am_sdr0.am0.multA[7] ),
    .X(_01801_));
 sg13g2_nand2_1 _09608_ (.Y(_01802_),
    .A(_01801_),
    .B(net39));
 sg13g2_nand3_1 _09609_ (.B(_01800_),
    .C(_01802_),
    .A(net23),
    .Y(_00133_));
 sg13g2_nand3_1 _09610_ (.B(_01801_),
    .C(net185),
    .A(_01760_),
    .Y(_01803_));
 sg13g2_buf_1 _09611_ (.A(\am_sdr0.am0.multA[8] ),
    .X(_01804_));
 sg13g2_nand2_1 _09612_ (.Y(_01805_),
    .A(_01804_),
    .B(net39));
 sg13g2_nand3_1 _09613_ (.B(_01803_),
    .C(_01805_),
    .A(net23),
    .Y(_00134_));
 sg13g2_nand3_1 _09614_ (.B(_01804_),
    .C(net185),
    .A(_01760_),
    .Y(_01806_));
 sg13g2_nand2_1 _09615_ (.Y(_01807_),
    .A(_01744_),
    .B(_01721_));
 sg13g2_nand3_1 _09616_ (.B(_01806_),
    .C(_01807_),
    .A(_01741_),
    .Y(_00135_));
 sg13g2_inv_1 _09617_ (.Y(_01808_),
    .A(\am_sdr0.am0.multB[1] ));
 sg13g2_o21ai_1 _09618_ (.B1(_01735_),
    .Y(_01809_),
    .A1(_01808_),
    .A2(net255));
 sg13g2_mux2_1 _09619_ (.A0(_01809_),
    .A1(\am_sdr0.am0.multB[0] ),
    .S(net40),
    .X(_00136_));
 sg13g2_a21oi_1 _09620_ (.A1(\am_sdr0.am0.multB[2] ),
    .A2(net256),
    .Y(_01810_),
    .B1(_01768_));
 sg13g2_nand2_1 _09621_ (.Y(_01811_),
    .A(\am_sdr0.am0.multB[1] ),
    .B(net38));
 sg13g2_o21ai_1 _09622_ (.B1(_01811_),
    .Y(_00137_),
    .A1(_01733_),
    .A2(_01810_));
 sg13g2_a21oi_1 _09623_ (.A1(\am_sdr0.am0.multB[3] ),
    .A2(net256),
    .Y(_01812_),
    .B1(_01774_));
 sg13g2_nand2_1 _09624_ (.Y(_01813_),
    .A(\am_sdr0.am0.multB[2] ),
    .B(net38));
 sg13g2_o21ai_1 _09625_ (.B1(_01813_),
    .Y(_00138_),
    .A1(_01733_),
    .A2(_01812_));
 sg13g2_a21oi_1 _09626_ (.A1(\am_sdr0.am0.multB[4] ),
    .A2(net256),
    .Y(_01814_),
    .B1(_01780_));
 sg13g2_nand2_1 _09627_ (.Y(_01815_),
    .A(\am_sdr0.am0.multB[3] ),
    .B(net38));
 sg13g2_o21ai_1 _09628_ (.B1(_01815_),
    .Y(_00139_),
    .A1(net40),
    .A2(_01814_));
 sg13g2_a21oi_1 _09629_ (.A1(\am_sdr0.am0.multB[5] ),
    .A2(_01710_),
    .Y(_01816_),
    .B1(_01786_));
 sg13g2_nand2_1 _09630_ (.Y(_01817_),
    .A(\am_sdr0.am0.multB[4] ),
    .B(_01729_));
 sg13g2_o21ai_1 _09631_ (.B1(_01817_),
    .Y(_00140_),
    .A1(_01714_),
    .A2(_01816_));
 sg13g2_inv_1 _09632_ (.Y(_01818_),
    .A(\am_sdr0.am0.multB[5] ));
 sg13g2_nand2_1 _09633_ (.Y(_01819_),
    .A(\am_sdr0.am0.multB[6] ),
    .B(net186));
 sg13g2_a22oi_1 _09634_ (.Y(_00141_),
    .B1(_01792_),
    .B2(_01819_),
    .A2(net37),
    .A1(_01818_));
 sg13g2_a21oi_1 _09635_ (.A1(\am_sdr0.am0.multB[7] ),
    .A2(_01710_),
    .Y(_01820_),
    .B1(_01796_));
 sg13g2_nand2_1 _09636_ (.Y(_01821_),
    .A(\am_sdr0.am0.multB[6] ),
    .B(_01729_));
 sg13g2_o21ai_1 _09637_ (.B1(_01821_),
    .Y(_00142_),
    .A1(_01714_),
    .A2(_01820_));
 sg13g2_nand2_1 _09638_ (.Y(_01822_),
    .A(\am_sdr0.am0.multB[7] ),
    .B(net40));
 sg13g2_nand2_1 _09639_ (.Y(_00143_),
    .A(_01742_),
    .B(_01822_));
 sg13g2_a22oi_1 _09640_ (.Y(_01823_),
    .B1(_01665_),
    .B2(_00022_),
    .A2(net13),
    .A1(\am_sdr0.am0.q[0] ));
 sg13g2_inv_1 _09641_ (.Y(_00144_),
    .A(_01823_));
 sg13g2_nand2_1 _09642_ (.Y(_01824_),
    .A(\am_sdr0.am0.q[0] ),
    .B(_01580_));
 sg13g2_nand2_1 _09643_ (.Y(_01825_),
    .A(\am_sdr0.am0.q[1] ),
    .B(net12));
 sg13g2_o21ai_1 _09644_ (.B1(_01825_),
    .Y(_00145_),
    .A1(net12),
    .A2(_01824_));
 sg13g2_nand2_1 _09645_ (.Y(_01826_),
    .A(\am_sdr0.am0.q[1] ),
    .B(_01580_));
 sg13g2_nand2_1 _09646_ (.Y(_01827_),
    .A(\am_sdr0.am0.q[2] ),
    .B(net12));
 sg13g2_o21ai_1 _09647_ (.B1(_01827_),
    .Y(_00146_),
    .A1(net12),
    .A2(_01826_));
 sg13g2_nand2_1 _09648_ (.Y(_01828_),
    .A(\am_sdr0.am0.q[2] ),
    .B(net188));
 sg13g2_nand2_1 _09649_ (.Y(_01829_),
    .A(\am_sdr0.am0.q[3] ),
    .B(net13));
 sg13g2_o21ai_1 _09650_ (.B1(_01829_),
    .Y(_00147_),
    .A1(_01667_),
    .A2(_01828_));
 sg13g2_nand2_1 _09651_ (.Y(_01830_),
    .A(\am_sdr0.am0.q[3] ),
    .B(net188));
 sg13g2_nand2_1 _09652_ (.Y(_01831_),
    .A(\am_sdr0.am0.q[4] ),
    .B(net13));
 sg13g2_o21ai_1 _09653_ (.B1(_01831_),
    .Y(_00148_),
    .A1(_01667_),
    .A2(_01830_));
 sg13g2_nand2_1 _09654_ (.Y(_01832_),
    .A(\am_sdr0.am0.q[4] ),
    .B(net188));
 sg13g2_nand2_1 _09655_ (.Y(_01833_),
    .A(\am_sdr0.am0.q[5] ),
    .B(_01662_));
 sg13g2_o21ai_1 _09656_ (.B1(_01833_),
    .Y(_00149_),
    .A1(net12),
    .A2(_01832_));
 sg13g2_nand2_1 _09657_ (.Y(_01834_),
    .A(\am_sdr0.am0.q[5] ),
    .B(_01580_));
 sg13g2_nand2_1 _09658_ (.Y(_01835_),
    .A(\am_sdr0.am0.q[6] ),
    .B(_01662_));
 sg13g2_o21ai_1 _09659_ (.B1(_01835_),
    .Y(_00150_),
    .A1(net12),
    .A2(_01834_));
 sg13g2_nand2_1 _09660_ (.Y(_01836_),
    .A(\am_sdr0.am0.q[6] ),
    .B(net188));
 sg13g2_nand2_1 _09661_ (.Y(_01837_),
    .A(\am_sdr0.am0.q[7] ),
    .B(net13));
 sg13g2_o21ai_1 _09662_ (.B1(_01837_),
    .Y(_00151_),
    .A1(net12),
    .A2(_01836_));
 sg13g2_buf_1 _09663_ (.A(\am_sdr0.am0.right[0] ),
    .X(_01838_));
 sg13g2_xnor2_1 _09664_ (.Y(_01839_),
    .A(_01685_),
    .B(_01838_));
 sg13g2_o21ai_1 _09665_ (.B1(_01580_),
    .Y(_01840_),
    .A1(_01577_),
    .A2(_01680_));
 sg13g2_nand2_1 _09666_ (.Y(_01841_),
    .A(net41),
    .B(_01840_));
 sg13g2_buf_1 _09667_ (.A(_01841_),
    .X(_01842_));
 sg13g2_nand2_1 _09668_ (.Y(_01843_),
    .A(\am_sdr0.am0.r[0] ),
    .B(net22));
 sg13g2_o21ai_1 _09669_ (.B1(_01843_),
    .Y(_00152_),
    .A1(net24),
    .A2(_01839_));
 sg13g2_inv_1 _09670_ (.Y(_01844_),
    .A(_01838_));
 sg13g2_buf_1 _09671_ (.A(\am_sdr0.am0.r[9] ),
    .X(_01845_));
 sg13g2_buf_1 _09672_ (.A(_01845_),
    .X(_01846_));
 sg13g2_buf_1 _09673_ (.A(net300),
    .X(_01847_));
 sg13g2_buf_1 _09674_ (.A(\am_sdr0.am0.right[1] ),
    .X(_01848_));
 sg13g2_nor2_1 _09675_ (.A(_01848_),
    .B(_01845_),
    .Y(_01849_));
 sg13g2_a21o_1 _09676_ (.A2(net252),
    .A1(_00041_),
    .B1(_01849_),
    .X(_01850_));
 sg13g2_nor2b_1 _09677_ (.A(_00041_),
    .B_N(_01845_),
    .Y(_01851_));
 sg13g2_a21oi_1 _09678_ (.A1(_01838_),
    .A2(_01851_),
    .Y(_01852_),
    .B1(_01849_));
 sg13g2_nor2b_1 _09679_ (.A(_01845_),
    .B_N(_01848_),
    .Y(_01853_));
 sg13g2_a221oi_1 _09680_ (.B2(_01838_),
    .C1(_01685_),
    .B1(_01853_),
    .A1(_00041_),
    .Y(_01854_),
    .A2(net252));
 sg13g2_a21oi_1 _09681_ (.A1(_01685_),
    .A2(_01852_),
    .Y(_01855_),
    .B1(_01854_));
 sg13g2_a21oi_1 _09682_ (.A1(_01844_),
    .A2(_01850_),
    .Y(_01856_),
    .B1(_01855_));
 sg13g2_xnor2_1 _09683_ (.Y(_01857_),
    .A(_01689_),
    .B(_01856_));
 sg13g2_nand2_1 _09684_ (.Y(_01858_),
    .A(\am_sdr0.am0.r[1] ),
    .B(net22));
 sg13g2_o21ai_1 _09685_ (.B1(_01858_),
    .Y(_00153_),
    .A1(net24),
    .A2(_01857_));
 sg13g2_o21ai_1 _09686_ (.B1(_01685_),
    .Y(_01859_),
    .A1(_01689_),
    .A2(_01851_));
 sg13g2_o21ai_1 _09687_ (.B1(_01849_),
    .Y(_01860_),
    .A1(_01685_),
    .A2(_01689_));
 sg13g2_a21oi_1 _09688_ (.A1(_01859_),
    .A2(_01860_),
    .Y(_01861_),
    .B1(_01844_));
 sg13g2_a21oi_1 _09689_ (.A1(_01844_),
    .A2(_01853_),
    .Y(_01862_),
    .B1(_01851_));
 sg13g2_nor2_1 _09690_ (.A(_01690_),
    .B(_01862_),
    .Y(_01863_));
 sg13g2_nor2_1 _09691_ (.A(_01861_),
    .B(_01863_),
    .Y(_01864_));
 sg13g2_inv_1 _09692_ (.Y(_01865_),
    .A(\am_sdr0.am0.right[2] ));
 sg13g2_nor2_1 _09693_ (.A(_01838_),
    .B(_01848_),
    .Y(_01866_));
 sg13g2_xnor2_1 _09694_ (.Y(_01867_),
    .A(_01865_),
    .B(_01866_));
 sg13g2_nand2b_1 _09695_ (.Y(_01868_),
    .B(net300),
    .A_N(_00043_));
 sg13g2_o21ai_1 _09696_ (.B1(_01868_),
    .Y(_01869_),
    .A1(net300),
    .A2(_01867_));
 sg13g2_buf_1 _09697_ (.A(_01869_),
    .X(_01870_));
 sg13g2_xor2_1 _09698_ (.B(_01870_),
    .A(_00042_),
    .X(_01871_));
 sg13g2_xnor2_1 _09699_ (.Y(_01872_),
    .A(_01864_),
    .B(_01871_));
 sg13g2_nand2_1 _09700_ (.Y(_01873_),
    .A(\am_sdr0.am0.r[2] ),
    .B(net22));
 sg13g2_o21ai_1 _09701_ (.B1(_01873_),
    .Y(_00154_),
    .A1(net24),
    .A2(_01872_));
 sg13g2_o21ai_1 _09702_ (.B1(_01870_),
    .Y(_01874_),
    .A1(_01861_),
    .A2(_01863_));
 sg13g2_nor3_1 _09703_ (.A(_01861_),
    .B(_01863_),
    .C(_01870_),
    .Y(_01875_));
 sg13g2_a21oi_2 _09704_ (.B1(_01875_),
    .Y(_01876_),
    .A2(_01874_),
    .A1(_00042_));
 sg13g2_buf_1 _09705_ (.A(\am_sdr0.am0.right[3] ),
    .X(_01877_));
 sg13g2_inv_1 _09706_ (.Y(_01878_),
    .A(_01877_));
 sg13g2_nor2_1 _09707_ (.A(_01848_),
    .B(\am_sdr0.am0.right[2] ),
    .Y(_01879_));
 sg13g2_nand2_1 _09708_ (.Y(_01880_),
    .A(_00045_),
    .B(_01879_));
 sg13g2_xnor2_1 _09709_ (.Y(_01881_),
    .A(_01878_),
    .B(_01880_));
 sg13g2_nand2_1 _09710_ (.Y(_01882_),
    .A(net300),
    .B(_00044_));
 sg13g2_o21ai_1 _09711_ (.B1(_01882_),
    .Y(_01883_),
    .A1(_01846_),
    .A2(_01881_));
 sg13g2_xnor2_1 _09712_ (.Y(_01884_),
    .A(\am_sdr0.am0.left[3] ),
    .B(_01883_));
 sg13g2_xnor2_1 _09713_ (.Y(_01885_),
    .A(_01876_),
    .B(_01884_));
 sg13g2_nand2_1 _09714_ (.Y(_01886_),
    .A(\am_sdr0.am0.r[3] ),
    .B(_01842_));
 sg13g2_o21ai_1 _09715_ (.B1(_01886_),
    .Y(_00155_),
    .A1(net24),
    .A2(_01885_));
 sg13g2_inv_1 _09716_ (.Y(_01887_),
    .A(_01883_));
 sg13g2_nand2_1 _09717_ (.Y(_01888_),
    .A(_01876_),
    .B(_01887_));
 sg13g2_o21ai_1 _09718_ (.B1(\am_sdr0.am0.left[3] ),
    .Y(_01889_),
    .A1(_01876_),
    .A2(_01887_));
 sg13g2_nand2_1 _09719_ (.Y(_01890_),
    .A(_01888_),
    .B(_01889_));
 sg13g2_buf_1 _09720_ (.A(\am_sdr0.am0.right[4] ),
    .X(_01891_));
 sg13g2_nand2_1 _09721_ (.Y(_01892_),
    .A(_01865_),
    .B(_01866_));
 sg13g2_nor2_1 _09722_ (.A(_01877_),
    .B(_01892_),
    .Y(_01893_));
 sg13g2_xnor2_1 _09723_ (.Y(_01894_),
    .A(_01891_),
    .B(_01893_));
 sg13g2_nand2_1 _09724_ (.Y(_01895_),
    .A(net300),
    .B(_00046_));
 sg13g2_o21ai_1 _09725_ (.B1(_01895_),
    .Y(_01896_),
    .A1(_01846_),
    .A2(_01894_));
 sg13g2_xnor2_1 _09726_ (.Y(_01897_),
    .A(\am_sdr0.am0.left[4] ),
    .B(_01896_));
 sg13g2_xnor2_1 _09727_ (.Y(_01898_),
    .A(_01890_),
    .B(_01897_));
 sg13g2_nand2_1 _09728_ (.Y(_01899_),
    .A(\am_sdr0.am0.r[4] ),
    .B(net22));
 sg13g2_o21ai_1 _09729_ (.B1(_01899_),
    .Y(_00156_),
    .A1(net24),
    .A2(_01898_));
 sg13g2_a21oi_1 _09730_ (.A1(_01888_),
    .A2(_01889_),
    .Y(_01900_),
    .B1(_01896_));
 sg13g2_nand3_1 _09731_ (.B(_01889_),
    .C(_01896_),
    .A(_01888_),
    .Y(_01901_));
 sg13g2_o21ai_1 _09732_ (.B1(_01901_),
    .Y(_01902_),
    .A1(\am_sdr0.am0.left[4] ),
    .A2(_01900_));
 sg13g2_buf_1 _09733_ (.A(_01902_),
    .X(_01903_));
 sg13g2_buf_1 _09734_ (.A(\am_sdr0.am0.right[5] ),
    .X(_01904_));
 sg13g2_nor3_1 _09735_ (.A(_01877_),
    .B(_01891_),
    .C(_01880_),
    .Y(_01905_));
 sg13g2_xnor2_1 _09736_ (.Y(_01906_),
    .A(_01904_),
    .B(_01905_));
 sg13g2_nand2_1 _09737_ (.Y(_01907_),
    .A(net300),
    .B(_00047_));
 sg13g2_o21ai_1 _09738_ (.B1(_01907_),
    .Y(_01908_),
    .A1(net300),
    .A2(_01906_));
 sg13g2_xnor2_1 _09739_ (.Y(_01909_),
    .A(_01698_),
    .B(_01908_));
 sg13g2_xnor2_1 _09740_ (.Y(_01910_),
    .A(_01903_),
    .B(_01909_));
 sg13g2_nand2_1 _09741_ (.Y(_01911_),
    .A(\am_sdr0.am0.r[5] ),
    .B(net22));
 sg13g2_o21ai_1 _09742_ (.B1(_01911_),
    .Y(_00157_),
    .A1(net24),
    .A2(_01910_));
 sg13g2_or2_1 _09743_ (.X(_01912_),
    .B(_01908_),
    .A(_01903_));
 sg13g2_buf_1 _09744_ (.A(_01912_),
    .X(_01913_));
 sg13g2_a21o_1 _09745_ (.A2(_01908_),
    .A1(_01903_),
    .B1(_01698_),
    .X(_01914_));
 sg13g2_buf_1 _09746_ (.A(_01914_),
    .X(_01915_));
 sg13g2_nand2_1 _09747_ (.Y(_01916_),
    .A(_01913_),
    .B(_01915_));
 sg13g2_nor4_1 _09748_ (.A(_01877_),
    .B(_01891_),
    .C(_01904_),
    .D(_01892_),
    .Y(_01917_));
 sg13g2_xnor2_1 _09749_ (.Y(_01918_),
    .A(\am_sdr0.am0.right[6] ),
    .B(_01917_));
 sg13g2_nand2_1 _09750_ (.Y(_01919_),
    .A(net300),
    .B(_00048_));
 sg13g2_o21ai_1 _09751_ (.B1(_01919_),
    .Y(_01920_),
    .A1(net252),
    .A2(_01918_));
 sg13g2_xnor2_1 _09752_ (.Y(_01921_),
    .A(\am_sdr0.am0.left[6] ),
    .B(_01920_));
 sg13g2_xnor2_1 _09753_ (.Y(_01922_),
    .A(_01916_),
    .B(_01921_));
 sg13g2_nand2_1 _09754_ (.Y(_01923_),
    .A(\am_sdr0.am0.r[6] ),
    .B(net22));
 sg13g2_o21ai_1 _09755_ (.B1(_01923_),
    .Y(_00158_),
    .A1(_01684_),
    .A2(_01922_));
 sg13g2_a21oi_1 _09756_ (.A1(_01913_),
    .A2(_01915_),
    .Y(_01924_),
    .B1(_01920_));
 sg13g2_nand3_1 _09757_ (.B(_01915_),
    .C(_01920_),
    .A(_01913_),
    .Y(_01925_));
 sg13g2_o21ai_1 _09758_ (.B1(_01925_),
    .Y(_01926_),
    .A1(\am_sdr0.am0.left[6] ),
    .A2(_01924_));
 sg13g2_buf_1 _09759_ (.A(_01926_),
    .X(_01927_));
 sg13g2_inv_1 _09760_ (.Y(_01928_),
    .A(\am_sdr0.am0.right[7] ));
 sg13g2_nor4_2 _09761_ (.A(_01877_),
    .B(_01891_),
    .C(_01904_),
    .Y(_01929_),
    .D(\am_sdr0.am0.right[6] ));
 sg13g2_nand3_1 _09762_ (.B(_01879_),
    .C(_01929_),
    .A(_00045_),
    .Y(_01930_));
 sg13g2_xnor2_1 _09763_ (.Y(_01931_),
    .A(_01928_),
    .B(_01930_));
 sg13g2_nand2_1 _09764_ (.Y(_01932_),
    .A(net252),
    .B(_00049_));
 sg13g2_o21ai_1 _09765_ (.B1(_01932_),
    .Y(_01933_),
    .A1(_01847_),
    .A2(_01931_));
 sg13g2_buf_1 _09766_ (.A(_01933_),
    .X(_01934_));
 sg13g2_xnor2_1 _09767_ (.Y(_01935_),
    .A(_01703_),
    .B(_01934_));
 sg13g2_xnor2_1 _09768_ (.Y(_01936_),
    .A(_01927_),
    .B(_01935_));
 sg13g2_nand2_1 _09769_ (.Y(_01937_),
    .A(\am_sdr0.am0.r[7] ),
    .B(net22));
 sg13g2_o21ai_1 _09770_ (.B1(_01937_),
    .Y(_00159_),
    .A1(_01684_),
    .A2(_01936_));
 sg13g2_inv_1 _09771_ (.Y(_01938_),
    .A(\am_sdr0.am0.right[9] ));
 sg13g2_nand2_1 _09772_ (.Y(_01939_),
    .A(_01928_),
    .B(_01929_));
 sg13g2_nor3_1 _09773_ (.A(\am_sdr0.am0.right[8] ),
    .B(_01880_),
    .C(_01939_),
    .Y(_01940_));
 sg13g2_xnor2_1 _09774_ (.Y(_01941_),
    .A(_01938_),
    .B(_01940_));
 sg13g2_mux2_1 _09775_ (.A0(_01941_),
    .A1(_00050_),
    .S(net252),
    .X(_01942_));
 sg13g2_xnor2_1 _09776_ (.Y(_01943_),
    .A(\am_sdr0.am0.left[9] ),
    .B(_01942_));
 sg13g2_nand4_1 _09777_ (.B(_01928_),
    .C(_01879_),
    .A(_01844_),
    .Y(_01944_),
    .D(_01929_));
 sg13g2_xnor2_1 _09778_ (.Y(_01945_),
    .A(\am_sdr0.am0.right[8] ),
    .B(_01944_));
 sg13g2_nand2b_1 _09779_ (.Y(_01946_),
    .B(net252),
    .A_N(_00051_));
 sg13g2_o21ai_1 _09780_ (.B1(_01946_),
    .Y(_01947_),
    .A1(_01847_),
    .A2(_01945_));
 sg13g2_o21ai_1 _09781_ (.B1(_01703_),
    .Y(_01948_),
    .A1(_01927_),
    .A2(_01934_));
 sg13g2_nand2_1 _09782_ (.Y(_01949_),
    .A(_01927_),
    .B(_01934_));
 sg13g2_a22oi_1 _09783_ (.Y(_01950_),
    .B1(_01948_),
    .B2(_01949_),
    .A2(_01947_),
    .A1(\am_sdr0.am0.left[8] ));
 sg13g2_nor2_1 _09784_ (.A(\am_sdr0.am0.left[8] ),
    .B(_01947_),
    .Y(_01951_));
 sg13g2_nor2_1 _09785_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sg13g2_xnor2_1 _09786_ (.Y(_01953_),
    .A(_01943_),
    .B(_01952_));
 sg13g2_nand2_1 _09787_ (.Y(_01954_),
    .A(net252),
    .B(net22));
 sg13g2_o21ai_1 _09788_ (.B1(_01954_),
    .Y(_00160_),
    .A1(net24),
    .A2(_01953_));
 sg13g2_nand2_1 _09789_ (.Y(_01955_),
    .A(net136),
    .B(net14));
 sg13g2_o21ai_1 _09790_ (.B1(_01955_),
    .Y(_00161_),
    .A1(_01844_),
    .A2(net7));
 sg13g2_inv_1 _09791_ (.Y(_01956_),
    .A(_01848_));
 sg13g2_nand3_1 _09792_ (.B(net189),
    .C(net16),
    .A(net252),
    .Y(_01957_));
 sg13g2_o21ai_1 _09793_ (.B1(_01957_),
    .Y(_00162_),
    .A1(_01956_),
    .A2(net7));
 sg13g2_or2_1 _09794_ (.X(_01958_),
    .B(_01824_),
    .A(_01582_));
 sg13g2_o21ai_1 _09795_ (.B1(_01958_),
    .Y(_00163_),
    .A1(_01865_),
    .A2(net7));
 sg13g2_or2_1 _09796_ (.X(_01959_),
    .B(_01826_),
    .A(_01582_));
 sg13g2_o21ai_1 _09797_ (.B1(_01959_),
    .Y(_00164_),
    .A1(_01878_),
    .A2(net7));
 sg13g2_nand2_1 _09798_ (.Y(_01960_),
    .A(_01891_),
    .B(net25));
 sg13g2_o21ai_1 _09799_ (.B1(_01960_),
    .Y(_00165_),
    .A1(net25),
    .A2(_01828_));
 sg13g2_nand2_1 _09800_ (.Y(_01961_),
    .A(_01904_),
    .B(net25));
 sg13g2_o21ai_1 _09801_ (.B1(_01961_),
    .Y(_00166_),
    .A1(net25),
    .A2(_01830_));
 sg13g2_nand2_1 _09802_ (.Y(_01962_),
    .A(\am_sdr0.am0.right[6] ),
    .B(net25));
 sg13g2_o21ai_1 _09803_ (.B1(_01962_),
    .Y(_00167_),
    .A1(net25),
    .A2(_01832_));
 sg13g2_or2_1 _09804_ (.X(_01963_),
    .B(_01834_),
    .A(_01582_));
 sg13g2_o21ai_1 _09805_ (.B1(_01963_),
    .Y(_00168_),
    .A1(_01928_),
    .A2(net7));
 sg13g2_nand2_1 _09806_ (.Y(_01964_),
    .A(\am_sdr0.am0.right[8] ),
    .B(net25));
 sg13g2_o21ai_1 _09807_ (.B1(_01964_),
    .Y(_00169_),
    .A1(net25),
    .A2(_01836_));
 sg13g2_nand3_1 _09808_ (.B(net189),
    .C(net16),
    .A(\am_sdr0.am0.q[7] ),
    .Y(_01965_));
 sg13g2_o21ai_1 _09809_ (.B1(_01965_),
    .Y(_00170_),
    .A1(_01938_),
    .A2(net7));
 sg13g2_buf_1 _09810_ (.A(_01570_),
    .X(_01966_));
 sg13g2_a21oi_1 _09811_ (.A1(net301),
    .A2(_01966_),
    .Y(_01967_),
    .B1(_01458_));
 sg13g2_buf_1 _09812_ (.A(net310),
    .X(_01968_));
 sg13g2_o21ai_1 _09813_ (.B1(_01458_),
    .Y(_01969_),
    .A1(net251),
    .A2(_01966_));
 sg13g2_o21ai_1 _09814_ (.B1(_01969_),
    .Y(_00171_),
    .A1(_01569_),
    .A2(_01967_));
 sg13g2_buf_1 _09815_ (.A(\am_sdr0.am0.sum[0] ),
    .X(_01970_));
 sg13g2_nand2_1 _09816_ (.Y(_01971_),
    .A(\am_sdr0.am0.multB[0] ),
    .B(net256));
 sg13g2_nor2_1 _09817_ (.A(_01467_),
    .B(_01971_),
    .Y(_01972_));
 sg13g2_buf_1 _09818_ (.A(_01972_),
    .X(_01973_));
 sg13g2_nand2_1 _09819_ (.Y(_01974_),
    .A(net363),
    .B(_01973_));
 sg13g2_nand2_1 _09820_ (.Y(_01975_),
    .A(\am_sdr0.am0.state[0] ),
    .B(_01722_));
 sg13g2_a21o_1 _09821_ (.A2(_01971_),
    .A1(_01975_),
    .B1(_01467_),
    .X(_01976_));
 sg13g2_buf_2 _09822_ (.A(_01976_),
    .X(_01977_));
 sg13g2_buf_1 _09823_ (.A(_01977_),
    .X(_01978_));
 sg13g2_or2_1 _09824_ (.X(_01979_),
    .B(_01971_),
    .A(_01467_));
 sg13g2_buf_1 _09825_ (.A(_01979_),
    .X(_01980_));
 sg13g2_buf_1 _09826_ (.A(_01980_),
    .X(_01981_));
 sg13g2_nor2_1 _09827_ (.A(net363),
    .B(net31),
    .Y(_01982_));
 sg13g2_o21ai_1 _09828_ (.B1(_01970_),
    .Y(_01983_),
    .A1(_01978_),
    .A2(_01982_));
 sg13g2_o21ai_1 _09829_ (.B1(_01983_),
    .Y(_00174_),
    .A1(_01970_),
    .A2(_01974_));
 sg13g2_buf_1 _09830_ (.A(net36),
    .X(_01984_));
 sg13g2_or2_1 _09831_ (.X(_01985_),
    .B(_01770_),
    .A(\am_sdr0.am0.multA[0] ));
 sg13g2_buf_1 _09832_ (.A(_01985_),
    .X(_01986_));
 sg13g2_or4_1 _09833_ (.A(_01776_),
    .B(_01782_),
    .C(_01788_),
    .D(\am_sdr0.am0.multA[5] ),
    .X(_01987_));
 sg13g2_buf_2 _09834_ (.A(_01987_),
    .X(_01988_));
 sg13g2_or3_1 _09835_ (.A(_01801_),
    .B(_01804_),
    .C(_01744_),
    .X(_01989_));
 sg13g2_nor4_1 _09836_ (.A(_01798_),
    .B(_01986_),
    .C(_01988_),
    .D(_01989_),
    .Y(_01990_));
 sg13g2_xnor2_1 _09837_ (.Y(_01991_),
    .A(_01746_),
    .B(_01990_));
 sg13g2_nand2_1 _09838_ (.Y(_01992_),
    .A(_00062_),
    .B(net42));
 sg13g2_o21ai_1 _09839_ (.B1(_01992_),
    .Y(_01993_),
    .A1(_01565_),
    .A2(_01991_));
 sg13g2_buf_1 _09840_ (.A(_01993_),
    .X(_01994_));
 sg13g2_or2_1 _09841_ (.X(_01995_),
    .B(_01804_),
    .A(_01801_));
 sg13g2_nand2b_1 _09842_ (.Y(_01996_),
    .B(_00055_),
    .A_N(_01770_));
 sg13g2_buf_1 _09843_ (.A(_01996_),
    .X(_01997_));
 sg13g2_nor4_1 _09844_ (.A(_01798_),
    .B(_01988_),
    .C(_01995_),
    .D(_01997_),
    .Y(_01998_));
 sg13g2_xnor2_1 _09845_ (.Y(_01999_),
    .A(_01744_),
    .B(_01998_));
 sg13g2_nand2_1 _09846_ (.Y(_02000_),
    .A(_00061_),
    .B(net138));
 sg13g2_o21ai_1 _09847_ (.B1(_02000_),
    .Y(_02001_),
    .A1(net138),
    .A2(_01999_));
 sg13g2_buf_1 _09848_ (.A(_02001_),
    .X(_02002_));
 sg13g2_or2_1 _09849_ (.X(_02003_),
    .B(_02002_),
    .A(_01648_));
 sg13g2_buf_2 _09850_ (.A(_02003_),
    .X(_02004_));
 sg13g2_nor2_1 _09851_ (.A(_00054_),
    .B(net190),
    .Y(_02005_));
 sg13g2_or3_1 _09852_ (.A(_01776_),
    .B(_01782_),
    .C(_01997_),
    .X(_02006_));
 sg13g2_o21ai_1 _09853_ (.B1(_01782_),
    .Y(_02007_),
    .A1(_01776_),
    .A2(_01997_));
 sg13g2_and3_1 _09854_ (.X(_02008_),
    .A(_01455_),
    .B(_02006_),
    .C(_02007_));
 sg13g2_buf_1 _09855_ (.A(_02008_),
    .X(_02009_));
 sg13g2_nor2_1 _09856_ (.A(_02005_),
    .B(_02009_),
    .Y(_02010_));
 sg13g2_or3_1 _09857_ (.A(_01449_),
    .B(_00052_),
    .C(_01562_),
    .X(_02011_));
 sg13g2_a21oi_1 _09858_ (.A1(_01567_),
    .A2(_02011_),
    .Y(_02012_),
    .B1(_01970_));
 sg13g2_a221oi_1 _09859_ (.B2(_01450_),
    .C1(_01770_),
    .B1(_01454_),
    .A1(_01970_),
    .Y(_02013_),
    .A2(_01567_));
 sg13g2_o21ai_1 _09860_ (.B1(_01736_),
    .Y(_02014_),
    .A1(_02012_),
    .A2(_02013_));
 sg13g2_buf_1 _09861_ (.A(_02014_),
    .X(_02015_));
 sg13g2_nor2_1 _09862_ (.A(_00052_),
    .B(net190),
    .Y(_02016_));
 sg13g2_inv_1 _09863_ (.Y(_02017_),
    .A(_01770_));
 sg13g2_nor3_1 _09864_ (.A(net363),
    .B(_02017_),
    .C(net138),
    .Y(_02018_));
 sg13g2_inv_1 _09865_ (.Y(_02019_),
    .A(_01567_));
 sg13g2_o21ai_1 _09866_ (.B1(_02019_),
    .Y(_02020_),
    .A1(_02016_),
    .A2(_02018_));
 sg13g2_buf_1 _09867_ (.A(_02020_),
    .X(_02021_));
 sg13g2_xnor2_1 _09868_ (.Y(_02022_),
    .A(_01776_),
    .B(_01986_));
 sg13g2_mux2_1 _09869_ (.A0(_00053_),
    .A1(_02022_),
    .S(net190),
    .X(_02023_));
 sg13g2_buf_1 _09870_ (.A(_02023_),
    .X(_02024_));
 sg13g2_a221oi_1 _09871_ (.B2(_02021_),
    .C1(_02024_),
    .B1(_02015_),
    .A1(_01620_),
    .Y(_02025_),
    .A2(_02010_));
 sg13g2_buf_1 _09872_ (.A(_02025_),
    .X(_02026_));
 sg13g2_a221oi_1 _09873_ (.B2(_02021_),
    .C1(_01618_),
    .B1(_02015_),
    .A1(_01620_),
    .Y(_02027_),
    .A2(_02010_));
 sg13g2_buf_1 _09874_ (.A(_02027_),
    .X(_02028_));
 sg13g2_nor3_1 _09875_ (.A(_01621_),
    .B(_02005_),
    .C(_02009_),
    .Y(_02029_));
 sg13g2_or2_1 _09876_ (.X(_02030_),
    .B(_02024_),
    .A(_01618_));
 sg13g2_o21ai_1 _09877_ (.B1(_01621_),
    .Y(_02031_),
    .A1(_02005_),
    .A2(_02009_));
 sg13g2_o21ai_1 _09878_ (.B1(_02031_),
    .Y(_02032_),
    .A1(_02029_),
    .A2(_02030_));
 sg13g2_nor2_1 _09879_ (.A(_01986_),
    .B(_01988_),
    .Y(_02033_));
 sg13g2_xnor2_1 _09880_ (.Y(_02034_),
    .A(_01798_),
    .B(_02033_));
 sg13g2_nand2_1 _09881_ (.Y(_02035_),
    .A(_00058_),
    .B(net138));
 sg13g2_o21ai_1 _09882_ (.B1(_02035_),
    .Y(_02036_),
    .A1(net138),
    .A2(_02034_));
 sg13g2_buf_1 _09883_ (.A(_02036_),
    .X(_02037_));
 sg13g2_nand2b_1 _09884_ (.Y(_02038_),
    .B(_01564_),
    .A_N(_00057_));
 sg13g2_nor3_1 _09885_ (.A(_01776_),
    .B(_01782_),
    .C(_01788_),
    .Y(_02039_));
 sg13g2_nor2b_1 _09886_ (.A(_01770_),
    .B_N(_00055_),
    .Y(_02040_));
 sg13g2_a21oi_1 _09887_ (.A1(_02039_),
    .A2(_02040_),
    .Y(_02041_),
    .B1(_01790_));
 sg13g2_and3_1 _09888_ (.X(_02042_),
    .A(_01790_),
    .B(_02039_),
    .C(_02040_));
 sg13g2_buf_1 _09889_ (.A(_02042_),
    .X(_02043_));
 sg13g2_or3_1 _09890_ (.A(_01564_),
    .B(_02041_),
    .C(_02043_),
    .X(_02044_));
 sg13g2_nand3_1 _09891_ (.B(_02038_),
    .C(_02044_),
    .A(_01629_),
    .Y(_02045_));
 sg13g2_buf_1 _09892_ (.A(_02045_),
    .X(_02046_));
 sg13g2_a21o_1 _09893_ (.A2(_02044_),
    .A1(_02038_),
    .B1(_01629_),
    .X(_02047_));
 sg13g2_buf_1 _09894_ (.A(_02047_),
    .X(_02048_));
 sg13g2_nor4_1 _09895_ (.A(net363),
    .B(_01770_),
    .C(_01776_),
    .D(_01782_),
    .Y(_02049_));
 sg13g2_xnor2_1 _09896_ (.Y(_02050_),
    .A(_01788_),
    .B(_02049_));
 sg13g2_nor3_1 _09897_ (.A(_01449_),
    .B(_00056_),
    .C(_01562_),
    .Y(_02051_));
 sg13g2_a21oi_2 _09898_ (.B1(_02051_),
    .Y(_02052_),
    .A2(_02050_),
    .A1(net190));
 sg13g2_xor2_1 _09899_ (.B(_02052_),
    .A(_01625_),
    .X(_02053_));
 sg13g2_nand4_1 _09900_ (.B(_02046_),
    .C(_02048_),
    .A(_02037_),
    .Y(_02054_),
    .D(_02053_));
 sg13g2_or4_1 _09901_ (.A(_02026_),
    .B(_02028_),
    .C(_02032_),
    .D(_02054_),
    .X(_02055_));
 sg13g2_nand4_1 _09902_ (.B(_02046_),
    .C(_02048_),
    .A(_01633_),
    .Y(_02056_),
    .D(_02053_));
 sg13g2_or4_1 _09903_ (.A(_02026_),
    .B(_02028_),
    .C(_02032_),
    .D(_02056_),
    .X(_02057_));
 sg13g2_o21ai_1 _09904_ (.B1(_01629_),
    .Y(_02058_),
    .A1(_02041_),
    .A2(_02043_));
 sg13g2_nand2b_1 _09905_ (.Y(_02059_),
    .B(_01625_),
    .A_N(_02050_));
 sg13g2_nor3_1 _09906_ (.A(_01629_),
    .B(_02041_),
    .C(_02043_),
    .Y(_02060_));
 sg13g2_a21oi_1 _09907_ (.A1(_02058_),
    .A2(_02059_),
    .Y(_02061_),
    .B1(_02060_));
 sg13g2_and2_1 _09908_ (.A(_01625_),
    .B(_00056_),
    .X(_02062_));
 sg13g2_o21ai_1 _09909_ (.B1(_02062_),
    .Y(_02063_),
    .A1(_01629_),
    .A2(_00057_));
 sg13g2_nand2_1 _09910_ (.Y(_02064_),
    .A(_01629_),
    .B(_00057_));
 sg13g2_a21oi_1 _09911_ (.A1(_02063_),
    .A2(_02064_),
    .Y(_02065_),
    .B1(net190));
 sg13g2_a21o_1 _09912_ (.A2(_02061_),
    .A1(_01456_),
    .B1(_02065_),
    .X(_02066_));
 sg13g2_buf_1 _09913_ (.A(_02066_),
    .X(_02067_));
 sg13g2_o21ai_1 _09914_ (.B1(_02067_),
    .Y(_02068_),
    .A1(_01633_),
    .A2(_02037_));
 sg13g2_nand2_1 _09915_ (.Y(_02069_),
    .A(_01633_),
    .B(_02037_));
 sg13g2_and4_1 _09916_ (.A(_02055_),
    .B(_02057_),
    .C(_02068_),
    .D(_02069_),
    .X(_02070_));
 sg13g2_buf_2 _09917_ (.A(_02070_),
    .X(_02071_));
 sg13g2_nor3_1 _09918_ (.A(_01798_),
    .B(_01988_),
    .C(_01997_),
    .Y(_02072_));
 sg13g2_xnor2_1 _09919_ (.Y(_02073_),
    .A(_01801_),
    .B(_02072_));
 sg13g2_nand2_1 _09920_ (.Y(_02074_),
    .A(_00059_),
    .B(_01565_));
 sg13g2_o21ai_1 _09921_ (.B1(_02074_),
    .Y(_02075_),
    .A1(net42),
    .A2(_02073_));
 sg13g2_buf_1 _09922_ (.A(_02075_),
    .X(_02076_));
 sg13g2_nand2_1 _09923_ (.Y(_02077_),
    .A(_01648_),
    .B(_02002_));
 sg13g2_buf_2 _09924_ (.A(_02077_),
    .X(_02078_));
 sg13g2_nor4_1 _09925_ (.A(_01798_),
    .B(_01801_),
    .C(_01986_),
    .D(_01988_),
    .Y(_02079_));
 sg13g2_xnor2_1 _09926_ (.Y(_02080_),
    .A(_01804_),
    .B(_02079_));
 sg13g2_nand2_1 _09927_ (.Y(_02081_),
    .A(_00060_),
    .B(net138));
 sg13g2_o21ai_1 _09928_ (.B1(_02081_),
    .Y(_02082_),
    .A1(net138),
    .A2(_02080_));
 sg13g2_buf_2 _09929_ (.A(_02082_),
    .X(_02083_));
 sg13g2_nand2_1 _09930_ (.Y(_02084_),
    .A(_01643_),
    .B(_02083_));
 sg13g2_nand2_1 _09931_ (.Y(_02085_),
    .A(_02078_),
    .B(_02084_));
 sg13g2_a21oi_2 _09932_ (.B1(_02085_),
    .Y(_02086_),
    .A2(_02076_),
    .A1(\am_sdr0.am0.sum[7] ));
 sg13g2_nand3b_1 _09933_ (.B(_02084_),
    .C(_01638_),
    .Y(_02087_),
    .A_N(_02076_));
 sg13g2_o21ai_1 _09934_ (.B1(_02087_),
    .Y(_02088_),
    .A1(_01643_),
    .A2(_02083_));
 sg13g2_buf_1 _09935_ (.A(_02088_),
    .X(_02089_));
 sg13g2_a22oi_1 _09936_ (.Y(_02090_),
    .B1(_02089_),
    .B2(_02078_),
    .A2(_02086_),
    .A1(_02071_));
 sg13g2_nand2_1 _09937_ (.Y(_02091_),
    .A(_02004_),
    .B(_02090_));
 sg13g2_xnor2_1 _09938_ (.Y(_02092_),
    .A(_01994_),
    .B(_02091_));
 sg13g2_nand2_1 _09939_ (.Y(_02093_),
    .A(net30),
    .B(_02092_));
 sg13g2_nor2_1 _09940_ (.A(_01981_),
    .B(_02092_),
    .Y(_02094_));
 sg13g2_o21ai_1 _09941_ (.B1(_01652_),
    .Y(_02095_),
    .A1(net32),
    .A2(_02094_));
 sg13g2_o21ai_1 _09942_ (.B1(_02095_),
    .Y(_00175_),
    .A1(_01652_),
    .A2(_02093_));
 sg13g2_or2_1 _09943_ (.X(_02096_),
    .B(_01989_),
    .A(_01746_));
 sg13g2_nor2b_1 _09944_ (.A(_02096_),
    .B_N(_02072_),
    .Y(_02097_));
 sg13g2_xnor2_1 _09945_ (.Y(_02098_),
    .A(_01749_),
    .B(_02097_));
 sg13g2_nand2_1 _09946_ (.Y(_02099_),
    .A(_00063_),
    .B(net42));
 sg13g2_o21ai_1 _09947_ (.B1(_02099_),
    .Y(_02100_),
    .A1(net42),
    .A2(_02098_));
 sg13g2_buf_1 _09948_ (.A(_02100_),
    .X(_02101_));
 sg13g2_nand3_1 _09949_ (.B(_02004_),
    .C(_02090_),
    .A(_01994_),
    .Y(_02102_));
 sg13g2_a21oi_1 _09950_ (.A1(_02004_),
    .A2(_02090_),
    .Y(_02103_),
    .B1(_01994_));
 sg13g2_a21oi_1 _09951_ (.A1(_01653_),
    .A2(_02102_),
    .Y(_02104_),
    .B1(_02103_));
 sg13g2_xnor2_1 _09952_ (.Y(_02105_),
    .A(_02101_),
    .B(_02104_));
 sg13g2_a21oi_1 _09953_ (.A1(net36),
    .A2(_02105_),
    .Y(_02106_),
    .B1(net32));
 sg13g2_nand3b_1 _09954_ (.B(_01591_),
    .C(net30),
    .Y(_02107_),
    .A_N(_02105_));
 sg13g2_o21ai_1 _09955_ (.B1(_02107_),
    .Y(_00176_),
    .A1(_01591_),
    .A2(_02106_));
 sg13g2_nor2b_1 _09956_ (.A(_01746_),
    .B_N(_01990_),
    .Y(_02108_));
 sg13g2_nor2b_1 _09957_ (.A(_01749_),
    .B_N(_02108_),
    .Y(_02109_));
 sg13g2_xnor2_1 _09958_ (.Y(_02110_),
    .A(_01752_),
    .B(_02109_));
 sg13g2_nand2_1 _09959_ (.Y(_02111_),
    .A(_00064_),
    .B(net42));
 sg13g2_o21ai_1 _09960_ (.B1(_02111_),
    .Y(_02112_),
    .A1(net33),
    .A2(_02110_));
 sg13g2_and2_1 _09961_ (.A(_01994_),
    .B(_02101_),
    .X(_02113_));
 sg13g2_nand2_1 _09962_ (.Y(_02114_),
    .A(_02004_),
    .B(_02113_));
 sg13g2_a221oi_1 _09963_ (.B2(_02078_),
    .C1(_02114_),
    .B1(_02089_),
    .A1(_02071_),
    .Y(_02115_),
    .A2(_02086_));
 sg13g2_nand3_1 _09964_ (.B(_02004_),
    .C(_02101_),
    .A(_01652_),
    .Y(_02116_));
 sg13g2_a221oi_1 _09965_ (.B2(_02078_),
    .C1(_02116_),
    .B1(_02089_),
    .A1(_02071_),
    .Y(_02117_),
    .A2(_02086_));
 sg13g2_nand3_1 _09966_ (.B(_01994_),
    .C(_02004_),
    .A(_01590_),
    .Y(_02118_));
 sg13g2_a221oi_1 _09967_ (.B2(_02078_),
    .C1(_02118_),
    .B1(_02089_),
    .A1(_02071_),
    .Y(_02119_),
    .A2(_02086_));
 sg13g2_nand3_1 _09968_ (.B(_01590_),
    .C(_02004_),
    .A(_01652_),
    .Y(_02120_));
 sg13g2_a221oi_1 _09969_ (.B2(_02078_),
    .C1(_02120_),
    .B1(_02089_),
    .A1(_02071_),
    .Y(_02121_),
    .A2(_02086_));
 sg13g2_nor4_2 _09970_ (.A(_02115_),
    .B(_02117_),
    .C(_02119_),
    .Y(_02122_),
    .D(_02121_));
 sg13g2_and3_1 _09971_ (.X(_02123_),
    .A(_01652_),
    .B(_01590_),
    .C(_01994_));
 sg13g2_a221oi_1 _09972_ (.B2(_01652_),
    .C1(_02123_),
    .B1(_02113_),
    .A1(_01590_),
    .Y(_02124_),
    .A2(_02101_));
 sg13g2_buf_1 _09973_ (.A(_02124_),
    .X(_02125_));
 sg13g2_nand2_1 _09974_ (.Y(_02126_),
    .A(_02122_),
    .B(_02125_));
 sg13g2_xnor2_1 _09975_ (.Y(_02127_),
    .A(_02112_),
    .B(_02126_));
 sg13g2_a21o_1 _09976_ (.A2(_02127_),
    .A1(net36),
    .B1(_01977_),
    .X(_02128_));
 sg13g2_nor3_1 _09977_ (.A(_01597_),
    .B(net31),
    .C(_02127_),
    .Y(_02129_));
 sg13g2_a21o_1 _09978_ (.A2(_02128_),
    .A1(_01597_),
    .B1(_02129_),
    .X(_00177_));
 sg13g2_nor2_1 _09979_ (.A(_01749_),
    .B(_01752_),
    .Y(_02130_));
 sg13g2_nand2_1 _09980_ (.Y(_02131_),
    .A(_02097_),
    .B(_02130_));
 sg13g2_xor2_1 _09981_ (.B(_02131_),
    .A(_01755_),
    .X(_02132_));
 sg13g2_nand2_1 _09982_ (.Y(_02133_),
    .A(_00065_),
    .B(net42));
 sg13g2_o21ai_1 _09983_ (.B1(_02133_),
    .Y(_02134_),
    .A1(net33),
    .A2(_02132_));
 sg13g2_buf_1 _09984_ (.A(_02134_),
    .X(_02135_));
 sg13g2_or2_1 _09985_ (.X(_02136_),
    .B(_02112_),
    .A(_01597_));
 sg13g2_buf_1 _09986_ (.A(_02136_),
    .X(_02137_));
 sg13g2_and2_1 _09987_ (.A(_01597_),
    .B(_02112_),
    .X(_02138_));
 sg13g2_nand3b_1 _09988_ (.B(_02125_),
    .C(_02122_),
    .Y(_02139_),
    .A_N(_02138_));
 sg13g2_nand2_1 _09989_ (.Y(_02140_),
    .A(_02137_),
    .B(_02139_));
 sg13g2_xnor2_1 _09990_ (.Y(_02141_),
    .A(_02135_),
    .B(_02140_));
 sg13g2_nand2_1 _09991_ (.Y(_02142_),
    .A(net30),
    .B(_02141_));
 sg13g2_nor2_1 _09992_ (.A(net31),
    .B(_02141_),
    .Y(_02143_));
 sg13g2_o21ai_1 _09993_ (.B1(_01603_),
    .Y(_02144_),
    .A1(net32),
    .A2(_02143_));
 sg13g2_o21ai_1 _09994_ (.B1(_02144_),
    .Y(_00178_),
    .A1(_01603_),
    .A2(_02142_));
 sg13g2_nor3_1 _09995_ (.A(_01749_),
    .B(_01752_),
    .C(_01755_),
    .Y(_02145_));
 sg13g2_nand2_1 _09996_ (.Y(_02146_),
    .A(_02108_),
    .B(_02145_));
 sg13g2_xor2_1 _09997_ (.B(_02146_),
    .A(_01758_),
    .X(_02147_));
 sg13g2_nor2_1 _09998_ (.A(net42),
    .B(_02147_),
    .Y(_02148_));
 sg13g2_a21oi_1 _09999_ (.A1(_00066_),
    .A2(net33),
    .Y(_02149_),
    .B1(_02148_));
 sg13g2_inv_1 _10000_ (.Y(_02150_),
    .A(_02149_));
 sg13g2_and2_1 _10001_ (.A(_02135_),
    .B(_02150_),
    .X(_02151_));
 sg13g2_buf_1 _10002_ (.A(_02151_),
    .X(_02152_));
 sg13g2_nand2_1 _10003_ (.Y(_02153_),
    .A(_02137_),
    .B(_02152_));
 sg13g2_nor2b_1 _10004_ (.A(_02149_),
    .B_N(_01603_),
    .Y(_02154_));
 sg13g2_nand2_1 _10005_ (.Y(_02155_),
    .A(_02137_),
    .B(_02154_));
 sg13g2_a22oi_1 _10006_ (.Y(_02156_),
    .B1(_02153_),
    .B2(_02155_),
    .A2(_02125_),
    .A1(_02122_));
 sg13g2_o21ai_1 _10007_ (.B1(_02138_),
    .Y(_02157_),
    .A1(_02152_),
    .A2(_02154_));
 sg13g2_nand2_1 _10008_ (.Y(_02158_),
    .A(_01603_),
    .B(_02152_));
 sg13g2_nand2_1 _10009_ (.Y(_02159_),
    .A(_02157_),
    .B(_02158_));
 sg13g2_and2_1 _10010_ (.A(_01603_),
    .B(_02135_),
    .X(_02160_));
 sg13g2_or2_1 _10011_ (.X(_02161_),
    .B(_02135_),
    .A(_01603_));
 sg13g2_and3_1 _10012_ (.X(_02162_),
    .A(_02137_),
    .B(_02139_),
    .C(_02161_));
 sg13g2_nor3_1 _10013_ (.A(_02150_),
    .B(_02160_),
    .C(_02162_),
    .Y(_02163_));
 sg13g2_or3_1 _10014_ (.A(_02156_),
    .B(_02159_),
    .C(_02163_),
    .X(_02164_));
 sg13g2_a21oi_1 _10015_ (.A1(net36),
    .A2(_02164_),
    .Y(_02165_),
    .B1(_01978_));
 sg13g2_nand3b_1 _10016_ (.B(_01607_),
    .C(_01984_),
    .Y(_02166_),
    .A_N(_02164_));
 sg13g2_o21ai_1 _10017_ (.B1(_02166_),
    .Y(_00179_),
    .A1(_01607_),
    .A2(_02165_));
 sg13g2_nor2b_1 _10018_ (.A(_01758_),
    .B_N(_02145_),
    .Y(_02167_));
 sg13g2_nand2_1 _10019_ (.Y(_02168_),
    .A(_02097_),
    .B(_02167_));
 sg13g2_xor2_1 _10020_ (.B(_02168_),
    .A(_01762_),
    .X(_02169_));
 sg13g2_nand2_1 _10021_ (.Y(_02170_),
    .A(_00067_),
    .B(net33));
 sg13g2_o21ai_1 _10022_ (.B1(_02170_),
    .Y(_02171_),
    .A1(_01566_),
    .A2(_02169_));
 sg13g2_buf_2 _10023_ (.A(_02171_),
    .X(_02172_));
 sg13g2_nor2_1 _10024_ (.A(_02156_),
    .B(_02159_),
    .Y(_02173_));
 sg13g2_a21oi_1 _10025_ (.A1(_01607_),
    .A2(_02173_),
    .Y(_02174_),
    .B1(_02163_));
 sg13g2_xnor2_1 _10026_ (.Y(_02175_),
    .A(_02172_),
    .B(_02174_));
 sg13g2_a21o_1 _10027_ (.A2(_02175_),
    .A1(_01973_),
    .B1(_01977_),
    .X(_02176_));
 sg13g2_nor3_1 _10028_ (.A(_01611_),
    .B(net31),
    .C(_02175_),
    .Y(_02177_));
 sg13g2_a21o_1 _10029_ (.A2(_02176_),
    .A1(_01611_),
    .B1(_02177_),
    .X(_00180_));
 sg13g2_xnor2_1 _10030_ (.Y(_02178_),
    .A(\am_sdr0.am0.sum[16] ),
    .B(\am_sdr0.am0.multA[16] ));
 sg13g2_nor2b_1 _10031_ (.A(_01762_),
    .B_N(_02167_),
    .Y(_02179_));
 sg13g2_a21oi_1 _10032_ (.A1(_02108_),
    .A2(_02179_),
    .Y(_02180_),
    .B1(net33));
 sg13g2_xnor2_1 _10033_ (.Y(_02181_),
    .A(_02178_),
    .B(_02180_));
 sg13g2_o21ai_1 _10034_ (.B1(\am_sdr0.am0.sum[14] ),
    .Y(_02182_),
    .A1(_01611_),
    .A2(_02172_));
 sg13g2_nor2b_1 _10035_ (.A(_02149_),
    .B_N(_02172_),
    .Y(_02183_));
 sg13g2_o21ai_1 _10036_ (.B1(_02183_),
    .Y(_02184_),
    .A1(_02160_),
    .A2(_02162_));
 sg13g2_o21ai_1 _10037_ (.B1(_02184_),
    .Y(_02185_),
    .A1(_02163_),
    .A2(_02182_));
 sg13g2_nor3_1 _10038_ (.A(_02156_),
    .B(_02159_),
    .C(_02172_),
    .Y(_02186_));
 sg13g2_nand2_1 _10039_ (.Y(_02187_),
    .A(_01611_),
    .B(_02181_));
 sg13g2_or3_1 _10040_ (.A(_01611_),
    .B(_02172_),
    .C(_02181_),
    .X(_02188_));
 sg13g2_o21ai_1 _10041_ (.B1(_02188_),
    .Y(_02189_),
    .A1(_02186_),
    .A2(_02187_));
 sg13g2_a21oi_1 _10042_ (.A1(_02181_),
    .A2(_02185_),
    .Y(_02190_),
    .B1(_02189_));
 sg13g2_and2_1 _10043_ (.A(_01611_),
    .B(_02172_),
    .X(_02191_));
 sg13g2_nor4_1 _10044_ (.A(_01980_),
    .B(_02174_),
    .C(_02181_),
    .D(_02191_),
    .Y(_02192_));
 sg13g2_a21oi_1 _10045_ (.A1(\am_sdr0.am0.sum[16] ),
    .A2(net32),
    .Y(_02193_),
    .B1(_02192_));
 sg13g2_o21ai_1 _10046_ (.B1(_02193_),
    .Y(_00181_),
    .A1(net31),
    .A2(_02190_));
 sg13g2_nor2_1 _10047_ (.A(_02017_),
    .B(net33),
    .Y(_02194_));
 sg13g2_nor3_1 _10048_ (.A(net363),
    .B(_02016_),
    .C(_02194_),
    .Y(_02195_));
 sg13g2_a22oi_1 _10049_ (.Y(_02196_),
    .B1(_02194_),
    .B2(net363),
    .A2(_01566_),
    .A1(_00052_));
 sg13g2_a221oi_1 _10050_ (.B2(net363),
    .C1(_01970_),
    .B1(_02016_),
    .A1(_02017_),
    .Y(_02197_),
    .A2(_01456_));
 sg13g2_a21oi_1 _10051_ (.A1(_01970_),
    .A2(_02196_),
    .Y(_02198_),
    .B1(_02197_));
 sg13g2_nor2_1 _10052_ (.A(_02195_),
    .B(_02198_),
    .Y(_02199_));
 sg13g2_nand2_1 _10053_ (.Y(_02200_),
    .A(_01984_),
    .B(_02199_));
 sg13g2_nor2_1 _10054_ (.A(net31),
    .B(_02199_),
    .Y(_02201_));
 sg13g2_o21ai_1 _10055_ (.B1(_01567_),
    .Y(_02202_),
    .A1(net32),
    .A2(_02201_));
 sg13g2_o21ai_1 _10056_ (.B1(_02202_),
    .Y(_00182_),
    .A1(_01567_),
    .A2(_02200_));
 sg13g2_nand2_1 _10057_ (.Y(_02203_),
    .A(_02015_),
    .B(_02021_));
 sg13g2_xnor2_1 _10058_ (.Y(_02204_),
    .A(_02203_),
    .B(_02024_));
 sg13g2_nand2_1 _10059_ (.Y(_02205_),
    .A(net30),
    .B(_02204_));
 sg13g2_nor2_1 _10060_ (.A(net31),
    .B(_02204_),
    .Y(_02206_));
 sg13g2_o21ai_1 _10061_ (.B1(_01618_),
    .Y(_02207_),
    .A1(_01977_),
    .A2(_02206_));
 sg13g2_o21ai_1 _10062_ (.B1(_02207_),
    .Y(_00183_),
    .A1(_01618_),
    .A2(_02205_));
 sg13g2_nand2b_1 _10063_ (.Y(_02208_),
    .B(_02203_),
    .A_N(_02024_));
 sg13g2_nor2b_1 _10064_ (.A(_02203_),
    .B_N(_02024_),
    .Y(_02209_));
 sg13g2_a21oi_1 _10065_ (.A1(_01618_),
    .A2(_02208_),
    .Y(_02210_),
    .B1(_02209_));
 sg13g2_xnor2_1 _10066_ (.Y(_02211_),
    .A(_02010_),
    .B(_02210_));
 sg13g2_nand2_1 _10067_ (.Y(_02212_),
    .A(net30),
    .B(_02211_));
 sg13g2_nor2_1 _10068_ (.A(_01980_),
    .B(_02211_),
    .Y(_02213_));
 sg13g2_o21ai_1 _10069_ (.B1(_01620_),
    .Y(_02214_),
    .A1(_01977_),
    .A2(_02213_));
 sg13g2_o21ai_1 _10070_ (.B1(_02214_),
    .Y(_00184_),
    .A1(_01620_),
    .A2(_02212_));
 sg13g2_nor3_2 _10071_ (.A(_02026_),
    .B(_02028_),
    .C(_02032_),
    .Y(_02215_));
 sg13g2_xnor2_1 _10072_ (.Y(_02216_),
    .A(_02215_),
    .B(_02052_));
 sg13g2_a21o_1 _10073_ (.A2(_02216_),
    .A1(net36),
    .B1(_01977_),
    .X(_02217_));
 sg13g2_nor3_1 _10074_ (.A(_01625_),
    .B(net31),
    .C(_02216_),
    .Y(_02218_));
 sg13g2_a21o_1 _10075_ (.A2(_02217_),
    .A1(_01625_),
    .B1(_02218_),
    .X(_00185_));
 sg13g2_nand2_1 _10076_ (.Y(_02219_),
    .A(_02046_),
    .B(_02048_));
 sg13g2_a21o_1 _10077_ (.A2(_02052_),
    .A1(_02215_),
    .B1(_01625_),
    .X(_02220_));
 sg13g2_o21ai_1 _10078_ (.B1(_02220_),
    .Y(_02221_),
    .A1(_02215_),
    .A2(_02052_));
 sg13g2_xnor2_1 _10079_ (.Y(_02222_),
    .A(_02219_),
    .B(_02221_));
 sg13g2_nand2_1 _10080_ (.Y(_02223_),
    .A(_01629_),
    .B(net32));
 sg13g2_o21ai_1 _10081_ (.B1(_02223_),
    .Y(_00186_),
    .A1(_01981_),
    .A2(_02222_));
 sg13g2_and4_1 _10082_ (.A(_02215_),
    .B(_02046_),
    .C(_02048_),
    .D(_02053_),
    .X(_02224_));
 sg13g2_nor3_1 _10083_ (.A(_02037_),
    .B(_02067_),
    .C(_02224_),
    .Y(_02225_));
 sg13g2_inv_1 _10084_ (.Y(_02226_),
    .A(_02225_));
 sg13g2_o21ai_1 _10085_ (.B1(_02037_),
    .Y(_02227_),
    .A1(_02067_),
    .A2(_02224_));
 sg13g2_nand3_1 _10086_ (.B(_02226_),
    .C(_02227_),
    .A(net36),
    .Y(_02228_));
 sg13g2_a21oi_1 _10087_ (.A1(_02226_),
    .A2(_02227_),
    .Y(_02229_),
    .B1(_01980_));
 sg13g2_o21ai_1 _10088_ (.B1(_01633_),
    .Y(_02230_),
    .A1(_01977_),
    .A2(_02229_));
 sg13g2_o21ai_1 _10089_ (.B1(_02230_),
    .Y(_00187_),
    .A1(_01633_),
    .A2(_02228_));
 sg13g2_nor2b_1 _10090_ (.A(_02076_),
    .B_N(_02071_),
    .Y(_02231_));
 sg13g2_nand2b_1 _10091_ (.Y(_02232_),
    .B(_02076_),
    .A_N(_02071_));
 sg13g2_nand2b_1 _10092_ (.Y(_02233_),
    .B(_02232_),
    .A_N(_02231_));
 sg13g2_a21oi_1 _10093_ (.A1(net36),
    .A2(_02233_),
    .Y(_02234_),
    .B1(net32));
 sg13g2_nand3b_1 _10094_ (.B(_01638_),
    .C(net30),
    .Y(_02235_),
    .A_N(_02233_));
 sg13g2_o21ai_1 _10095_ (.B1(_02235_),
    .Y(_00188_),
    .A1(_01638_),
    .A2(_02234_));
 sg13g2_a21oi_1 _10096_ (.A1(_01638_),
    .A2(_02232_),
    .Y(_02236_),
    .B1(_02231_));
 sg13g2_xnor2_1 _10097_ (.Y(_02237_),
    .A(_02083_),
    .B(_02236_));
 sg13g2_a21oi_1 _10098_ (.A1(net36),
    .A2(_02237_),
    .Y(_02238_),
    .B1(net32));
 sg13g2_nand3b_1 _10099_ (.B(_01644_),
    .C(net30),
    .Y(_02239_),
    .A_N(_02237_));
 sg13g2_o21ai_1 _10100_ (.B1(_02239_),
    .Y(_00189_),
    .A1(_01644_),
    .A2(_02238_));
 sg13g2_a21o_1 _10101_ (.A2(_02236_),
    .A1(_02083_),
    .B1(_01643_),
    .X(_02240_));
 sg13g2_o21ai_1 _10102_ (.B1(_02240_),
    .Y(_02241_),
    .A1(_02083_),
    .A2(_02236_));
 sg13g2_xnor2_1 _10103_ (.Y(_02242_),
    .A(_02002_),
    .B(_02241_));
 sg13g2_nand2_1 _10104_ (.Y(_02243_),
    .A(net30),
    .B(_02242_));
 sg13g2_nor2_1 _10105_ (.A(_01980_),
    .B(_02242_),
    .Y(_02244_));
 sg13g2_o21ai_1 _10106_ (.B1(_01648_),
    .Y(_02245_),
    .A1(_01977_),
    .A2(_02244_));
 sg13g2_o21ai_1 _10107_ (.B1(_02245_),
    .Y(_00190_),
    .A1(_01648_),
    .A2(_02243_));
 sg13g2_buf_2 _10108_ (.A(\am_sdr0.cic0.integ_sample[0] ),
    .X(_02246_));
 sg13g2_buf_2 _10109_ (.A(\am_sdr0.cic0.integ3[0] ),
    .X(_02247_));
 sg13g2_buf_1 _10110_ (.A(\am_sdr0.cic0.count[4] ),
    .X(_02248_));
 sg13g2_inv_1 _10111_ (.Y(_02249_),
    .A(\am_sdr0.cic0.count[3] ));
 sg13g2_nand3_1 _10112_ (.B(\am_sdr0.cic0.count[0] ),
    .C(\am_sdr0.cic0.count[2] ),
    .A(\am_sdr0.cic0.count[1] ),
    .Y(_02250_));
 sg13g2_nor2_2 _10113_ (.A(_02249_),
    .B(_02250_),
    .Y(_02251_));
 sg13g2_nand3_1 _10114_ (.B(_02248_),
    .C(_02251_),
    .A(\am_sdr0.cic0.count[5] ),
    .Y(_02252_));
 sg13g2_or3_1 _10115_ (.A(\am_sdr0.cic0.count[7] ),
    .B(\am_sdr0.cic0.count[6] ),
    .C(_02252_),
    .X(_02253_));
 sg13g2_buf_1 _10116_ (.A(_02253_),
    .X(_02254_));
 sg13g2_nor2_1 _10117_ (.A(net310),
    .B(_02254_),
    .Y(_02255_));
 sg13g2_buf_2 _10118_ (.A(_02255_),
    .X(_02256_));
 sg13g2_buf_1 _10119_ (.A(_02256_),
    .X(_00397_));
 sg13g2_mux2_1 _10120_ (.A0(_02246_),
    .A1(_02247_),
    .S(net21),
    .X(_00376_));
 sg13g2_buf_1 _10121_ (.A(\am_sdr0.cic0.integ_sample[10] ),
    .X(_02257_));
 sg13g2_buf_2 _10122_ (.A(\am_sdr0.cic0.integ3[10] ),
    .X(_02258_));
 sg13g2_mux2_1 _10123_ (.A0(_02257_),
    .A1(_02258_),
    .S(net21),
    .X(_00377_));
 sg13g2_buf_1 _10124_ (.A(\am_sdr0.cic0.integ_sample[11] ),
    .X(_02259_));
 sg13g2_buf_1 _10125_ (.A(\am_sdr0.cic0.integ3[11] ),
    .X(_02260_));
 sg13g2_mux2_1 _10126_ (.A0(_02259_),
    .A1(_02260_),
    .S(net21),
    .X(_00378_));
 sg13g2_inv_1 _10127_ (.Y(_02261_),
    .A(\am_sdr0.cic0.integ_sample[12] ));
 sg13g2_buf_1 _10128_ (.A(\am_sdr0.cic0.integ3[12] ),
    .X(_02262_));
 sg13g2_nand2_1 _10129_ (.Y(_02263_),
    .A(_02262_),
    .B(_02256_));
 sg13g2_o21ai_1 _10130_ (.B1(_02263_),
    .Y(_00379_),
    .A1(_02261_),
    .A2(_00397_));
 sg13g2_buf_1 _10131_ (.A(\am_sdr0.cic0.integ_sample[13] ),
    .X(_02264_));
 sg13g2_buf_1 _10132_ (.A(\am_sdr0.cic0.integ3[13] ),
    .X(_02265_));
 sg13g2_mux2_1 _10133_ (.A0(_02264_),
    .A1(_02265_),
    .S(net21),
    .X(_00380_));
 sg13g2_buf_1 _10134_ (.A(\am_sdr0.cic0.integ_sample[14] ),
    .X(_02266_));
 sg13g2_mux2_1 _10135_ (.A0(_02266_),
    .A1(\am_sdr0.cic0.integ3[14] ),
    .S(net21),
    .X(_00381_));
 sg13g2_buf_2 _10136_ (.A(\am_sdr0.cic0.integ_sample[15] ),
    .X(_02267_));
 sg13g2_buf_1 _10137_ (.A(\am_sdr0.cic0.integ3[15] ),
    .X(_02268_));
 sg13g2_buf_1 _10138_ (.A(_02256_),
    .X(_02269_));
 sg13g2_mux2_1 _10139_ (.A0(_02267_),
    .A1(_02268_),
    .S(net20),
    .X(_00382_));
 sg13g2_buf_1 _10140_ (.A(\am_sdr0.cic0.integ_sample[16] ),
    .X(_02270_));
 sg13g2_inv_1 _10141_ (.Y(_02271_),
    .A(_02270_));
 sg13g2_buf_2 _10142_ (.A(\am_sdr0.cic0.integ3[16] ),
    .X(_02272_));
 sg13g2_nand2_1 _10143_ (.Y(_02273_),
    .A(_02272_),
    .B(_02256_));
 sg13g2_o21ai_1 _10144_ (.B1(_02273_),
    .Y(_00383_),
    .A1(_02271_),
    .A2(_00397_));
 sg13g2_buf_1 _10145_ (.A(\am_sdr0.cic0.integ_sample[17] ),
    .X(_02274_));
 sg13g2_buf_2 _10146_ (.A(\am_sdr0.cic0.integ3[17] ),
    .X(_02275_));
 sg13g2_mux2_1 _10147_ (.A0(_02274_),
    .A1(_02275_),
    .S(net20),
    .X(_00384_));
 sg13g2_buf_1 _10148_ (.A(\am_sdr0.cic0.integ_sample[18] ),
    .X(_02276_));
 sg13g2_buf_1 _10149_ (.A(\am_sdr0.cic0.integ3[18] ),
    .X(_02277_));
 sg13g2_mux2_1 _10150_ (.A0(_02276_),
    .A1(_02277_),
    .S(_02269_),
    .X(_00385_));
 sg13g2_mux2_1 _10151_ (.A0(\am_sdr0.cic0.integ_sample[19] ),
    .A1(\am_sdr0.cic0.integ3[19] ),
    .S(_02269_),
    .X(_00386_));
 sg13g2_buf_2 _10152_ (.A(\am_sdr0.cic0.integ_sample[1] ),
    .X(_02278_));
 sg13g2_buf_2 _10153_ (.A(\am_sdr0.cic0.integ3[1] ),
    .X(_02279_));
 sg13g2_mux2_1 _10154_ (.A0(_02278_),
    .A1(_02279_),
    .S(net20),
    .X(_00387_));
 sg13g2_inv_1 _10155_ (.Y(_02280_),
    .A(\am_sdr0.cic0.integ_sample[2] ));
 sg13g2_buf_1 _10156_ (.A(\am_sdr0.cic0.integ3[2] ),
    .X(_02281_));
 sg13g2_nand2_1 _10157_ (.Y(_02282_),
    .A(_02281_),
    .B(_02256_));
 sg13g2_o21ai_1 _10158_ (.B1(_02282_),
    .Y(_00388_),
    .A1(_02280_),
    .A2(net21));
 sg13g2_inv_1 _10159_ (.Y(_02283_),
    .A(\am_sdr0.cic0.integ_sample[3] ));
 sg13g2_buf_1 _10160_ (.A(\am_sdr0.cic0.integ3[3] ),
    .X(_02284_));
 sg13g2_nand2_1 _10161_ (.Y(_02285_),
    .A(_02284_),
    .B(_02256_));
 sg13g2_o21ai_1 _10162_ (.B1(_02285_),
    .Y(_00389_),
    .A1(_02283_),
    .A2(net21));
 sg13g2_buf_1 _10163_ (.A(\am_sdr0.cic0.integ_sample[4] ),
    .X(_02286_));
 sg13g2_buf_1 _10164_ (.A(\am_sdr0.cic0.integ3[4] ),
    .X(_02287_));
 sg13g2_mux2_1 _10165_ (.A0(_02286_),
    .A1(_02287_),
    .S(net20),
    .X(_00390_));
 sg13g2_buf_2 _10166_ (.A(\am_sdr0.cic0.integ_sample[5] ),
    .X(_02288_));
 sg13g2_mux2_1 _10167_ (.A0(_02288_),
    .A1(\am_sdr0.cic0.integ3[5] ),
    .S(net20),
    .X(_00391_));
 sg13g2_buf_1 _10168_ (.A(\am_sdr0.cic0.integ_sample[6] ),
    .X(_02289_));
 sg13g2_buf_2 _10169_ (.A(\am_sdr0.cic0.integ3[6] ),
    .X(_02290_));
 sg13g2_mux2_1 _10170_ (.A0(_02289_),
    .A1(_02290_),
    .S(net20),
    .X(_00392_));
 sg13g2_buf_1 _10171_ (.A(\am_sdr0.cic0.integ_sample[7] ),
    .X(_02291_));
 sg13g2_buf_2 _10172_ (.A(\am_sdr0.cic0.integ3[7] ),
    .X(_02292_));
 sg13g2_mux2_1 _10173_ (.A0(_02291_),
    .A1(_02292_),
    .S(net20),
    .X(_00393_));
 sg13g2_buf_1 _10174_ (.A(\am_sdr0.cic0.integ_sample[8] ),
    .X(_02293_));
 sg13g2_buf_1 _10175_ (.A(\am_sdr0.cic0.integ3[8] ),
    .X(_02294_));
 sg13g2_mux2_1 _10176_ (.A0(_02293_),
    .A1(_02294_),
    .S(net20),
    .X(_00394_));
 sg13g2_buf_1 _10177_ (.A(\am_sdr0.cic0.integ_sample[9] ),
    .X(_02295_));
 sg13g2_buf_2 _10178_ (.A(\am_sdr0.cic0.integ3[9] ),
    .X(_02296_));
 sg13g2_mux2_1 _10179_ (.A0(_02295_),
    .A1(_02296_),
    .S(_02256_),
    .X(_00395_));
 sg13g2_buf_1 _10180_ (.A(\am_sdr0.cic1.integ3[0] ),
    .X(_02297_));
 sg13g2_buf_2 _10181_ (.A(\am_sdr0.cic1.integ_sample[0] ),
    .X(_02298_));
 sg13g2_buf_1 _10182_ (.A(\am_sdr0.cic1.count[4] ),
    .X(_02299_));
 sg13g2_inv_1 _10183_ (.Y(_02300_),
    .A(\am_sdr0.cic1.count[3] ));
 sg13g2_nand3_1 _10184_ (.B(\am_sdr0.cic1.count[0] ),
    .C(\am_sdr0.cic1.count[2] ),
    .A(\am_sdr0.cic1.count[1] ),
    .Y(_02301_));
 sg13g2_nor2_2 _10185_ (.A(_02300_),
    .B(_02301_),
    .Y(_02302_));
 sg13g2_nand3_1 _10186_ (.B(_02299_),
    .C(_02302_),
    .A(\am_sdr0.cic1.count[5] ),
    .Y(_02303_));
 sg13g2_nor3_1 _10187_ (.A(\am_sdr0.cic1.count[7] ),
    .B(\am_sdr0.cic1.count[6] ),
    .C(_02303_),
    .Y(_02304_));
 sg13g2_nand2_1 _10188_ (.Y(_02305_),
    .A(net364),
    .B(_02304_));
 sg13g2_buf_1 _10189_ (.A(_02305_),
    .X(_02306_));
 sg13g2_buf_1 _10190_ (.A(_02306_),
    .X(_02307_));
 sg13g2_mux2_1 _10191_ (.A0(_02297_),
    .A1(_02298_),
    .S(net29),
    .X(_00591_));
 sg13g2_buf_2 _10192_ (.A(\am_sdr0.cic1.integ3[10] ),
    .X(_02308_));
 sg13g2_inv_1 _10193_ (.Y(_02309_),
    .A(_02308_));
 sg13g2_buf_1 _10194_ (.A(\am_sdr0.cic1.integ_sample[10] ),
    .X(_02310_));
 sg13g2_buf_1 _10195_ (.A(_02306_),
    .X(_02311_));
 sg13g2_nand2_1 _10196_ (.Y(_02312_),
    .A(_02310_),
    .B(net28));
 sg13g2_o21ai_1 _10197_ (.B1(_02312_),
    .Y(_00592_),
    .A1(_02309_),
    .A2(_02307_));
 sg13g2_buf_1 _10198_ (.A(\am_sdr0.cic1.integ3[11] ),
    .X(_02313_));
 sg13g2_inv_1 _10199_ (.Y(_02314_),
    .A(_02313_));
 sg13g2_buf_1 _10200_ (.A(\am_sdr0.cic1.integ_sample[11] ),
    .X(_02315_));
 sg13g2_nand2_1 _10201_ (.Y(_02316_),
    .A(_02315_),
    .B(net28));
 sg13g2_o21ai_1 _10202_ (.B1(_02316_),
    .Y(_00593_),
    .A1(_02314_),
    .A2(net29));
 sg13g2_buf_1 _10203_ (.A(\am_sdr0.cic1.integ3[12] ),
    .X(_02317_));
 sg13g2_inv_1 _10204_ (.Y(_02318_),
    .A(_02317_));
 sg13g2_buf_1 _10205_ (.A(\am_sdr0.cic1.integ_sample[12] ),
    .X(_02319_));
 sg13g2_nand2_1 _10206_ (.Y(_02320_),
    .A(_02319_),
    .B(net28));
 sg13g2_o21ai_1 _10207_ (.B1(_02320_),
    .Y(_00594_),
    .A1(_02318_),
    .A2(net29));
 sg13g2_buf_1 _10208_ (.A(\am_sdr0.cic1.integ3[13] ),
    .X(_02321_));
 sg13g2_buf_2 _10209_ (.A(\am_sdr0.cic1.integ_sample[13] ),
    .X(_02322_));
 sg13g2_mux2_1 _10210_ (.A0(_02321_),
    .A1(_02322_),
    .S(_02307_),
    .X(_00595_));
 sg13g2_buf_1 _10211_ (.A(\am_sdr0.cic1.integ3[14] ),
    .X(_02323_));
 sg13g2_buf_1 _10212_ (.A(\am_sdr0.cic1.integ_sample[14] ),
    .X(_02324_));
 sg13g2_mux2_1 _10213_ (.A0(_02323_),
    .A1(_02324_),
    .S(net29),
    .X(_00596_));
 sg13g2_buf_1 _10214_ (.A(\am_sdr0.cic1.integ_sample[15] ),
    .X(_02325_));
 sg13g2_inv_1 _10215_ (.Y(_02326_),
    .A(_02325_));
 sg13g2_inv_1 _10216_ (.Y(_00612_),
    .A(_02306_));
 sg13g2_buf_1 _10217_ (.A(\am_sdr0.cic1.integ3[15] ),
    .X(_02327_));
 sg13g2_nand2_1 _10218_ (.Y(_02328_),
    .A(_02327_),
    .B(net27));
 sg13g2_o21ai_1 _10219_ (.B1(_02328_),
    .Y(_00597_),
    .A1(_02326_),
    .A2(_00612_));
 sg13g2_buf_1 _10220_ (.A(\am_sdr0.cic1.integ3[16] ),
    .X(_02329_));
 sg13g2_buf_1 _10221_ (.A(\am_sdr0.cic1.integ_sample[16] ),
    .X(_02330_));
 sg13g2_mux2_1 _10222_ (.A0(_02329_),
    .A1(_02330_),
    .S(net28),
    .X(_00598_));
 sg13g2_buf_1 _10223_ (.A(\am_sdr0.cic1.integ3[17] ),
    .X(_02331_));
 sg13g2_buf_2 _10224_ (.A(\am_sdr0.cic1.integ_sample[17] ),
    .X(_02332_));
 sg13g2_mux2_1 _10225_ (.A0(_02331_),
    .A1(_02332_),
    .S(net28),
    .X(_00599_));
 sg13g2_buf_1 _10226_ (.A(\am_sdr0.cic1.integ3[18] ),
    .X(_02333_));
 sg13g2_buf_1 _10227_ (.A(\am_sdr0.cic1.integ_sample[18] ),
    .X(_02334_));
 sg13g2_mux2_1 _10228_ (.A0(_02333_),
    .A1(_02334_),
    .S(_02311_),
    .X(_00600_));
 sg13g2_mux2_1 _10229_ (.A0(\am_sdr0.cic1.integ3[19] ),
    .A1(\am_sdr0.cic1.integ_sample[19] ),
    .S(_02311_),
    .X(_00601_));
 sg13g2_buf_1 _10230_ (.A(\am_sdr0.cic1.integ3[1] ),
    .X(_02335_));
 sg13g2_buf_2 _10231_ (.A(\am_sdr0.cic1.integ_sample[1] ),
    .X(_02336_));
 sg13g2_mux2_1 _10232_ (.A0(_02335_),
    .A1(_02336_),
    .S(net28),
    .X(_00602_));
 sg13g2_inv_1 _10233_ (.Y(_02337_),
    .A(\am_sdr0.cic1.integ_sample[2] ));
 sg13g2_buf_1 _10234_ (.A(\am_sdr0.cic1.integ3[2] ),
    .X(_02338_));
 sg13g2_nand2_1 _10235_ (.Y(_02339_),
    .A(_02338_),
    .B(net27));
 sg13g2_o21ai_1 _10236_ (.B1(_02339_),
    .Y(_00603_),
    .A1(_02337_),
    .A2(net27));
 sg13g2_inv_1 _10237_ (.Y(_02340_),
    .A(\am_sdr0.cic1.integ3[3] ));
 sg13g2_buf_1 _10238_ (.A(\am_sdr0.cic1.integ_sample[3] ),
    .X(_02341_));
 sg13g2_nand2_1 _10239_ (.Y(_02342_),
    .A(_02341_),
    .B(net28));
 sg13g2_o21ai_1 _10240_ (.B1(_02342_),
    .Y(_00604_),
    .A1(_02340_),
    .A2(net29));
 sg13g2_buf_1 _10241_ (.A(\am_sdr0.cic1.integ3[4] ),
    .X(_02343_));
 sg13g2_inv_1 _10242_ (.Y(_02344_),
    .A(_02343_));
 sg13g2_buf_1 _10243_ (.A(\am_sdr0.cic1.integ_sample[4] ),
    .X(_02345_));
 sg13g2_nand2_1 _10244_ (.Y(_02346_),
    .A(_02345_),
    .B(_02306_));
 sg13g2_o21ai_1 _10245_ (.B1(_02346_),
    .Y(_00605_),
    .A1(_02344_),
    .A2(net29));
 sg13g2_inv_1 _10246_ (.Y(_02347_),
    .A(\am_sdr0.cic1.integ3[5] ));
 sg13g2_buf_2 _10247_ (.A(\am_sdr0.cic1.integ_sample[5] ),
    .X(_02348_));
 sg13g2_nand2_1 _10248_ (.Y(_02349_),
    .A(_02348_),
    .B(_02306_));
 sg13g2_o21ai_1 _10249_ (.B1(_02349_),
    .Y(_00606_),
    .A1(_02347_),
    .A2(net29));
 sg13g2_buf_1 _10250_ (.A(\am_sdr0.cic1.integ3[6] ),
    .X(_02350_));
 sg13g2_buf_2 _10251_ (.A(\am_sdr0.cic1.integ_sample[6] ),
    .X(_02351_));
 sg13g2_mux2_1 _10252_ (.A0(_02350_),
    .A1(_02351_),
    .S(net28),
    .X(_00607_));
 sg13g2_inv_1 _10253_ (.Y(_02352_),
    .A(\am_sdr0.cic1.integ3[7] ));
 sg13g2_buf_1 _10254_ (.A(\am_sdr0.cic1.integ_sample[7] ),
    .X(_02353_));
 sg13g2_nand2_1 _10255_ (.Y(_02354_),
    .A(_02353_),
    .B(_02306_));
 sg13g2_o21ai_1 _10256_ (.B1(_02354_),
    .Y(_00608_),
    .A1(_02352_),
    .A2(net29));
 sg13g2_buf_1 _10257_ (.A(\am_sdr0.cic1.integ_sample[8] ),
    .X(_02355_));
 sg13g2_inv_1 _10258_ (.Y(_02356_),
    .A(_02355_));
 sg13g2_buf_1 _10259_ (.A(\am_sdr0.cic1.integ3[8] ),
    .X(_02357_));
 sg13g2_nand2_1 _10260_ (.Y(_02358_),
    .A(_02357_),
    .B(net27));
 sg13g2_o21ai_1 _10261_ (.B1(_02358_),
    .Y(_00609_),
    .A1(_02356_),
    .A2(net27));
 sg13g2_buf_1 _10262_ (.A(\am_sdr0.cic1.integ_sample[9] ),
    .X(_02359_));
 sg13g2_inv_1 _10263_ (.Y(_02360_),
    .A(_02359_));
 sg13g2_buf_1 _10264_ (.A(\am_sdr0.cic1.integ3[9] ),
    .X(_02361_));
 sg13g2_nand2_1 _10265_ (.Y(_02362_),
    .A(_02361_),
    .B(net27));
 sg13g2_o21ai_1 _10266_ (.B1(_02362_),
    .Y(_00610_),
    .A1(_02360_),
    .A2(net27));
 sg13g2_buf_1 _10267_ (.A(\am_sdr0.cic2.integ_sample[0] ),
    .X(_02363_));
 sg13g2_buf_1 _10268_ (.A(\am_sdr0.cic2.count[6] ),
    .X(_02364_));
 sg13g2_buf_1 _10269_ (.A(\am_sdr0.cic2.count[3] ),
    .X(_02365_));
 sg13g2_inv_1 _10270_ (.Y(_02366_),
    .A(\am_sdr0.cic2.count[2] ));
 sg13g2_nand3_1 _10271_ (.B(\am_sdr0.cic2.count[1] ),
    .C(\am_sdr0.cic2.count[0] ),
    .A(\am_sdr0.cic0.out_tick ),
    .Y(_02367_));
 sg13g2_nor2_2 _10272_ (.A(_02366_),
    .B(_02367_),
    .Y(_02368_));
 sg13g2_nand4_1 _10273_ (.B(\am_sdr0.cic2.count[5] ),
    .C(\am_sdr0.cic2.count[4] ),
    .A(_02365_),
    .Y(_02369_),
    .D(_02368_));
 sg13g2_buf_1 _10274_ (.A(_02369_),
    .X(_02370_));
 sg13g2_or4_1 _10275_ (.A(_01444_),
    .B(\am_sdr0.cic2.count[7] ),
    .C(_02364_),
    .D(_02370_),
    .X(_02371_));
 sg13g2_buf_1 _10276_ (.A(_02371_),
    .X(_02372_));
 sg13g2_buf_1 _10277_ (.A(_02372_),
    .X(_02373_));
 sg13g2_buf_1 _10278_ (.A(_02373_),
    .X(_02374_));
 sg13g2_mux2_1 _10279_ (.A0(\am_sdr0.cic2.integ3[0] ),
    .A1(_02363_),
    .S(net19),
    .X(_00806_));
 sg13g2_buf_1 _10280_ (.A(\am_sdr0.cic2.integ3[10] ),
    .X(_02375_));
 sg13g2_buf_1 _10281_ (.A(\am_sdr0.cic2.integ_sample[10] ),
    .X(_02376_));
 sg13g2_mux2_1 _10282_ (.A0(_02375_),
    .A1(_02376_),
    .S(net19),
    .X(_00807_));
 sg13g2_buf_1 _10283_ (.A(\am_sdr0.cic2.integ3[11] ),
    .X(_02377_));
 sg13g2_buf_1 _10284_ (.A(\am_sdr0.cic2.integ_sample[11] ),
    .X(_02378_));
 sg13g2_mux2_1 _10285_ (.A0(_02377_),
    .A1(_02378_),
    .S(net19),
    .X(_00808_));
 sg13g2_buf_1 _10286_ (.A(\am_sdr0.cic2.integ3[12] ),
    .X(_02379_));
 sg13g2_buf_1 _10287_ (.A(\am_sdr0.cic2.integ_sample[12] ),
    .X(_02380_));
 sg13g2_mux2_1 _10288_ (.A0(_02379_),
    .A1(_02380_),
    .S(net19),
    .X(_00809_));
 sg13g2_buf_1 _10289_ (.A(\am_sdr0.cic2.integ3[13] ),
    .X(_02381_));
 sg13g2_buf_1 _10290_ (.A(\am_sdr0.cic2.integ_sample[13] ),
    .X(_02382_));
 sg13g2_mux2_1 _10291_ (.A0(_02381_),
    .A1(_02382_),
    .S(net19),
    .X(_00810_));
 sg13g2_buf_2 _10292_ (.A(\am_sdr0.cic2.integ3[14] ),
    .X(_02383_));
 sg13g2_buf_1 _10293_ (.A(\am_sdr0.cic2.integ_sample[14] ),
    .X(_02384_));
 sg13g2_mux2_1 _10294_ (.A0(_02383_),
    .A1(_02384_),
    .S(_02374_),
    .X(_00811_));
 sg13g2_buf_2 _10295_ (.A(\am_sdr0.cic2.integ3[15] ),
    .X(_02385_));
 sg13g2_buf_1 _10296_ (.A(\am_sdr0.cic2.integ_sample[15] ),
    .X(_02386_));
 sg13g2_mux2_1 _10297_ (.A0(_02385_),
    .A1(_02386_),
    .S(net19),
    .X(_00812_));
 sg13g2_buf_1 _10298_ (.A(\am_sdr0.cic2.integ3[16] ),
    .X(_02387_));
 sg13g2_buf_1 _10299_ (.A(\am_sdr0.cic2.integ_sample[16] ),
    .X(_02388_));
 sg13g2_mux2_1 _10300_ (.A0(_02387_),
    .A1(_02388_),
    .S(net19),
    .X(_00813_));
 sg13g2_buf_1 _10301_ (.A(\am_sdr0.cic2.integ3[17] ),
    .X(_02389_));
 sg13g2_buf_1 _10302_ (.A(\am_sdr0.cic2.integ_sample[17] ),
    .X(_02390_));
 sg13g2_mux2_1 _10303_ (.A0(_02389_),
    .A1(_02390_),
    .S(net26),
    .X(_00814_));
 sg13g2_buf_1 _10304_ (.A(\am_sdr0.cic2.integ3[18] ),
    .X(_02391_));
 sg13g2_buf_1 _10305_ (.A(\am_sdr0.cic2.integ_sample[18] ),
    .X(_02392_));
 sg13g2_mux2_1 _10306_ (.A0(_02391_),
    .A1(_02392_),
    .S(net26),
    .X(_00815_));
 sg13g2_inv_1 _10307_ (.Y(_02393_),
    .A(\am_sdr0.cic2.integ3[19] ));
 sg13g2_nand2_1 _10308_ (.Y(_02394_),
    .A(\am_sdr0.cic2.integ_sample[19] ),
    .B(_02373_));
 sg13g2_o21ai_1 _10309_ (.B1(_02394_),
    .Y(_00816_),
    .A1(_02393_),
    .A2(_02374_));
 sg13g2_buf_1 _10310_ (.A(\am_sdr0.cic2.integ3[1] ),
    .X(_02395_));
 sg13g2_buf_2 _10311_ (.A(\am_sdr0.cic2.integ_sample[1] ),
    .X(_02396_));
 sg13g2_mux2_1 _10312_ (.A0(_02395_),
    .A1(_02396_),
    .S(net26),
    .X(_00817_));
 sg13g2_buf_1 _10313_ (.A(\am_sdr0.cic2.integ3[2] ),
    .X(_02397_));
 sg13g2_buf_1 _10314_ (.A(\am_sdr0.cic2.integ_sample[2] ),
    .X(_02398_));
 sg13g2_mux2_1 _10315_ (.A0(_02397_),
    .A1(_02398_),
    .S(net26),
    .X(_00818_));
 sg13g2_inv_1 _10316_ (.Y(_02399_),
    .A(\am_sdr0.cic2.integ3[3] ));
 sg13g2_buf_2 _10317_ (.A(\am_sdr0.cic2.integ_sample[3] ),
    .X(_02400_));
 sg13g2_nand2_1 _10318_ (.Y(_02401_),
    .A(_02400_),
    .B(net26));
 sg13g2_o21ai_1 _10319_ (.B1(_02401_),
    .Y(_00819_),
    .A1(_02399_),
    .A2(net19));
 sg13g2_buf_1 _10320_ (.A(\am_sdr0.cic2.integ3[4] ),
    .X(_02402_));
 sg13g2_buf_2 _10321_ (.A(\am_sdr0.cic2.integ_sample[4] ),
    .X(_02403_));
 sg13g2_mux2_1 _10322_ (.A0(_02402_),
    .A1(_02403_),
    .S(net26),
    .X(_00820_));
 sg13g2_buf_2 _10323_ (.A(\am_sdr0.cic2.integ_sample[5] ),
    .X(_02404_));
 sg13g2_inv_1 _10324_ (.Y(_02405_),
    .A(_02404_));
 sg13g2_inv_2 _10325_ (.Y(_00827_),
    .A(_02372_));
 sg13g2_buf_1 _10326_ (.A(\am_sdr0.cic2.integ3[5] ),
    .X(_02406_));
 sg13g2_nand2_1 _10327_ (.Y(_02407_),
    .A(_02406_),
    .B(_00827_));
 sg13g2_o21ai_1 _10328_ (.B1(_02407_),
    .Y(_00821_),
    .A1(_02405_),
    .A2(_00827_));
 sg13g2_buf_1 _10329_ (.A(\am_sdr0.cic2.integ3[6] ),
    .X(_02408_));
 sg13g2_buf_2 _10330_ (.A(\am_sdr0.cic2.integ_sample[6] ),
    .X(_02409_));
 sg13g2_mux2_1 _10331_ (.A0(_02408_),
    .A1(_02409_),
    .S(net26),
    .X(_00822_));
 sg13g2_buf_1 _10332_ (.A(\am_sdr0.cic2.integ_sample[7] ),
    .X(_02410_));
 sg13g2_inv_1 _10333_ (.Y(_02411_),
    .A(_02410_));
 sg13g2_buf_1 _10334_ (.A(\am_sdr0.cic2.integ3[7] ),
    .X(_02412_));
 sg13g2_nand2_1 _10335_ (.Y(_02413_),
    .A(_02412_),
    .B(_00827_));
 sg13g2_o21ai_1 _10336_ (.B1(_02413_),
    .Y(_00823_),
    .A1(_02411_),
    .A2(_00827_));
 sg13g2_buf_1 _10337_ (.A(\am_sdr0.cic2.integ3[8] ),
    .X(_02414_));
 sg13g2_buf_2 _10338_ (.A(\am_sdr0.cic2.integ_sample[8] ),
    .X(_02415_));
 sg13g2_mux2_1 _10339_ (.A0(_02414_),
    .A1(_02415_),
    .S(net26),
    .X(_00824_));
 sg13g2_buf_1 _10340_ (.A(\am_sdr0.cic2.integ_sample[9] ),
    .X(_02416_));
 sg13g2_inv_1 _10341_ (.Y(_02417_),
    .A(_02416_));
 sg13g2_buf_1 _10342_ (.A(\am_sdr0.cic2.integ3[9] ),
    .X(_02418_));
 sg13g2_nand2_1 _10343_ (.Y(_02419_),
    .A(_02418_),
    .B(_00827_));
 sg13g2_o21ai_1 _10344_ (.B1(_02419_),
    .Y(_00825_),
    .A1(_02417_),
    .A2(_00827_));
 sg13g2_buf_1 _10345_ (.A(\am_sdr0.cic3.integ3[0] ),
    .X(_02420_));
 sg13g2_buf_2 _10346_ (.A(\am_sdr0.cic3.integ_sample[0] ),
    .X(_02421_));
 sg13g2_buf_1 _10347_ (.A(\am_sdr0.cic3.count[6] ),
    .X(_02422_));
 sg13g2_buf_1 _10348_ (.A(\am_sdr0.cic3.count[3] ),
    .X(_02423_));
 sg13g2_inv_1 _10349_ (.Y(_02424_),
    .A(\am_sdr0.cic3.count[2] ));
 sg13g2_buf_1 _10350_ (.A(\am_sdr0.cic1.out_tick ),
    .X(_02425_));
 sg13g2_nand3_1 _10351_ (.B(\am_sdr0.cic3.count[0] ),
    .C(_02425_),
    .A(\am_sdr0.cic3.count[1] ),
    .Y(_02426_));
 sg13g2_nor2_2 _10352_ (.A(_02424_),
    .B(_02426_),
    .Y(_02427_));
 sg13g2_nand4_1 _10353_ (.B(\am_sdr0.cic3.count[5] ),
    .C(\am_sdr0.cic3.count[4] ),
    .A(_02423_),
    .Y(_02428_),
    .D(_02427_));
 sg13g2_buf_1 _10354_ (.A(_02428_),
    .X(_02429_));
 sg13g2_or4_1 _10355_ (.A(net310),
    .B(\am_sdr0.cic3.count[7] ),
    .C(_02422_),
    .D(_02429_),
    .X(_02430_));
 sg13g2_buf_1 _10356_ (.A(_02430_),
    .X(_02431_));
 sg13g2_buf_1 _10357_ (.A(_02431_),
    .X(_02432_));
 sg13g2_mux2_1 _10358_ (.A0(_02420_),
    .A1(_02421_),
    .S(net18),
    .X(_01021_));
 sg13g2_buf_1 _10359_ (.A(\am_sdr0.cic3.integ_sample[10] ),
    .X(_02433_));
 sg13g2_inv_1 _10360_ (.Y(_02434_),
    .A(_02433_));
 sg13g2_inv_1 _10361_ (.Y(_02435_),
    .A(_02431_));
 sg13g2_buf_1 _10362_ (.A(_02435_),
    .X(_01041_));
 sg13g2_buf_1 _10363_ (.A(\am_sdr0.cic3.integ3[10] ),
    .X(_02436_));
 sg13g2_nand2_1 _10364_ (.Y(_02437_),
    .A(_02436_),
    .B(net11));
 sg13g2_o21ai_1 _10365_ (.B1(_02437_),
    .Y(_01022_),
    .A1(_02434_),
    .A2(net11));
 sg13g2_buf_2 _10366_ (.A(\am_sdr0.cic3.integ3[11] ),
    .X(_02438_));
 sg13g2_buf_1 _10367_ (.A(\am_sdr0.cic3.integ_sample[11] ),
    .X(_02439_));
 sg13g2_mux2_1 _10368_ (.A0(_02438_),
    .A1(_02439_),
    .S(net18),
    .X(_01023_));
 sg13g2_buf_2 _10369_ (.A(\am_sdr0.cic3.integ3[12] ),
    .X(_02440_));
 sg13g2_buf_1 _10370_ (.A(\am_sdr0.cic3.integ_sample[12] ),
    .X(_02441_));
 sg13g2_mux2_1 _10371_ (.A0(_02440_),
    .A1(_02441_),
    .S(net18),
    .X(_01024_));
 sg13g2_buf_1 _10372_ (.A(\am_sdr0.cic3.integ_sample[13] ),
    .X(_02442_));
 sg13g2_inv_1 _10373_ (.Y(_02443_),
    .A(_02442_));
 sg13g2_buf_1 _10374_ (.A(\am_sdr0.cic3.integ3[13] ),
    .X(_02444_));
 sg13g2_nand2_1 _10375_ (.Y(_02445_),
    .A(_02444_),
    .B(_01041_));
 sg13g2_o21ai_1 _10376_ (.B1(_02445_),
    .Y(_01025_),
    .A1(_02443_),
    .A2(_01041_));
 sg13g2_buf_1 _10377_ (.A(\am_sdr0.cic3.integ3[14] ),
    .X(_02446_));
 sg13g2_inv_1 _10378_ (.Y(_02447_),
    .A(_02446_));
 sg13g2_buf_1 _10379_ (.A(\am_sdr0.cic3.integ_sample[14] ),
    .X(_02448_));
 sg13g2_buf_1 _10380_ (.A(_02431_),
    .X(_02449_));
 sg13g2_nand2_1 _10381_ (.Y(_02450_),
    .A(_02448_),
    .B(net17));
 sg13g2_o21ai_1 _10382_ (.B1(_02450_),
    .Y(_01026_),
    .A1(_02447_),
    .A2(net18));
 sg13g2_buf_1 _10383_ (.A(\am_sdr0.cic3.integ3[15] ),
    .X(_02451_));
 sg13g2_buf_2 _10384_ (.A(\am_sdr0.cic3.integ_sample[15] ),
    .X(_02452_));
 sg13g2_mux2_1 _10385_ (.A0(_02451_),
    .A1(_02452_),
    .S(net18),
    .X(_01027_));
 sg13g2_inv_1 _10386_ (.Y(_02453_),
    .A(\am_sdr0.cic3.integ3[16] ));
 sg13g2_buf_1 _10387_ (.A(\am_sdr0.cic3.integ_sample[16] ),
    .X(_02454_));
 sg13g2_nand2_1 _10388_ (.Y(_02455_),
    .A(_02454_),
    .B(net17));
 sg13g2_o21ai_1 _10389_ (.B1(_02455_),
    .Y(_01028_),
    .A1(_02453_),
    .A2(net18));
 sg13g2_buf_1 _10390_ (.A(\am_sdr0.cic3.integ3[17] ),
    .X(_02456_));
 sg13g2_inv_1 _10391_ (.Y(_02457_),
    .A(_02456_));
 sg13g2_buf_1 _10392_ (.A(\am_sdr0.cic3.integ_sample[17] ),
    .X(_02458_));
 sg13g2_nand2_1 _10393_ (.Y(_02459_),
    .A(_02458_),
    .B(_02449_));
 sg13g2_o21ai_1 _10394_ (.B1(_02459_),
    .Y(_01029_),
    .A1(_02457_),
    .A2(_02432_));
 sg13g2_buf_1 _10395_ (.A(\am_sdr0.cic3.integ3[18] ),
    .X(_02460_));
 sg13g2_buf_1 _10396_ (.A(\am_sdr0.cic3.integ_sample[18] ),
    .X(_02461_));
 sg13g2_mux2_1 _10397_ (.A0(_02460_),
    .A1(_02461_),
    .S(_02432_),
    .X(_01030_));
 sg13g2_mux2_1 _10398_ (.A0(\am_sdr0.cic3.integ3[19] ),
    .A1(\am_sdr0.cic3.integ_sample[19] ),
    .S(_02449_),
    .X(_01031_));
 sg13g2_buf_1 _10399_ (.A(\am_sdr0.cic3.integ3[1] ),
    .X(_02462_));
 sg13g2_buf_2 _10400_ (.A(\am_sdr0.cic3.integ_sample[1] ),
    .X(_02463_));
 sg13g2_mux2_1 _10401_ (.A0(_02462_),
    .A1(_02463_),
    .S(net17),
    .X(_01032_));
 sg13g2_inv_1 _10402_ (.Y(_02464_),
    .A(\am_sdr0.cic3.integ_sample[2] ));
 sg13g2_buf_1 _10403_ (.A(\am_sdr0.cic3.integ3[2] ),
    .X(_02465_));
 sg13g2_nand2_1 _10404_ (.Y(_02466_),
    .A(_02465_),
    .B(net11));
 sg13g2_o21ai_1 _10405_ (.B1(_02466_),
    .Y(_01033_),
    .A1(_02464_),
    .A2(net11));
 sg13g2_inv_1 _10406_ (.Y(_02467_),
    .A(\am_sdr0.cic3.integ3[3] ));
 sg13g2_buf_1 _10407_ (.A(\am_sdr0.cic3.integ_sample[3] ),
    .X(_02468_));
 sg13g2_nand2_1 _10408_ (.Y(_02469_),
    .A(_02468_),
    .B(net17));
 sg13g2_o21ai_1 _10409_ (.B1(_02469_),
    .Y(_01034_),
    .A1(_02467_),
    .A2(net18));
 sg13g2_buf_1 _10410_ (.A(\am_sdr0.cic3.integ3[4] ),
    .X(_02470_));
 sg13g2_buf_1 _10411_ (.A(\am_sdr0.cic3.integ_sample[4] ),
    .X(_02471_));
 sg13g2_mux2_1 _10412_ (.A0(_02470_),
    .A1(_02471_),
    .S(net17),
    .X(_01035_));
 sg13g2_inv_1 _10413_ (.Y(_02472_),
    .A(\am_sdr0.cic3.integ3[5] ));
 sg13g2_buf_2 _10414_ (.A(\am_sdr0.cic3.integ_sample[5] ),
    .X(_02473_));
 sg13g2_nand2_1 _10415_ (.Y(_02474_),
    .A(_02473_),
    .B(net17));
 sg13g2_o21ai_1 _10416_ (.B1(_02474_),
    .Y(_01036_),
    .A1(_02472_),
    .A2(net18));
 sg13g2_buf_1 _10417_ (.A(\am_sdr0.cic3.integ3[6] ),
    .X(_02475_));
 sg13g2_buf_2 _10418_ (.A(\am_sdr0.cic3.integ_sample[6] ),
    .X(_02476_));
 sg13g2_mux2_1 _10419_ (.A0(_02475_),
    .A1(_02476_),
    .S(net17),
    .X(_01037_));
 sg13g2_buf_2 _10420_ (.A(\am_sdr0.cic3.integ3[7] ),
    .X(_02477_));
 sg13g2_buf_1 _10421_ (.A(\am_sdr0.cic3.integ_sample[7] ),
    .X(_02478_));
 sg13g2_mux2_1 _10422_ (.A0(_02477_),
    .A1(_02478_),
    .S(net17),
    .X(_01038_));
 sg13g2_buf_1 _10423_ (.A(\am_sdr0.cic3.integ_sample[8] ),
    .X(_02479_));
 sg13g2_inv_1 _10424_ (.Y(_02480_),
    .A(_02479_));
 sg13g2_buf_2 _10425_ (.A(\am_sdr0.cic3.integ3[8] ),
    .X(_02481_));
 sg13g2_nand2_1 _10426_ (.Y(_02482_),
    .A(_02481_),
    .B(net11));
 sg13g2_o21ai_1 _10427_ (.B1(_02482_),
    .Y(_01039_),
    .A1(_02480_),
    .A2(net11));
 sg13g2_buf_1 _10428_ (.A(\am_sdr0.cic3.integ_sample[9] ),
    .X(_02483_));
 sg13g2_inv_1 _10429_ (.Y(_02484_),
    .A(_02483_));
 sg13g2_buf_2 _10430_ (.A(\am_sdr0.cic3.integ3[9] ),
    .X(_02485_));
 sg13g2_nand2_1 _10431_ (.Y(_02486_),
    .A(_02485_),
    .B(_02435_));
 sg13g2_o21ai_1 _10432_ (.B1(_02486_),
    .Y(_01040_),
    .A1(_02484_),
    .A2(net11));
 sg13g2_inv_1 _10433_ (.Y(_02487_),
    .A(\am_sdr0.spi0.shift_reg[0] ));
 sg13g2_buf_1 _10434_ (.A(\am_sdr0.spi0.state[0] ),
    .X(_02488_));
 sg13g2_nand3b_1 _10435_ (.B(_02488_),
    .C(\am_sdr0.spi0.SCK_qq ),
    .Y(_02489_),
    .A_N(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_inv_1 _10436_ (.Y(_02490_),
    .A(\am_sdr0.spi0.CS_qq ));
 sg13g2_nand3b_1 _10437_ (.B(\am_sdr0.spi0.CS_qqq ),
    .C(_02490_),
    .Y(_02491_),
    .A_N(_02488_));
 sg13g2_buf_1 _10438_ (.A(\am_sdr0.spi0.state[1] ),
    .X(_02492_));
 sg13g2_nand2b_1 _10439_ (.Y(_02493_),
    .B(net364),
    .A_N(_02492_));
 sg13g2_a21oi_1 _10440_ (.A1(_02489_),
    .A2(_02491_),
    .Y(_02494_),
    .B1(_02493_));
 sg13g2_buf_1 _10441_ (.A(_02494_),
    .X(_02495_));
 sg13g2_buf_1 _10442_ (.A(_02495_),
    .X(_02496_));
 sg13g2_buf_1 _10443_ (.A(_02496_),
    .X(_02497_));
 sg13g2_buf_1 _10444_ (.A(_02495_),
    .X(_02498_));
 sg13g2_nor2b_1 _10445_ (.A(_02492_),
    .B_N(_02488_),
    .Y(_02499_));
 sg13g2_buf_1 _10446_ (.A(_02499_),
    .X(_02500_));
 sg13g2_buf_1 _10447_ (.A(_02500_),
    .X(_02501_));
 sg13g2_nand3_1 _10448_ (.B(net134),
    .C(net184),
    .A(\am_sdr0.spi0.MOSI_qq ),
    .Y(_02502_));
 sg13g2_o21ai_1 _10449_ (.B1(_02502_),
    .Y(_01141_),
    .A1(_02487_),
    .A2(net35));
 sg13g2_inv_1 _10450_ (.Y(_02503_),
    .A(\am_sdr0.spi0.shift_reg[10] ));
 sg13g2_buf_1 _10451_ (.A(_02495_),
    .X(_02504_));
 sg13g2_nand3_1 _10452_ (.B(_02504_),
    .C(_02501_),
    .A(\am_sdr0.spi0.shift_reg[9] ),
    .Y(_02505_));
 sg13g2_o21ai_1 _10453_ (.B1(_02505_),
    .Y(_01142_),
    .A1(_02503_),
    .A2(net35));
 sg13g2_inv_1 _10454_ (.Y(_02506_),
    .A(\am_sdr0.spi0.shift_reg[11] ));
 sg13g2_nand3_1 _10455_ (.B(_02504_),
    .C(_02501_),
    .A(\am_sdr0.spi0.shift_reg[10] ),
    .Y(_02507_));
 sg13g2_o21ai_1 _10456_ (.B1(_02507_),
    .Y(_01143_),
    .A1(_02506_),
    .A2(_02497_));
 sg13g2_inv_1 _10457_ (.Y(_02508_),
    .A(\am_sdr0.spi0.shift_reg[12] ));
 sg13g2_nand3_1 _10458_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[11] ),
    .Y(_02509_));
 sg13g2_o21ai_1 _10459_ (.B1(_02509_),
    .Y(_01144_),
    .A1(_02508_),
    .A2(_02497_));
 sg13g2_inv_1 _10460_ (.Y(_02510_),
    .A(\am_sdr0.spi0.shift_reg[13] ));
 sg13g2_nand3_1 _10461_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[12] ),
    .Y(_02511_));
 sg13g2_o21ai_1 _10462_ (.B1(_02511_),
    .Y(_01145_),
    .A1(_02510_),
    .A2(net35));
 sg13g2_inv_1 _10463_ (.Y(_02512_),
    .A(\am_sdr0.spi0.shift_reg[14] ));
 sg13g2_nand3_1 _10464_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[13] ),
    .Y(_02513_));
 sg13g2_o21ai_1 _10465_ (.B1(_02513_),
    .Y(_01146_),
    .A1(_02512_),
    .A2(net35));
 sg13g2_inv_1 _10466_ (.Y(_02514_),
    .A(\am_sdr0.spi0.shift_reg[15] ));
 sg13g2_nand3_1 _10467_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[14] ),
    .Y(_02515_));
 sg13g2_o21ai_1 _10468_ (.B1(_02515_),
    .Y(_01147_),
    .A1(_02514_),
    .A2(net35));
 sg13g2_inv_1 _10469_ (.Y(_02516_),
    .A(\am_sdr0.spi0.shift_reg[16] ));
 sg13g2_nand3_1 _10470_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[15] ),
    .Y(_02517_));
 sg13g2_o21ai_1 _10471_ (.B1(_02517_),
    .Y(_01148_),
    .A1(_02516_),
    .A2(net35));
 sg13g2_inv_1 _10472_ (.Y(_02518_),
    .A(\am_sdr0.spi0.shift_reg[17] ));
 sg13g2_nand3_1 _10473_ (.B(net133),
    .C(net184),
    .A(\am_sdr0.spi0.shift_reg[16] ),
    .Y(_02519_));
 sg13g2_o21ai_1 _10474_ (.B1(_02519_),
    .Y(_01149_),
    .A1(_02518_),
    .A2(net35));
 sg13g2_inv_1 _10475_ (.Y(_02520_),
    .A(\am_sdr0.spi0.shift_reg[18] ));
 sg13g2_buf_1 _10476_ (.A(_02500_),
    .X(_02521_));
 sg13g2_nand3_1 _10477_ (.B(net133),
    .C(_02521_),
    .A(\am_sdr0.spi0.shift_reg[17] ),
    .Y(_02522_));
 sg13g2_o21ai_1 _10478_ (.B1(_02522_),
    .Y(_01150_),
    .A1(_02520_),
    .A2(net35));
 sg13g2_inv_1 _10479_ (.Y(_02523_),
    .A(\am_sdr0.spi0.shift_reg[19] ));
 sg13g2_buf_1 _10480_ (.A(net135),
    .X(_02524_));
 sg13g2_nand3_1 _10481_ (.B(net133),
    .C(_02521_),
    .A(\am_sdr0.spi0.shift_reg[18] ),
    .Y(_02525_));
 sg13g2_o21ai_1 _10482_ (.B1(_02525_),
    .Y(_01151_),
    .A1(_02523_),
    .A2(net34));
 sg13g2_inv_1 _10483_ (.Y(_02526_),
    .A(\am_sdr0.spi0.shift_reg[1] ));
 sg13g2_buf_1 _10484_ (.A(_02495_),
    .X(_02527_));
 sg13g2_nand3_1 _10485_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[0] ),
    .Y(_02528_));
 sg13g2_o21ai_1 _10486_ (.B1(_02528_),
    .Y(_01152_),
    .A1(_02526_),
    .A2(net34));
 sg13g2_inv_1 _10487_ (.Y(_02529_),
    .A(\am_sdr0.spi0.shift_reg[20] ));
 sg13g2_nand3_1 _10488_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[19] ),
    .Y(_02530_));
 sg13g2_o21ai_1 _10489_ (.B1(_02530_),
    .Y(_01153_),
    .A1(_02529_),
    .A2(_02524_));
 sg13g2_inv_1 _10490_ (.Y(_02531_),
    .A(\am_sdr0.spi0.shift_reg[21] ));
 sg13g2_nand3_1 _10491_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[20] ),
    .Y(_02532_));
 sg13g2_o21ai_1 _10492_ (.B1(_02532_),
    .Y(_01154_),
    .A1(_02531_),
    .A2(_02524_));
 sg13g2_inv_1 _10493_ (.Y(_02533_),
    .A(\am_sdr0.spi0.shift_reg[22] ));
 sg13g2_nand3_1 _10494_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[21] ),
    .Y(_02534_));
 sg13g2_o21ai_1 _10495_ (.B1(_02534_),
    .Y(_01155_),
    .A1(_02533_),
    .A2(net34));
 sg13g2_inv_1 _10496_ (.Y(_02535_),
    .A(\am_sdr0.spi0.shift_reg[23] ));
 sg13g2_nand3_1 _10497_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[22] ),
    .Y(_02536_));
 sg13g2_o21ai_1 _10498_ (.B1(_02536_),
    .Y(_01156_),
    .A1(_02535_),
    .A2(net34));
 sg13g2_inv_1 _10499_ (.Y(_02537_),
    .A(\am_sdr0.spi0.shift_reg[24] ));
 sg13g2_nand3_1 _10500_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[23] ),
    .Y(_02538_));
 sg13g2_o21ai_1 _10501_ (.B1(_02538_),
    .Y(_01157_),
    .A1(_02537_),
    .A2(net34));
 sg13g2_inv_1 _10502_ (.Y(_02539_),
    .A(\am_sdr0.spi0.shift_reg[25] ));
 sg13g2_nand3_1 _10503_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[24] ),
    .Y(_02540_));
 sg13g2_o21ai_1 _10504_ (.B1(_02540_),
    .Y(_01158_),
    .A1(_02539_),
    .A2(net34));
 sg13g2_inv_1 _10505_ (.Y(_02541_),
    .A(\am_sdr0.spi0.shift_reg[26] ));
 sg13g2_nand3_1 _10506_ (.B(net132),
    .C(net183),
    .A(\am_sdr0.spi0.shift_reg[25] ),
    .Y(_02542_));
 sg13g2_o21ai_1 _10507_ (.B1(_02542_),
    .Y(_01159_),
    .A1(_02541_),
    .A2(net34));
 sg13g2_inv_1 _10508_ (.Y(_02543_),
    .A(\am_sdr0.spi0.shift_reg[27] ));
 sg13g2_buf_1 _10509_ (.A(_02500_),
    .X(_02544_));
 sg13g2_nand3_1 _10510_ (.B(_02527_),
    .C(_02544_),
    .A(\am_sdr0.spi0.shift_reg[26] ),
    .Y(_02545_));
 sg13g2_o21ai_1 _10511_ (.B1(_02545_),
    .Y(_01160_),
    .A1(_02543_),
    .A2(net34));
 sg13g2_inv_1 _10512_ (.Y(_02546_),
    .A(\am_sdr0.spi0.shift_reg[28] ));
 sg13g2_nand3_1 _10513_ (.B(_02527_),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[27] ),
    .Y(_02547_));
 sg13g2_o21ai_1 _10514_ (.B1(_02547_),
    .Y(_01161_),
    .A1(_02546_),
    .A2(net134));
 sg13g2_inv_1 _10515_ (.Y(_02548_),
    .A(\am_sdr0.spi0.shift_reg[2] ));
 sg13g2_nand3_1 _10516_ (.B(_02496_),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[1] ),
    .Y(_02549_));
 sg13g2_o21ai_1 _10517_ (.B1(_02549_),
    .Y(_01162_),
    .A1(_02548_),
    .A2(net134));
 sg13g2_inv_1 _10518_ (.Y(_02550_),
    .A(\am_sdr0.spi0.shift_reg[3] ));
 sg13g2_nand3_1 _10519_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[2] ),
    .Y(_02551_));
 sg13g2_o21ai_1 _10520_ (.B1(_02551_),
    .Y(_01163_),
    .A1(_02550_),
    .A2(net134));
 sg13g2_inv_1 _10521_ (.Y(_02552_),
    .A(\am_sdr0.spi0.shift_reg[4] ));
 sg13g2_nand3_1 _10522_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[3] ),
    .Y(_02553_));
 sg13g2_o21ai_1 _10523_ (.B1(_02553_),
    .Y(_01164_),
    .A1(_02552_),
    .A2(net134));
 sg13g2_inv_1 _10524_ (.Y(_02554_),
    .A(\am_sdr0.spi0.shift_reg[5] ));
 sg13g2_nand3_1 _10525_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[4] ),
    .Y(_02555_));
 sg13g2_o21ai_1 _10526_ (.B1(_02555_),
    .Y(_01165_),
    .A1(_02554_),
    .A2(net134));
 sg13g2_inv_1 _10527_ (.Y(_02556_),
    .A(\am_sdr0.spi0.shift_reg[6] ));
 sg13g2_nand3_1 _10528_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[5] ),
    .Y(_02557_));
 sg13g2_o21ai_1 _10529_ (.B1(_02557_),
    .Y(_01166_),
    .A1(_02556_),
    .A2(net134));
 sg13g2_inv_1 _10530_ (.Y(_02558_),
    .A(\am_sdr0.spi0.shift_reg[7] ));
 sg13g2_nand3_1 _10531_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[6] ),
    .Y(_02559_));
 sg13g2_o21ai_1 _10532_ (.B1(_02559_),
    .Y(_01167_),
    .A1(_02558_),
    .A2(net134));
 sg13g2_inv_1 _10533_ (.Y(_02560_),
    .A(\am_sdr0.spi0.shift_reg[8] ));
 sg13g2_nand3_1 _10534_ (.B(net135),
    .C(_02544_),
    .A(\am_sdr0.spi0.shift_reg[7] ),
    .Y(_02561_));
 sg13g2_o21ai_1 _10535_ (.B1(_02561_),
    .Y(_01168_),
    .A1(_02560_),
    .A2(_02498_));
 sg13g2_inv_1 _10536_ (.Y(_02562_),
    .A(\am_sdr0.spi0.shift_reg[9] ));
 sg13g2_nand3_1 _10537_ (.B(net135),
    .C(net182),
    .A(\am_sdr0.spi0.shift_reg[8] ),
    .Y(_02563_));
 sg13g2_o21ai_1 _10538_ (.B1(_02563_),
    .Y(_01169_),
    .A1(_02562_),
    .A2(_02498_));
 sg13g2_and3_1 _10539_ (.X(_00299_),
    .A(net257),
    .B(_00072_),
    .C(_02254_));
 sg13g2_nand2_1 _10540_ (.Y(_02564_),
    .A(net301),
    .B(_02254_));
 sg13g2_xnor2_1 _10541_ (.Y(_02565_),
    .A(\am_sdr0.cic0.count[1] ),
    .B(\am_sdr0.cic0.count[0] ));
 sg13g2_nor2_1 _10542_ (.A(_02564_),
    .B(_02565_),
    .Y(_00300_));
 sg13g2_nand2_1 _10543_ (.Y(_02566_),
    .A(\am_sdr0.cic0.count[1] ),
    .B(\am_sdr0.cic0.count[0] ));
 sg13g2_xor2_1 _10544_ (.B(_02566_),
    .A(\am_sdr0.cic0.count[2] ),
    .X(_02567_));
 sg13g2_nor2_1 _10545_ (.A(_02564_),
    .B(_02567_),
    .Y(_00301_));
 sg13g2_xnor2_1 _10546_ (.Y(_02568_),
    .A(_02249_),
    .B(_02250_));
 sg13g2_nor2_1 _10547_ (.A(_02564_),
    .B(_02568_),
    .Y(_00302_));
 sg13g2_xnor2_1 _10548_ (.Y(_02569_),
    .A(_02248_),
    .B(_02251_));
 sg13g2_nor2_1 _10549_ (.A(net139),
    .B(_02569_),
    .Y(_00303_));
 sg13g2_nand2_1 _10550_ (.Y(_02570_),
    .A(_02248_),
    .B(_02251_));
 sg13g2_xor2_1 _10551_ (.B(_02570_),
    .A(\am_sdr0.cic0.count[5] ),
    .X(_02571_));
 sg13g2_nor2_1 _10552_ (.A(net139),
    .B(_02571_),
    .Y(_00304_));
 sg13g2_xor2_1 _10553_ (.B(_02252_),
    .A(\am_sdr0.cic0.count[6] ),
    .X(_02572_));
 sg13g2_nor2_1 _10554_ (.A(_02564_),
    .B(_02572_),
    .Y(_00305_));
 sg13g2_nand4_1 _10555_ (.B(_02248_),
    .C(\am_sdr0.cic0.count[6] ),
    .A(\am_sdr0.cic0.count[5] ),
    .Y(_02573_),
    .D(_02251_));
 sg13g2_xor2_1 _10556_ (.B(_02573_),
    .A(\am_sdr0.cic0.count[7] ),
    .X(_02574_));
 sg13g2_nor2_1 _10557_ (.A(net139),
    .B(_02574_),
    .Y(_00306_));
 sg13g2_inv_1 _10558_ (.Y(_02575_),
    .A(_00073_));
 sg13g2_nand2b_1 _10559_ (.Y(_02576_),
    .B(net303),
    .A_N(_02304_));
 sg13g2_buf_1 _10560_ (.A(_02576_),
    .X(_02577_));
 sg13g2_nor2_1 _10561_ (.A(_02575_),
    .B(_02577_),
    .Y(_00514_));
 sg13g2_xnor2_1 _10562_ (.Y(_02578_),
    .A(\am_sdr0.cic1.count[1] ),
    .B(\am_sdr0.cic1.count[0] ));
 sg13g2_nor2_1 _10563_ (.A(_02577_),
    .B(_02578_),
    .Y(_00515_));
 sg13g2_nand2_1 _10564_ (.Y(_02579_),
    .A(\am_sdr0.cic1.count[1] ),
    .B(\am_sdr0.cic1.count[0] ));
 sg13g2_xor2_1 _10565_ (.B(_02579_),
    .A(\am_sdr0.cic1.count[2] ),
    .X(_02580_));
 sg13g2_nor2_1 _10566_ (.A(_02577_),
    .B(_02580_),
    .Y(_00516_));
 sg13g2_xnor2_1 _10567_ (.Y(_02581_),
    .A(_02300_),
    .B(_02301_));
 sg13g2_nor2_1 _10568_ (.A(net139),
    .B(_02581_),
    .Y(_00517_));
 sg13g2_xnor2_1 _10569_ (.Y(_02582_),
    .A(_02299_),
    .B(_02302_));
 sg13g2_nor2_1 _10570_ (.A(net139),
    .B(_02582_),
    .Y(_00518_));
 sg13g2_nand2_1 _10571_ (.Y(_02583_),
    .A(_02299_),
    .B(_02302_));
 sg13g2_xor2_1 _10572_ (.B(_02583_),
    .A(\am_sdr0.cic1.count[5] ),
    .X(_02584_));
 sg13g2_nor2_1 _10573_ (.A(net139),
    .B(_02584_),
    .Y(_00519_));
 sg13g2_xor2_1 _10574_ (.B(_02303_),
    .A(\am_sdr0.cic1.count[6] ),
    .X(_02585_));
 sg13g2_nor2_1 _10575_ (.A(_02577_),
    .B(_02585_),
    .Y(_00520_));
 sg13g2_nand4_1 _10576_ (.B(_02299_),
    .C(\am_sdr0.cic1.count[6] ),
    .A(\am_sdr0.cic1.count[5] ),
    .Y(_02586_),
    .D(_02302_));
 sg13g2_xor2_1 _10577_ (.B(_02586_),
    .A(\am_sdr0.cic1.count[7] ),
    .X(_02587_));
 sg13g2_nor2_1 _10578_ (.A(net139),
    .B(_02587_),
    .Y(_00521_));
 sg13g2_buf_1 _10579_ (.A(\am_sdr0.gain_spi[0] ),
    .X(_02588_));
 sg13g2_buf_2 _10580_ (.A(\am_sdr0.am0.demod_out[13] ),
    .X(_02589_));
 sg13g2_buf_1 _10581_ (.A(\am_sdr0.count[6] ),
    .X(_02590_));
 sg13g2_buf_1 _10582_ (.A(\am_sdr0.am0.demod_out[12] ),
    .X(_02591_));
 sg13g2_inv_1 _10583_ (.Y(_02592_),
    .A(_02591_));
 sg13g2_inv_2 _10584_ (.Y(_02593_),
    .A(_02590_));
 sg13g2_buf_2 _10585_ (.A(\am_sdr0.am0.demod_out[10] ),
    .X(_02594_));
 sg13g2_inv_2 _10586_ (.Y(_02595_),
    .A(_02594_));
 sg13g2_buf_1 _10587_ (.A(\am_sdr0.count[4] ),
    .X(_02596_));
 sg13g2_buf_1 _10588_ (.A(_02596_),
    .X(_02597_));
 sg13g2_inv_1 _10589_ (.Y(_02598_),
    .A(_02596_));
 sg13g2_buf_1 _10590_ (.A(\am_sdr0.am0.demod_out[8] ),
    .X(_02599_));
 sg13g2_inv_1 _10591_ (.Y(_02600_),
    .A(_02599_));
 sg13g2_buf_2 _10592_ (.A(\am_sdr0.count[2] ),
    .X(_02601_));
 sg13g2_buf_1 _10593_ (.A(\am_sdr0.count[3] ),
    .X(_02602_));
 sg13g2_o21ai_1 _10594_ (.B1(_02602_),
    .Y(_02603_),
    .A1(_02600_),
    .A2(_02601_));
 sg13g2_buf_1 _10595_ (.A(\am_sdr0.am0.demod_out[9] ),
    .X(_02604_));
 sg13g2_inv_1 _10596_ (.Y(_02605_),
    .A(_02602_));
 sg13g2_nand2_1 _10597_ (.Y(_02606_),
    .A(_02599_),
    .B(_02605_));
 sg13g2_nor2_1 _10598_ (.A(_02601_),
    .B(_02606_),
    .Y(_02607_));
 sg13g2_a221oi_1 _10599_ (.B2(_02604_),
    .C1(_02607_),
    .B1(_02603_),
    .A1(_02594_),
    .Y(_02608_),
    .A2(_02598_));
 sg13g2_a21oi_1 _10600_ (.A1(_02595_),
    .A2(_02597_),
    .Y(_02609_),
    .B1(_02608_));
 sg13g2_buf_2 _10601_ (.A(\am_sdr0.am0.demod_out[11] ),
    .X(_02610_));
 sg13g2_buf_1 _10602_ (.A(\am_sdr0.count[5] ),
    .X(_02611_));
 sg13g2_nor2_1 _10603_ (.A(_02610_),
    .B(_02609_),
    .Y(_02612_));
 sg13g2_nor2_1 _10604_ (.A(_02611_),
    .B(_02612_),
    .Y(_02613_));
 sg13g2_a221oi_1 _10605_ (.B2(_02610_),
    .C1(_02613_),
    .B1(_02609_),
    .A1(_02593_),
    .Y(_02614_),
    .A2(_02591_));
 sg13g2_a21oi_1 _10606_ (.A1(_02590_),
    .A2(_02592_),
    .Y(_02615_),
    .B1(_02614_));
 sg13g2_buf_1 _10607_ (.A(\am_sdr0.count[7] ),
    .X(_02616_));
 sg13g2_inv_1 _10608_ (.Y(_02617_),
    .A(_02616_));
 sg13g2_a21oi_1 _10609_ (.A1(_02589_),
    .A2(_02615_),
    .Y(_02618_),
    .B1(_02617_));
 sg13g2_buf_2 _10610_ (.A(\am_sdr0.gain_spi[1] ),
    .X(_02619_));
 sg13g2_o21ai_1 _10611_ (.B1(_02619_),
    .Y(_02620_),
    .A1(_02589_),
    .A2(_02615_));
 sg13g2_nor3_1 _10612_ (.A(_02588_),
    .B(_02618_),
    .C(_02620_),
    .Y(_02621_));
 sg13g2_inv_1 _10613_ (.Y(_02622_),
    .A(_02588_));
 sg13g2_buf_1 _10614_ (.A(\am_sdr0.am0.demod_out[14] ),
    .X(_02623_));
 sg13g2_inv_1 _10615_ (.Y(_02624_),
    .A(_02589_));
 sg13g2_inv_1 _10616_ (.Y(_02625_),
    .A(_02611_));
 sg13g2_buf_1 _10617_ (.A(\am_sdr0.count[1] ),
    .X(_02626_));
 sg13g2_nand2b_1 _10618_ (.Y(_02627_),
    .B(_02599_),
    .A_N(_02626_));
 sg13g2_nor2_1 _10619_ (.A(_02601_),
    .B(_02627_),
    .Y(_02628_));
 sg13g2_nor2_1 _10620_ (.A(_02604_),
    .B(_02628_),
    .Y(_02629_));
 sg13g2_a221oi_1 _10621_ (.B2(_02627_),
    .C1(_02629_),
    .B1(_02601_),
    .A1(_02595_),
    .Y(_02630_),
    .A2(_02602_));
 sg13g2_a21oi_1 _10622_ (.A1(_02594_),
    .A2(_02605_),
    .Y(_02631_),
    .B1(_02630_));
 sg13g2_nand2_1 _10623_ (.Y(_02632_),
    .A(_02597_),
    .B(_02631_));
 sg13g2_inv_1 _10624_ (.Y(_02633_),
    .A(_02610_));
 sg13g2_o21ai_1 _10625_ (.B1(_02633_),
    .Y(_02634_),
    .A1(net298),
    .A2(_02631_));
 sg13g2_a22oi_1 _10626_ (.Y(_02635_),
    .B1(_02632_),
    .B2(_02634_),
    .A2(_02591_),
    .A1(_02625_));
 sg13g2_a221oi_1 _10627_ (.B2(_02590_),
    .C1(_02635_),
    .B1(_02624_),
    .A1(_02611_),
    .Y(_02636_),
    .A2(_02592_));
 sg13g2_a221oi_1 _10628_ (.B2(_02617_),
    .C1(_02636_),
    .B1(_02623_),
    .A1(_02593_),
    .Y(_02637_),
    .A2(_02589_));
 sg13g2_nor2_1 _10629_ (.A(_02617_),
    .B(_02623_),
    .Y(_02638_));
 sg13g2_nor4_1 _10630_ (.A(_02622_),
    .B(_02619_),
    .C(_02637_),
    .D(_02638_),
    .Y(_02639_));
 sg13g2_buf_1 _10631_ (.A(_00040_),
    .X(_02640_));
 sg13g2_o21ai_1 _10632_ (.B1(_02640_),
    .Y(_02641_),
    .A1(_02621_),
    .A2(_02639_));
 sg13g2_inv_1 _10633_ (.Y(_02642_),
    .A(_02619_));
 sg13g2_buf_1 _10634_ (.A(\am_sdr0.gain_spi[2] ),
    .X(_02643_));
 sg13g2_nand2_1 _10635_ (.Y(_02644_),
    .A(net298),
    .B(_02606_));
 sg13g2_nor2_1 _10636_ (.A(net298),
    .B(_02606_),
    .Y(_02645_));
 sg13g2_a221oi_1 _10637_ (.B2(_02604_),
    .C1(_02645_),
    .B1(_02644_),
    .A1(_02594_),
    .Y(_02646_),
    .A2(_02625_));
 sg13g2_a21oi_1 _10638_ (.A1(_02595_),
    .A2(_02611_),
    .Y(_02647_),
    .B1(_02646_));
 sg13g2_nand2_1 _10639_ (.Y(_02648_),
    .A(_02610_),
    .B(_02647_));
 sg13g2_o21ai_1 _10640_ (.B1(_02593_),
    .Y(_02649_),
    .A1(_02610_),
    .A2(_02647_));
 sg13g2_a22oi_1 _10641_ (.Y(_02650_),
    .B1(_02648_),
    .B2(_02649_),
    .A2(_02592_),
    .A1(_02616_));
 sg13g2_nor2_1 _10642_ (.A(_02616_),
    .B(_02592_),
    .Y(_02651_));
 sg13g2_nor4_1 _10643_ (.A(_02642_),
    .B(_02643_),
    .C(_02650_),
    .D(_02651_),
    .Y(_02652_));
 sg13g2_a21oi_1 _10644_ (.A1(_02642_),
    .A2(_02640_),
    .Y(_02653_),
    .B1(_02652_));
 sg13g2_o21ai_1 _10645_ (.B1(_02611_),
    .Y(_02654_),
    .A1(_02600_),
    .A2(net298));
 sg13g2_nor2_1 _10646_ (.A(_02600_),
    .B(_02611_),
    .Y(_02655_));
 sg13g2_a21o_1 _10647_ (.A2(_02655_),
    .A1(_02598_),
    .B1(_02604_),
    .X(_02656_));
 sg13g2_a22oi_1 _10648_ (.Y(_02657_),
    .B1(_02654_),
    .B2(_02656_),
    .A2(_02593_),
    .A1(_02594_));
 sg13g2_a21oi_1 _10649_ (.A1(_02595_),
    .A2(_02590_),
    .Y(_02658_),
    .B1(_02657_));
 sg13g2_a21oi_1 _10650_ (.A1(_02610_),
    .A2(_02658_),
    .Y(_02659_),
    .B1(_02617_));
 sg13g2_nor2_1 _10651_ (.A(_02610_),
    .B(_02658_),
    .Y(_02660_));
 sg13g2_nor2_1 _10652_ (.A(_02659_),
    .B(_02660_),
    .Y(_02661_));
 sg13g2_nor2_1 _10653_ (.A(_02619_),
    .B(_02661_),
    .Y(_02662_));
 sg13g2_nor2_1 _10654_ (.A(_02640_),
    .B(_02662_),
    .Y(_02663_));
 sg13g2_nand2b_1 _10655_ (.Y(_02664_),
    .B(_02590_),
    .A_N(_02623_));
 sg13g2_inv_1 _10656_ (.Y(_02665_),
    .A(_02601_));
 sg13g2_buf_1 _10657_ (.A(\am_sdr0.count[0] ),
    .X(_02666_));
 sg13g2_o21ai_1 _10658_ (.B1(_02626_),
    .Y(_02667_),
    .A1(_02600_),
    .A2(_02666_));
 sg13g2_nor2_1 _10659_ (.A(_02666_),
    .B(_02627_),
    .Y(_02668_));
 sg13g2_a21oi_1 _10660_ (.A1(_02604_),
    .A2(_02667_),
    .Y(_02669_),
    .B1(_02668_));
 sg13g2_o21ai_1 _10661_ (.B1(_02669_),
    .Y(_02670_),
    .A1(_02595_),
    .A2(_02601_));
 sg13g2_o21ai_1 _10662_ (.B1(_02670_),
    .Y(_02671_),
    .A1(_02594_),
    .A2(_02665_));
 sg13g2_nand2_1 _10663_ (.Y(_02672_),
    .A(_02602_),
    .B(_02671_));
 sg13g2_o21ai_1 _10664_ (.B1(_02633_),
    .Y(_02673_),
    .A1(_02602_),
    .A2(_02671_));
 sg13g2_a22oi_1 _10665_ (.Y(_02674_),
    .B1(_02672_),
    .B2(_02673_),
    .A2(_02591_),
    .A1(_02598_));
 sg13g2_a21oi_1 _10666_ (.A1(net298),
    .A2(_02592_),
    .Y(_02675_),
    .B1(_02674_));
 sg13g2_nor2_1 _10667_ (.A(_02589_),
    .B(_02675_),
    .Y(_02676_));
 sg13g2_a21oi_1 _10668_ (.A1(_02589_),
    .A2(_02675_),
    .Y(_02677_),
    .B1(_02625_));
 sg13g2_nor2_1 _10669_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sg13g2_nor2b_1 _10670_ (.A(_02590_),
    .B_N(_02623_),
    .Y(_02679_));
 sg13g2_a21o_1 _10671_ (.A2(_02678_),
    .A1(_02664_),
    .B1(_02679_),
    .X(_02680_));
 sg13g2_o21ai_1 _10672_ (.B1(_02617_),
    .Y(_02681_),
    .A1(\am_sdr0.am0.demod_out[15] ),
    .A2(_02680_));
 sg13g2_nand2_1 _10673_ (.Y(_02682_),
    .A(\am_sdr0.am0.demod_out[15] ),
    .B(_02680_));
 sg13g2_or2_1 _10674_ (.X(_02683_),
    .B(_02643_),
    .A(_02619_));
 sg13g2_a21oi_1 _10675_ (.A1(_02681_),
    .A2(_02682_),
    .Y(_02684_),
    .B1(_02683_));
 sg13g2_or3_1 _10676_ (.A(_02588_),
    .B(_02663_),
    .C(_02684_),
    .X(_02685_));
 sg13g2_o21ai_1 _10677_ (.B1(_02685_),
    .Y(_02686_),
    .A1(_02622_),
    .A2(_02653_));
 sg13g2_xnor2_1 _10678_ (.Y(_02687_),
    .A(_02588_),
    .B(_02619_));
 sg13g2_nand3_1 _10679_ (.B(_02619_),
    .C(_02643_),
    .A(_02588_),
    .Y(_02688_));
 sg13g2_o21ai_1 _10680_ (.B1(_02688_),
    .Y(_02689_),
    .A1(_02640_),
    .A2(_02687_));
 sg13g2_o21ai_1 _10681_ (.B1(_02689_),
    .Y(_02690_),
    .A1(_02595_),
    .A2(_02616_));
 sg13g2_o21ai_1 _10682_ (.B1(_02604_),
    .Y(_02691_),
    .A1(_02593_),
    .A2(_02655_));
 sg13g2_nand2_1 _10683_ (.Y(_02692_),
    .A(_02593_),
    .B(_02655_));
 sg13g2_a22oi_1 _10684_ (.Y(_02693_),
    .B1(_02691_),
    .B2(_02692_),
    .A2(_02616_),
    .A1(_02595_));
 sg13g2_o21ai_1 _10685_ (.B1(net257),
    .Y(_02694_),
    .A1(_02690_),
    .A2(_02693_));
 sg13g2_a21oi_1 _10686_ (.A1(_02641_),
    .A2(_02686_),
    .Y(_00074_),
    .B1(_02694_));
 sg13g2_nand3_1 _10687_ (.B(net299),
    .C(\am_sdr0.am0.q[2] ),
    .A(net302),
    .Y(_02695_));
 sg13g2_nand2_1 _10688_ (.Y(_02696_),
    .A(_01574_),
    .B(_01570_));
 sg13g2_buf_2 _10689_ (.A(_02696_),
    .X(_02697_));
 sg13g2_nand2_1 _10690_ (.Y(_02698_),
    .A(_02594_),
    .B(_02697_));
 sg13g2_buf_1 _10691_ (.A(net251),
    .X(_02699_));
 sg13g2_a21oi_1 _10692_ (.A1(_02695_),
    .A2(_02698_),
    .Y(_00097_),
    .B1(net181));
 sg13g2_nand3_1 _10693_ (.B(net299),
    .C(\am_sdr0.am0.q[3] ),
    .A(net302),
    .Y(_02700_));
 sg13g2_nand2_1 _10694_ (.Y(_02701_),
    .A(_02610_),
    .B(_02697_));
 sg13g2_a21oi_1 _10695_ (.A1(_02700_),
    .A2(_02701_),
    .Y(_00098_),
    .B1(net181));
 sg13g2_nand3_1 _10696_ (.B(net299),
    .C(\am_sdr0.am0.q[4] ),
    .A(net302),
    .Y(_02702_));
 sg13g2_nand2_1 _10697_ (.Y(_02703_),
    .A(_02591_),
    .B(_02697_));
 sg13g2_a21oi_1 _10698_ (.A1(_02702_),
    .A2(_02703_),
    .Y(_00099_),
    .B1(net181));
 sg13g2_nand3_1 _10699_ (.B(net299),
    .C(\am_sdr0.am0.q[5] ),
    .A(net302),
    .Y(_02704_));
 sg13g2_nand2_1 _10700_ (.Y(_02705_),
    .A(_02589_),
    .B(_02697_));
 sg13g2_a21oi_1 _10701_ (.A1(_02704_),
    .A2(_02705_),
    .Y(_00100_),
    .B1(net181));
 sg13g2_nand3_1 _10702_ (.B(net299),
    .C(\am_sdr0.am0.q[6] ),
    .A(net302),
    .Y(_02706_));
 sg13g2_nand2_1 _10703_ (.Y(_02707_),
    .A(_02623_),
    .B(_02697_));
 sg13g2_a21oi_1 _10704_ (.A1(_02706_),
    .A2(_02707_),
    .Y(_00101_),
    .B1(_02699_));
 sg13g2_nand3_1 _10705_ (.B(net299),
    .C(\am_sdr0.am0.q[7] ),
    .A(net302),
    .Y(_02708_));
 sg13g2_nand2_1 _10706_ (.Y(_02709_),
    .A(\am_sdr0.am0.demod_out[15] ),
    .B(_02697_));
 sg13g2_a21oi_1 _10707_ (.A1(_02708_),
    .A2(_02709_),
    .Y(_00102_),
    .B1(net181));
 sg13g2_nand3_1 _10708_ (.B(net299),
    .C(\am_sdr0.am0.q[0] ),
    .A(net302),
    .Y(_02710_));
 sg13g2_nand2_1 _10709_ (.Y(_02711_),
    .A(_02599_),
    .B(_02697_));
 sg13g2_a21oi_1 _10710_ (.A1(_02710_),
    .A2(_02711_),
    .Y(_00103_),
    .B1(net181));
 sg13g2_nand3_1 _10711_ (.B(net299),
    .C(\am_sdr0.am0.q[1] ),
    .A(net302),
    .Y(_02712_));
 sg13g2_nand2_1 _10712_ (.Y(_02713_),
    .A(_02604_),
    .B(_02697_));
 sg13g2_a21oi_1 _10713_ (.A1(_02712_),
    .A2(_02713_),
    .Y(_00104_),
    .B1(_02699_));
 sg13g2_nand2b_1 _10714_ (.Y(_02714_),
    .B(\am_sdr0.am0.state[3] ),
    .A_N(_01570_));
 sg13g2_a221oi_1 _10715_ (.B2(_01664_),
    .C1(_01663_),
    .B1(_02714_),
    .A1(_01687_),
    .Y(_00172_),
    .A2(_01678_));
 sg13g2_buf_1 _10716_ (.A(\am_sdr0.cic0.sample ),
    .X(_02715_));
 sg13g2_buf_2 _10717_ (.A(_02715_),
    .X(_02716_));
 sg13g2_buf_1 _10718_ (.A(_02716_),
    .X(_02717_));
 sg13g2_buf_1 _10719_ (.A(net250),
    .X(_02718_));
 sg13g2_xnor2_1 _10720_ (.Y(_02719_),
    .A(_02246_),
    .B(\am_sdr0.cic0.comb1_in_del[0] ));
 sg13g2_buf_2 _10721_ (.A(\am_sdr0.cic0.comb1[0] ),
    .X(_02720_));
 sg13g2_buf_1 _10722_ (.A(_02716_),
    .X(_02721_));
 sg13g2_o21ai_1 _10723_ (.B1(net257),
    .Y(_02722_),
    .A1(_02720_),
    .A2(net249));
 sg13g2_a21oi_1 _10724_ (.A1(net180),
    .A2(_02719_),
    .Y(_00191_),
    .B1(_02722_));
 sg13g2_buf_1 _10725_ (.A(\am_sdr0.cic0.comb1[10] ),
    .X(_02723_));
 sg13g2_inv_1 _10726_ (.Y(_02724_),
    .A(_02715_));
 sg13g2_buf_1 _10727_ (.A(_02724_),
    .X(_02725_));
 sg13g2_buf_1 _10728_ (.A(net248),
    .X(_02726_));
 sg13g2_nand2_1 _10729_ (.Y(_02727_),
    .A(_02723_),
    .B(net179));
 sg13g2_buf_1 _10730_ (.A(_02716_),
    .X(_02728_));
 sg13g2_buf_1 _10731_ (.A(_02728_),
    .X(_02729_));
 sg13g2_buf_1 _10732_ (.A(\am_sdr0.cic0.comb1_in_del[8] ),
    .X(_02730_));
 sg13g2_buf_1 _10733_ (.A(\am_sdr0.cic0.comb1_in_del[9] ),
    .X(_02731_));
 sg13g2_nor2_1 _10734_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sg13g2_nor2b_1 _10735_ (.A(_02731_),
    .B_N(_02293_),
    .Y(_02733_));
 sg13g2_buf_1 _10736_ (.A(\am_sdr0.cic0.comb1_in_del[5] ),
    .X(_02734_));
 sg13g2_inv_1 _10737_ (.Y(_02735_),
    .A(_02734_));
 sg13g2_buf_1 _10738_ (.A(\am_sdr0.cic0.comb1_in_del[4] ),
    .X(_02736_));
 sg13g2_nand2b_1 _10739_ (.Y(_02737_),
    .B(_02736_),
    .A_N(_02286_));
 sg13g2_inv_1 _10740_ (.Y(_02738_),
    .A(\am_sdr0.cic0.comb1_in_del[3] ));
 sg13g2_buf_1 _10741_ (.A(\am_sdr0.cic0.comb1_in_del[2] ),
    .X(_02739_));
 sg13g2_nor2_1 _10742_ (.A(_02280_),
    .B(_02739_),
    .Y(_02740_));
 sg13g2_nor2b_1 _10743_ (.A(_02246_),
    .B_N(\am_sdr0.cic0.comb1_in_del[0] ),
    .Y(_02741_));
 sg13g2_buf_1 _10744_ (.A(\am_sdr0.cic0.comb1_in_del[1] ),
    .X(_02742_));
 sg13g2_nand2b_1 _10745_ (.Y(_02743_),
    .B(_02278_),
    .A_N(_02742_));
 sg13g2_nor2b_1 _10746_ (.A(_02278_),
    .B_N(_02742_),
    .Y(_02744_));
 sg13g2_a221oi_1 _10747_ (.B2(_02743_),
    .C1(_02744_),
    .B1(_02741_),
    .A1(_02280_),
    .Y(_02745_),
    .A2(_02739_));
 sg13g2_buf_1 _10748_ (.A(_02745_),
    .X(_02746_));
 sg13g2_nor3_1 _10749_ (.A(_02738_),
    .B(_02740_),
    .C(_02746_),
    .Y(_02747_));
 sg13g2_o21ai_1 _10750_ (.B1(_02738_),
    .Y(_02748_),
    .A1(_02740_),
    .A2(_02746_));
 sg13g2_o21ai_1 _10751_ (.B1(_02748_),
    .Y(_02749_),
    .A1(_02283_),
    .A2(_02747_));
 sg13g2_buf_2 _10752_ (.A(_02749_),
    .X(_02750_));
 sg13g2_nor2b_1 _10753_ (.A(\am_sdr0.cic0.comb1_in_del[6] ),
    .B_N(_02289_),
    .Y(_02751_));
 sg13g2_nor2b_1 _10754_ (.A(_02736_),
    .B_N(_02286_),
    .Y(_02752_));
 sg13g2_or2_1 _10755_ (.X(_02753_),
    .B(_02752_),
    .A(_02751_));
 sg13g2_a221oi_1 _10756_ (.B2(_02750_),
    .C1(_02753_),
    .B1(_02737_),
    .A1(_02288_),
    .Y(_02754_),
    .A2(_02735_));
 sg13g2_buf_1 _10757_ (.A(_02754_),
    .X(_02755_));
 sg13g2_nand2b_1 _10758_ (.Y(_02756_),
    .B(_02734_),
    .A_N(_02288_));
 sg13g2_nand2b_1 _10759_ (.Y(_02757_),
    .B(\am_sdr0.cic0.comb1_in_del[6] ),
    .A_N(_02289_));
 sg13g2_o21ai_1 _10760_ (.B1(_02757_),
    .Y(_02758_),
    .A1(_02751_),
    .A2(_02756_));
 sg13g2_buf_1 _10761_ (.A(\am_sdr0.cic0.comb1_in_del[7] ),
    .X(_02759_));
 sg13g2_o21ai_1 _10762_ (.B1(_02759_),
    .Y(_02760_),
    .A1(_02755_),
    .A2(_02758_));
 sg13g2_nor3_1 _10763_ (.A(_02759_),
    .B(_02755_),
    .C(_02758_),
    .Y(_02761_));
 sg13g2_a21o_1 _10764_ (.A2(_02760_),
    .A1(_02291_),
    .B1(_02761_),
    .X(_02762_));
 sg13g2_buf_2 _10765_ (.A(_02762_),
    .X(_02763_));
 sg13g2_o21ai_1 _10766_ (.B1(_02763_),
    .Y(_02764_),
    .A1(_02732_),
    .A2(_02733_));
 sg13g2_inv_1 _10767_ (.Y(_02765_),
    .A(_02731_));
 sg13g2_nor2b_1 _10768_ (.A(_02730_),
    .B_N(_02293_),
    .Y(_02766_));
 sg13g2_a21oi_1 _10769_ (.A1(_02765_),
    .A2(_02766_),
    .Y(_02767_),
    .B1(_02295_));
 sg13g2_inv_1 _10770_ (.Y(_02768_),
    .A(_02730_));
 sg13g2_a21oi_1 _10771_ (.A1(_02768_),
    .A2(_02763_),
    .Y(_02769_),
    .B1(_02765_));
 sg13g2_o21ai_1 _10772_ (.B1(_02293_),
    .Y(_02770_),
    .A1(_02768_),
    .A2(_02763_));
 sg13g2_buf_1 _10773_ (.A(_02770_),
    .X(_02771_));
 sg13g2_a22oi_1 _10774_ (.Y(_02772_),
    .B1(_02769_),
    .B2(_02771_),
    .A2(_02767_),
    .A1(_02764_));
 sg13g2_buf_2 _10775_ (.A(_02772_),
    .X(_02773_));
 sg13g2_buf_1 _10776_ (.A(\am_sdr0.cic0.comb1_in_del[10] ),
    .X(_02774_));
 sg13g2_xor2_1 _10777_ (.B(_02774_),
    .A(_02257_),
    .X(_02775_));
 sg13g2_xnor2_1 _10778_ (.Y(_02776_),
    .A(_02773_),
    .B(_02775_));
 sg13g2_nand2_1 _10779_ (.Y(_02777_),
    .A(net178),
    .B(_02776_));
 sg13g2_buf_2 _10780_ (.A(net310),
    .X(_02778_));
 sg13g2_buf_2 _10781_ (.A(_02778_),
    .X(_02779_));
 sg13g2_buf_1 _10782_ (.A(_02779_),
    .X(_02780_));
 sg13g2_a21oi_1 _10783_ (.A1(_02727_),
    .A2(_02777_),
    .Y(_00192_),
    .B1(net131));
 sg13g2_buf_1 _10784_ (.A(net251),
    .X(_02781_));
 sg13g2_buf_1 _10785_ (.A(\am_sdr0.cic0.comb1[11] ),
    .X(_02782_));
 sg13g2_buf_1 _10786_ (.A(_02716_),
    .X(_02783_));
 sg13g2_nor2_1 _10787_ (.A(_02782_),
    .B(net247),
    .Y(_02784_));
 sg13g2_buf_2 _10788_ (.A(_02724_),
    .X(_02785_));
 sg13g2_buf_1 _10789_ (.A(_02785_),
    .X(_02786_));
 sg13g2_inv_1 _10790_ (.Y(_02787_),
    .A(_02774_));
 sg13g2_a21oi_1 _10791_ (.A1(_02787_),
    .A2(_02773_),
    .Y(_02788_),
    .B1(_02257_));
 sg13g2_nor2_1 _10792_ (.A(_02787_),
    .B(_02773_),
    .Y(_02789_));
 sg13g2_nor2_1 _10793_ (.A(_02788_),
    .B(_02789_),
    .Y(_02790_));
 sg13g2_buf_1 _10794_ (.A(\am_sdr0.cic0.comb1_in_del[11] ),
    .X(_02791_));
 sg13g2_nor2b_1 _10795_ (.A(_02791_),
    .B_N(_02259_),
    .Y(_02792_));
 sg13g2_nand2b_1 _10796_ (.Y(_02793_),
    .B(_02791_),
    .A_N(_02259_));
 sg13g2_nor2b_1 _10797_ (.A(_02792_),
    .B_N(_02793_),
    .Y(_02794_));
 sg13g2_xor2_1 _10798_ (.B(_02794_),
    .A(_02790_),
    .X(_02795_));
 sg13g2_nor2_1 _10799_ (.A(net176),
    .B(_02795_),
    .Y(_02796_));
 sg13g2_nor3_1 _10800_ (.A(net177),
    .B(_02784_),
    .C(_02796_),
    .Y(_00193_));
 sg13g2_buf_1 _10801_ (.A(\am_sdr0.cic0.comb1[12] ),
    .X(_02797_));
 sg13g2_nor2_1 _10802_ (.A(_02797_),
    .B(net247),
    .Y(_02798_));
 sg13g2_o21ai_1 _10803_ (.B1(_02791_),
    .Y(_02799_),
    .A1(_02788_),
    .A2(_02789_));
 sg13g2_nor3_1 _10804_ (.A(_02791_),
    .B(_02788_),
    .C(_02789_),
    .Y(_02800_));
 sg13g2_a21oi_2 _10805_ (.B1(_02800_),
    .Y(_02801_),
    .A2(_02799_),
    .A1(_02259_));
 sg13g2_buf_2 _10806_ (.A(\am_sdr0.cic0.comb1_in_del[12] ),
    .X(_02802_));
 sg13g2_nor2_1 _10807_ (.A(_02261_),
    .B(_02802_),
    .Y(_02803_));
 sg13g2_nand2_1 _10808_ (.Y(_02804_),
    .A(_02261_),
    .B(_02802_));
 sg13g2_nor2b_1 _10809_ (.A(_02803_),
    .B_N(_02804_),
    .Y(_02805_));
 sg13g2_xnor2_1 _10810_ (.Y(_02806_),
    .A(_02801_),
    .B(_02805_));
 sg13g2_nor2_1 _10811_ (.A(net176),
    .B(_02806_),
    .Y(_02807_));
 sg13g2_nor3_1 _10812_ (.A(net177),
    .B(_02798_),
    .C(_02807_),
    .Y(_00194_));
 sg13g2_buf_1 _10813_ (.A(net364),
    .X(_02808_));
 sg13g2_buf_1 _10814_ (.A(net297),
    .X(_02809_));
 sg13g2_buf_2 _10815_ (.A(\am_sdr0.cic0.comb1[13] ),
    .X(_02810_));
 sg13g2_nand2_1 _10816_ (.Y(_02811_),
    .A(_02810_),
    .B(net248));
 sg13g2_nand2_1 _10817_ (.Y(_02812_),
    .A(_02802_),
    .B(_02801_));
 sg13g2_o21ai_1 _10818_ (.B1(_02261_),
    .Y(_02813_),
    .A1(_02802_),
    .A2(_02801_));
 sg13g2_nand2b_1 _10819_ (.Y(_02814_),
    .B(_02264_),
    .A_N(\am_sdr0.cic0.comb1_in_del[13] ));
 sg13g2_buf_1 _10820_ (.A(_02814_),
    .X(_02815_));
 sg13g2_nand2b_1 _10821_ (.Y(_02816_),
    .B(\am_sdr0.cic0.comb1_in_del[13] ),
    .A_N(_02264_));
 sg13g2_buf_1 _10822_ (.A(_02816_),
    .X(_02817_));
 sg13g2_a21oi_1 _10823_ (.A1(_02815_),
    .A2(_02817_),
    .Y(_02818_),
    .B1(_02785_));
 sg13g2_nand3_1 _10824_ (.B(_02813_),
    .C(_02818_),
    .A(_02812_),
    .Y(_02819_));
 sg13g2_nand3_1 _10825_ (.B(_02815_),
    .C(_02817_),
    .A(_02716_),
    .Y(_02820_));
 sg13g2_a21o_1 _10826_ (.A2(_02813_),
    .A1(_02812_),
    .B1(_02820_),
    .X(_02821_));
 sg13g2_nand3_1 _10827_ (.B(_02819_),
    .C(_02821_),
    .A(_02811_),
    .Y(_02822_));
 sg13g2_and2_1 _10828_ (.A(net246),
    .B(_02822_),
    .X(_00195_));
 sg13g2_buf_1 _10829_ (.A(\am_sdr0.cic0.comb1[14] ),
    .X(_02823_));
 sg13g2_nand2_1 _10830_ (.Y(_02824_),
    .A(_02823_),
    .B(net179));
 sg13g2_and4_1 _10831_ (.A(_02794_),
    .B(_02805_),
    .C(_02815_),
    .D(_02817_),
    .X(_02825_));
 sg13g2_buf_1 _10832_ (.A(_02825_),
    .X(_02826_));
 sg13g2_nor2b_1 _10833_ (.A(_02775_),
    .B_N(_02826_),
    .Y(_02827_));
 sg13g2_nor2b_1 _10834_ (.A(_02774_),
    .B_N(_02257_),
    .Y(_02828_));
 sg13g2_a21oi_1 _10835_ (.A1(_02828_),
    .A2(_02793_),
    .Y(_02829_),
    .B1(_02792_));
 sg13g2_nand2_1 _10836_ (.Y(_02830_),
    .A(_02802_),
    .B(_02829_));
 sg13g2_o21ai_1 _10837_ (.B1(_02261_),
    .Y(_02831_),
    .A1(_02802_),
    .A2(_02829_));
 sg13g2_nand3_1 _10838_ (.B(_02830_),
    .C(_02831_),
    .A(_02817_),
    .Y(_02832_));
 sg13g2_nand2_1 _10839_ (.Y(_02833_),
    .A(_02815_),
    .B(_02832_));
 sg13g2_a21oi_1 _10840_ (.A1(_02773_),
    .A2(_02827_),
    .Y(_02834_),
    .B1(_02833_));
 sg13g2_buf_1 _10841_ (.A(\am_sdr0.cic0.comb1_in_del[14] ),
    .X(_02835_));
 sg13g2_xnor2_1 _10842_ (.Y(_02836_),
    .A(_02266_),
    .B(_02835_));
 sg13g2_xnor2_1 _10843_ (.Y(_02837_),
    .A(_02834_),
    .B(_02836_));
 sg13g2_nand2_1 _10844_ (.Y(_02838_),
    .A(net178),
    .B(_02837_));
 sg13g2_a21oi_1 _10845_ (.A1(_02824_),
    .A2(_02838_),
    .Y(_00196_),
    .B1(net131));
 sg13g2_buf_1 _10846_ (.A(net191),
    .X(_02839_));
 sg13g2_buf_1 _10847_ (.A(\am_sdr0.cic0.comb1[15] ),
    .X(_02840_));
 sg13g2_inv_1 _10848_ (.Y(_02841_),
    .A(_02835_));
 sg13g2_a21oi_1 _10849_ (.A1(_02841_),
    .A2(_02833_),
    .Y(_02842_),
    .B1(_02266_));
 sg13g2_nand3_1 _10850_ (.B(_02773_),
    .C(_02827_),
    .A(_02841_),
    .Y(_02843_));
 sg13g2_buf_1 _10851_ (.A(_02843_),
    .X(_02844_));
 sg13g2_nand2_1 _10852_ (.Y(_02845_),
    .A(_02828_),
    .B(_02826_));
 sg13g2_a21oi_1 _10853_ (.A1(_02792_),
    .A2(_02804_),
    .Y(_02846_),
    .B1(_02803_));
 sg13g2_nand2b_1 _10854_ (.Y(_02847_),
    .B(_02817_),
    .A_N(_02846_));
 sg13g2_nand4_1 _10855_ (.B(_02815_),
    .C(_02845_),
    .A(_02835_),
    .Y(_02848_),
    .D(_02847_));
 sg13g2_nand2_1 _10856_ (.Y(_02849_),
    .A(_02787_),
    .B(_02826_));
 sg13g2_a221oi_1 _10857_ (.B2(_02771_),
    .C1(_02849_),
    .B1(_02769_),
    .A1(_02764_),
    .Y(_02850_),
    .A2(_02767_));
 sg13g2_nand2_1 _10858_ (.Y(_02851_),
    .A(_02257_),
    .B(_02826_));
 sg13g2_a221oi_1 _10859_ (.B2(_02771_),
    .C1(_02851_),
    .B1(_02769_),
    .A1(_02764_),
    .Y(_02852_),
    .A2(_02767_));
 sg13g2_nor3_1 _10860_ (.A(_02848_),
    .B(_02850_),
    .C(_02852_),
    .Y(_02853_));
 sg13g2_a21o_1 _10861_ (.A2(_02844_),
    .A1(_02842_),
    .B1(_02853_),
    .X(_02854_));
 sg13g2_buf_1 _10862_ (.A(_02854_),
    .X(_02855_));
 sg13g2_buf_2 _10863_ (.A(\am_sdr0.cic0.comb1_in_del[15] ),
    .X(_02856_));
 sg13g2_xor2_1 _10864_ (.B(_02856_),
    .A(_02267_),
    .X(_02857_));
 sg13g2_xnor2_1 _10865_ (.Y(_02858_),
    .A(_02855_),
    .B(_02857_));
 sg13g2_nor2_1 _10866_ (.A(net248),
    .B(_02858_),
    .Y(_02859_));
 sg13g2_a21oi_1 _10867_ (.A1(_02840_),
    .A2(_02726_),
    .Y(_02860_),
    .B1(_02859_));
 sg13g2_nor2_1 _10868_ (.A(net130),
    .B(_02860_),
    .Y(_00197_));
 sg13g2_nor2_1 _10869_ (.A(_02856_),
    .B(_02855_),
    .Y(_02861_));
 sg13g2_nand2_1 _10870_ (.Y(_02862_),
    .A(_02856_),
    .B(_02855_));
 sg13g2_o21ai_1 _10871_ (.B1(_02862_),
    .Y(_02863_),
    .A1(_02267_),
    .A2(_02861_));
 sg13g2_buf_1 _10872_ (.A(\am_sdr0.cic0.comb1_in_del[16] ),
    .X(_02864_));
 sg13g2_xor2_1 _10873_ (.B(_02864_),
    .A(_02270_),
    .X(_02865_));
 sg13g2_xnor2_1 _10874_ (.Y(_02866_),
    .A(_02863_),
    .B(_02865_));
 sg13g2_buf_1 _10875_ (.A(\am_sdr0.cic0.comb1[16] ),
    .X(_02867_));
 sg13g2_o21ai_1 _10876_ (.B1(net257),
    .Y(_02868_),
    .A1(_02867_),
    .A2(net249));
 sg13g2_a21oi_1 _10877_ (.A1(net180),
    .A2(_02866_),
    .Y(_00198_),
    .B1(_02868_));
 sg13g2_buf_1 _10878_ (.A(\am_sdr0.cic0.comb1[17] ),
    .X(_02869_));
 sg13g2_buf_1 _10879_ (.A(_02716_),
    .X(_02870_));
 sg13g2_nor2_1 _10880_ (.A(_02271_),
    .B(_02864_),
    .Y(_02871_));
 sg13g2_or2_1 _10881_ (.X(_02872_),
    .B(_02864_),
    .A(_02856_));
 sg13g2_nand2b_1 _10882_ (.Y(_02873_),
    .B(_02267_),
    .A_N(_02864_));
 sg13g2_a221oi_1 _10883_ (.B2(_02873_),
    .C1(_02853_),
    .B1(_02872_),
    .A1(_02842_),
    .Y(_02874_),
    .A2(_02844_));
 sg13g2_nand2b_1 _10884_ (.Y(_02875_),
    .B(_02270_),
    .A_N(_02856_));
 sg13g2_nand2_1 _10885_ (.Y(_02876_),
    .A(_02267_),
    .B(_02270_));
 sg13g2_a221oi_1 _10886_ (.B2(_02876_),
    .C1(_02853_),
    .B1(_02875_),
    .A1(_02842_),
    .Y(_02877_),
    .A2(_02844_));
 sg13g2_nand2b_1 _10887_ (.Y(_02878_),
    .B(_02267_),
    .A_N(_02856_));
 sg13g2_a21oi_1 _10888_ (.A1(_02271_),
    .A2(_02864_),
    .Y(_02879_),
    .B1(_02878_));
 sg13g2_nor4_2 _10889_ (.A(_02871_),
    .B(_02874_),
    .C(_02877_),
    .Y(_02880_),
    .D(_02879_));
 sg13g2_nor2b_1 _10890_ (.A(_02274_),
    .B_N(\am_sdr0.cic0.comb1_in_del[17] ),
    .Y(_02881_));
 sg13g2_nand2b_1 _10891_ (.Y(_02882_),
    .B(_02274_),
    .A_N(\am_sdr0.cic0.comb1_in_del[17] ));
 sg13g2_nand2b_1 _10892_ (.Y(_02883_),
    .B(_02882_),
    .A_N(_02881_));
 sg13g2_xnor2_1 _10893_ (.Y(_02884_),
    .A(_02880_),
    .B(_02883_));
 sg13g2_nand2_1 _10894_ (.Y(_02885_),
    .A(net245),
    .B(_02884_));
 sg13g2_o21ai_1 _10895_ (.B1(_02885_),
    .Y(_02886_),
    .A1(_02869_),
    .A2(net178));
 sg13g2_nor2_1 _10896_ (.A(net130),
    .B(_02886_),
    .Y(_00199_));
 sg13g2_buf_1 _10897_ (.A(\am_sdr0.cic0.comb1[18] ),
    .X(_02887_));
 sg13g2_nor2_1 _10898_ (.A(_02887_),
    .B(net247),
    .Y(_02888_));
 sg13g2_buf_1 _10899_ (.A(\am_sdr0.cic0.comb1_in_del[18] ),
    .X(_02889_));
 sg13g2_xor2_1 _10900_ (.B(_02889_),
    .A(_02276_),
    .X(_02890_));
 sg13g2_a21oi_1 _10901_ (.A1(_02880_),
    .A2(_02882_),
    .Y(_02891_),
    .B1(_02881_));
 sg13g2_xnor2_1 _10902_ (.Y(_02892_),
    .A(_02890_),
    .B(_02891_));
 sg13g2_nor2_1 _10903_ (.A(net176),
    .B(_02892_),
    .Y(_02893_));
 sg13g2_nor3_1 _10904_ (.A(net177),
    .B(_02888_),
    .C(_02893_),
    .Y(_00200_));
 sg13g2_nand2b_1 _10905_ (.Y(_02894_),
    .B(_02889_),
    .A_N(_02276_));
 sg13g2_nor2b_1 _10906_ (.A(_02889_),
    .B_N(_02276_),
    .Y(_02895_));
 sg13g2_a21oi_1 _10907_ (.A1(_02894_),
    .A2(_02891_),
    .Y(_02896_),
    .B1(_02895_));
 sg13g2_xor2_1 _10908_ (.B(\am_sdr0.cic0.comb1_in_del[19] ),
    .A(\am_sdr0.cic0.integ_sample[19] ),
    .X(_02897_));
 sg13g2_and3_1 _10909_ (.X(_02898_),
    .A(net245),
    .B(_02896_),
    .C(_02897_));
 sg13g2_nor3_1 _10910_ (.A(_02725_),
    .B(_02896_),
    .C(_02897_),
    .Y(_02899_));
 sg13g2_o21ai_1 _10911_ (.B1(net253),
    .Y(_02900_),
    .A1(\am_sdr0.cic0.comb1[19] ),
    .A2(net249));
 sg13g2_nor3_1 _10912_ (.A(_02898_),
    .B(_02899_),
    .C(_02900_),
    .Y(_00201_));
 sg13g2_buf_2 _10913_ (.A(\am_sdr0.cic0.comb1[1] ),
    .X(_02901_));
 sg13g2_nand2_1 _10914_ (.Y(_02902_),
    .A(_02901_),
    .B(net179));
 sg13g2_xnor2_1 _10915_ (.Y(_02903_),
    .A(_02278_),
    .B(_02742_));
 sg13g2_xnor2_1 _10916_ (.Y(_02904_),
    .A(_02741_),
    .B(_02903_));
 sg13g2_nand2_1 _10917_ (.Y(_02905_),
    .A(net178),
    .B(_02904_));
 sg13g2_a21oi_1 _10918_ (.A1(_02902_),
    .A2(_02905_),
    .Y(_00202_),
    .B1(net131));
 sg13g2_buf_1 _10919_ (.A(\am_sdr0.cic0.comb1[2] ),
    .X(_02906_));
 sg13g2_a21oi_1 _10920_ (.A1(_02741_),
    .A2(_02743_),
    .Y(_02907_),
    .B1(_02744_));
 sg13g2_xnor2_1 _10921_ (.Y(_02908_),
    .A(\am_sdr0.cic0.integ_sample[2] ),
    .B(_02739_));
 sg13g2_xnor2_1 _10922_ (.Y(_02909_),
    .A(_02907_),
    .B(_02908_));
 sg13g2_nor2_1 _10923_ (.A(net248),
    .B(_02909_),
    .Y(_02910_));
 sg13g2_a21oi_1 _10924_ (.A1(_02906_),
    .A2(net179),
    .Y(_02911_),
    .B1(_02910_));
 sg13g2_nor2_1 _10925_ (.A(net130),
    .B(_02911_),
    .Y(_00203_));
 sg13g2_buf_1 _10926_ (.A(\am_sdr0.cic0.comb1[3] ),
    .X(_02912_));
 sg13g2_nand2_1 _10927_ (.Y(_02913_),
    .A(_02912_),
    .B(net179));
 sg13g2_nor2_1 _10928_ (.A(_02740_),
    .B(_02746_),
    .Y(_02914_));
 sg13g2_xnor2_1 _10929_ (.Y(_02915_),
    .A(\am_sdr0.cic0.integ_sample[3] ),
    .B(\am_sdr0.cic0.comb1_in_del[3] ));
 sg13g2_xnor2_1 _10930_ (.Y(_02916_),
    .A(_02914_),
    .B(_02915_));
 sg13g2_nand2_1 _10931_ (.Y(_02917_),
    .A(net178),
    .B(_02916_));
 sg13g2_a21oi_1 _10932_ (.A1(_02913_),
    .A2(_02917_),
    .Y(_00204_),
    .B1(net131));
 sg13g2_buf_1 _10933_ (.A(\am_sdr0.cic0.comb1[4] ),
    .X(_02918_));
 sg13g2_nor2_1 _10934_ (.A(_02918_),
    .B(net249),
    .Y(_02919_));
 sg13g2_xor2_1 _10935_ (.B(_02736_),
    .A(_02286_),
    .X(_02920_));
 sg13g2_xnor2_1 _10936_ (.Y(_02921_),
    .A(_02750_),
    .B(_02920_));
 sg13g2_nor2_1 _10937_ (.A(net248),
    .B(_02921_),
    .Y(_02922_));
 sg13g2_nor3_1 _10938_ (.A(net177),
    .B(_02919_),
    .C(_02922_),
    .Y(_00205_));
 sg13g2_buf_2 _10939_ (.A(\am_sdr0.cic0.comb1[5] ),
    .X(_02923_));
 sg13g2_a21oi_2 _10940_ (.B1(_02752_),
    .Y(_02924_),
    .A2(_02750_),
    .A1(_02737_));
 sg13g2_xor2_1 _10941_ (.B(_02734_),
    .A(_02288_),
    .X(_02925_));
 sg13g2_xnor2_1 _10942_ (.Y(_02926_),
    .A(_02924_),
    .B(_02925_));
 sg13g2_nand2_1 _10943_ (.Y(_02927_),
    .A(net245),
    .B(_02926_));
 sg13g2_o21ai_1 _10944_ (.B1(_02927_),
    .Y(_02928_),
    .A1(_02923_),
    .A2(net178));
 sg13g2_nor2_1 _10945_ (.A(net130),
    .B(_02928_),
    .Y(_00206_));
 sg13g2_buf_2 _10946_ (.A(\am_sdr0.cic0.comb1[6] ),
    .X(_02929_));
 sg13g2_nand2_1 _10947_ (.Y(_02930_),
    .A(_02929_),
    .B(net179));
 sg13g2_nand2_1 _10948_ (.Y(_02931_),
    .A(_02734_),
    .B(_02924_));
 sg13g2_nor2_1 _10949_ (.A(_02734_),
    .B(_02924_),
    .Y(_02932_));
 sg13g2_a21oi_1 _10950_ (.A1(_02288_),
    .A2(_02931_),
    .Y(_02933_),
    .B1(_02932_));
 sg13g2_nor2b_1 _10951_ (.A(_02751_),
    .B_N(_02757_),
    .Y(_02934_));
 sg13g2_xnor2_1 _10952_ (.Y(_02935_),
    .A(_02933_),
    .B(_02934_));
 sg13g2_nand2_1 _10953_ (.Y(_02936_),
    .A(net178),
    .B(_02935_));
 sg13g2_a21oi_1 _10954_ (.A1(_02930_),
    .A2(_02936_),
    .Y(_00207_),
    .B1(net131));
 sg13g2_buf_1 _10955_ (.A(\am_sdr0.cic0.comb1[7] ),
    .X(_02937_));
 sg13g2_nor2_1 _10956_ (.A(_02755_),
    .B(_02758_),
    .Y(_02938_));
 sg13g2_xnor2_1 _10957_ (.Y(_02939_),
    .A(_02291_),
    .B(_02759_));
 sg13g2_xnor2_1 _10958_ (.Y(_02940_),
    .A(_02938_),
    .B(_02939_));
 sg13g2_nor2_1 _10959_ (.A(net248),
    .B(_02940_),
    .Y(_02941_));
 sg13g2_a21oi_1 _10960_ (.A1(_02937_),
    .A2(net179),
    .Y(_02942_),
    .B1(_02941_));
 sg13g2_nor2_1 _10961_ (.A(net130),
    .B(_02942_),
    .Y(_00208_));
 sg13g2_buf_2 _10962_ (.A(\am_sdr0.cic0.comb1[8] ),
    .X(_02943_));
 sg13g2_xnor2_1 _10963_ (.Y(_02944_),
    .A(_02293_),
    .B(_02730_));
 sg13g2_xnor2_1 _10964_ (.Y(_02945_),
    .A(_02763_),
    .B(_02944_));
 sg13g2_nand2_1 _10965_ (.Y(_02946_),
    .A(net245),
    .B(_02945_));
 sg13g2_o21ai_1 _10966_ (.B1(_02946_),
    .Y(_02947_),
    .A1(_02943_),
    .A2(net178));
 sg13g2_nor2_1 _10967_ (.A(net130),
    .B(_02947_),
    .Y(_00209_));
 sg13g2_buf_1 _10968_ (.A(\am_sdr0.cic0.comb1[9] ),
    .X(_02948_));
 sg13g2_inv_1 _10969_ (.Y(_02949_),
    .A(_02948_));
 sg13g2_inv_1 _10970_ (.Y(_02950_),
    .A(_02763_));
 sg13g2_o21ai_1 _10971_ (.B1(_02771_),
    .Y(_02951_),
    .A1(_02730_),
    .A2(_02950_));
 sg13g2_xnor2_1 _10972_ (.Y(_02952_),
    .A(_02295_),
    .B(_02731_));
 sg13g2_xnor2_1 _10973_ (.Y(_02953_),
    .A(_02951_),
    .B(_02952_));
 sg13g2_mux2_1 _10974_ (.A0(_02949_),
    .A1(_02953_),
    .S(net245),
    .X(_02954_));
 sg13g2_nor2_1 _10975_ (.A(net130),
    .B(_02954_),
    .Y(_00210_));
 sg13g2_buf_1 _10976_ (.A(_02728_),
    .X(_02955_));
 sg13g2_nand2_1 _10977_ (.Y(_02956_),
    .A(_02246_),
    .B(net175));
 sg13g2_nand2_1 _10978_ (.Y(_02957_),
    .A(\am_sdr0.cic0.comb1_in_del[0] ),
    .B(net179));
 sg13g2_a21oi_1 _10979_ (.A1(_02956_),
    .A2(_02957_),
    .Y(_00211_),
    .B1(_02780_));
 sg13g2_nand2_1 _10980_ (.Y(_02958_),
    .A(_02257_),
    .B(net175));
 sg13g2_buf_1 _10981_ (.A(_02725_),
    .X(_02959_));
 sg13g2_nand2_1 _10982_ (.Y(_02960_),
    .A(_02774_),
    .B(net174));
 sg13g2_a21oi_1 _10983_ (.A1(_02958_),
    .A2(_02960_),
    .Y(_00212_),
    .B1(net131));
 sg13g2_nand2_1 _10984_ (.Y(_02961_),
    .A(_02259_),
    .B(net175));
 sg13g2_nand2_1 _10985_ (.Y(_02962_),
    .A(_02791_),
    .B(net174));
 sg13g2_a21oi_1 _10986_ (.A1(_02961_),
    .A2(_02962_),
    .Y(_00213_),
    .B1(net131));
 sg13g2_nand2_1 _10987_ (.Y(_02963_),
    .A(\am_sdr0.cic0.integ_sample[12] ),
    .B(net175));
 sg13g2_nand2_1 _10988_ (.Y(_02964_),
    .A(_02802_),
    .B(net174));
 sg13g2_a21oi_1 _10989_ (.A1(_02963_),
    .A2(_02964_),
    .Y(_00214_),
    .B1(_02780_));
 sg13g2_nand2_1 _10990_ (.Y(_02965_),
    .A(_02264_),
    .B(net175));
 sg13g2_nand2_1 _10991_ (.Y(_02966_),
    .A(\am_sdr0.cic0.comb1_in_del[13] ),
    .B(net174));
 sg13g2_a21oi_1 _10992_ (.A1(_02965_),
    .A2(_02966_),
    .Y(_00215_),
    .B1(net131));
 sg13g2_nand2_1 _10993_ (.Y(_02967_),
    .A(_02266_),
    .B(_02955_));
 sg13g2_nand2_1 _10994_ (.Y(_02968_),
    .A(_02835_),
    .B(net174));
 sg13g2_buf_1 _10995_ (.A(_02779_),
    .X(_02969_));
 sg13g2_a21oi_1 _10996_ (.A1(_02967_),
    .A2(_02968_),
    .Y(_00216_),
    .B1(net129));
 sg13g2_nand2_1 _10997_ (.Y(_02970_),
    .A(_02267_),
    .B(net175));
 sg13g2_nand2_1 _10998_ (.Y(_02971_),
    .A(_02856_),
    .B(net174));
 sg13g2_a21oi_1 _10999_ (.A1(_02970_),
    .A2(_02971_),
    .Y(_00217_),
    .B1(net129));
 sg13g2_nand2_1 _11000_ (.Y(_02972_),
    .A(_02270_),
    .B(net175));
 sg13g2_nand2_1 _11001_ (.Y(_02973_),
    .A(_02864_),
    .B(net174));
 sg13g2_a21oi_1 _11002_ (.A1(_02972_),
    .A2(_02973_),
    .Y(_00218_),
    .B1(net129));
 sg13g2_nand2_1 _11003_ (.Y(_02974_),
    .A(_02274_),
    .B(_02955_));
 sg13g2_nand2_1 _11004_ (.Y(_02975_),
    .A(\am_sdr0.cic0.comb1_in_del[17] ),
    .B(net174));
 sg13g2_a21oi_1 _11005_ (.A1(_02974_),
    .A2(_02975_),
    .Y(_00219_),
    .B1(net129));
 sg13g2_nand2_1 _11006_ (.Y(_02976_),
    .A(_02276_),
    .B(net175));
 sg13g2_nand2_1 _11007_ (.Y(_02977_),
    .A(_02889_),
    .B(_02959_));
 sg13g2_a21oi_1 _11008_ (.A1(_02976_),
    .A2(_02977_),
    .Y(_00220_),
    .B1(_02969_));
 sg13g2_buf_1 _11009_ (.A(_02728_),
    .X(_02978_));
 sg13g2_nand2_1 _11010_ (.Y(_02979_),
    .A(\am_sdr0.cic0.integ_sample[19] ),
    .B(_02978_));
 sg13g2_nand2_1 _11011_ (.Y(_02980_),
    .A(\am_sdr0.cic0.comb1_in_del[19] ),
    .B(_02959_));
 sg13g2_a21oi_1 _11012_ (.A1(_02979_),
    .A2(_02980_),
    .Y(_00221_),
    .B1(_02969_));
 sg13g2_nand2_1 _11013_ (.Y(_02981_),
    .A(_02278_),
    .B(net173));
 sg13g2_buf_1 _11014_ (.A(_02785_),
    .X(_02982_));
 sg13g2_nand2_1 _11015_ (.Y(_02983_),
    .A(_02742_),
    .B(_02982_));
 sg13g2_a21oi_1 _11016_ (.A1(_02981_),
    .A2(_02983_),
    .Y(_00222_),
    .B1(net129));
 sg13g2_nand2_1 _11017_ (.Y(_02984_),
    .A(\am_sdr0.cic0.integ_sample[2] ),
    .B(_02978_));
 sg13g2_nand2_1 _11018_ (.Y(_02985_),
    .A(_02739_),
    .B(_02982_));
 sg13g2_a21oi_1 _11019_ (.A1(_02984_),
    .A2(_02985_),
    .Y(_00223_),
    .B1(net129));
 sg13g2_nand2_1 _11020_ (.Y(_02986_),
    .A(\am_sdr0.cic0.integ_sample[3] ),
    .B(net173));
 sg13g2_nand2_1 _11021_ (.Y(_02987_),
    .A(\am_sdr0.cic0.comb1_in_del[3] ),
    .B(net172));
 sg13g2_a21oi_1 _11022_ (.A1(_02986_),
    .A2(_02987_),
    .Y(_00224_),
    .B1(net129));
 sg13g2_nand2_1 _11023_ (.Y(_02988_),
    .A(_02286_),
    .B(net173));
 sg13g2_nand2_1 _11024_ (.Y(_02989_),
    .A(_02736_),
    .B(net172));
 sg13g2_a21oi_1 _11025_ (.A1(_02988_),
    .A2(_02989_),
    .Y(_00225_),
    .B1(net129));
 sg13g2_nand2_1 _11026_ (.Y(_02990_),
    .A(_02288_),
    .B(net173));
 sg13g2_nand2_1 _11027_ (.Y(_02991_),
    .A(_02734_),
    .B(net172));
 sg13g2_buf_1 _11028_ (.A(_02779_),
    .X(_02992_));
 sg13g2_a21oi_1 _11029_ (.A1(_02990_),
    .A2(_02991_),
    .Y(_00226_),
    .B1(net128));
 sg13g2_nand2_1 _11030_ (.Y(_02993_),
    .A(_02289_),
    .B(net173));
 sg13g2_nand2_1 _11031_ (.Y(_02994_),
    .A(\am_sdr0.cic0.comb1_in_del[6] ),
    .B(net172));
 sg13g2_a21oi_1 _11032_ (.A1(_02993_),
    .A2(_02994_),
    .Y(_00227_),
    .B1(net128));
 sg13g2_nand2_1 _11033_ (.Y(_02995_),
    .A(_02291_),
    .B(net173));
 sg13g2_nand2_1 _11034_ (.Y(_02996_),
    .A(_02759_),
    .B(net172));
 sg13g2_a21oi_1 _11035_ (.A1(_02995_),
    .A2(_02996_),
    .Y(_00228_),
    .B1(net128));
 sg13g2_nand2_1 _11036_ (.Y(_02997_),
    .A(_02293_),
    .B(net173));
 sg13g2_nand2_1 _11037_ (.Y(_02998_),
    .A(_02730_),
    .B(net172));
 sg13g2_a21oi_1 _11038_ (.A1(_02997_),
    .A2(_02998_),
    .Y(_00229_),
    .B1(net128));
 sg13g2_nand2_1 _11039_ (.Y(_02999_),
    .A(_02295_),
    .B(net173));
 sg13g2_nand2_1 _11040_ (.Y(_03000_),
    .A(_02731_),
    .B(net172));
 sg13g2_a21oi_1 _11041_ (.A1(_02999_),
    .A2(_03000_),
    .Y(_00230_),
    .B1(net128));
 sg13g2_xnor2_1 _11042_ (.Y(_03001_),
    .A(_02720_),
    .B(\am_sdr0.cic0.comb2_in_del[0] ));
 sg13g2_buf_1 _11043_ (.A(net303),
    .X(_03002_));
 sg13g2_o21ai_1 _11044_ (.B1(net244),
    .Y(_03003_),
    .A1(\am_sdr0.cic0.comb2[0] ),
    .A2(net249));
 sg13g2_a21oi_1 _11045_ (.A1(net180),
    .A2(_03001_),
    .Y(_00231_),
    .B1(_03003_));
 sg13g2_buf_1 _11046_ (.A(net250),
    .X(_03004_));
 sg13g2_inv_1 _11047_ (.Y(_03005_),
    .A(_02912_));
 sg13g2_inv_1 _11048_ (.Y(_03006_),
    .A(_02906_));
 sg13g2_buf_1 _11049_ (.A(\am_sdr0.cic0.comb2_in_del[2] ),
    .X(_03007_));
 sg13g2_nor2_1 _11050_ (.A(_03006_),
    .B(_03007_),
    .Y(_03008_));
 sg13g2_nor2b_1 _11051_ (.A(_02720_),
    .B_N(\am_sdr0.cic0.comb2_in_del[0] ),
    .Y(_03009_));
 sg13g2_buf_1 _11052_ (.A(\am_sdr0.cic0.comb2_in_del[1] ),
    .X(_03010_));
 sg13g2_nand2b_1 _11053_ (.Y(_03011_),
    .B(_02901_),
    .A_N(_03010_));
 sg13g2_nor2b_1 _11054_ (.A(_02901_),
    .B_N(_03010_),
    .Y(_03012_));
 sg13g2_a221oi_1 _11055_ (.B2(_03011_),
    .C1(_03012_),
    .B1(_03009_),
    .A1(_03006_),
    .Y(_03013_),
    .A2(_03007_));
 sg13g2_buf_1 _11056_ (.A(_03013_),
    .X(_03014_));
 sg13g2_inv_1 _11057_ (.Y(_03015_),
    .A(\am_sdr0.cic0.comb2_in_del[3] ));
 sg13g2_o21ai_1 _11058_ (.B1(_03015_),
    .Y(_03016_),
    .A1(_03008_),
    .A2(_03014_));
 sg13g2_nor3_1 _11059_ (.A(_03015_),
    .B(_03008_),
    .C(_03014_),
    .Y(_03017_));
 sg13g2_a21o_1 _11060_ (.A2(_03016_),
    .A1(_03005_),
    .B1(_03017_),
    .X(_03018_));
 sg13g2_buf_1 _11061_ (.A(_03018_),
    .X(_03019_));
 sg13g2_nand2b_1 _11062_ (.Y(_03020_),
    .B(_02918_),
    .A_N(\am_sdr0.cic0.comb2_in_del[4] ));
 sg13g2_buf_1 _11063_ (.A(\am_sdr0.cic0.comb2_in_del[5] ),
    .X(_03021_));
 sg13g2_nand2b_1 _11064_ (.Y(_03022_),
    .B(\am_sdr0.cic0.comb2_in_del[4] ),
    .A_N(_02918_));
 sg13g2_buf_1 _11065_ (.A(_03022_),
    .X(_03023_));
 sg13g2_nand2b_1 _11066_ (.Y(_03024_),
    .B(_03023_),
    .A_N(_03021_));
 sg13g2_nand2_1 _11067_ (.Y(_03025_),
    .A(_02923_),
    .B(_03023_));
 sg13g2_buf_1 _11068_ (.A(\am_sdr0.cic0.comb2_in_del[7] ),
    .X(_03026_));
 sg13g2_nand2b_1 _11069_ (.Y(_03027_),
    .B(_03026_),
    .A_N(_02937_));
 sg13g2_buf_1 _11070_ (.A(_03027_),
    .X(_03028_));
 sg13g2_buf_1 _11071_ (.A(\am_sdr0.cic0.comb2_in_del[8] ),
    .X(_03029_));
 sg13g2_inv_1 _11072_ (.Y(_03030_),
    .A(_03029_));
 sg13g2_o21ai_1 _11073_ (.B1(_03030_),
    .Y(_03031_),
    .A1(_02943_),
    .A2(_03028_));
 sg13g2_nand2_1 _11074_ (.Y(_03032_),
    .A(_02943_),
    .B(_03028_));
 sg13g2_buf_1 _11075_ (.A(\am_sdr0.cic0.comb2_in_del[6] ),
    .X(_03033_));
 sg13g2_nor2b_1 _11076_ (.A(_02929_),
    .B_N(_03033_),
    .Y(_03034_));
 sg13g2_a21o_1 _11077_ (.A2(_03032_),
    .A1(_03031_),
    .B1(_03034_),
    .X(_03035_));
 sg13g2_a221oi_1 _11078_ (.B2(_03025_),
    .C1(_03035_),
    .B1(_03024_),
    .A1(_03019_),
    .Y(_03036_),
    .A2(_03020_));
 sg13g2_buf_2 _11079_ (.A(_03036_),
    .X(_03037_));
 sg13g2_nand2b_1 _11080_ (.Y(_03038_),
    .B(_02923_),
    .A_N(_03021_));
 sg13g2_inv_1 _11081_ (.Y(_03039_),
    .A(_02943_));
 sg13g2_nand2b_1 _11082_ (.Y(_03040_),
    .B(_02937_),
    .A_N(_03026_));
 sg13g2_nand3b_1 _11083_ (.B(_03028_),
    .C(_02929_),
    .Y(_03041_),
    .A_N(_03033_));
 sg13g2_a22oi_1 _11084_ (.Y(_03042_),
    .B1(_03040_),
    .B2(_03041_),
    .A2(_03029_),
    .A1(_03039_));
 sg13g2_a21oi_1 _11085_ (.A1(_02943_),
    .A2(_03030_),
    .Y(_03043_),
    .B1(_03042_));
 sg13g2_o21ai_1 _11086_ (.B1(_03043_),
    .Y(_03044_),
    .A1(_03035_),
    .A2(_03038_));
 sg13g2_buf_1 _11087_ (.A(_03044_),
    .X(_03045_));
 sg13g2_buf_1 _11088_ (.A(\am_sdr0.cic0.comb2_in_del[9] ),
    .X(_03046_));
 sg13g2_inv_1 _11089_ (.Y(_03047_),
    .A(_03046_));
 sg13g2_o21ai_1 _11090_ (.B1(_03047_),
    .Y(_03048_),
    .A1(_03037_),
    .A2(_03045_));
 sg13g2_nor3_1 _11091_ (.A(_03047_),
    .B(_03037_),
    .C(_03045_),
    .Y(_03049_));
 sg13g2_a21oi_1 _11092_ (.A1(_02949_),
    .A2(_03048_),
    .Y(_03050_),
    .B1(_03049_));
 sg13g2_buf_1 _11093_ (.A(\am_sdr0.cic0.comb2_in_del[10] ),
    .X(_03051_));
 sg13g2_nor2b_1 _11094_ (.A(_03051_),
    .B_N(_02723_),
    .Y(_03052_));
 sg13g2_nand2b_1 _11095_ (.Y(_03053_),
    .B(_03051_),
    .A_N(_02723_));
 sg13g2_nand2b_1 _11096_ (.Y(_03054_),
    .B(_03053_),
    .A_N(_03052_));
 sg13g2_xnor2_1 _11097_ (.Y(_03055_),
    .A(_03050_),
    .B(_03054_));
 sg13g2_buf_1 _11098_ (.A(\am_sdr0.cic0.comb2[10] ),
    .X(_03056_));
 sg13g2_nor2b_1 _11099_ (.A(net250),
    .B_N(_03056_),
    .Y(_03057_));
 sg13g2_a21oi_1 _11100_ (.A1(net171),
    .A2(_03055_),
    .Y(_03058_),
    .B1(_03057_));
 sg13g2_nor2_1 _11101_ (.A(net130),
    .B(_03058_),
    .Y(_00232_));
 sg13g2_buf_2 _11102_ (.A(\am_sdr0.cic0.comb2[11] ),
    .X(_03059_));
 sg13g2_o21ai_1 _11103_ (.B1(_03053_),
    .Y(_03060_),
    .A1(_03050_),
    .A2(_03052_));
 sg13g2_buf_2 _11104_ (.A(\am_sdr0.cic0.comb2_in_del[11] ),
    .X(_03061_));
 sg13g2_xor2_1 _11105_ (.B(_03061_),
    .A(_02782_),
    .X(_03062_));
 sg13g2_xnor2_1 _11106_ (.Y(_03063_),
    .A(_03060_),
    .B(_03062_));
 sg13g2_nand2_1 _11107_ (.Y(_03064_),
    .A(net245),
    .B(_03063_));
 sg13g2_o21ai_1 _11108_ (.B1(_03064_),
    .Y(_03065_),
    .A1(_03059_),
    .A2(_02729_));
 sg13g2_nor2_1 _11109_ (.A(_02839_),
    .B(_03065_),
    .Y(_00233_));
 sg13g2_buf_1 _11110_ (.A(\am_sdr0.cic0.comb2[12] ),
    .X(_03066_));
 sg13g2_or2_1 _11111_ (.X(_03067_),
    .B(_03061_),
    .A(_03051_));
 sg13g2_inv_1 _11112_ (.Y(_03068_),
    .A(_03061_));
 sg13g2_nand2_1 _11113_ (.Y(_03069_),
    .A(_02723_),
    .B(_03068_));
 sg13g2_a221oi_1 _11114_ (.B2(_03069_),
    .C1(_03049_),
    .B1(_03067_),
    .A1(_02949_),
    .Y(_03070_),
    .A2(_03048_));
 sg13g2_a21oi_1 _11115_ (.A1(_03068_),
    .A2(_03052_),
    .Y(_03071_),
    .B1(_02782_));
 sg13g2_nand2b_1 _11116_ (.Y(_03072_),
    .B(_03071_),
    .A_N(_03070_));
 sg13g2_nand3_1 _11117_ (.B(_03051_),
    .C(_03061_),
    .A(_03046_),
    .Y(_03073_));
 sg13g2_nor3_1 _11118_ (.A(_03037_),
    .B(_03045_),
    .C(_03073_),
    .Y(_03074_));
 sg13g2_nand2_1 _11119_ (.Y(_03075_),
    .A(_02949_),
    .B(_03051_));
 sg13g2_nor4_1 _11120_ (.A(_03068_),
    .B(_03037_),
    .C(_03045_),
    .D(_03075_),
    .Y(_03076_));
 sg13g2_nand2b_1 _11121_ (.Y(_03077_),
    .B(_03046_),
    .A_N(_02723_));
 sg13g2_nor4_1 _11122_ (.A(_03068_),
    .B(_03037_),
    .C(_03045_),
    .D(_03077_),
    .Y(_03078_));
 sg13g2_or2_1 _11123_ (.X(_03079_),
    .B(_02723_),
    .A(_02948_));
 sg13g2_nor4_1 _11124_ (.A(_03068_),
    .B(_03037_),
    .C(_03045_),
    .D(_03079_),
    .Y(_03080_));
 sg13g2_or4_1 _11125_ (.A(_03074_),
    .B(_03076_),
    .C(_03078_),
    .D(_03080_),
    .X(_03081_));
 sg13g2_buf_1 _11126_ (.A(_03081_),
    .X(_03082_));
 sg13g2_nor2_1 _11127_ (.A(_03068_),
    .B(_03053_),
    .Y(_03083_));
 sg13g2_nor2_1 _11128_ (.A(_02948_),
    .B(_03047_),
    .Y(_03084_));
 sg13g2_nand3_1 _11129_ (.B(_03061_),
    .C(_03084_),
    .A(_03051_),
    .Y(_03085_));
 sg13g2_nand3b_1 _11130_ (.B(_03061_),
    .C(_03084_),
    .Y(_03086_),
    .A_N(_02723_));
 sg13g2_nand3b_1 _11131_ (.B(_03085_),
    .C(_03086_),
    .Y(_03087_),
    .A_N(_03083_));
 sg13g2_buf_1 _11132_ (.A(_03087_),
    .X(_03088_));
 sg13g2_nor2_1 _11133_ (.A(_03082_),
    .B(_03088_),
    .Y(_03089_));
 sg13g2_and2_1 _11134_ (.A(_03072_),
    .B(_03089_),
    .X(_03090_));
 sg13g2_buf_1 _11135_ (.A(\am_sdr0.cic0.comb2_in_del[12] ),
    .X(_03091_));
 sg13g2_xnor2_1 _11136_ (.Y(_03092_),
    .A(_02797_),
    .B(_03091_));
 sg13g2_xnor2_1 _11137_ (.Y(_03093_),
    .A(_03090_),
    .B(_03092_));
 sg13g2_nand2_1 _11138_ (.Y(_03094_),
    .A(net245),
    .B(_03093_));
 sg13g2_o21ai_1 _11139_ (.B1(_03094_),
    .Y(_03095_),
    .A1(_03066_),
    .A2(_02729_));
 sg13g2_nor2_1 _11140_ (.A(_02839_),
    .B(_03095_),
    .Y(_00234_));
 sg13g2_buf_1 _11141_ (.A(net191),
    .X(_03096_));
 sg13g2_buf_1 _11142_ (.A(\am_sdr0.cic0.comb2[13] ),
    .X(_03097_));
 sg13g2_buf_1 _11143_ (.A(_02716_),
    .X(_03098_));
 sg13g2_nor2b_1 _11144_ (.A(_03091_),
    .B_N(_02797_),
    .Y(_03099_));
 sg13g2_nand2b_1 _11145_ (.Y(_03100_),
    .B(_03091_),
    .A_N(_02797_));
 sg13g2_o21ai_1 _11146_ (.B1(_03100_),
    .Y(_03101_),
    .A1(_03090_),
    .A2(_03099_));
 sg13g2_xor2_1 _11147_ (.B(\am_sdr0.cic0.comb2_in_del[13] ),
    .A(_02810_),
    .X(_03102_));
 sg13g2_xnor2_1 _11148_ (.Y(_03103_),
    .A(_03101_),
    .B(_03102_));
 sg13g2_nand2_1 _11149_ (.Y(_03104_),
    .A(net243),
    .B(_03103_));
 sg13g2_o21ai_1 _11150_ (.B1(_03104_),
    .Y(_03105_),
    .A1(_03097_),
    .A2(_02783_));
 sg13g2_nor2_1 _11151_ (.A(_03096_),
    .B(_03105_),
    .Y(_00235_));
 sg13g2_buf_1 _11152_ (.A(\am_sdr0.cic0.comb2[14] ),
    .X(_03106_));
 sg13g2_nand2_1 _11153_ (.Y(_03107_),
    .A(_02810_),
    .B(_03100_));
 sg13g2_nor3_1 _11154_ (.A(_03082_),
    .B(_03088_),
    .C(_03107_),
    .Y(_03108_));
 sg13g2_inv_1 _11155_ (.Y(_03109_),
    .A(\am_sdr0.cic0.comb2_in_del[13] ));
 sg13g2_nand2_1 _11156_ (.Y(_03110_),
    .A(_03109_),
    .B(_03100_));
 sg13g2_nor3_1 _11157_ (.A(_03082_),
    .B(_03088_),
    .C(_03110_),
    .Y(_03111_));
 sg13g2_o21ai_1 _11158_ (.B1(_03072_),
    .Y(_03112_),
    .A1(_03108_),
    .A2(_03111_));
 sg13g2_nand2_1 _11159_ (.Y(_03113_),
    .A(_02810_),
    .B(_03109_));
 sg13g2_o21ai_1 _11160_ (.B1(_03099_),
    .Y(_03114_),
    .A1(_02810_),
    .A2(_03109_));
 sg13g2_and2_1 _11161_ (.A(_03113_),
    .B(_03114_),
    .X(_03115_));
 sg13g2_buf_1 _11162_ (.A(_03115_),
    .X(_03116_));
 sg13g2_and2_1 _11163_ (.A(_03112_),
    .B(_03116_),
    .X(_03117_));
 sg13g2_nor2b_1 _11164_ (.A(_02823_),
    .B_N(\am_sdr0.cic0.comb2_in_del[14] ),
    .Y(_03118_));
 sg13g2_nand2b_1 _11165_ (.Y(_03119_),
    .B(_02823_),
    .A_N(\am_sdr0.cic0.comb2_in_del[14] ));
 sg13g2_buf_1 _11166_ (.A(_03119_),
    .X(_03120_));
 sg13g2_nor2b_1 _11167_ (.A(_03118_),
    .B_N(_03120_),
    .Y(_03121_));
 sg13g2_xor2_1 _11168_ (.B(_03121_),
    .A(_03117_),
    .X(_03122_));
 sg13g2_nand2_1 _11169_ (.Y(_03123_),
    .A(net243),
    .B(_03122_));
 sg13g2_o21ai_1 _11170_ (.B1(_03123_),
    .Y(_03124_),
    .A1(_03106_),
    .A2(_02783_));
 sg13g2_nor2_1 _11171_ (.A(_03096_),
    .B(_03124_),
    .Y(_00236_));
 sg13g2_buf_1 _11172_ (.A(\am_sdr0.cic0.comb2[15] ),
    .X(_03125_));
 sg13g2_inv_1 _11173_ (.Y(_03126_),
    .A(_03125_));
 sg13g2_a21oi_1 _11174_ (.A1(_03117_),
    .A2(_03120_),
    .Y(_03127_),
    .B1(_03118_));
 sg13g2_buf_1 _11175_ (.A(\am_sdr0.cic0.comb2_in_del[15] ),
    .X(_03128_));
 sg13g2_xnor2_1 _11176_ (.Y(_03129_),
    .A(_02840_),
    .B(_03128_));
 sg13g2_xnor2_1 _11177_ (.Y(_03130_),
    .A(_03127_),
    .B(_03129_));
 sg13g2_mux2_1 _11178_ (.A0(_03126_),
    .A1(_03130_),
    .S(net245),
    .X(_03131_));
 sg13g2_nor2_1 _11179_ (.A(net127),
    .B(_03131_),
    .Y(_00237_));
 sg13g2_inv_1 _11180_ (.Y(_03132_),
    .A(\am_sdr0.cic0.comb2[16] ));
 sg13g2_inv_1 _11181_ (.Y(_03133_),
    .A(_02840_));
 sg13g2_nand2_1 _11182_ (.Y(_03134_),
    .A(_03133_),
    .B(_03128_));
 sg13g2_nand4_1 _11183_ (.B(_03112_),
    .C(_03116_),
    .A(_03128_),
    .Y(_03135_),
    .D(_03120_));
 sg13g2_nand4_1 _11184_ (.B(_03112_),
    .C(_03116_),
    .A(_03133_),
    .Y(_03136_),
    .D(_03120_));
 sg13g2_o21ai_1 _11185_ (.B1(_03118_),
    .Y(_03137_),
    .A1(_03133_),
    .A2(_03128_));
 sg13g2_and4_1 _11186_ (.A(_03134_),
    .B(_03135_),
    .C(_03136_),
    .D(_03137_),
    .X(_03138_));
 sg13g2_buf_2 _11187_ (.A(_03138_),
    .X(_03139_));
 sg13g2_buf_1 _11188_ (.A(\am_sdr0.cic0.comb2_in_del[16] ),
    .X(_03140_));
 sg13g2_xnor2_1 _11189_ (.Y(_03141_),
    .A(_02867_),
    .B(_03140_));
 sg13g2_xnor2_1 _11190_ (.Y(_03142_),
    .A(_03139_),
    .B(_03141_));
 sg13g2_mux2_1 _11191_ (.A0(_03132_),
    .A1(_03142_),
    .S(_02870_),
    .X(_03143_));
 sg13g2_nor2_1 _11192_ (.A(net127),
    .B(_03143_),
    .Y(_00238_));
 sg13g2_inv_1 _11193_ (.Y(_03144_),
    .A(\am_sdr0.cic0.comb2[17] ));
 sg13g2_inv_1 _11194_ (.Y(_03145_),
    .A(_03140_));
 sg13g2_a21o_1 _11195_ (.A2(_03139_),
    .A1(_03145_),
    .B1(_02867_),
    .X(_03146_));
 sg13g2_o21ai_1 _11196_ (.B1(_03146_),
    .Y(_03147_),
    .A1(_03145_),
    .A2(_03139_));
 sg13g2_xor2_1 _11197_ (.B(\am_sdr0.cic0.comb2_in_del[17] ),
    .A(_02869_),
    .X(_03148_));
 sg13g2_xnor2_1 _11198_ (.Y(_03149_),
    .A(_03147_),
    .B(_03148_));
 sg13g2_mux2_1 _11199_ (.A0(_03144_),
    .A1(_03149_),
    .S(_02870_),
    .X(_03150_));
 sg13g2_nor2_1 _11200_ (.A(net127),
    .B(_03150_),
    .Y(_00239_));
 sg13g2_inv_1 _11201_ (.Y(_03151_),
    .A(\am_sdr0.cic0.comb2_in_del[17] ));
 sg13g2_nor2_1 _11202_ (.A(_02869_),
    .B(_03151_),
    .Y(_03152_));
 sg13g2_a221oi_1 _11203_ (.B2(_03151_),
    .C1(_03139_),
    .B1(_02869_),
    .A1(_02867_),
    .Y(_03153_),
    .A2(_03145_));
 sg13g2_nand2b_1 _11204_ (.Y(_03154_),
    .B(_03140_),
    .A_N(_02867_));
 sg13g2_a21oi_1 _11205_ (.A1(_02869_),
    .A2(_03151_),
    .Y(_03155_),
    .B1(_03154_));
 sg13g2_nor3_1 _11206_ (.A(_03152_),
    .B(_03153_),
    .C(_03155_),
    .Y(_03156_));
 sg13g2_buf_1 _11207_ (.A(\am_sdr0.cic0.comb2_in_del[18] ),
    .X(_03157_));
 sg13g2_xnor2_1 _11208_ (.Y(_03158_),
    .A(_02887_),
    .B(_03157_));
 sg13g2_xnor2_1 _11209_ (.Y(_03159_),
    .A(_03156_),
    .B(_03158_));
 sg13g2_o21ai_1 _11210_ (.B1(net244),
    .Y(_03160_),
    .A1(\am_sdr0.cic0.comb2[18] ),
    .A2(net249));
 sg13g2_a21oi_1 _11211_ (.A1(net180),
    .A2(_03159_),
    .Y(_00240_),
    .B1(_03160_));
 sg13g2_nor2b_1 _11212_ (.A(_03157_),
    .B_N(_02887_),
    .Y(_03161_));
 sg13g2_nand2b_1 _11213_ (.Y(_03162_),
    .B(_03157_),
    .A_N(_02887_));
 sg13g2_o21ai_1 _11214_ (.B1(_03162_),
    .Y(_03163_),
    .A1(_03156_),
    .A2(_03161_));
 sg13g2_xor2_1 _11215_ (.B(\am_sdr0.cic0.comb2_in_del[19] ),
    .A(\am_sdr0.cic0.comb1[19] ),
    .X(_03164_));
 sg13g2_xnor2_1 _11216_ (.Y(_03165_),
    .A(_03163_),
    .B(_03164_));
 sg13g2_o21ai_1 _11217_ (.B1(net244),
    .Y(_03166_),
    .A1(\am_sdr0.cic0.comb2[19] ),
    .A2(_02721_));
 sg13g2_a21oi_1 _11218_ (.A1(_02718_),
    .A2(_03165_),
    .Y(_00241_),
    .B1(_03166_));
 sg13g2_xnor2_1 _11219_ (.Y(_03167_),
    .A(_02901_),
    .B(_03010_));
 sg13g2_xnor2_1 _11220_ (.Y(_03168_),
    .A(_03009_),
    .B(_03167_));
 sg13g2_buf_1 _11221_ (.A(\am_sdr0.cic0.comb2[1] ),
    .X(_03169_));
 sg13g2_nor2b_1 _11222_ (.A(net250),
    .B_N(_03169_),
    .Y(_03170_));
 sg13g2_a21oi_1 _11223_ (.A1(net171),
    .A2(_03168_),
    .Y(_03171_),
    .B1(_03170_));
 sg13g2_nor2_1 _11224_ (.A(net127),
    .B(_03171_),
    .Y(_00242_));
 sg13g2_a21oi_1 _11225_ (.A1(_03009_),
    .A2(_03011_),
    .Y(_03172_),
    .B1(_03012_));
 sg13g2_xor2_1 _11226_ (.B(_03007_),
    .A(_02906_),
    .X(_03173_));
 sg13g2_xnor2_1 _11227_ (.Y(_03174_),
    .A(_03172_),
    .B(_03173_));
 sg13g2_buf_1 _11228_ (.A(\am_sdr0.cic0.comb2[2] ),
    .X(_03175_));
 sg13g2_nor2b_1 _11229_ (.A(net250),
    .B_N(_03175_),
    .Y(_03176_));
 sg13g2_a21oi_1 _11230_ (.A1(net171),
    .A2(_03174_),
    .Y(_03177_),
    .B1(_03176_));
 sg13g2_nor2_1 _11231_ (.A(net127),
    .B(_03177_),
    .Y(_00243_));
 sg13g2_nor2_1 _11232_ (.A(_03008_),
    .B(_03014_),
    .Y(_03178_));
 sg13g2_xnor2_1 _11233_ (.Y(_03179_),
    .A(_02912_),
    .B(\am_sdr0.cic0.comb2_in_del[3] ));
 sg13g2_xnor2_1 _11234_ (.Y(_03180_),
    .A(_03178_),
    .B(_03179_));
 sg13g2_buf_1 _11235_ (.A(\am_sdr0.cic0.comb2[3] ),
    .X(_03181_));
 sg13g2_nor2b_1 _11236_ (.A(net250),
    .B_N(_03181_),
    .Y(_03182_));
 sg13g2_a21oi_1 _11237_ (.A1(net171),
    .A2(_03180_),
    .Y(_03183_),
    .B1(_03182_));
 sg13g2_nor2_1 _11238_ (.A(net127),
    .B(_03183_),
    .Y(_00244_));
 sg13g2_buf_1 _11239_ (.A(\am_sdr0.cic0.comb2[4] ),
    .X(_03184_));
 sg13g2_nand2_1 _11240_ (.Y(_03185_),
    .A(_03020_),
    .B(_03023_));
 sg13g2_xnor2_1 _11241_ (.Y(_03186_),
    .A(_03019_),
    .B(_03185_));
 sg13g2_nand2_1 _11242_ (.Y(_03187_),
    .A(net243),
    .B(_03186_));
 sg13g2_o21ai_1 _11243_ (.B1(_03187_),
    .Y(_03188_),
    .A1(_03184_),
    .A2(net247));
 sg13g2_nor2_1 _11244_ (.A(net127),
    .B(_03188_),
    .Y(_00245_));
 sg13g2_nand2_1 _11245_ (.Y(_03189_),
    .A(_03019_),
    .B(_03020_));
 sg13g2_nand2_1 _11246_ (.Y(_03190_),
    .A(_03189_),
    .B(_03023_));
 sg13g2_xor2_1 _11247_ (.B(_03021_),
    .A(_02923_),
    .X(_03191_));
 sg13g2_xnor2_1 _11248_ (.Y(_03192_),
    .A(_03190_),
    .B(_03191_));
 sg13g2_nand2_1 _11249_ (.Y(_03193_),
    .A(net243),
    .B(_03192_));
 sg13g2_o21ai_1 _11250_ (.B1(_03193_),
    .Y(_03194_),
    .A1(\am_sdr0.cic0.comb2[5] ),
    .A2(net247));
 sg13g2_nor2_1 _11251_ (.A(net127),
    .B(_03194_),
    .Y(_00246_));
 sg13g2_buf_1 _11252_ (.A(net259),
    .X(_03195_));
 sg13g2_buf_1 _11253_ (.A(_03195_),
    .X(_03196_));
 sg13g2_buf_1 _11254_ (.A(\am_sdr0.cic0.comb2[6] ),
    .X(_03197_));
 sg13g2_nor2_1 _11255_ (.A(_03021_),
    .B(_03190_),
    .Y(_03198_));
 sg13g2_nand2_1 _11256_ (.Y(_03199_),
    .A(_03021_),
    .B(_03190_));
 sg13g2_o21ai_1 _11257_ (.B1(_03199_),
    .Y(_03200_),
    .A1(_02923_),
    .A2(_03198_));
 sg13g2_buf_1 _11258_ (.A(_03200_),
    .X(_03201_));
 sg13g2_xor2_1 _11259_ (.B(_03033_),
    .A(_02929_),
    .X(_03202_));
 sg13g2_xnor2_1 _11260_ (.Y(_03203_),
    .A(_03201_),
    .B(_03202_));
 sg13g2_nand2_1 _11261_ (.Y(_03204_),
    .A(net243),
    .B(_03203_));
 sg13g2_o21ai_1 _11262_ (.B1(_03204_),
    .Y(_03205_),
    .A1(_03197_),
    .A2(net247));
 sg13g2_nor2_1 _11263_ (.A(net126),
    .B(_03205_),
    .Y(_00247_));
 sg13g2_nor2_1 _11264_ (.A(_03033_),
    .B(_03201_),
    .Y(_03206_));
 sg13g2_nand2_1 _11265_ (.Y(_03207_),
    .A(_03033_),
    .B(_03201_));
 sg13g2_o21ai_1 _11266_ (.B1(_03207_),
    .Y(_03208_),
    .A1(_02929_),
    .A2(_03206_));
 sg13g2_buf_1 _11267_ (.A(_03208_),
    .X(_03209_));
 sg13g2_nand2_1 _11268_ (.Y(_03210_),
    .A(_03028_),
    .B(_03040_));
 sg13g2_xnor2_1 _11269_ (.Y(_03211_),
    .A(_03209_),
    .B(_03210_));
 sg13g2_nand2_1 _11270_ (.Y(_03212_),
    .A(net243),
    .B(_03211_));
 sg13g2_o21ai_1 _11271_ (.B1(_03212_),
    .Y(_03213_),
    .A1(\am_sdr0.cic0.comb2[7] ),
    .A2(net247));
 sg13g2_nor2_1 _11272_ (.A(net126),
    .B(_03213_),
    .Y(_00248_));
 sg13g2_nand2_1 _11273_ (.Y(_03214_),
    .A(_03026_),
    .B(_03209_));
 sg13g2_nor2_1 _11274_ (.A(_03026_),
    .B(_03209_),
    .Y(_03215_));
 sg13g2_a21oi_1 _11275_ (.A1(_02937_),
    .A2(_03214_),
    .Y(_03216_),
    .B1(_03215_));
 sg13g2_xor2_1 _11276_ (.B(_03029_),
    .A(_02943_),
    .X(_03217_));
 sg13g2_xnor2_1 _11277_ (.Y(_03218_),
    .A(_03216_),
    .B(_03217_));
 sg13g2_nand2_1 _11278_ (.Y(_03219_),
    .A(net243),
    .B(_03218_));
 sg13g2_o21ai_1 _11279_ (.B1(_03219_),
    .Y(_03220_),
    .A1(\am_sdr0.cic0.comb2[8] ),
    .A2(net247));
 sg13g2_nor2_1 _11280_ (.A(net126),
    .B(_03220_),
    .Y(_00249_));
 sg13g2_nor2_1 _11281_ (.A(_03037_),
    .B(_03045_),
    .Y(_03221_));
 sg13g2_xnor2_1 _11282_ (.Y(_03222_),
    .A(_02948_),
    .B(_03046_));
 sg13g2_xnor2_1 _11283_ (.Y(_03223_),
    .A(_03221_),
    .B(_03222_));
 sg13g2_buf_1 _11284_ (.A(\am_sdr0.cic0.comb2[9] ),
    .X(_03224_));
 sg13g2_nor2b_1 _11285_ (.A(net250),
    .B_N(_03224_),
    .Y(_03225_));
 sg13g2_a21oi_1 _11286_ (.A1(net171),
    .A2(_03223_),
    .Y(_03226_),
    .B1(_03225_));
 sg13g2_nor2_1 _11287_ (.A(net126),
    .B(_03226_),
    .Y(_00250_));
 sg13g2_buf_1 _11288_ (.A(_02728_),
    .X(_03227_));
 sg13g2_nand2_1 _11289_ (.Y(_03228_),
    .A(_02720_),
    .B(net170));
 sg13g2_nand2_1 _11290_ (.Y(_03229_),
    .A(\am_sdr0.cic0.comb2_in_del[0] ),
    .B(net172));
 sg13g2_a21oi_1 _11291_ (.A1(_03228_),
    .A2(_03229_),
    .Y(_00251_),
    .B1(net128));
 sg13g2_nand2_1 _11292_ (.Y(_03230_),
    .A(_02723_),
    .B(net170));
 sg13g2_buf_1 _11293_ (.A(_02785_),
    .X(_03231_));
 sg13g2_nand2_1 _11294_ (.Y(_03232_),
    .A(_03051_),
    .B(net169));
 sg13g2_a21oi_1 _11295_ (.A1(_03230_),
    .A2(_03232_),
    .Y(_00252_),
    .B1(net128));
 sg13g2_nand2_1 _11296_ (.Y(_03233_),
    .A(_02782_),
    .B(net170));
 sg13g2_nand2_1 _11297_ (.Y(_03234_),
    .A(_03061_),
    .B(net169));
 sg13g2_a21oi_1 _11298_ (.A1(_03233_),
    .A2(_03234_),
    .Y(_00253_),
    .B1(net128));
 sg13g2_nand2_1 _11299_ (.Y(_03235_),
    .A(_02797_),
    .B(net170));
 sg13g2_nand2_1 _11300_ (.Y(_03236_),
    .A(_03091_),
    .B(net169));
 sg13g2_a21oi_1 _11301_ (.A1(_03235_),
    .A2(_03236_),
    .Y(_00254_),
    .B1(_02992_));
 sg13g2_nand2_1 _11302_ (.Y(_03237_),
    .A(_02810_),
    .B(net170));
 sg13g2_nand2_1 _11303_ (.Y(_03238_),
    .A(\am_sdr0.cic0.comb2_in_del[13] ),
    .B(net169));
 sg13g2_a21oi_1 _11304_ (.A1(_03237_),
    .A2(_03238_),
    .Y(_00255_),
    .B1(_02992_));
 sg13g2_nand2_1 _11305_ (.Y(_03239_),
    .A(_02823_),
    .B(net170));
 sg13g2_nand2_1 _11306_ (.Y(_03240_),
    .A(\am_sdr0.cic0.comb2_in_del[14] ),
    .B(net169));
 sg13g2_buf_1 _11307_ (.A(_02779_),
    .X(_03241_));
 sg13g2_a21oi_1 _11308_ (.A1(_03239_),
    .A2(_03240_),
    .Y(_00256_),
    .B1(_03241_));
 sg13g2_nand2_1 _11309_ (.Y(_03242_),
    .A(_02840_),
    .B(net170));
 sg13g2_nand2_1 _11310_ (.Y(_03243_),
    .A(_03128_),
    .B(net169));
 sg13g2_a21oi_1 _11311_ (.A1(_03242_),
    .A2(_03243_),
    .Y(_00257_),
    .B1(net125));
 sg13g2_nand2_1 _11312_ (.Y(_03244_),
    .A(_02867_),
    .B(net170));
 sg13g2_nand2_1 _11313_ (.Y(_03245_),
    .A(_03140_),
    .B(net169));
 sg13g2_a21oi_1 _11314_ (.A1(_03244_),
    .A2(_03245_),
    .Y(_00258_),
    .B1(net125));
 sg13g2_nand2_1 _11315_ (.Y(_03246_),
    .A(_02869_),
    .B(_03227_));
 sg13g2_nand2_1 _11316_ (.Y(_03247_),
    .A(\am_sdr0.cic0.comb2_in_del[17] ),
    .B(net169));
 sg13g2_a21oi_1 _11317_ (.A1(_03246_),
    .A2(_03247_),
    .Y(_00259_),
    .B1(net125));
 sg13g2_nand2_1 _11318_ (.Y(_03248_),
    .A(_02887_),
    .B(_03227_));
 sg13g2_nand2_1 _11319_ (.Y(_03249_),
    .A(_03157_),
    .B(_03231_));
 sg13g2_a21oi_1 _11320_ (.A1(_03248_),
    .A2(_03249_),
    .Y(_00260_),
    .B1(_03241_));
 sg13g2_buf_1 _11321_ (.A(_02728_),
    .X(_03250_));
 sg13g2_nand2_1 _11322_ (.Y(_03251_),
    .A(\am_sdr0.cic0.comb1[19] ),
    .B(_03250_));
 sg13g2_nand2_1 _11323_ (.Y(_03252_),
    .A(\am_sdr0.cic0.comb2_in_del[19] ),
    .B(_03231_));
 sg13g2_a21oi_1 _11324_ (.A1(_03251_),
    .A2(_03252_),
    .Y(_00261_),
    .B1(net125));
 sg13g2_nand2_1 _11325_ (.Y(_03253_),
    .A(_02901_),
    .B(_03250_));
 sg13g2_buf_1 _11326_ (.A(_02785_),
    .X(_03254_));
 sg13g2_nand2_1 _11327_ (.Y(_03255_),
    .A(_03010_),
    .B(net167));
 sg13g2_a21oi_1 _11328_ (.A1(_03253_),
    .A2(_03255_),
    .Y(_00262_),
    .B1(net125));
 sg13g2_nand2_1 _11329_ (.Y(_03256_),
    .A(_02906_),
    .B(net168));
 sg13g2_nand2_1 _11330_ (.Y(_03257_),
    .A(_03007_),
    .B(_03254_));
 sg13g2_a21oi_1 _11331_ (.A1(_03256_),
    .A2(_03257_),
    .Y(_00263_),
    .B1(net125));
 sg13g2_nand2_1 _11332_ (.Y(_03258_),
    .A(_02912_),
    .B(net168));
 sg13g2_nand2_1 _11333_ (.Y(_03259_),
    .A(\am_sdr0.cic0.comb2_in_del[3] ),
    .B(_03254_));
 sg13g2_a21oi_1 _11334_ (.A1(_03258_),
    .A2(_03259_),
    .Y(_00264_),
    .B1(net125));
 sg13g2_nand2_1 _11335_ (.Y(_03260_),
    .A(_02918_),
    .B(net168));
 sg13g2_nand2_1 _11336_ (.Y(_03261_),
    .A(\am_sdr0.cic0.comb2_in_del[4] ),
    .B(net167));
 sg13g2_a21oi_1 _11337_ (.A1(_03260_),
    .A2(_03261_),
    .Y(_00265_),
    .B1(net125));
 sg13g2_nand2_1 _11338_ (.Y(_03262_),
    .A(_02923_),
    .B(net168));
 sg13g2_nand2_1 _11339_ (.Y(_03263_),
    .A(_03021_),
    .B(net167));
 sg13g2_buf_1 _11340_ (.A(_02779_),
    .X(_03264_));
 sg13g2_a21oi_1 _11341_ (.A1(_03262_),
    .A2(_03263_),
    .Y(_00266_),
    .B1(net124));
 sg13g2_nand2_1 _11342_ (.Y(_03265_),
    .A(_02929_),
    .B(net168));
 sg13g2_nand2_1 _11343_ (.Y(_03266_),
    .A(_03033_),
    .B(net167));
 sg13g2_a21oi_1 _11344_ (.A1(_03265_),
    .A2(_03266_),
    .Y(_00267_),
    .B1(net124));
 sg13g2_nand2_1 _11345_ (.Y(_03267_),
    .A(_02937_),
    .B(net168));
 sg13g2_nand2_1 _11346_ (.Y(_03268_),
    .A(_03026_),
    .B(net167));
 sg13g2_a21oi_1 _11347_ (.A1(_03267_),
    .A2(_03268_),
    .Y(_00268_),
    .B1(net124));
 sg13g2_nand2_1 _11348_ (.Y(_03269_),
    .A(_02943_),
    .B(net168));
 sg13g2_nand2_1 _11349_ (.Y(_03270_),
    .A(_03029_),
    .B(net167));
 sg13g2_a21oi_1 _11350_ (.A1(_03269_),
    .A2(_03270_),
    .Y(_00269_),
    .B1(net124));
 sg13g2_nand2_1 _11351_ (.Y(_03271_),
    .A(_02948_),
    .B(net168));
 sg13g2_nand2_1 _11352_ (.Y(_03272_),
    .A(_03046_),
    .B(net167));
 sg13g2_a21oi_1 _11353_ (.A1(_03271_),
    .A2(_03272_),
    .Y(_00270_),
    .B1(_03264_));
 sg13g2_inv_1 _11354_ (.Y(_03273_),
    .A(\am_sdr0.cic0.comb3_in_del[9] ));
 sg13g2_inv_1 _11355_ (.Y(_03274_),
    .A(\am_sdr0.cic0.comb2[7] ));
 sg13g2_inv_1 _11356_ (.Y(_03275_),
    .A(\am_sdr0.cic0.comb2[5] ));
 sg13g2_xnor2_1 _11357_ (.Y(_03276_),
    .A(\am_sdr0.cic0.comb3_in_del[3] ),
    .B(_03181_));
 sg13g2_nand2b_1 _11358_ (.Y(_03277_),
    .B(\am_sdr0.cic0.comb3_in_del[4] ),
    .A_N(_03184_));
 sg13g2_xnor2_1 _11359_ (.Y(_03278_),
    .A(\am_sdr0.cic0.comb3_in_del[2] ),
    .B(_03175_));
 sg13g2_nand2b_1 _11360_ (.Y(_03279_),
    .B(\am_sdr0.cic0.comb3_in_del[0] ),
    .A_N(\am_sdr0.cic0.comb2[0] ));
 sg13g2_nor2_1 _11361_ (.A(_03169_),
    .B(_03279_),
    .Y(_03280_));
 sg13g2_nand2_1 _11362_ (.Y(_03281_),
    .A(_03169_),
    .B(_03279_));
 sg13g2_o21ai_1 _11363_ (.B1(_03281_),
    .Y(_03282_),
    .A1(\am_sdr0.cic0.comb3_in_del[1] ),
    .A2(_03280_));
 sg13g2_nand4_1 _11364_ (.B(_03277_),
    .C(_03278_),
    .A(_03276_),
    .Y(_03283_),
    .D(_03282_));
 sg13g2_nor2b_1 _11365_ (.A(\am_sdr0.cic0.comb3_in_del[4] ),
    .B_N(_03184_),
    .Y(_03284_));
 sg13g2_nor2b_1 _11366_ (.A(\am_sdr0.cic0.comb3_in_del[2] ),
    .B_N(_03175_),
    .Y(_03285_));
 sg13g2_nor2_1 _11367_ (.A(_03181_),
    .B(_03285_),
    .Y(_03286_));
 sg13g2_nand2_1 _11368_ (.Y(_03287_),
    .A(_03181_),
    .B(_03285_));
 sg13g2_o21ai_1 _11369_ (.B1(_03287_),
    .Y(_03288_),
    .A1(\am_sdr0.cic0.comb3_in_del[3] ),
    .A2(_03286_));
 sg13g2_o21ai_1 _11370_ (.B1(_03277_),
    .Y(_03289_),
    .A1(_03284_),
    .A2(_03288_));
 sg13g2_a22oi_1 _11371_ (.Y(_03290_),
    .B1(_03283_),
    .B2(_03289_),
    .A2(_03275_),
    .A1(\am_sdr0.cic0.comb3_in_del[5] ));
 sg13g2_nand2b_1 _11372_ (.Y(_03291_),
    .B(_03197_),
    .A_N(\am_sdr0.cic0.comb3_in_del[6] ));
 sg13g2_o21ai_1 _11373_ (.B1(_03291_),
    .Y(_03292_),
    .A1(\am_sdr0.cic0.comb3_in_del[5] ),
    .A2(_03275_));
 sg13g2_nand2b_1 _11374_ (.Y(_03293_),
    .B(\am_sdr0.cic0.comb3_in_del[6] ),
    .A_N(_03197_));
 sg13g2_o21ai_1 _11375_ (.B1(_03293_),
    .Y(_03294_),
    .A1(_03290_),
    .A2(_03292_));
 sg13g2_o21ai_1 _11376_ (.B1(_03294_),
    .Y(_03295_),
    .A1(\am_sdr0.cic0.comb3_in_del[7] ),
    .A2(_03274_));
 sg13g2_inv_1 _11377_ (.Y(_03296_),
    .A(\am_sdr0.cic0.comb2[8] ));
 sg13g2_a22oi_1 _11378_ (.Y(_03297_),
    .B1(\am_sdr0.cic0.comb3_in_del[7] ),
    .B2(_03274_),
    .A2(_03296_),
    .A1(\am_sdr0.cic0.comb3_in_del[8] ));
 sg13g2_nor2_1 _11379_ (.A(\am_sdr0.cic0.comb3_in_del[8] ),
    .B(_03296_),
    .Y(_03298_));
 sg13g2_a221oi_1 _11380_ (.B2(_03297_),
    .C1(_03298_),
    .B1(_03295_),
    .A1(_03273_),
    .Y(_03299_),
    .A2(_03224_));
 sg13g2_nand2b_1 _11381_ (.Y(_03300_),
    .B(\am_sdr0.cic0.comb3_in_del[10] ),
    .A_N(_03056_));
 sg13g2_o21ai_1 _11382_ (.B1(_03300_),
    .Y(_03301_),
    .A1(_03273_),
    .A2(_03224_));
 sg13g2_nand2b_1 _11383_ (.Y(_03302_),
    .B(_03056_),
    .A_N(\am_sdr0.cic0.comb3_in_del[10] ));
 sg13g2_o21ai_1 _11384_ (.B1(_03302_),
    .Y(_03303_),
    .A1(_03299_),
    .A2(_03301_));
 sg13g2_buf_1 _11385_ (.A(_03303_),
    .X(_03304_));
 sg13g2_inv_1 _11386_ (.Y(_03305_),
    .A(\am_sdr0.cic0.comb3_in_del[11] ));
 sg13g2_o21ai_1 _11387_ (.B1(_03305_),
    .Y(_03306_),
    .A1(_03059_),
    .A2(_03304_));
 sg13g2_nand2_1 _11388_ (.Y(_03307_),
    .A(_03059_),
    .B(_03304_));
 sg13g2_nand2_1 _11389_ (.Y(_03308_),
    .A(_03306_),
    .B(_03307_));
 sg13g2_buf_1 _11390_ (.A(\am_sdr0.cic0.comb3_in_del[12] ),
    .X(_03309_));
 sg13g2_xor2_1 _11391_ (.B(_03309_),
    .A(_03066_),
    .X(_03310_));
 sg13g2_xor2_1 _11392_ (.B(_03310_),
    .A(_03308_),
    .X(_03311_));
 sg13g2_nor2_1 _11393_ (.A(net248),
    .B(_03311_),
    .Y(_03312_));
 sg13g2_a21oi_1 _11394_ (.A1(_02726_),
    .A2(\am_sdr0.cic0.comb3[12] ),
    .Y(_03313_),
    .B1(_03312_));
 sg13g2_nor2_1 _11395_ (.A(_03196_),
    .B(_03313_),
    .Y(_00271_));
 sg13g2_nand3_1 _11396_ (.B(_03306_),
    .C(_03307_),
    .A(_03309_),
    .Y(_03314_));
 sg13g2_a21oi_1 _11397_ (.A1(_03306_),
    .A2(_03307_),
    .Y(_03315_),
    .B1(_03309_));
 sg13g2_a21oi_2 _11398_ (.B1(_03315_),
    .Y(_03316_),
    .A2(_03314_),
    .A1(_03066_));
 sg13g2_buf_2 _11399_ (.A(\am_sdr0.cic0.comb3_in_del[13] ),
    .X(_03317_));
 sg13g2_xnor2_1 _11400_ (.Y(_03318_),
    .A(_03097_),
    .B(_03317_));
 sg13g2_xnor2_1 _11401_ (.Y(_03319_),
    .A(_03316_),
    .B(_03318_));
 sg13g2_nor2b_1 _11402_ (.A(net250),
    .B_N(\am_sdr0.cic0.comb3[13] ),
    .Y(_03320_));
 sg13g2_a21oi_1 _11403_ (.A1(net171),
    .A2(_03319_),
    .Y(_03321_),
    .B1(_03320_));
 sg13g2_nor2_1 _11404_ (.A(net126),
    .B(_03321_),
    .Y(_00272_));
 sg13g2_nor2b_1 _11405_ (.A(_02717_),
    .B_N(\am_sdr0.cic0.comb3[14] ),
    .Y(_03322_));
 sg13g2_nand2_1 _11406_ (.Y(_03323_),
    .A(_03317_),
    .B(_03316_));
 sg13g2_inv_1 _11407_ (.Y(_03324_),
    .A(_03097_));
 sg13g2_o21ai_1 _11408_ (.B1(_03324_),
    .Y(_03325_),
    .A1(_03317_),
    .A2(_03316_));
 sg13g2_buf_1 _11409_ (.A(\am_sdr0.cic0.comb3_in_del[14] ),
    .X(_03326_));
 sg13g2_xnor2_1 _11410_ (.Y(_03327_),
    .A(_03106_),
    .B(_03326_));
 sg13g2_nor2_1 _11411_ (.A(_02785_),
    .B(_03327_),
    .Y(_03328_));
 sg13g2_and3_1 _11412_ (.X(_03329_),
    .A(_03323_),
    .B(_03325_),
    .C(_03328_));
 sg13g2_nand2_1 _11413_ (.Y(_03330_),
    .A(_02716_),
    .B(_03327_));
 sg13g2_a21oi_1 _11414_ (.A1(_03323_),
    .A2(_03325_),
    .Y(_03331_),
    .B1(_03330_));
 sg13g2_nor3_1 _11415_ (.A(_03322_),
    .B(_03329_),
    .C(_03331_),
    .Y(_03332_));
 sg13g2_nor2_1 _11416_ (.A(net126),
    .B(_03332_),
    .Y(_00273_));
 sg13g2_inv_1 _11417_ (.Y(_03333_),
    .A(_03326_));
 sg13g2_nand2_1 _11418_ (.Y(_03334_),
    .A(_03305_),
    .B(_03059_));
 sg13g2_inv_1 _11419_ (.Y(_03335_),
    .A(_03066_));
 sg13g2_o21ai_1 _11420_ (.B1(_03335_),
    .Y(_03336_),
    .A1(_03309_),
    .A2(_03334_));
 sg13g2_nand2_1 _11421_ (.Y(_03337_),
    .A(_03309_),
    .B(_03334_));
 sg13g2_a22oi_1 _11422_ (.Y(_03338_),
    .B1(_03336_),
    .B2(_03337_),
    .A2(_03333_),
    .A1(_03106_));
 sg13g2_o21ai_1 _11423_ (.B1(_03338_),
    .Y(_03339_),
    .A1(_03324_),
    .A2(_03317_));
 sg13g2_xor2_1 _11424_ (.B(_03059_),
    .A(\am_sdr0.cic0.comb3_in_del[11] ),
    .X(_03340_));
 sg13g2_o21ai_1 _11425_ (.B1(_03338_),
    .Y(_03341_),
    .A1(_03310_),
    .A2(_03340_));
 sg13g2_inv_1 _11426_ (.Y(_03342_),
    .A(_03341_));
 sg13g2_a21o_1 _11427_ (.A2(_03317_),
    .A1(_03324_),
    .B1(_03326_),
    .X(_03343_));
 sg13g2_inv_1 _11428_ (.Y(_03344_),
    .A(_03106_));
 sg13g2_nand2_1 _11429_ (.Y(_03345_),
    .A(_03317_),
    .B(_03326_));
 sg13g2_a21oi_1 _11430_ (.A1(_03341_),
    .A2(_03345_),
    .Y(_03346_),
    .B1(_03097_));
 sg13g2_a221oi_1 _11431_ (.B2(_03344_),
    .C1(_03346_),
    .B1(_03343_),
    .A1(_03317_),
    .Y(_03347_),
    .A2(_03342_));
 sg13g2_o21ai_1 _11432_ (.B1(_03347_),
    .Y(_03348_),
    .A1(_03304_),
    .A2(_03339_));
 sg13g2_buf_1 _11433_ (.A(_03348_),
    .X(_03349_));
 sg13g2_buf_1 _11434_ (.A(\am_sdr0.cic0.comb3_in_del[15] ),
    .X(_03350_));
 sg13g2_xor2_1 _11435_ (.B(_03350_),
    .A(_03125_),
    .X(_03351_));
 sg13g2_xnor2_1 _11436_ (.Y(_03352_),
    .A(_03349_),
    .B(_03351_));
 sg13g2_nand2_1 _11437_ (.Y(_03353_),
    .A(_03098_),
    .B(_03352_));
 sg13g2_o21ai_1 _11438_ (.B1(_03353_),
    .Y(_03354_),
    .A1(_02721_),
    .A2(\am_sdr0.cic0.comb3[15] ));
 sg13g2_nor2_1 _11439_ (.A(net126),
    .B(_03354_),
    .Y(_00274_));
 sg13g2_nand2_1 _11440_ (.Y(_03355_),
    .A(_03350_),
    .B(_03349_));
 sg13g2_o21ai_1 _11441_ (.B1(_03126_),
    .Y(_03356_),
    .A1(_03350_),
    .A2(_03349_));
 sg13g2_nand2_1 _11442_ (.Y(_03357_),
    .A(_03355_),
    .B(_03356_));
 sg13g2_buf_1 _11443_ (.A(\am_sdr0.cic0.comb3_in_del[16] ),
    .X(_03358_));
 sg13g2_xor2_1 _11444_ (.B(_03358_),
    .A(\am_sdr0.cic0.comb2[16] ),
    .X(_03359_));
 sg13g2_xnor2_1 _11445_ (.Y(_03360_),
    .A(_03357_),
    .B(_03359_));
 sg13g2_nand2_1 _11446_ (.Y(_03361_),
    .A(_03098_),
    .B(_03360_));
 sg13g2_o21ai_1 _11447_ (.B1(_03361_),
    .Y(_03362_),
    .A1(net249),
    .A2(\am_sdr0.cic0.comb3[16] ));
 sg13g2_nor2_1 _11448_ (.A(_03196_),
    .B(_03362_),
    .Y(_00275_));
 sg13g2_a221oi_1 _11449_ (.B2(_03358_),
    .C1(_03349_),
    .B1(_03132_),
    .A1(_03126_),
    .Y(_03363_),
    .A2(_03350_));
 sg13g2_buf_1 _11450_ (.A(_03363_),
    .X(_03364_));
 sg13g2_nand2b_1 _11451_ (.Y(_03365_),
    .B(_03125_),
    .A_N(_03350_));
 sg13g2_a21o_1 _11452_ (.A2(_03358_),
    .A1(_03132_),
    .B1(_03365_),
    .X(_03366_));
 sg13g2_o21ai_1 _11453_ (.B1(_03366_),
    .Y(_03367_),
    .A1(_03132_),
    .A2(_03358_));
 sg13g2_nor2_1 _11454_ (.A(_03364_),
    .B(_03367_),
    .Y(_03368_));
 sg13g2_xor2_1 _11455_ (.B(\am_sdr0.cic0.comb3_in_del[17] ),
    .A(\am_sdr0.cic0.comb2[17] ),
    .X(_03369_));
 sg13g2_xnor2_1 _11456_ (.Y(_03370_),
    .A(_03368_),
    .B(_03369_));
 sg13g2_nand2_1 _11457_ (.Y(_03371_),
    .A(net243),
    .B(_03370_));
 sg13g2_o21ai_1 _11458_ (.B1(_03371_),
    .Y(_03372_),
    .A1(net249),
    .A2(\am_sdr0.cic0.comb3[17] ));
 sg13g2_nor2_1 _11459_ (.A(net126),
    .B(_03372_),
    .Y(_00276_));
 sg13g2_buf_1 _11460_ (.A(_03195_),
    .X(_03373_));
 sg13g2_inv_1 _11461_ (.Y(_03374_),
    .A(\am_sdr0.cic0.comb3_in_del[17] ));
 sg13g2_o21ai_1 _11462_ (.B1(_03374_),
    .Y(_03375_),
    .A1(_03364_),
    .A2(_03367_));
 sg13g2_nor3_1 _11463_ (.A(_03374_),
    .B(_03364_),
    .C(_03367_),
    .Y(_03376_));
 sg13g2_a21oi_1 _11464_ (.A1(_03144_),
    .A2(_03375_),
    .Y(_03377_),
    .B1(_03376_));
 sg13g2_inv_1 _11465_ (.Y(_03378_),
    .A(\am_sdr0.cic0.comb2[18] ));
 sg13g2_nor2_1 _11466_ (.A(_03378_),
    .B(\am_sdr0.cic0.comb3_in_del[18] ),
    .Y(_03379_));
 sg13g2_nand2_1 _11467_ (.Y(_03380_),
    .A(_03378_),
    .B(\am_sdr0.cic0.comb3_in_del[18] ));
 sg13g2_nand2b_1 _11468_ (.Y(_03381_),
    .B(_03380_),
    .A_N(_03379_));
 sg13g2_xnor2_1 _11469_ (.Y(_03382_),
    .A(_03377_),
    .B(_03381_));
 sg13g2_nor2b_1 _11470_ (.A(_02717_),
    .B_N(\am_sdr0.cic0.comb3[18] ),
    .Y(_03383_));
 sg13g2_a21oi_1 _11471_ (.A1(net171),
    .A2(_03382_),
    .Y(_03384_),
    .B1(_03383_));
 sg13g2_nor2_1 _11472_ (.A(_03373_),
    .B(_03384_),
    .Y(_00277_));
 sg13g2_xnor2_1 _11473_ (.Y(_03385_),
    .A(\am_sdr0.cic0.comb2[19] ),
    .B(\am_sdr0.cic0.comb3_in_del[19] ));
 sg13g2_nor2_1 _11474_ (.A(net310),
    .B(_02724_),
    .Y(_00396_));
 sg13g2_a21o_1 _11475_ (.A2(_03380_),
    .A1(_03377_),
    .B1(_03379_),
    .X(_03386_));
 sg13g2_nand3b_1 _11476_ (.B(_00396_),
    .C(_03386_),
    .Y(_03387_),
    .A_N(_03385_));
 sg13g2_nand2_1 _11477_ (.Y(_03388_),
    .A(_00396_),
    .B(_03385_));
 sg13g2_or2_1 _11478_ (.X(_03389_),
    .B(_03388_),
    .A(_03386_));
 sg13g2_nand3_1 _11479_ (.B(net248),
    .C(\am_sdr0.cic0.comb3[19] ),
    .A(net253),
    .Y(_03390_));
 sg13g2_nand3_1 _11480_ (.B(_03389_),
    .C(_03390_),
    .A(_03387_),
    .Y(_00278_));
 sg13g2_buf_1 _11481_ (.A(_02728_),
    .X(_03391_));
 sg13g2_nand2_1 _11482_ (.Y(_03392_),
    .A(\am_sdr0.cic0.comb2[0] ),
    .B(net166));
 sg13g2_nand2_1 _11483_ (.Y(_03393_),
    .A(\am_sdr0.cic0.comb3_in_del[0] ),
    .B(net167));
 sg13g2_a21oi_1 _11484_ (.A1(_03392_),
    .A2(_03393_),
    .Y(_00279_),
    .B1(net124));
 sg13g2_nand2_1 _11485_ (.Y(_03394_),
    .A(_03056_),
    .B(net166));
 sg13g2_buf_1 _11486_ (.A(_02785_),
    .X(_03395_));
 sg13g2_nand2_1 _11487_ (.Y(_03396_),
    .A(\am_sdr0.cic0.comb3_in_del[10] ),
    .B(net165));
 sg13g2_a21oi_1 _11488_ (.A1(_03394_),
    .A2(_03396_),
    .Y(_00280_),
    .B1(net124));
 sg13g2_nand2_1 _11489_ (.Y(_03397_),
    .A(_03059_),
    .B(net166));
 sg13g2_nand2_1 _11490_ (.Y(_03398_),
    .A(\am_sdr0.cic0.comb3_in_del[11] ),
    .B(net165));
 sg13g2_a21oi_1 _11491_ (.A1(_03397_),
    .A2(_03398_),
    .Y(_00281_),
    .B1(net124));
 sg13g2_nand2_1 _11492_ (.Y(_03399_),
    .A(_03066_),
    .B(net166));
 sg13g2_nand2_1 _11493_ (.Y(_03400_),
    .A(_03309_),
    .B(net165));
 sg13g2_a21oi_1 _11494_ (.A1(_03399_),
    .A2(_03400_),
    .Y(_00282_),
    .B1(_03264_));
 sg13g2_nand2_1 _11495_ (.Y(_03401_),
    .A(_03097_),
    .B(net166));
 sg13g2_nand2_1 _11496_ (.Y(_03402_),
    .A(_03317_),
    .B(net165));
 sg13g2_a21oi_1 _11497_ (.A1(_03401_),
    .A2(_03402_),
    .Y(_00283_),
    .B1(net124));
 sg13g2_nand2_1 _11498_ (.Y(_03403_),
    .A(_03106_),
    .B(net166));
 sg13g2_nand2_1 _11499_ (.Y(_03404_),
    .A(_03326_),
    .B(_03395_));
 sg13g2_buf_1 _11500_ (.A(_02779_),
    .X(_03405_));
 sg13g2_a21oi_1 _11501_ (.A1(_03403_),
    .A2(_03404_),
    .Y(_00284_),
    .B1(net122));
 sg13g2_nand2_1 _11502_ (.Y(_03406_),
    .A(_03125_),
    .B(net166));
 sg13g2_nand2_1 _11503_ (.Y(_03407_),
    .A(_03350_),
    .B(net165));
 sg13g2_a21oi_1 _11504_ (.A1(_03406_),
    .A2(_03407_),
    .Y(_00285_),
    .B1(net122));
 sg13g2_nand2_1 _11505_ (.Y(_03408_),
    .A(\am_sdr0.cic0.comb2[16] ),
    .B(net166));
 sg13g2_nand2_1 _11506_ (.Y(_03409_),
    .A(_03358_),
    .B(net165));
 sg13g2_a21oi_1 _11507_ (.A1(_03408_),
    .A2(_03409_),
    .Y(_00286_),
    .B1(net122));
 sg13g2_nand2_1 _11508_ (.Y(_03410_),
    .A(\am_sdr0.cic0.comb2[17] ),
    .B(_03391_));
 sg13g2_nand2_1 _11509_ (.Y(_03411_),
    .A(\am_sdr0.cic0.comb3_in_del[17] ),
    .B(net165));
 sg13g2_a21oi_1 _11510_ (.A1(_03410_),
    .A2(_03411_),
    .Y(_00287_),
    .B1(net122));
 sg13g2_nand2_1 _11511_ (.Y(_03412_),
    .A(\am_sdr0.cic0.comb2[18] ),
    .B(_03391_));
 sg13g2_nand2_1 _11512_ (.Y(_03413_),
    .A(\am_sdr0.cic0.comb3_in_del[18] ),
    .B(_03395_));
 sg13g2_a21oi_1 _11513_ (.A1(_03412_),
    .A2(_03413_),
    .Y(_00288_),
    .B1(_03405_));
 sg13g2_buf_1 _11514_ (.A(_02728_),
    .X(_03414_));
 sg13g2_nand2_1 _11515_ (.Y(_03415_),
    .A(\am_sdr0.cic0.comb2[19] ),
    .B(_03414_));
 sg13g2_nand2_1 _11516_ (.Y(_03416_),
    .A(\am_sdr0.cic0.comb3_in_del[19] ),
    .B(net165));
 sg13g2_a21oi_1 _11517_ (.A1(_03415_),
    .A2(_03416_),
    .Y(_00289_),
    .B1(_03405_));
 sg13g2_nand2_1 _11518_ (.Y(_03417_),
    .A(_03169_),
    .B(net164));
 sg13g2_buf_1 _11519_ (.A(_02785_),
    .X(_03418_));
 sg13g2_nand2_1 _11520_ (.Y(_03419_),
    .A(\am_sdr0.cic0.comb3_in_del[1] ),
    .B(net163));
 sg13g2_a21oi_1 _11521_ (.A1(_03417_),
    .A2(_03419_),
    .Y(_00290_),
    .B1(net122));
 sg13g2_nand2_1 _11522_ (.Y(_03420_),
    .A(_03175_),
    .B(_03414_));
 sg13g2_nand2_1 _11523_ (.Y(_03421_),
    .A(\am_sdr0.cic0.comb3_in_del[2] ),
    .B(_03418_));
 sg13g2_a21oi_1 _11524_ (.A1(_03420_),
    .A2(_03421_),
    .Y(_00291_),
    .B1(net122));
 sg13g2_nand2_1 _11525_ (.Y(_03422_),
    .A(_03181_),
    .B(net164));
 sg13g2_nand2_1 _11526_ (.Y(_03423_),
    .A(\am_sdr0.cic0.comb3_in_del[3] ),
    .B(net163));
 sg13g2_a21oi_1 _11527_ (.A1(_03422_),
    .A2(_03423_),
    .Y(_00292_),
    .B1(net122));
 sg13g2_nand2_1 _11528_ (.Y(_03424_),
    .A(_03184_),
    .B(net164));
 sg13g2_nand2_1 _11529_ (.Y(_03425_),
    .A(\am_sdr0.cic0.comb3_in_del[4] ),
    .B(net163));
 sg13g2_a21oi_1 _11530_ (.A1(_03424_),
    .A2(_03425_),
    .Y(_00293_),
    .B1(net122));
 sg13g2_nand2_1 _11531_ (.Y(_03426_),
    .A(\am_sdr0.cic0.comb2[5] ),
    .B(net164));
 sg13g2_nand2_1 _11532_ (.Y(_03427_),
    .A(\am_sdr0.cic0.comb3_in_del[5] ),
    .B(net163));
 sg13g2_buf_1 _11533_ (.A(_02778_),
    .X(_03428_));
 sg13g2_buf_1 _11534_ (.A(_03428_),
    .X(_03429_));
 sg13g2_a21oi_1 _11535_ (.A1(_03426_),
    .A2(_03427_),
    .Y(_00294_),
    .B1(net121));
 sg13g2_nand2_1 _11536_ (.Y(_03430_),
    .A(_03197_),
    .B(net164));
 sg13g2_nand2_1 _11537_ (.Y(_03431_),
    .A(\am_sdr0.cic0.comb3_in_del[6] ),
    .B(net163));
 sg13g2_a21oi_1 _11538_ (.A1(_03430_),
    .A2(_03431_),
    .Y(_00295_),
    .B1(net121));
 sg13g2_nand2_1 _11539_ (.Y(_03432_),
    .A(\am_sdr0.cic0.comb2[7] ),
    .B(net164));
 sg13g2_nand2_1 _11540_ (.Y(_03433_),
    .A(\am_sdr0.cic0.comb3_in_del[7] ),
    .B(net163));
 sg13g2_a21oi_1 _11541_ (.A1(_03432_),
    .A2(_03433_),
    .Y(_00296_),
    .B1(net121));
 sg13g2_nand2_1 _11542_ (.Y(_03434_),
    .A(\am_sdr0.cic0.comb2[8] ),
    .B(net164));
 sg13g2_nand2_1 _11543_ (.Y(_03435_),
    .A(\am_sdr0.cic0.comb3_in_del[8] ),
    .B(net163));
 sg13g2_a21oi_1 _11544_ (.A1(_03434_),
    .A2(_03435_),
    .Y(_00297_),
    .B1(net121));
 sg13g2_nand2_1 _11545_ (.Y(_03436_),
    .A(_03224_),
    .B(net164));
 sg13g2_nand2_1 _11546_ (.Y(_03437_),
    .A(\am_sdr0.cic0.comb3_in_del[9] ),
    .B(net163));
 sg13g2_a21oi_1 _11547_ (.A1(_03436_),
    .A2(_03437_),
    .Y(_00298_),
    .B1(net121));
 sg13g2_xnor2_1 _11548_ (.Y(_03438_),
    .A(\am_sdr0.I_out[0] ),
    .B(\am_sdr0.cic0.integ1[0] ));
 sg13g2_nor2_1 _11549_ (.A(_03373_),
    .B(_03438_),
    .Y(_00307_));
 sg13g2_buf_1 _11550_ (.A(\am_sdr0.cic0.integ1[10] ),
    .X(_03439_));
 sg13g2_buf_1 _11551_ (.A(_03439_),
    .X(_03440_));
 sg13g2_buf_1 _11552_ (.A(\am_sdr0.I_out[7] ),
    .X(_03441_));
 sg13g2_buf_1 _11553_ (.A(_03441_),
    .X(_03442_));
 sg13g2_buf_1 _11554_ (.A(net295),
    .X(_03443_));
 sg13g2_buf_1 _11555_ (.A(\am_sdr0.cic0.integ1[7] ),
    .X(_03444_));
 sg13g2_inv_1 _11556_ (.Y(_03445_),
    .A(net362));
 sg13g2_nor2_1 _11557_ (.A(net242),
    .B(_03445_),
    .Y(_03446_));
 sg13g2_buf_2 _11558_ (.A(\am_sdr0.cic0.integ1[8] ),
    .X(_03447_));
 sg13g2_inv_1 _11559_ (.Y(_03448_),
    .A(_03447_));
 sg13g2_inv_1 _11560_ (.Y(_03449_),
    .A(\am_sdr0.cic0.integ1[9] ));
 sg13g2_buf_1 _11561_ (.A(\am_sdr0.cic0.integ1[6] ),
    .X(_03450_));
 sg13g2_buf_2 _11562_ (.A(\am_sdr0.cic0.integ1[5] ),
    .X(_03451_));
 sg13g2_inv_1 _11563_ (.Y(_03452_),
    .A(_03451_));
 sg13g2_buf_2 _11564_ (.A(\am_sdr0.cic0.integ1[4] ),
    .X(_03453_));
 sg13g2_inv_1 _11565_ (.Y(_03454_),
    .A(\am_sdr0.I_out[3] ));
 sg13g2_nor2_1 _11566_ (.A(\am_sdr0.I_out[1] ),
    .B(\am_sdr0.cic0.integ1[1] ),
    .Y(_03455_));
 sg13g2_a22oi_1 _11567_ (.Y(_03456_),
    .B1(\am_sdr0.I_out[1] ),
    .B2(\am_sdr0.cic0.integ1[1] ),
    .A2(\am_sdr0.cic0.integ1[0] ),
    .A1(\am_sdr0.I_out[0] ));
 sg13g2_nand2_1 _11568_ (.Y(_03457_),
    .A(\am_sdr0.I_out[2] ),
    .B(\am_sdr0.cic0.integ1[2] ));
 sg13g2_o21ai_1 _11569_ (.B1(_03457_),
    .Y(_03458_),
    .A1(_03455_),
    .A2(_03456_));
 sg13g2_or2_1 _11570_ (.X(_03459_),
    .B(\am_sdr0.cic0.integ1[2] ),
    .A(\am_sdr0.I_out[2] ));
 sg13g2_buf_1 _11571_ (.A(_03459_),
    .X(_03460_));
 sg13g2_buf_2 _11572_ (.A(\am_sdr0.cic0.integ1[3] ),
    .X(_03461_));
 sg13g2_a21oi_1 _11573_ (.A1(_03458_),
    .A2(_03460_),
    .Y(_03462_),
    .B1(_03461_));
 sg13g2_nand3_1 _11574_ (.B(_03458_),
    .C(_03460_),
    .A(_03461_),
    .Y(_03463_));
 sg13g2_o21ai_1 _11575_ (.B1(_03463_),
    .Y(_03464_),
    .A1(_03454_),
    .A2(_03462_));
 sg13g2_buf_1 _11576_ (.A(_03464_),
    .X(_03465_));
 sg13g2_nand2_1 _11577_ (.Y(_03466_),
    .A(_03453_),
    .B(_03465_));
 sg13g2_o21ai_1 _11578_ (.B1(\am_sdr0.I_out[4] ),
    .Y(_03467_),
    .A1(_03453_),
    .A2(_03465_));
 sg13g2_buf_1 _11579_ (.A(_03467_),
    .X(_03468_));
 sg13g2_nand3_1 _11580_ (.B(_03466_),
    .C(_03468_),
    .A(_03452_),
    .Y(_03469_));
 sg13g2_a21oi_1 _11581_ (.A1(_03466_),
    .A2(_03468_),
    .Y(_03470_),
    .B1(_03452_));
 sg13g2_a21o_1 _11582_ (.A2(_03469_),
    .A1(\am_sdr0.I_out[5] ),
    .B1(_03470_),
    .X(_03471_));
 sg13g2_buf_2 _11583_ (.A(_03471_),
    .X(_03472_));
 sg13g2_nor2_1 _11584_ (.A(net361),
    .B(_03472_),
    .Y(_03473_));
 sg13g2_a21oi_1 _11585_ (.A1(net361),
    .A2(_03472_),
    .Y(_03474_),
    .B1(\am_sdr0.I_out[6] ));
 sg13g2_nor4_2 _11586_ (.A(_03448_),
    .B(_03449_),
    .C(_03473_),
    .Y(_03475_),
    .D(_03474_));
 sg13g2_inv_2 _11587_ (.Y(_03476_),
    .A(_03441_));
 sg13g2_nor2_2 _11588_ (.A(_03476_),
    .B(net362),
    .Y(_03477_));
 sg13g2_nor2_2 _11589_ (.A(_03473_),
    .B(_03474_),
    .Y(_03478_));
 sg13g2_nor3_1 _11590_ (.A(_03447_),
    .B(\am_sdr0.cic0.integ1[9] ),
    .C(_03478_),
    .Y(_03479_));
 sg13g2_a22oi_1 _11591_ (.Y(_03480_),
    .B1(_03477_),
    .B2(_03479_),
    .A2(_03475_),
    .A1(_03446_));
 sg13g2_xor2_1 _11592_ (.B(_03480_),
    .A(net296),
    .X(_03481_));
 sg13g2_nor2_1 _11593_ (.A(net123),
    .B(_03481_),
    .Y(_00308_));
 sg13g2_a21oi_1 _11594_ (.A1(net296),
    .A2(_03475_),
    .Y(_03482_),
    .B1(_03441_));
 sg13g2_nand2_1 _11595_ (.Y(_03483_),
    .A(net361),
    .B(_03472_));
 sg13g2_o21ai_1 _11596_ (.B1(\am_sdr0.I_out[6] ),
    .Y(_03484_),
    .A1(net361),
    .A2(_03472_));
 sg13g2_nand4_1 _11597_ (.B(_03449_),
    .C(_03483_),
    .A(_03448_),
    .Y(_03485_),
    .D(_03484_));
 sg13g2_buf_1 _11598_ (.A(_03485_),
    .X(_03486_));
 sg13g2_o21ai_1 _11599_ (.B1(_03441_),
    .Y(_03487_),
    .A1(net296),
    .A2(_03486_));
 sg13g2_o21ai_1 _11600_ (.B1(_03487_),
    .Y(_03488_),
    .A1(_03445_),
    .A2(_03482_));
 sg13g2_buf_2 _11601_ (.A(_03488_),
    .X(_03489_));
 sg13g2_buf_1 _11602_ (.A(\am_sdr0.cic0.integ1[11] ),
    .X(_03490_));
 sg13g2_xor2_1 _11603_ (.B(net360),
    .A(net242),
    .X(_03491_));
 sg13g2_xnor2_1 _11604_ (.Y(_03492_),
    .A(_03489_),
    .B(_03491_));
 sg13g2_nor2_1 _11605_ (.A(net123),
    .B(_03492_),
    .Y(_00309_));
 sg13g2_or4_1 _11606_ (.A(net362),
    .B(net296),
    .C(net360),
    .D(_03486_),
    .X(_03493_));
 sg13g2_and4_1 _11607_ (.A(net362),
    .B(_03440_),
    .C(net360),
    .D(_03475_),
    .X(_03494_));
 sg13g2_buf_2 _11608_ (.A(_03494_),
    .X(_03495_));
 sg13g2_a21oi_2 _11609_ (.B1(_03495_),
    .Y(_03496_),
    .A2(_03493_),
    .A1(net295));
 sg13g2_buf_1 _11610_ (.A(\am_sdr0.cic0.integ1[12] ),
    .X(_03497_));
 sg13g2_buf_1 _11611_ (.A(_03497_),
    .X(_03498_));
 sg13g2_xnor2_1 _11612_ (.Y(_03499_),
    .A(net242),
    .B(net294));
 sg13g2_xnor2_1 _11613_ (.Y(_03500_),
    .A(_03496_),
    .B(_03499_));
 sg13g2_nor2_1 _11614_ (.A(net123),
    .B(_03500_),
    .Y(_00310_));
 sg13g2_buf_1 _11615_ (.A(\am_sdr0.cic0.integ1[13] ),
    .X(_03501_));
 sg13g2_buf_1 _11616_ (.A(_03501_),
    .X(_03502_));
 sg13g2_nor4_1 _11617_ (.A(_03476_),
    .B(net360),
    .C(net294),
    .D(_03489_),
    .Y(_03503_));
 sg13g2_nand4_1 _11618_ (.B(net360),
    .C(net294),
    .A(_03476_),
    .Y(_03504_),
    .D(_03489_));
 sg13g2_nor2b_1 _11619_ (.A(_03503_),
    .B_N(_03504_),
    .Y(_03505_));
 sg13g2_xor2_1 _11620_ (.B(_03505_),
    .A(net293),
    .X(_03506_));
 sg13g2_nor2_1 _11621_ (.A(net123),
    .B(_03506_),
    .Y(_00311_));
 sg13g2_buf_2 _11622_ (.A(\am_sdr0.cic0.integ1[14] ),
    .X(_03507_));
 sg13g2_nand2_1 _11623_ (.Y(_03508_),
    .A(net294),
    .B(net293));
 sg13g2_or2_1 _11624_ (.X(_03509_),
    .B(_03508_),
    .A(_03496_));
 sg13g2_nor2_1 _11625_ (.A(_03497_),
    .B(_03501_),
    .Y(_03510_));
 sg13g2_nand3_1 _11626_ (.B(_03496_),
    .C(_03510_),
    .A(net242),
    .Y(_03511_));
 sg13g2_o21ai_1 _11627_ (.B1(_03511_),
    .Y(_03512_),
    .A1(net242),
    .A2(_03509_));
 sg13g2_xnor2_1 _11628_ (.Y(_03513_),
    .A(_03507_),
    .B(_03512_));
 sg13g2_nor2_1 _11629_ (.A(net123),
    .B(_03513_),
    .Y(_00312_));
 sg13g2_and3_1 _11630_ (.X(_03514_),
    .A(_03497_),
    .B(_03501_),
    .C(_03507_));
 sg13g2_a21o_1 _11631_ (.A2(_03514_),
    .A1(_03489_),
    .B1(net295),
    .X(_03515_));
 sg13g2_or4_1 _11632_ (.A(_03498_),
    .B(net293),
    .C(_03507_),
    .D(_03489_),
    .X(_03516_));
 sg13g2_a22oi_1 _11633_ (.Y(_03517_),
    .B1(_03516_),
    .B2(net295),
    .A2(_03515_),
    .A1(_03490_));
 sg13g2_buf_1 _11634_ (.A(_03517_),
    .X(_03518_));
 sg13g2_buf_1 _11635_ (.A(\am_sdr0.cic0.integ1[15] ),
    .X(_03519_));
 sg13g2_xnor2_1 _11636_ (.Y(_03520_),
    .A(net242),
    .B(net359));
 sg13g2_xnor2_1 _11637_ (.Y(_03521_),
    .A(_03518_),
    .B(_03520_));
 sg13g2_nor2_1 _11638_ (.A(net123),
    .B(_03521_),
    .Y(_00313_));
 sg13g2_nor4_2 _11639_ (.A(_03444_),
    .B(_03440_),
    .C(_03490_),
    .Y(_03522_),
    .D(_03486_));
 sg13g2_nor2_1 _11640_ (.A(_03507_),
    .B(net359),
    .Y(_03523_));
 sg13g2_nand3_1 _11641_ (.B(_03510_),
    .C(_03523_),
    .A(_03522_),
    .Y(_03524_));
 sg13g2_and2_1 _11642_ (.A(_03507_),
    .B(net359),
    .X(_03525_));
 sg13g2_buf_1 _11643_ (.A(_03525_),
    .X(_03526_));
 sg13g2_and4_1 _11644_ (.A(net294),
    .B(net293),
    .C(_03495_),
    .D(_03526_),
    .X(_03527_));
 sg13g2_a21oi_2 _11645_ (.B1(_03527_),
    .Y(_03528_),
    .A2(_03524_),
    .A1(net295));
 sg13g2_buf_1 _11646_ (.A(\am_sdr0.cic0.integ1[16] ),
    .X(_03529_));
 sg13g2_xnor2_1 _11647_ (.Y(_03530_),
    .A(_03443_),
    .B(net358));
 sg13g2_xnor2_1 _11648_ (.Y(_03531_),
    .A(_03528_),
    .B(_03530_));
 sg13g2_nor2_1 _11649_ (.A(net123),
    .B(_03531_),
    .Y(_00314_));
 sg13g2_inv_1 _11650_ (.Y(_03532_),
    .A(net358));
 sg13g2_nand4_1 _11651_ (.B(_03522_),
    .C(_03510_),
    .A(_03532_),
    .Y(_03533_),
    .D(_03523_));
 sg13g2_a22oi_1 _11652_ (.Y(_03534_),
    .B1(_03533_),
    .B2(net295),
    .A2(_03527_),
    .A1(net358));
 sg13g2_buf_2 _11653_ (.A(\am_sdr0.cic0.integ1[17] ),
    .X(_03535_));
 sg13g2_nor2b_1 _11654_ (.A(_03441_),
    .B_N(_03535_),
    .Y(_03536_));
 sg13g2_buf_1 _11655_ (.A(_03536_),
    .X(_03537_));
 sg13g2_nor2_1 _11656_ (.A(_03476_),
    .B(_03535_),
    .Y(_03538_));
 sg13g2_nor2_1 _11657_ (.A(_03537_),
    .B(_03538_),
    .Y(_03539_));
 sg13g2_xnor2_1 _11658_ (.Y(_03540_),
    .A(_03534_),
    .B(_03539_));
 sg13g2_nor2_1 _11659_ (.A(net123),
    .B(_03540_),
    .Y(_00315_));
 sg13g2_buf_1 _11660_ (.A(_03195_),
    .X(_03541_));
 sg13g2_buf_1 _11661_ (.A(\am_sdr0.cic0.integ1[18] ),
    .X(_03542_));
 sg13g2_nand3_1 _11662_ (.B(_03523_),
    .C(_03538_),
    .A(_03532_),
    .Y(_03543_));
 sg13g2_a21oi_1 _11663_ (.A1(net293),
    .A2(_03495_),
    .Y(_03544_),
    .B1(net295));
 sg13g2_nand2b_1 _11664_ (.Y(_03545_),
    .B(net294),
    .A_N(_03544_));
 sg13g2_o21ai_1 _11665_ (.B1(net295),
    .Y(_03546_),
    .A1(net293),
    .A2(_03493_));
 sg13g2_nand3_1 _11666_ (.B(_03526_),
    .C(_03537_),
    .A(net358),
    .Y(_03547_));
 sg13g2_a22oi_1 _11667_ (.Y(_03548_),
    .B1(_03547_),
    .B2(_03543_),
    .A2(_03546_),
    .A1(_03545_));
 sg13g2_mux2_1 _11668_ (.A0(_03543_),
    .A1(net242),
    .S(_03548_),
    .X(_03549_));
 sg13g2_xor2_1 _11669_ (.B(_03549_),
    .A(net357),
    .X(_03550_));
 sg13g2_nor2_1 _11670_ (.A(net120),
    .B(_03550_),
    .Y(_00316_));
 sg13g2_buf_1 _11671_ (.A(\am_sdr0.cic0.integ1[19] ),
    .X(_03551_));
 sg13g2_nand4_1 _11672_ (.B(_03529_),
    .C(net357),
    .A(net359),
    .Y(_03552_),
    .D(_03537_));
 sg13g2_nor2_1 _11673_ (.A(_03519_),
    .B(net357),
    .Y(_03553_));
 sg13g2_nand3_1 _11674_ (.B(_03538_),
    .C(_03553_),
    .A(_03532_),
    .Y(_03554_));
 sg13g2_mux2_1 _11675_ (.A0(_03552_),
    .A1(_03554_),
    .S(_03518_),
    .X(_03555_));
 sg13g2_xor2_1 _11676_ (.B(_03555_),
    .A(net356),
    .X(_03556_));
 sg13g2_nor2_1 _11677_ (.A(net120),
    .B(_03556_),
    .Y(_00317_));
 sg13g2_nand2_1 _11678_ (.Y(_03557_),
    .A(\am_sdr0.I_out[0] ),
    .B(\am_sdr0.cic0.integ1[0] ));
 sg13g2_xnor2_1 _11679_ (.Y(_03558_),
    .A(\am_sdr0.I_out[1] ),
    .B(\am_sdr0.cic0.integ1[1] ));
 sg13g2_xnor2_1 _11680_ (.Y(_03559_),
    .A(_03557_),
    .B(_03558_));
 sg13g2_nor2_1 _11681_ (.A(_03541_),
    .B(_03559_),
    .Y(_00318_));
 sg13g2_buf_1 _11682_ (.A(\am_sdr0.cic0.integ1[20] ),
    .X(_03560_));
 sg13g2_nor4_2 _11683_ (.A(_03476_),
    .B(_03535_),
    .C(net357),
    .Y(_03561_),
    .D(net356));
 sg13g2_and2_1 _11684_ (.A(_03532_),
    .B(_03561_),
    .X(_03562_));
 sg13g2_buf_1 _11685_ (.A(_03562_),
    .X(_03563_));
 sg13g2_and4_1 _11686_ (.A(_03529_),
    .B(net357),
    .C(net356),
    .D(_03537_),
    .X(_03564_));
 sg13g2_buf_1 _11687_ (.A(_03564_),
    .X(_03565_));
 sg13g2_nand2_1 _11688_ (.Y(_03566_),
    .A(_03507_),
    .B(net359));
 sg13g2_nor3_1 _11689_ (.A(_03496_),
    .B(_03508_),
    .C(_03566_),
    .Y(_03567_));
 sg13g2_a22oi_1 _11690_ (.Y(_03568_),
    .B1(_03565_),
    .B2(_03567_),
    .A2(_03563_),
    .A1(_03528_));
 sg13g2_xor2_1 _11691_ (.B(_03568_),
    .A(net355),
    .X(_03569_));
 sg13g2_nor2_1 _11692_ (.A(net120),
    .B(_03569_),
    .Y(_00319_));
 sg13g2_buf_2 _11693_ (.A(\am_sdr0.cic0.integ1[21] ),
    .X(_03570_));
 sg13g2_and4_1 _11694_ (.A(_03502_),
    .B(net355),
    .C(_03526_),
    .D(_03565_),
    .X(_03571_));
 sg13g2_nand2_1 _11695_ (.Y(_03572_),
    .A(_03523_),
    .B(_03563_));
 sg13g2_nor3_1 _11696_ (.A(_03502_),
    .B(net355),
    .C(_03572_),
    .Y(_03573_));
 sg13g2_nand2b_1 _11697_ (.Y(_03574_),
    .B(_03522_),
    .A_N(net294));
 sg13g2_a22oi_1 _11698_ (.Y(_03575_),
    .B1(_03574_),
    .B2(net242),
    .A2(_03495_),
    .A1(net294));
 sg13g2_mux2_1 _11699_ (.A0(_03571_),
    .A1(_03573_),
    .S(_03575_),
    .X(_03576_));
 sg13g2_xnor2_1 _11700_ (.Y(_03577_),
    .A(_03570_),
    .B(_03576_));
 sg13g2_nor2_1 _11701_ (.A(net120),
    .B(_03577_),
    .Y(_00320_));
 sg13g2_buf_2 _11702_ (.A(\am_sdr0.cic0.integ1[22] ),
    .X(_03578_));
 sg13g2_or2_1 _11703_ (.X(_03579_),
    .B(_03570_),
    .A(net355));
 sg13g2_buf_1 _11704_ (.A(_03579_),
    .X(_03580_));
 sg13g2_or2_1 _11705_ (.X(_03581_),
    .B(_03580_),
    .A(_03572_));
 sg13g2_nand4_1 _11706_ (.B(_03570_),
    .C(_03567_),
    .A(net355),
    .Y(_03582_),
    .D(_03565_));
 sg13g2_o21ai_1 _11707_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_03548_),
    .A2(_03581_));
 sg13g2_xnor2_1 _11708_ (.Y(_03584_),
    .A(_03578_),
    .B(_03583_));
 sg13g2_nor2_1 _11709_ (.A(net120),
    .B(_03584_),
    .Y(_00321_));
 sg13g2_buf_2 _11710_ (.A(\am_sdr0.cic0.integ1[23] ),
    .X(_03585_));
 sg13g2_inv_1 _11711_ (.Y(_03586_),
    .A(_03578_));
 sg13g2_nor2_1 _11712_ (.A(_03442_),
    .B(_03586_),
    .Y(_03587_));
 sg13g2_and3_1 _11713_ (.X(_03588_),
    .A(net355),
    .B(_03570_),
    .C(_03587_));
 sg13g2_nand2_1 _11714_ (.Y(_03589_),
    .A(net356),
    .B(_03588_));
 sg13g2_a21oi_1 _11715_ (.A1(_03552_),
    .A2(_03554_),
    .Y(_03590_),
    .B1(_03589_));
 sg13g2_nor4_1 _11716_ (.A(net356),
    .B(_03578_),
    .C(_03554_),
    .D(_03580_),
    .Y(_03591_));
 sg13g2_mux2_1 _11717_ (.A0(_03590_),
    .A1(_03591_),
    .S(_03518_),
    .X(_03592_));
 sg13g2_xnor2_1 _11718_ (.Y(_03593_),
    .A(_03585_),
    .B(_03592_));
 sg13g2_nor2_1 _11719_ (.A(net120),
    .B(_03593_),
    .Y(_00322_));
 sg13g2_buf_2 _11720_ (.A(\am_sdr0.cic0.integ1[24] ),
    .X(_03594_));
 sg13g2_and2_1 _11721_ (.A(_03585_),
    .B(_03588_),
    .X(_03595_));
 sg13g2_o21ai_1 _11722_ (.B1(_03595_),
    .Y(_03596_),
    .A1(_03563_),
    .A2(_03565_));
 sg13g2_nor3_1 _11723_ (.A(_03578_),
    .B(_03585_),
    .C(_03580_),
    .Y(_03597_));
 sg13g2_nand2_1 _11724_ (.Y(_03598_),
    .A(_03563_),
    .B(_03597_));
 sg13g2_mux2_1 _11725_ (.A0(_03596_),
    .A1(_03598_),
    .S(_03528_),
    .X(_03599_));
 sg13g2_xor2_1 _11726_ (.B(_03599_),
    .A(_03594_),
    .X(_03600_));
 sg13g2_nor2_1 _11727_ (.A(net120),
    .B(_03600_),
    .Y(_00323_));
 sg13g2_nand3b_1 _11728_ (.B(_03561_),
    .C(_03597_),
    .Y(_03601_),
    .A_N(_03594_));
 sg13g2_nand4_1 _11729_ (.B(_03585_),
    .C(_03594_),
    .A(_03570_),
    .Y(_03602_),
    .D(_03587_));
 sg13g2_inv_1 _11730_ (.Y(_03603_),
    .A(_03585_));
 sg13g2_nor2_1 _11731_ (.A(_03570_),
    .B(_03594_),
    .Y(_03604_));
 sg13g2_nand4_1 _11732_ (.B(_03586_),
    .C(_03603_),
    .A(_03442_),
    .Y(_03605_),
    .D(_03604_));
 sg13g2_nand2b_1 _11733_ (.Y(_03606_),
    .B(_03561_),
    .A_N(net355));
 sg13g2_nand4_1 _11734_ (.B(net356),
    .C(net355),
    .A(net357),
    .Y(_03607_),
    .D(_03537_));
 sg13g2_a221oi_1 _11735_ (.B2(_03607_),
    .C1(_03534_),
    .B1(_03606_),
    .A1(_03602_),
    .Y(_03608_),
    .A2(_03605_));
 sg13g2_mux2_1 _11736_ (.A0(_03601_),
    .A1(_03443_),
    .S(_03608_),
    .X(_03609_));
 sg13g2_xor2_1 _11737_ (.B(_03609_),
    .A(\am_sdr0.cic0.integ1[25] ),
    .X(_03610_));
 sg13g2_nor2_1 _11738_ (.A(net120),
    .B(_03610_),
    .Y(_00324_));
 sg13g2_nor2_1 _11739_ (.A(_03455_),
    .B(_03456_),
    .Y(_03611_));
 sg13g2_xor2_1 _11740_ (.B(\am_sdr0.cic0.integ1[2] ),
    .A(\am_sdr0.I_out[2] ),
    .X(_03612_));
 sg13g2_xnor2_1 _11741_ (.Y(_03613_),
    .A(_03611_),
    .B(_03612_));
 sg13g2_nor2_1 _11742_ (.A(_03541_),
    .B(_03613_),
    .Y(_00325_));
 sg13g2_buf_1 _11743_ (.A(_03195_),
    .X(_03614_));
 sg13g2_nand2_1 _11744_ (.Y(_03615_),
    .A(_03458_),
    .B(_03460_));
 sg13g2_xnor2_1 _11745_ (.Y(_03616_),
    .A(\am_sdr0.I_out[3] ),
    .B(_03461_));
 sg13g2_xnor2_1 _11746_ (.Y(_03617_),
    .A(_03615_),
    .B(_03616_));
 sg13g2_nor2_1 _11747_ (.A(_03614_),
    .B(_03617_),
    .Y(_00326_));
 sg13g2_xor2_1 _11748_ (.B(_03453_),
    .A(\am_sdr0.I_out[4] ),
    .X(_03618_));
 sg13g2_xnor2_1 _11749_ (.Y(_03619_),
    .A(_03465_),
    .B(_03618_));
 sg13g2_nor2_1 _11750_ (.A(net119),
    .B(_03619_),
    .Y(_00327_));
 sg13g2_xnor2_1 _11751_ (.Y(_03620_),
    .A(\am_sdr0.I_out[5] ),
    .B(_03451_));
 sg13g2_and3_1 _11752_ (.X(_03621_),
    .A(_03466_),
    .B(_03468_),
    .C(_03620_));
 sg13g2_a21oi_1 _11753_ (.A1(_03466_),
    .A2(_03468_),
    .Y(_03622_),
    .B1(_03620_));
 sg13g2_nor3_1 _11754_ (.A(net177),
    .B(_03621_),
    .C(_03622_),
    .Y(_00328_));
 sg13g2_xor2_1 _11755_ (.B(_03450_),
    .A(\am_sdr0.I_out[6] ),
    .X(_03623_));
 sg13g2_xnor2_1 _11756_ (.Y(_03624_),
    .A(_03472_),
    .B(_03623_));
 sg13g2_nor2_1 _11757_ (.A(_03614_),
    .B(_03624_),
    .Y(_00329_));
 sg13g2_nor2_1 _11758_ (.A(_03446_),
    .B(_03477_),
    .Y(_03625_));
 sg13g2_xor2_1 _11759_ (.B(_03625_),
    .A(_03478_),
    .X(_03626_));
 sg13g2_nor2_1 _11760_ (.A(net119),
    .B(_03626_),
    .Y(_00330_));
 sg13g2_mux2_1 _11761_ (.A0(_03477_),
    .A1(_03446_),
    .S(_03478_),
    .X(_03627_));
 sg13g2_xnor2_1 _11762_ (.Y(_03628_),
    .A(_03447_),
    .B(_03627_));
 sg13g2_nor2_1 _11763_ (.A(net119),
    .B(_03628_),
    .Y(_00331_));
 sg13g2_a21oi_1 _11764_ (.A1(_03483_),
    .A2(_03484_),
    .Y(_03629_),
    .B1(_03448_));
 sg13g2_nor2_1 _11765_ (.A(_03447_),
    .B(_03478_),
    .Y(_03630_));
 sg13g2_a22oi_1 _11766_ (.Y(_03631_),
    .B1(_03477_),
    .B2(_03630_),
    .A2(_03629_),
    .A1(_03446_));
 sg13g2_xnor2_1 _11767_ (.Y(_03632_),
    .A(_03449_),
    .B(_03631_));
 sg13g2_nor2_1 _11768_ (.A(net119),
    .B(_03632_),
    .Y(_00332_));
 sg13g2_xnor2_1 _11769_ (.Y(_03633_),
    .A(_03461_),
    .B(\am_sdr0.cic0.integ2[0] ));
 sg13g2_nor2_1 _11770_ (.A(net119),
    .B(_03633_),
    .Y(_00333_));
 sg13g2_buf_1 _11771_ (.A(\am_sdr0.cic0.integ2[6] ),
    .X(_03634_));
 sg13g2_buf_2 _11772_ (.A(\am_sdr0.cic0.integ2[5] ),
    .X(_03635_));
 sg13g2_and2_1 _11773_ (.A(_03447_),
    .B(_03635_),
    .X(_03636_));
 sg13g2_buf_2 _11774_ (.A(_03636_),
    .X(_03637_));
 sg13g2_buf_2 _11775_ (.A(\am_sdr0.cic0.integ2[3] ),
    .X(_03638_));
 sg13g2_buf_1 _11776_ (.A(\am_sdr0.cic0.integ2[2] ),
    .X(_03639_));
 sg13g2_or2_1 _11777_ (.X(_03640_),
    .B(_03639_),
    .A(_03451_));
 sg13g2_o21ai_1 _11778_ (.B1(_03640_),
    .Y(_03641_),
    .A1(net361),
    .A2(_03638_));
 sg13g2_or2_1 _11779_ (.X(_03642_),
    .B(\am_sdr0.cic0.integ2[1] ),
    .A(_03453_));
 sg13g2_and2_1 _11780_ (.A(_03461_),
    .B(\am_sdr0.cic0.integ2[0] ),
    .X(_03643_));
 sg13g2_buf_1 _11781_ (.A(_03643_),
    .X(_03644_));
 sg13g2_and2_1 _11782_ (.A(_03453_),
    .B(\am_sdr0.cic0.integ2[1] ),
    .X(_03645_));
 sg13g2_a221oi_1 _11783_ (.B2(_03644_),
    .C1(_03645_),
    .B1(_03642_),
    .A1(_03451_),
    .Y(_03646_),
    .A2(_03639_));
 sg13g2_buf_2 _11784_ (.A(\am_sdr0.cic0.integ2[4] ),
    .X(_03647_));
 sg13g2_a22oi_1 _11785_ (.Y(_03648_),
    .B1(_03647_),
    .B2(net362),
    .A2(_03638_),
    .A1(net361));
 sg13g2_o21ai_1 _11786_ (.B1(_03648_),
    .Y(_03649_),
    .A1(_03641_),
    .A2(_03646_));
 sg13g2_buf_2 _11787_ (.A(_03649_),
    .X(_03650_));
 sg13g2_inv_1 _11788_ (.Y(_03651_),
    .A(net354));
 sg13g2_nor2_1 _11789_ (.A(_03447_),
    .B(_03635_),
    .Y(_03652_));
 sg13g2_nor2_1 _11790_ (.A(net362),
    .B(_03647_),
    .Y(_03653_));
 sg13g2_nor3_2 _11791_ (.A(_03651_),
    .B(_03652_),
    .C(_03653_),
    .Y(_03654_));
 sg13g2_buf_1 _11792_ (.A(\am_sdr0.cic0.integ2[7] ),
    .X(_03655_));
 sg13g2_buf_2 _11793_ (.A(\am_sdr0.cic0.integ2[8] ),
    .X(_03656_));
 sg13g2_or2_1 _11794_ (.X(_03657_),
    .B(_03656_),
    .A(net353));
 sg13g2_a221oi_1 _11795_ (.B2(_03654_),
    .C1(_03657_),
    .B1(_03650_),
    .A1(net354),
    .Y(_03658_),
    .A2(_03637_));
 sg13g2_or2_1 _11796_ (.X(_03659_),
    .B(_03656_),
    .A(_03439_));
 sg13g2_a221oi_1 _11797_ (.B2(_03654_),
    .C1(_03659_),
    .B1(_03650_),
    .A1(net354),
    .Y(_03660_),
    .A2(_03637_));
 sg13g2_a21o_1 _11798_ (.A2(_03635_),
    .A1(_03447_),
    .B1(net354),
    .X(_03661_));
 sg13g2_or2_1 _11799_ (.X(_03662_),
    .B(_03647_),
    .A(net362));
 sg13g2_or2_1 _11800_ (.X(_03663_),
    .B(_03635_),
    .A(_03447_));
 sg13g2_o21ai_1 _11801_ (.B1(_03663_),
    .Y(_03664_),
    .A1(_03662_),
    .A2(_03637_));
 sg13g2_a21oi_1 _11802_ (.A1(_03651_),
    .A2(_03664_),
    .Y(_03665_),
    .B1(_03449_));
 sg13g2_o21ai_1 _11803_ (.B1(_03665_),
    .Y(_03666_),
    .A1(_03650_),
    .A2(_03661_));
 sg13g2_o21ai_1 _11804_ (.B1(_03666_),
    .Y(_03667_),
    .A1(_03658_),
    .A2(_03660_));
 sg13g2_or2_1 _11805_ (.X(_03668_),
    .B(net353),
    .A(net360));
 sg13g2_a221oi_1 _11806_ (.B2(_03654_),
    .C1(_03668_),
    .B1(_03650_),
    .A1(net354),
    .Y(_03669_),
    .A2(_03637_));
 sg13g2_or2_1 _11807_ (.X(_03670_),
    .B(\am_sdr0.cic0.integ1[11] ),
    .A(_03439_));
 sg13g2_a221oi_1 _11808_ (.B2(_03654_),
    .C1(_03670_),
    .B1(_03650_),
    .A1(_03634_),
    .Y(_03671_),
    .A2(_03637_));
 sg13g2_o21ai_1 _11809_ (.B1(_03666_),
    .Y(_03672_),
    .A1(_03669_),
    .A2(_03671_));
 sg13g2_nor2_1 _11810_ (.A(net360),
    .B(_03656_),
    .Y(_03673_));
 sg13g2_nor3_1 _11811_ (.A(net296),
    .B(net353),
    .C(_03656_),
    .Y(_03674_));
 sg13g2_nor2_1 _11812_ (.A(net353),
    .B(_03670_),
    .Y(_03675_));
 sg13g2_nor3_1 _11813_ (.A(_03673_),
    .B(_03674_),
    .C(_03675_),
    .Y(_03676_));
 sg13g2_nand3_1 _11814_ (.B(_03672_),
    .C(_03676_),
    .A(_03667_),
    .Y(_03677_));
 sg13g2_buf_1 _11815_ (.A(_03677_),
    .X(_03678_));
 sg13g2_buf_2 _11816_ (.A(\am_sdr0.cic0.integ2[9] ),
    .X(_03679_));
 sg13g2_nand2_1 _11817_ (.Y(_03680_),
    .A(_03497_),
    .B(_03679_));
 sg13g2_nor2_1 _11818_ (.A(_03497_),
    .B(_03679_),
    .Y(_03681_));
 sg13g2_a21o_1 _11819_ (.A2(_03680_),
    .A1(_03678_),
    .B1(_03681_),
    .X(_03682_));
 sg13g2_buf_1 _11820_ (.A(\am_sdr0.cic0.integ2[10] ),
    .X(_03683_));
 sg13g2_xnor2_1 _11821_ (.Y(_03684_),
    .A(net293),
    .B(net352));
 sg13g2_xnor2_1 _11822_ (.Y(_03685_),
    .A(_03682_),
    .B(_03684_));
 sg13g2_nor2_1 _11823_ (.A(net119),
    .B(_03685_),
    .Y(_00334_));
 sg13g2_buf_1 _11824_ (.A(\am_sdr0.cic0.integ2[11] ),
    .X(_03686_));
 sg13g2_nand2_1 _11825_ (.Y(_03687_),
    .A(_03507_),
    .B(_03686_));
 sg13g2_or2_1 _11826_ (.X(_03688_),
    .B(_03686_),
    .A(_03507_));
 sg13g2_buf_1 _11827_ (.A(_03688_),
    .X(_03689_));
 sg13g2_nand2_1 _11828_ (.Y(_03690_),
    .A(_03687_),
    .B(_03689_));
 sg13g2_nor2_1 _11829_ (.A(_03501_),
    .B(net352),
    .Y(_03691_));
 sg13g2_nand2_1 _11830_ (.Y(_03692_),
    .A(net293),
    .B(net352));
 sg13g2_o21ai_1 _11831_ (.B1(_03692_),
    .Y(_03693_),
    .A1(_03682_),
    .A2(_03691_));
 sg13g2_xor2_1 _11832_ (.B(_03693_),
    .A(_03690_),
    .X(_03694_));
 sg13g2_nor2_1 _11833_ (.A(net119),
    .B(_03694_),
    .Y(_00335_));
 sg13g2_nand2_1 _11834_ (.Y(_03695_),
    .A(_03680_),
    .B(_03687_));
 sg13g2_nor2_1 _11835_ (.A(\am_sdr0.cic0.integ2[10] ),
    .B(_03695_),
    .Y(_03696_));
 sg13g2_nor2_1 _11836_ (.A(_03501_),
    .B(_03695_),
    .Y(_03697_));
 sg13g2_o21ai_1 _11837_ (.B1(_03678_),
    .Y(_03698_),
    .A1(_03696_),
    .A2(_03697_));
 sg13g2_nand2_1 _11838_ (.Y(_03699_),
    .A(_03681_),
    .B(_03687_));
 sg13g2_a21oi_1 _11839_ (.A1(_03501_),
    .A2(net352),
    .Y(_03700_),
    .B1(_03699_));
 sg13g2_a21oi_1 _11840_ (.A1(_03687_),
    .A2(_03691_),
    .Y(_03701_),
    .B1(_03700_));
 sg13g2_nand3_1 _11841_ (.B(_03698_),
    .C(_03701_),
    .A(_03689_),
    .Y(_03702_));
 sg13g2_buf_1 _11842_ (.A(\am_sdr0.cic0.integ2[12] ),
    .X(_03703_));
 sg13g2_xnor2_1 _11843_ (.Y(_03704_),
    .A(net359),
    .B(net351));
 sg13g2_xnor2_1 _11844_ (.Y(_03705_),
    .A(_03702_),
    .B(_03704_));
 sg13g2_nor2_1 _11845_ (.A(net119),
    .B(_03705_),
    .Y(_00336_));
 sg13g2_buf_1 _11846_ (.A(_03195_),
    .X(_03706_));
 sg13g2_nand4_1 _11847_ (.B(_03689_),
    .C(_03698_),
    .A(net351),
    .Y(_03707_),
    .D(_03701_));
 sg13g2_nand4_1 _11848_ (.B(_03689_),
    .C(_03698_),
    .A(net359),
    .Y(_03708_),
    .D(_03701_));
 sg13g2_buf_1 _11849_ (.A(_03708_),
    .X(_03709_));
 sg13g2_nand2_1 _11850_ (.Y(_03710_),
    .A(net359),
    .B(net351));
 sg13g2_and3_1 _11851_ (.X(_03711_),
    .A(_03707_),
    .B(_03709_),
    .C(_03710_));
 sg13g2_buf_1 _11852_ (.A(\am_sdr0.cic0.integ2[13] ),
    .X(_03712_));
 sg13g2_xnor2_1 _11853_ (.Y(_03713_),
    .A(net358),
    .B(net350));
 sg13g2_xnor2_1 _11854_ (.Y(_03714_),
    .A(_03711_),
    .B(_03713_));
 sg13g2_nor2_1 _11855_ (.A(net118),
    .B(_03714_),
    .Y(_00337_));
 sg13g2_buf_2 _11856_ (.A(\am_sdr0.cic0.integ2[14] ),
    .X(_03715_));
 sg13g2_xor2_1 _11857_ (.B(_03715_),
    .A(_03535_),
    .X(_03716_));
 sg13g2_nor2_1 _11858_ (.A(net358),
    .B(net350),
    .Y(_03717_));
 sg13g2_nand2_1 _11859_ (.Y(_03718_),
    .A(net358),
    .B(net350));
 sg13g2_o21ai_1 _11860_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_03711_),
    .A2(_03717_));
 sg13g2_xnor2_1 _11861_ (.Y(_03720_),
    .A(_03716_),
    .B(_03719_));
 sg13g2_nor2_1 _11862_ (.A(net118),
    .B(_03720_),
    .Y(_00338_));
 sg13g2_a21oi_1 _11863_ (.A1(_03535_),
    .A2(_03715_),
    .Y(_03721_),
    .B1(net350));
 sg13g2_nand4_1 _11864_ (.B(_03709_),
    .C(_03710_),
    .A(_03707_),
    .Y(_03722_),
    .D(_03721_));
 sg13g2_a21oi_1 _11865_ (.A1(_03535_),
    .A2(_03715_),
    .Y(_03723_),
    .B1(net358));
 sg13g2_nand4_1 _11866_ (.B(_03709_),
    .C(_03710_),
    .A(_03707_),
    .Y(_03724_),
    .D(_03723_));
 sg13g2_nand2_1 _11867_ (.Y(_03725_),
    .A(_03535_),
    .B(_03715_));
 sg13g2_nor2_1 _11868_ (.A(_03535_),
    .B(_03715_),
    .Y(_03726_));
 sg13g2_a21oi_1 _11869_ (.A1(_03725_),
    .A2(_03717_),
    .Y(_03727_),
    .B1(_03726_));
 sg13g2_nand3_1 _11870_ (.B(_03724_),
    .C(_03727_),
    .A(_03722_),
    .Y(_03728_));
 sg13g2_buf_2 _11871_ (.A(\am_sdr0.cic0.integ2[15] ),
    .X(_03729_));
 sg13g2_xnor2_1 _11872_ (.Y(_03730_),
    .A(net357),
    .B(_03729_));
 sg13g2_xnor2_1 _11873_ (.Y(_03731_),
    .A(_03728_),
    .B(_03730_));
 sg13g2_nor2_1 _11874_ (.A(net118),
    .B(_03731_),
    .Y(_00339_));
 sg13g2_buf_2 _11875_ (.A(\am_sdr0.cic0.integ2[16] ),
    .X(_03732_));
 sg13g2_xor2_1 _11876_ (.B(_03732_),
    .A(net356),
    .X(_03733_));
 sg13g2_nor2_1 _11877_ (.A(net357),
    .B(_03729_),
    .Y(_03734_));
 sg13g2_nand2_1 _11878_ (.Y(_03735_),
    .A(_03542_),
    .B(_03729_));
 sg13g2_o21ai_1 _11879_ (.B1(_03735_),
    .Y(_03736_),
    .A1(_03728_),
    .A2(_03734_));
 sg13g2_xnor2_1 _11880_ (.Y(_03737_),
    .A(_03733_),
    .B(_03736_));
 sg13g2_nor2_1 _11881_ (.A(net118),
    .B(_03737_),
    .Y(_00340_));
 sg13g2_nor2_1 _11882_ (.A(net356),
    .B(_03732_),
    .Y(_03738_));
 sg13g2_nand2_1 _11883_ (.Y(_03739_),
    .A(_03551_),
    .B(_03732_));
 sg13g2_nand2b_1 _11884_ (.Y(_03740_),
    .B(_03739_),
    .A_N(_03736_));
 sg13g2_nand2b_1 _11885_ (.Y(_03741_),
    .B(_03740_),
    .A_N(_03738_));
 sg13g2_buf_2 _11886_ (.A(\am_sdr0.cic0.integ2[17] ),
    .X(_03742_));
 sg13g2_xnor2_1 _11887_ (.Y(_03743_),
    .A(_03560_),
    .B(_03742_));
 sg13g2_xnor2_1 _11888_ (.Y(_03744_),
    .A(_03741_),
    .B(_03743_));
 sg13g2_nor2_1 _11889_ (.A(net118),
    .B(_03744_),
    .Y(_00341_));
 sg13g2_buf_1 _11890_ (.A(\am_sdr0.cic0.integ2[18] ),
    .X(_03745_));
 sg13g2_nand2_1 _11891_ (.Y(_03746_),
    .A(_03570_),
    .B(_03745_));
 sg13g2_or2_1 _11892_ (.X(_03747_),
    .B(_03745_),
    .A(_03570_));
 sg13g2_nand2_1 _11893_ (.Y(_03748_),
    .A(_03746_),
    .B(_03747_));
 sg13g2_nor2_1 _11894_ (.A(\am_sdr0.cic0.integ1[20] ),
    .B(_03742_),
    .Y(_03749_));
 sg13g2_nand2_1 _11895_ (.Y(_03750_),
    .A(_03560_),
    .B(_03742_));
 sg13g2_o21ai_1 _11896_ (.B1(_03750_),
    .Y(_03751_),
    .A1(_03741_),
    .A2(_03749_));
 sg13g2_xnor2_1 _11897_ (.Y(_03752_),
    .A(_03748_),
    .B(_03751_));
 sg13g2_and2_1 _11898_ (.A(net246),
    .B(_03752_),
    .X(_00342_));
 sg13g2_nand3_1 _11899_ (.B(_03746_),
    .C(_03750_),
    .A(_03739_),
    .Y(_03753_));
 sg13g2_o21ai_1 _11900_ (.B1(_03750_),
    .Y(_03754_),
    .A1(_03738_),
    .A2(_03749_));
 sg13g2_nand2_1 _11901_ (.Y(_03755_),
    .A(_03747_),
    .B(_03754_));
 sg13g2_nand2_1 _11902_ (.Y(_03756_),
    .A(_03746_),
    .B(_03755_));
 sg13g2_o21ai_1 _11903_ (.B1(_03756_),
    .Y(_03757_),
    .A1(_03736_),
    .A2(_03753_));
 sg13g2_buf_1 _11904_ (.A(_03757_),
    .X(_03758_));
 sg13g2_buf_1 _11905_ (.A(\am_sdr0.cic0.integ2[19] ),
    .X(_03759_));
 sg13g2_xnor2_1 _11906_ (.Y(_03760_),
    .A(_03578_),
    .B(net349));
 sg13g2_xnor2_1 _11907_ (.Y(_03761_),
    .A(_03758_),
    .B(_03760_));
 sg13g2_nor2_1 _11908_ (.A(net118),
    .B(_03761_),
    .Y(_00343_));
 sg13g2_xor2_1 _11909_ (.B(\am_sdr0.cic0.integ2[1] ),
    .A(_03453_),
    .X(_03762_));
 sg13g2_xnor2_1 _11910_ (.Y(_03763_),
    .A(_03644_),
    .B(_03762_));
 sg13g2_nor2_1 _11911_ (.A(net118),
    .B(_03763_),
    .Y(_00344_));
 sg13g2_inv_1 _11912_ (.Y(_03764_),
    .A(net349));
 sg13g2_o21ai_1 _11913_ (.B1(_03586_),
    .Y(_03765_),
    .A1(_03764_),
    .A2(_03758_));
 sg13g2_nand2_1 _11914_ (.Y(_03766_),
    .A(_03764_),
    .B(_03758_));
 sg13g2_nand2_1 _11915_ (.Y(_03767_),
    .A(_03765_),
    .B(_03766_));
 sg13g2_buf_1 _11916_ (.A(\am_sdr0.cic0.integ2[20] ),
    .X(_03768_));
 sg13g2_xnor2_1 _11917_ (.Y(_03769_),
    .A(_03585_),
    .B(net348));
 sg13g2_xnor2_1 _11918_ (.Y(_03770_),
    .A(_03767_),
    .B(_03769_));
 sg13g2_nor2_1 _11919_ (.A(_03706_),
    .B(_03770_),
    .Y(_00345_));
 sg13g2_inv_1 _11920_ (.Y(_03771_),
    .A(net348));
 sg13g2_a221oi_1 _11921_ (.B2(_03603_),
    .C1(_03758_),
    .B1(_03771_),
    .A1(_03586_),
    .Y(_03772_),
    .A2(_03764_));
 sg13g2_nand2_1 _11922_ (.Y(_03773_),
    .A(_03585_),
    .B(net348));
 sg13g2_nand3_1 _11923_ (.B(net349),
    .C(net348),
    .A(_03578_),
    .Y(_03774_));
 sg13g2_nand3_1 _11924_ (.B(_03585_),
    .C(net349),
    .A(_03578_),
    .Y(_03775_));
 sg13g2_nand3_1 _11925_ (.B(_03774_),
    .C(_03775_),
    .A(_03773_),
    .Y(_03776_));
 sg13g2_nor2_1 _11926_ (.A(_03772_),
    .B(_03776_),
    .Y(_03777_));
 sg13g2_buf_2 _11927_ (.A(\am_sdr0.cic0.integ2[21] ),
    .X(_03778_));
 sg13g2_xnor2_1 _11928_ (.Y(_03779_),
    .A(_03594_),
    .B(_03778_));
 sg13g2_xnor2_1 _11929_ (.Y(_03780_),
    .A(_03777_),
    .B(_03779_));
 sg13g2_nor2_1 _11930_ (.A(_03706_),
    .B(_03780_),
    .Y(_00346_));
 sg13g2_nand2_1 _11931_ (.Y(_03781_),
    .A(_03594_),
    .B(_03778_));
 sg13g2_xor2_1 _11932_ (.B(\am_sdr0.cic0.integ2[22] ),
    .A(\am_sdr0.cic0.integ1[25] ),
    .X(_03782_));
 sg13g2_nand4_1 _11933_ (.B(_03777_),
    .C(_03781_),
    .A(net301),
    .Y(_03783_),
    .D(_03782_));
 sg13g2_nor2_1 _11934_ (.A(_03594_),
    .B(_03778_),
    .Y(_03784_));
 sg13g2_or4_1 _11935_ (.A(net259),
    .B(_03777_),
    .C(_03784_),
    .D(_03782_),
    .X(_03785_));
 sg13g2_nand3_1 _11936_ (.B(_03784_),
    .C(_03782_),
    .A(net301),
    .Y(_03786_));
 sg13g2_or3_1 _11937_ (.A(net259),
    .B(_03781_),
    .C(_03782_),
    .X(_03787_));
 sg13g2_nand4_1 _11938_ (.B(_03785_),
    .C(_03786_),
    .A(_03783_),
    .Y(_00347_),
    .D(_03787_));
 sg13g2_a21o_1 _11939_ (.A2(_03644_),
    .A1(_03642_),
    .B1(_03645_),
    .X(_03788_));
 sg13g2_buf_1 _11940_ (.A(_03788_),
    .X(_03789_));
 sg13g2_xor2_1 _11941_ (.B(_03639_),
    .A(_03451_),
    .X(_03790_));
 sg13g2_xnor2_1 _11942_ (.Y(_03791_),
    .A(_03789_),
    .B(_03790_));
 sg13g2_nor2_1 _11943_ (.A(net118),
    .B(_03791_),
    .Y(_00348_));
 sg13g2_buf_1 _11944_ (.A(_03195_),
    .X(_03792_));
 sg13g2_a21oi_1 _11945_ (.A1(_03639_),
    .A2(_03789_),
    .Y(_03793_),
    .B1(_03451_));
 sg13g2_nor2_1 _11946_ (.A(_03639_),
    .B(_03789_),
    .Y(_03794_));
 sg13g2_nor2_1 _11947_ (.A(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sg13g2_xor2_1 _11948_ (.B(_03638_),
    .A(net361),
    .X(_03796_));
 sg13g2_xnor2_1 _11949_ (.Y(_03797_),
    .A(_03795_),
    .B(_03796_));
 sg13g2_nor2_1 _11950_ (.A(net117),
    .B(_03797_),
    .Y(_00349_));
 sg13g2_a21o_1 _11951_ (.A2(_03795_),
    .A1(_03638_),
    .B1(net361),
    .X(_03798_));
 sg13g2_o21ai_1 _11952_ (.B1(_03798_),
    .Y(_03799_),
    .A1(_03638_),
    .A2(_03795_));
 sg13g2_xnor2_1 _11953_ (.Y(_03800_),
    .A(net362),
    .B(_03647_));
 sg13g2_xnor2_1 _11954_ (.Y(_03801_),
    .A(_03799_),
    .B(_03800_));
 sg13g2_nor2_1 _11955_ (.A(net117),
    .B(_03801_),
    .Y(_00350_));
 sg13g2_and2_1 _11956_ (.A(_03662_),
    .B(_03650_),
    .X(_03802_));
 sg13g2_nor2_1 _11957_ (.A(_03652_),
    .B(_03637_),
    .Y(_03803_));
 sg13g2_xnor2_1 _11958_ (.Y(_03804_),
    .A(_03802_),
    .B(_03803_));
 sg13g2_nor2_1 _11959_ (.A(net117),
    .B(_03804_),
    .Y(_00351_));
 sg13g2_nor2_1 _11960_ (.A(_03652_),
    .B(_03653_),
    .Y(_03805_));
 sg13g2_a21oi_1 _11961_ (.A1(_03650_),
    .A2(_03805_),
    .Y(_03806_),
    .B1(_03637_));
 sg13g2_xnor2_1 _11962_ (.Y(_03807_),
    .A(\am_sdr0.cic0.integ1[9] ),
    .B(net354));
 sg13g2_xnor2_1 _11963_ (.Y(_03808_),
    .A(_03806_),
    .B(_03807_));
 sg13g2_nor2_1 _11964_ (.A(net117),
    .B(_03808_),
    .Y(_00352_));
 sg13g2_a22oi_1 _11965_ (.Y(_03809_),
    .B1(_03650_),
    .B2(_03654_),
    .A2(_03637_),
    .A1(net354));
 sg13g2_nand2_1 _11966_ (.Y(_03810_),
    .A(_03666_),
    .B(_03809_));
 sg13g2_xor2_1 _11967_ (.B(net353),
    .A(net296),
    .X(_03811_));
 sg13g2_xnor2_1 _11968_ (.Y(_03812_),
    .A(_03810_),
    .B(_03811_));
 sg13g2_nor2_1 _11969_ (.A(net117),
    .B(_03812_),
    .Y(_00353_));
 sg13g2_o21ai_1 _11970_ (.B1(_03810_),
    .Y(_03813_),
    .A1(net296),
    .A2(net353));
 sg13g2_inv_1 _11971_ (.Y(_03814_),
    .A(_03813_));
 sg13g2_a21oi_1 _11972_ (.A1(net296),
    .A2(net353),
    .Y(_03815_),
    .B1(_03814_));
 sg13g2_xnor2_1 _11973_ (.Y(_03816_),
    .A(net360),
    .B(_03656_));
 sg13g2_xnor2_1 _11974_ (.Y(_03817_),
    .A(_03815_),
    .B(_03816_));
 sg13g2_nor2_1 _11975_ (.A(net117),
    .B(_03817_),
    .Y(_00354_));
 sg13g2_xnor2_1 _11976_ (.Y(_03818_),
    .A(_03498_),
    .B(_03679_));
 sg13g2_xnor2_1 _11977_ (.Y(_03819_),
    .A(_03678_),
    .B(_03818_));
 sg13g2_nor2_1 _11978_ (.A(net117),
    .B(_03819_),
    .Y(_00355_));
 sg13g2_xnor2_1 _11979_ (.Y(_03820_),
    .A(_03638_),
    .B(_02247_));
 sg13g2_nor2_1 _11980_ (.A(_03792_),
    .B(_03820_),
    .Y(_00356_));
 sg13g2_xor2_1 _11981_ (.B(_02258_),
    .A(net350),
    .X(_03821_));
 sg13g2_inv_1 _11982_ (.Y(_03822_),
    .A(\am_sdr0.cic0.integ3[5] ));
 sg13g2_and2_1 _11983_ (.A(_03635_),
    .B(_02281_),
    .X(_03823_));
 sg13g2_buf_1 _11984_ (.A(_03823_),
    .X(_03824_));
 sg13g2_nor2_1 _11985_ (.A(_03635_),
    .B(_02281_),
    .Y(_03825_));
 sg13g2_nor2_1 _11986_ (.A(_03647_),
    .B(_02279_),
    .Y(_03826_));
 sg13g2_a22oi_1 _11987_ (.Y(_03827_),
    .B1(_03647_),
    .B2(_02279_),
    .A2(_02247_),
    .A1(_03638_));
 sg13g2_nor3_1 _11988_ (.A(_03825_),
    .B(_03826_),
    .C(_03827_),
    .Y(_03828_));
 sg13g2_nor3_1 _11989_ (.A(_02284_),
    .B(_03824_),
    .C(_03828_),
    .Y(_03829_));
 sg13g2_o21ai_1 _11990_ (.B1(_02284_),
    .Y(_03830_),
    .A1(_03824_),
    .A2(_03828_));
 sg13g2_o21ai_1 _11991_ (.B1(_03830_),
    .Y(_03831_),
    .A1(_03651_),
    .A2(_03829_));
 sg13g2_buf_1 _11992_ (.A(_03831_),
    .X(_03832_));
 sg13g2_nand2_1 _11993_ (.Y(_03833_),
    .A(_02287_),
    .B(_03832_));
 sg13g2_o21ai_1 _11994_ (.B1(net353),
    .Y(_03834_),
    .A1(_02287_),
    .A2(_03832_));
 sg13g2_buf_1 _11995_ (.A(_03834_),
    .X(_03835_));
 sg13g2_nand3_1 _11996_ (.B(_03833_),
    .C(_03835_),
    .A(_03822_),
    .Y(_03836_));
 sg13g2_a21oi_1 _11997_ (.A1(_03833_),
    .A2(_03835_),
    .Y(_03837_),
    .B1(_03822_));
 sg13g2_a21o_1 _11998_ (.A2(_03836_),
    .A1(_03656_),
    .B1(_03837_),
    .X(_03838_));
 sg13g2_buf_2 _11999_ (.A(_03838_),
    .X(_03839_));
 sg13g2_a21oi_1 _12000_ (.A1(_02290_),
    .A2(_03839_),
    .Y(_03840_),
    .B1(_02292_));
 sg13g2_a21oi_1 _12001_ (.A1(_02290_),
    .A2(_03839_),
    .Y(_03841_),
    .B1(net352));
 sg13g2_or2_1 _12002_ (.X(_03842_),
    .B(_03839_),
    .A(_02290_));
 sg13g2_nand2_1 _12003_ (.Y(_03843_),
    .A(_03679_),
    .B(_03842_));
 sg13g2_o21ai_1 _12004_ (.B1(_03843_),
    .Y(_03844_),
    .A1(_03840_),
    .A2(_03841_));
 sg13g2_buf_1 _12005_ (.A(_03844_),
    .X(_03845_));
 sg13g2_nor2_1 _12006_ (.A(net352),
    .B(_02292_),
    .Y(_03846_));
 sg13g2_nor2b_1 _12007_ (.A(_03846_),
    .B_N(_02294_),
    .Y(_03847_));
 sg13g2_inv_1 _12008_ (.Y(_03848_),
    .A(_03686_));
 sg13g2_a21o_1 _12009_ (.A2(_03839_),
    .A1(_02290_),
    .B1(_03679_),
    .X(_03849_));
 sg13g2_a221oi_1 _12010_ (.B2(_03849_),
    .C1(_02294_),
    .B1(_03842_),
    .A1(net352),
    .Y(_03850_),
    .A2(_02292_));
 sg13g2_nor3_1 _12011_ (.A(net352),
    .B(_02292_),
    .C(_02294_),
    .Y(_03851_));
 sg13g2_nor3_2 _12012_ (.A(_03848_),
    .B(_03850_),
    .C(_03851_),
    .Y(_03852_));
 sg13g2_a21o_1 _12013_ (.A2(_03847_),
    .A1(_03845_),
    .B1(_03852_),
    .X(_03853_));
 sg13g2_and2_1 _12014_ (.A(net351),
    .B(_02296_),
    .X(_03854_));
 sg13g2_or2_1 _12015_ (.X(_03855_),
    .B(_02296_),
    .A(net351));
 sg13g2_buf_1 _12016_ (.A(_03855_),
    .X(_03856_));
 sg13g2_o21ai_1 _12017_ (.B1(_03856_),
    .Y(_03857_),
    .A1(_03853_),
    .A2(_03854_));
 sg13g2_xor2_1 _12018_ (.B(_03857_),
    .A(_03821_),
    .X(_03858_));
 sg13g2_nor2_1 _12019_ (.A(_03792_),
    .B(_03858_),
    .Y(_00357_));
 sg13g2_or2_1 _12020_ (.X(_03859_),
    .B(_02258_),
    .A(_02296_));
 sg13g2_or2_1 _12021_ (.X(_03860_),
    .B(_02258_),
    .A(net351));
 sg13g2_a221oi_1 _12022_ (.B2(_03860_),
    .C1(_03852_),
    .B1(_03859_),
    .A1(_03845_),
    .Y(_03861_),
    .A2(_03847_));
 sg13g2_or2_1 _12023_ (.X(_03862_),
    .B(net350),
    .A(_02296_));
 sg13g2_or2_1 _12024_ (.X(_03863_),
    .B(net350),
    .A(net351));
 sg13g2_a221oi_1 _12025_ (.B2(_03863_),
    .C1(_03852_),
    .B1(_03862_),
    .A1(_03845_),
    .Y(_03864_),
    .A2(_03847_));
 sg13g2_nor2_1 _12026_ (.A(net350),
    .B(_02258_),
    .Y(_03865_));
 sg13g2_a21oi_1 _12027_ (.A1(_03712_),
    .A2(_02258_),
    .Y(_03866_),
    .B1(_03856_));
 sg13g2_nor2_1 _12028_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sg13g2_inv_1 _12029_ (.Y(_03868_),
    .A(_03867_));
 sg13g2_nor3_1 _12030_ (.A(_03861_),
    .B(_03864_),
    .C(_03868_),
    .Y(_03869_));
 sg13g2_xnor2_1 _12031_ (.Y(_03870_),
    .A(_03715_),
    .B(_02260_));
 sg13g2_xor2_1 _12032_ (.B(_03870_),
    .A(_03869_),
    .X(_03871_));
 sg13g2_nor2_1 _12033_ (.A(net117),
    .B(_03871_),
    .Y(_00358_));
 sg13g2_buf_1 _12034_ (.A(_03195_),
    .X(_03872_));
 sg13g2_xnor2_1 _12035_ (.Y(_03873_),
    .A(_03729_),
    .B(_02262_));
 sg13g2_or2_1 _12036_ (.X(_03874_),
    .B(_02260_),
    .A(_03715_));
 sg13g2_and2_1 _12037_ (.A(_03715_),
    .B(_02260_),
    .X(_03875_));
 sg13g2_buf_1 _12038_ (.A(_03875_),
    .X(_03876_));
 sg13g2_a21o_1 _12039_ (.A2(_03874_),
    .A1(_03869_),
    .B1(_03876_),
    .X(_03877_));
 sg13g2_xor2_1 _12040_ (.B(_03877_),
    .A(_03873_),
    .X(_03878_));
 sg13g2_nor2_1 _12041_ (.A(_03872_),
    .B(_03878_),
    .Y(_00359_));
 sg13g2_xor2_1 _12042_ (.B(_02265_),
    .A(_03732_),
    .X(_03879_));
 sg13g2_or2_1 _12043_ (.X(_03880_),
    .B(_02262_),
    .A(_03729_));
 sg13g2_buf_1 _12044_ (.A(_03880_),
    .X(_03881_));
 sg13g2_and2_1 _12045_ (.A(_03729_),
    .B(_02262_),
    .X(_03882_));
 sg13g2_buf_1 _12046_ (.A(_03882_),
    .X(_03883_));
 sg13g2_a21oi_1 _12047_ (.A1(_03877_),
    .A2(_03881_),
    .Y(_03884_),
    .B1(_03883_));
 sg13g2_xor2_1 _12048_ (.B(_03884_),
    .A(_03879_),
    .X(_03885_));
 sg13g2_nor2_1 _12049_ (.A(_03872_),
    .B(_03885_),
    .Y(_00360_));
 sg13g2_and2_1 _12050_ (.A(_03712_),
    .B(_02258_),
    .X(_03886_));
 sg13g2_a21o_1 _12051_ (.A2(_03874_),
    .A1(_03886_),
    .B1(_03876_),
    .X(_03887_));
 sg13g2_a21o_1 _12052_ (.A2(_03887_),
    .A1(_03881_),
    .B1(_03883_),
    .X(_03888_));
 sg13g2_nor2_1 _12053_ (.A(_02265_),
    .B(_03888_),
    .Y(_03889_));
 sg13g2_a21oi_1 _12054_ (.A1(_02265_),
    .A2(_03888_),
    .Y(_03890_),
    .B1(_03732_));
 sg13g2_nor2_1 _12055_ (.A(_03889_),
    .B(_03890_),
    .Y(_03891_));
 sg13g2_or2_1 _12056_ (.X(_03892_),
    .B(_03891_),
    .A(_02296_));
 sg13g2_or2_1 _12057_ (.X(_03893_),
    .B(_03891_),
    .A(net351));
 sg13g2_a221oi_1 _12058_ (.B2(_03893_),
    .C1(_03852_),
    .B1(_03892_),
    .A1(_03845_),
    .Y(_03894_),
    .A2(_03847_));
 sg13g2_nand2b_1 _12059_ (.Y(_03895_),
    .B(_03879_),
    .A_N(_03873_));
 sg13g2_nor2_1 _12060_ (.A(_03870_),
    .B(_03895_),
    .Y(_03896_));
 sg13g2_and2_1 _12061_ (.A(_03821_),
    .B(_03896_),
    .X(_03897_));
 sg13g2_a21oi_1 _12062_ (.A1(_03856_),
    .A2(_03897_),
    .Y(_03898_),
    .B1(_03891_));
 sg13g2_nor2_1 _12063_ (.A(_03894_),
    .B(_03898_),
    .Y(_03899_));
 sg13g2_xor2_1 _12064_ (.B(\am_sdr0.cic0.integ3[14] ),
    .A(_03742_),
    .X(_03900_));
 sg13g2_xnor2_1 _12065_ (.Y(_03901_),
    .A(_03899_),
    .B(_03900_));
 sg13g2_nor2_1 _12066_ (.A(net116),
    .B(_03901_),
    .Y(_00361_));
 sg13g2_inv_1 _12067_ (.Y(_03902_),
    .A(\am_sdr0.cic0.integ3[14] ));
 sg13g2_nor3_1 _12068_ (.A(_03902_),
    .B(_03894_),
    .C(_03898_),
    .Y(_03903_));
 sg13g2_nand2_1 _12069_ (.Y(_03904_),
    .A(_03742_),
    .B(_03896_));
 sg13g2_nor4_2 _12070_ (.A(_03861_),
    .B(_03864_),
    .C(_03868_),
    .Y(_03905_),
    .D(_03904_));
 sg13g2_nor2_1 _12071_ (.A(_03732_),
    .B(_02265_),
    .Y(_03906_));
 sg13g2_a221oi_1 _12072_ (.B2(_03881_),
    .C1(_03883_),
    .B1(_03876_),
    .A1(_03732_),
    .Y(_03907_),
    .A2(_02265_));
 sg13g2_o21ai_1 _12073_ (.B1(_03902_),
    .Y(_03908_),
    .A1(_03906_),
    .A2(_03907_));
 sg13g2_and2_1 _12074_ (.A(_03742_),
    .B(_03908_),
    .X(_03909_));
 sg13g2_nor3_2 _12075_ (.A(_03903_),
    .B(_03905_),
    .C(_03909_),
    .Y(_03910_));
 sg13g2_xnor2_1 _12076_ (.Y(_03911_),
    .A(_03745_),
    .B(_02268_));
 sg13g2_xnor2_1 _12077_ (.Y(_03912_),
    .A(_03910_),
    .B(_03911_));
 sg13g2_nor2_1 _12078_ (.A(net116),
    .B(_03912_),
    .Y(_00362_));
 sg13g2_xnor2_1 _12079_ (.Y(_03913_),
    .A(net349),
    .B(_02272_));
 sg13g2_or3_1 _12080_ (.A(_03903_),
    .B(_03905_),
    .C(_03909_),
    .X(_03914_));
 sg13g2_or2_1 _12081_ (.X(_03915_),
    .B(_02268_),
    .A(_03745_));
 sg13g2_and2_1 _12082_ (.A(_03745_),
    .B(_02268_),
    .X(_03916_));
 sg13g2_buf_1 _12083_ (.A(_03916_),
    .X(_03917_));
 sg13g2_a21oi_1 _12084_ (.A1(_03914_),
    .A2(_03915_),
    .Y(_03918_),
    .B1(_03917_));
 sg13g2_xnor2_1 _12085_ (.Y(_03919_),
    .A(_03913_),
    .B(_03918_));
 sg13g2_nor2_1 _12086_ (.A(net116),
    .B(_03919_),
    .Y(_00363_));
 sg13g2_o21ai_1 _12087_ (.B1(_02268_),
    .Y(_03920_),
    .A1(net349),
    .A2(_02272_));
 sg13g2_o21ai_1 _12088_ (.B1(_03745_),
    .Y(_03921_),
    .A1(net349),
    .A2(_02272_));
 sg13g2_a21oi_1 _12089_ (.A1(_03920_),
    .A2(_03921_),
    .Y(_03922_),
    .B1(_03910_));
 sg13g2_nor2_1 _12090_ (.A(net349),
    .B(_02272_),
    .Y(_03923_));
 sg13g2_a21oi_1 _12091_ (.A1(_03759_),
    .A2(_02272_),
    .Y(_03924_),
    .B1(_03917_));
 sg13g2_nor2_2 _12092_ (.A(_03923_),
    .B(_03924_),
    .Y(_03925_));
 sg13g2_xnor2_1 _12093_ (.Y(_03926_),
    .A(net348),
    .B(_02275_));
 sg13g2_or3_1 _12094_ (.A(_03922_),
    .B(_03925_),
    .C(_03926_),
    .X(_03927_));
 sg13g2_o21ai_1 _12095_ (.B1(_03926_),
    .Y(_03928_),
    .A1(_03922_),
    .A2(_03925_));
 sg13g2_a21oi_1 _12096_ (.A1(_03927_),
    .A2(_03928_),
    .Y(_00364_),
    .B1(_03429_));
 sg13g2_xnor2_1 _12097_ (.Y(_03929_),
    .A(_03778_),
    .B(_02277_));
 sg13g2_nand2_1 _12098_ (.Y(_03930_),
    .A(net348),
    .B(_02275_));
 sg13g2_nand2_1 _12099_ (.Y(_03931_),
    .A(net364),
    .B(_03930_));
 sg13g2_nor4_1 _12100_ (.A(_03922_),
    .B(_03925_),
    .C(_03929_),
    .D(_03931_),
    .Y(_03932_));
 sg13g2_a221oi_1 _12101_ (.B2(_03915_),
    .C1(_03917_),
    .B1(_03914_),
    .A1(_03759_),
    .Y(_03933_),
    .A2(_02272_));
 sg13g2_inv_1 _12102_ (.Y(_03934_),
    .A(_03929_));
 sg13g2_o21ai_1 _12103_ (.B1(net364),
    .Y(_03935_),
    .A1(net348),
    .A2(_02275_));
 sg13g2_nor4_1 _12104_ (.A(_03923_),
    .B(_03933_),
    .C(_03934_),
    .D(_03935_),
    .Y(_03936_));
 sg13g2_nor4_1 _12105_ (.A(net259),
    .B(net348),
    .C(_02275_),
    .D(_03929_),
    .Y(_03937_));
 sg13g2_nor3_1 _12106_ (.A(net259),
    .B(_03934_),
    .C(_03930_),
    .Y(_03938_));
 sg13g2_or4_1 _12107_ (.A(_03932_),
    .B(_03936_),
    .C(_03937_),
    .D(_03938_),
    .X(_00365_));
 sg13g2_xor2_1 _12108_ (.B(\am_sdr0.cic0.integ3[19] ),
    .A(\am_sdr0.cic0.integ2[22] ),
    .X(_03939_));
 sg13g2_or4_1 _12109_ (.A(_03911_),
    .B(_03913_),
    .C(_03926_),
    .D(_03929_),
    .X(_03940_));
 sg13g2_nand2_1 _12110_ (.Y(_03941_),
    .A(_03778_),
    .B(_02277_));
 sg13g2_nand2_1 _12111_ (.Y(_03942_),
    .A(_02275_),
    .B(_03925_));
 sg13g2_o21ai_1 _12112_ (.B1(_03768_),
    .Y(_03943_),
    .A1(_02275_),
    .A2(_03925_));
 sg13g2_nand3_1 _12113_ (.B(_03942_),
    .C(_03943_),
    .A(_03941_),
    .Y(_03944_));
 sg13g2_o21ai_1 _12114_ (.B1(_03944_),
    .Y(_03945_),
    .A1(_03778_),
    .A2(_02277_));
 sg13g2_o21ai_1 _12115_ (.B1(_03945_),
    .Y(_03946_),
    .A1(_03910_),
    .A2(_03940_));
 sg13g2_xnor2_1 _12116_ (.Y(_03947_),
    .A(_03939_),
    .B(_03946_));
 sg13g2_nor2_1 _12117_ (.A(net116),
    .B(_03947_),
    .Y(_00366_));
 sg13g2_nand2_1 _12118_ (.Y(_03948_),
    .A(_03638_),
    .B(_02247_));
 sg13g2_xnor2_1 _12119_ (.Y(_03949_),
    .A(_03647_),
    .B(_02279_));
 sg13g2_xnor2_1 _12120_ (.Y(_03950_),
    .A(_03948_),
    .B(_03949_));
 sg13g2_nor2_1 _12121_ (.A(net116),
    .B(_03950_),
    .Y(_00367_));
 sg13g2_nor2_1 _12122_ (.A(_03826_),
    .B(_03827_),
    .Y(_03951_));
 sg13g2_xor2_1 _12123_ (.B(_02281_),
    .A(_03635_),
    .X(_03952_));
 sg13g2_xnor2_1 _12124_ (.Y(_03953_),
    .A(_03951_),
    .B(_03952_));
 sg13g2_nor2_1 _12125_ (.A(net116),
    .B(_03953_),
    .Y(_00368_));
 sg13g2_nor2_1 _12126_ (.A(_03824_),
    .B(_03828_),
    .Y(_03954_));
 sg13g2_xnor2_1 _12127_ (.Y(_03955_),
    .A(net354),
    .B(_02284_));
 sg13g2_xnor2_1 _12128_ (.Y(_03956_),
    .A(_03954_),
    .B(_03955_));
 sg13g2_nor2_1 _12129_ (.A(net116),
    .B(_03956_),
    .Y(_00369_));
 sg13g2_xor2_1 _12130_ (.B(_02287_),
    .A(_03655_),
    .X(_03957_));
 sg13g2_xnor2_1 _12131_ (.Y(_03958_),
    .A(_03832_),
    .B(_03957_));
 sg13g2_nor2_1 _12132_ (.A(net116),
    .B(_03958_),
    .Y(_00370_));
 sg13g2_xnor2_1 _12133_ (.Y(_03959_),
    .A(_03656_),
    .B(\am_sdr0.cic0.integ3[5] ));
 sg13g2_and3_1 _12134_ (.X(_03960_),
    .A(_03833_),
    .B(_03835_),
    .C(_03959_));
 sg13g2_a21oi_1 _12135_ (.A1(_03833_),
    .A2(_03835_),
    .Y(_03961_),
    .B1(_03959_));
 sg13g2_nor3_1 _12136_ (.A(net177),
    .B(_03960_),
    .C(_03961_),
    .Y(_00371_));
 sg13g2_buf_1 _12137_ (.A(_01445_),
    .X(_03962_));
 sg13g2_buf_1 _12138_ (.A(_03962_),
    .X(_03963_));
 sg13g2_xor2_1 _12139_ (.B(_02290_),
    .A(_03679_),
    .X(_03964_));
 sg13g2_xnor2_1 _12140_ (.Y(_03965_),
    .A(_03839_),
    .B(_03964_));
 sg13g2_nor2_1 _12141_ (.A(net115),
    .B(_03965_),
    .Y(_00372_));
 sg13g2_nand2_1 _12142_ (.Y(_03966_),
    .A(_02290_),
    .B(_03839_));
 sg13g2_nand2_1 _12143_ (.Y(_03967_),
    .A(_03966_),
    .B(_03843_));
 sg13g2_xor2_1 _12144_ (.B(_02292_),
    .A(_03683_),
    .X(_03968_));
 sg13g2_xnor2_1 _12145_ (.Y(_03969_),
    .A(_03967_),
    .B(_03968_));
 sg13g2_nor2_1 _12146_ (.A(net115),
    .B(_03969_),
    .Y(_00373_));
 sg13g2_a21oi_1 _12147_ (.A1(_03966_),
    .A2(_03843_),
    .Y(_03970_),
    .B1(_03846_));
 sg13g2_a21oi_1 _12148_ (.A1(_03683_),
    .A2(_02292_),
    .Y(_03971_),
    .B1(_03970_));
 sg13g2_xnor2_1 _12149_ (.Y(_03972_),
    .A(_03686_),
    .B(_02294_));
 sg13g2_xnor2_1 _12150_ (.Y(_03973_),
    .A(_03971_),
    .B(_03972_));
 sg13g2_nor2_1 _12151_ (.A(net115),
    .B(_03973_),
    .Y(_00374_));
 sg13g2_xor2_1 _12152_ (.B(_02296_),
    .A(_03703_),
    .X(_03974_));
 sg13g2_xnor2_1 _12153_ (.Y(_03975_),
    .A(_03853_),
    .B(_03974_));
 sg13g2_nor2_1 _12154_ (.A(net115),
    .B(_03975_),
    .Y(_00375_));
 sg13g2_nand2_1 _12155_ (.Y(_03976_),
    .A(net180),
    .B(\am_sdr0.cic0.comb3[14] ));
 sg13g2_buf_1 _12156_ (.A(\am_sdr0.cic0.x_out[10] ),
    .X(_03977_));
 sg13g2_nand2_1 _12157_ (.Y(_03978_),
    .A(_03977_),
    .B(_03418_));
 sg13g2_a21oi_1 _12158_ (.A1(_03976_),
    .A2(_03978_),
    .Y(_00398_),
    .B1(net121));
 sg13g2_nand2_1 _12159_ (.Y(_03979_),
    .A(net180),
    .B(\am_sdr0.cic0.comb3[15] ));
 sg13g2_nand2_1 _12160_ (.Y(_03980_),
    .A(\am_sdr0.cic0.x_out[11] ),
    .B(net176));
 sg13g2_a21oi_1 _12161_ (.A1(_03979_),
    .A2(_03980_),
    .Y(_00399_),
    .B1(_03429_));
 sg13g2_nand2_1 _12162_ (.Y(_03981_),
    .A(net180),
    .B(\am_sdr0.cic0.comb3[16] ));
 sg13g2_buf_1 _12163_ (.A(\am_sdr0.cic0.x_out[12] ),
    .X(_03982_));
 sg13g2_nand2_1 _12164_ (.Y(_03983_),
    .A(_03982_),
    .B(net176));
 sg13g2_a21oi_1 _12165_ (.A1(_03981_),
    .A2(_03983_),
    .Y(_00400_),
    .B1(net121));
 sg13g2_nand2_1 _12166_ (.Y(_03984_),
    .A(net180),
    .B(\am_sdr0.cic0.comb3[17] ));
 sg13g2_nand2_1 _12167_ (.Y(_03985_),
    .A(\am_sdr0.cic0.x_out[13] ),
    .B(net176));
 sg13g2_a21oi_1 _12168_ (.A1(_03984_),
    .A2(_03985_),
    .Y(_00401_),
    .B1(net121));
 sg13g2_nand2_1 _12169_ (.Y(_03986_),
    .A(_02718_),
    .B(\am_sdr0.cic0.comb3[18] ));
 sg13g2_buf_1 _12170_ (.A(\am_sdr0.cic0.x_out[14] ),
    .X(_03987_));
 sg13g2_nand2_1 _12171_ (.Y(_03988_),
    .A(_03987_),
    .B(net176));
 sg13g2_buf_1 _12172_ (.A(_03428_),
    .X(_03989_));
 sg13g2_a21oi_1 _12173_ (.A1(_03986_),
    .A2(_03988_),
    .Y(_00402_),
    .B1(net114));
 sg13g2_nand2_1 _12174_ (.Y(_03990_),
    .A(net171),
    .B(\am_sdr0.cic0.comb3[19] ));
 sg13g2_buf_1 _12175_ (.A(\am_sdr0.cic0.x_out[15] ),
    .X(_03991_));
 sg13g2_buf_1 _12176_ (.A(_03991_),
    .X(_03992_));
 sg13g2_buf_1 _12177_ (.A(net292),
    .X(_03993_));
 sg13g2_nand2_1 _12178_ (.Y(_03994_),
    .A(_03993_),
    .B(net176));
 sg13g2_a21oi_1 _12179_ (.A1(_03990_),
    .A2(_03994_),
    .Y(_00403_),
    .B1(net114));
 sg13g2_nand2_1 _12180_ (.Y(_03995_),
    .A(_03004_),
    .B(\am_sdr0.cic0.comb3[12] ));
 sg13g2_nand2_1 _12181_ (.Y(_03996_),
    .A(\am_sdr0.cic0.x_out[8] ),
    .B(_02786_));
 sg13g2_a21oi_1 _12182_ (.A1(_03995_),
    .A2(_03996_),
    .Y(_00404_),
    .B1(net114));
 sg13g2_nand2_1 _12183_ (.Y(_03997_),
    .A(_03004_),
    .B(\am_sdr0.cic0.comb3[13] ));
 sg13g2_buf_1 _12184_ (.A(\am_sdr0.cic0.x_out[9] ),
    .X(_03998_));
 sg13g2_nand2_1 _12185_ (.Y(_03999_),
    .A(_03998_),
    .B(_02786_));
 sg13g2_a21oi_1 _12186_ (.A1(_03997_),
    .A2(_03999_),
    .Y(_00405_),
    .B1(net114));
 sg13g2_buf_1 _12187_ (.A(\am_sdr0.cic1.sample ),
    .X(_04000_));
 sg13g2_buf_1 _12188_ (.A(_04000_),
    .X(_04001_));
 sg13g2_buf_1 _12189_ (.A(net291),
    .X(_04002_));
 sg13g2_xnor2_1 _12190_ (.Y(_04003_),
    .A(_02298_),
    .B(\am_sdr0.cic1.comb1_in_del[0] ));
 sg13g2_buf_1 _12191_ (.A(\am_sdr0.cic1.comb1[0] ),
    .X(_04004_));
 sg13g2_buf_1 _12192_ (.A(_04000_),
    .X(_04005_));
 sg13g2_buf_1 _12193_ (.A(_04005_),
    .X(_04006_));
 sg13g2_o21ai_1 _12194_ (.B1(net244),
    .Y(_04007_),
    .A1(_04004_),
    .A2(net239));
 sg13g2_a21oi_1 _12195_ (.A1(net240),
    .A2(_04003_),
    .Y(_00406_),
    .B1(_04007_));
 sg13g2_buf_1 _12196_ (.A(\am_sdr0.cic1.comb1[10] ),
    .X(_04008_));
 sg13g2_inv_1 _12197_ (.Y(_04009_),
    .A(_04000_));
 sg13g2_buf_1 _12198_ (.A(_04009_),
    .X(_04010_));
 sg13g2_buf_1 _12199_ (.A(_04010_),
    .X(_04011_));
 sg13g2_buf_1 _12200_ (.A(net162),
    .X(_04012_));
 sg13g2_nand2_1 _12201_ (.Y(_04013_),
    .A(_04008_),
    .B(_04012_));
 sg13g2_buf_1 _12202_ (.A(_04005_),
    .X(_04014_));
 sg13g2_inv_1 _12203_ (.Y(_04015_),
    .A(_02341_));
 sg13g2_buf_1 _12204_ (.A(\am_sdr0.cic1.comb1_in_del[2] ),
    .X(_04016_));
 sg13g2_nor2_1 _12205_ (.A(_02337_),
    .B(_04016_),
    .Y(_04017_));
 sg13g2_nor2b_1 _12206_ (.A(_02298_),
    .B_N(\am_sdr0.cic1.comb1_in_del[0] ),
    .Y(_04018_));
 sg13g2_buf_1 _12207_ (.A(\am_sdr0.cic1.comb1_in_del[1] ),
    .X(_04019_));
 sg13g2_nand2b_1 _12208_ (.Y(_04020_),
    .B(_02336_),
    .A_N(_04019_));
 sg13g2_nor2b_1 _12209_ (.A(_02336_),
    .B_N(_04019_),
    .Y(_04021_));
 sg13g2_a221oi_1 _12210_ (.B2(_04020_),
    .C1(_04021_),
    .B1(_04018_),
    .A1(_02337_),
    .Y(_04022_),
    .A2(_04016_));
 sg13g2_buf_1 _12211_ (.A(_04022_),
    .X(_04023_));
 sg13g2_inv_1 _12212_ (.Y(_04024_),
    .A(\am_sdr0.cic1.comb1_in_del[3] ));
 sg13g2_o21ai_1 _12213_ (.B1(_04024_),
    .Y(_04025_),
    .A1(_04017_),
    .A2(_04023_));
 sg13g2_nor3_1 _12214_ (.A(_04024_),
    .B(_04017_),
    .C(_04023_),
    .Y(_04026_));
 sg13g2_a21o_1 _12215_ (.A2(_04025_),
    .A1(_04015_),
    .B1(_04026_),
    .X(_04027_));
 sg13g2_buf_1 _12216_ (.A(_04027_),
    .X(_04028_));
 sg13g2_nand2b_1 _12217_ (.Y(_04029_),
    .B(_02345_),
    .A_N(\am_sdr0.cic1.comb1_in_del[4] ));
 sg13g2_buf_1 _12218_ (.A(\am_sdr0.cic1.comb1_in_del[5] ),
    .X(_04030_));
 sg13g2_nand2b_1 _12219_ (.Y(_04031_),
    .B(\am_sdr0.cic1.comb1_in_del[4] ),
    .A_N(_02345_));
 sg13g2_buf_1 _12220_ (.A(_04031_),
    .X(_04032_));
 sg13g2_nand2b_1 _12221_ (.Y(_04033_),
    .B(_04032_),
    .A_N(_04030_));
 sg13g2_nand2_1 _12222_ (.Y(_04034_),
    .A(_02348_),
    .B(_04032_));
 sg13g2_buf_1 _12223_ (.A(\am_sdr0.cic1.comb1_in_del[7] ),
    .X(_04035_));
 sg13g2_nand2b_1 _12224_ (.Y(_04036_),
    .B(_04035_),
    .A_N(_02353_));
 sg13g2_buf_1 _12225_ (.A(_04036_),
    .X(_04037_));
 sg13g2_buf_1 _12226_ (.A(\am_sdr0.cic1.comb1_in_del[8] ),
    .X(_04038_));
 sg13g2_inv_1 _12227_ (.Y(_04039_),
    .A(_04038_));
 sg13g2_o21ai_1 _12228_ (.B1(_04039_),
    .Y(_04040_),
    .A1(_02355_),
    .A2(_04037_));
 sg13g2_nand2_1 _12229_ (.Y(_04041_),
    .A(_02355_),
    .B(_04037_));
 sg13g2_buf_1 _12230_ (.A(\am_sdr0.cic1.comb1_in_del[6] ),
    .X(_04042_));
 sg13g2_nor2b_1 _12231_ (.A(_02351_),
    .B_N(_04042_),
    .Y(_04043_));
 sg13g2_a21o_1 _12232_ (.A2(_04041_),
    .A1(_04040_),
    .B1(_04043_),
    .X(_04044_));
 sg13g2_a221oi_1 _12233_ (.B2(_04034_),
    .C1(_04044_),
    .B1(_04033_),
    .A1(_04028_),
    .Y(_04045_),
    .A2(_04029_));
 sg13g2_buf_2 _12234_ (.A(_04045_),
    .X(_04046_));
 sg13g2_nand2b_1 _12235_ (.Y(_04047_),
    .B(_02348_),
    .A_N(_04030_));
 sg13g2_nand2b_1 _12236_ (.Y(_04048_),
    .B(_02353_),
    .A_N(_04035_));
 sg13g2_nand3b_1 _12237_ (.B(_04037_),
    .C(_02351_),
    .Y(_04049_),
    .A_N(_04042_));
 sg13g2_a22oi_1 _12238_ (.Y(_04050_),
    .B1(_04048_),
    .B2(_04049_),
    .A2(_04038_),
    .A1(_02356_));
 sg13g2_a21oi_1 _12239_ (.A1(_02355_),
    .A2(_04039_),
    .Y(_04051_),
    .B1(_04050_));
 sg13g2_o21ai_1 _12240_ (.B1(_04051_),
    .Y(_04052_),
    .A1(_04044_),
    .A2(_04047_));
 sg13g2_buf_1 _12241_ (.A(_04052_),
    .X(_04053_));
 sg13g2_buf_1 _12242_ (.A(\am_sdr0.cic1.comb1_in_del[9] ),
    .X(_04054_));
 sg13g2_inv_1 _12243_ (.Y(_04055_),
    .A(_04054_));
 sg13g2_o21ai_1 _12244_ (.B1(_04055_),
    .Y(_04056_),
    .A1(_04046_),
    .A2(_04053_));
 sg13g2_nor3_1 _12245_ (.A(_04055_),
    .B(_04046_),
    .C(_04053_),
    .Y(_04057_));
 sg13g2_a21oi_1 _12246_ (.A1(_02360_),
    .A2(_04056_),
    .Y(_04058_),
    .B1(_04057_));
 sg13g2_buf_1 _12247_ (.A(\am_sdr0.cic1.comb1_in_del[10] ),
    .X(_04059_));
 sg13g2_nor2b_1 _12248_ (.A(_04059_),
    .B_N(_02310_),
    .Y(_04060_));
 sg13g2_nand2b_1 _12249_ (.Y(_04061_),
    .B(_04059_),
    .A_N(_02310_));
 sg13g2_nand2b_1 _12250_ (.Y(_04062_),
    .B(_04061_),
    .A_N(_04060_));
 sg13g2_xnor2_1 _12251_ (.Y(_04063_),
    .A(_04058_),
    .B(_04062_));
 sg13g2_nand2_1 _12252_ (.Y(_04064_),
    .A(_04014_),
    .B(_04063_));
 sg13g2_a21oi_1 _12253_ (.A1(_04013_),
    .A2(_04064_),
    .Y(_00407_),
    .B1(net114));
 sg13g2_buf_1 _12254_ (.A(\am_sdr0.cic1.comb1[11] ),
    .X(_04065_));
 sg13g2_buf_1 _12255_ (.A(_04005_),
    .X(_04066_));
 sg13g2_buf_1 _12256_ (.A(_04005_),
    .X(_04067_));
 sg13g2_o21ai_1 _12257_ (.B1(_04061_),
    .Y(_04068_),
    .A1(_04058_),
    .A2(_04060_));
 sg13g2_buf_2 _12258_ (.A(\am_sdr0.cic1.comb1_in_del[11] ),
    .X(_04069_));
 sg13g2_xor2_1 _12259_ (.B(_04069_),
    .A(_02315_),
    .X(_04070_));
 sg13g2_xnor2_1 _12260_ (.Y(_04071_),
    .A(_04068_),
    .B(_04070_));
 sg13g2_nand2_1 _12261_ (.Y(_04072_),
    .A(net236),
    .B(_04071_));
 sg13g2_o21ai_1 _12262_ (.B1(_04072_),
    .Y(_04073_),
    .A1(_04065_),
    .A2(net237));
 sg13g2_nor2_1 _12263_ (.A(net115),
    .B(_04073_),
    .Y(_00408_));
 sg13g2_nor2_1 _12264_ (.A(\am_sdr0.cic1.comb1[12] ),
    .B(net239),
    .Y(_04074_));
 sg13g2_buf_1 _12265_ (.A(_04010_),
    .X(_04075_));
 sg13g2_or2_1 _12266_ (.X(_04076_),
    .B(_04069_),
    .A(_04059_));
 sg13g2_inv_1 _12267_ (.Y(_04077_),
    .A(_04069_));
 sg13g2_nand2_1 _12268_ (.Y(_04078_),
    .A(_02310_),
    .B(_04077_));
 sg13g2_a221oi_1 _12269_ (.B2(_04078_),
    .C1(_04057_),
    .B1(_04076_),
    .A1(_02360_),
    .Y(_04079_),
    .A2(_04056_));
 sg13g2_a21oi_1 _12270_ (.A1(_04077_),
    .A2(_04060_),
    .Y(_04080_),
    .B1(_02315_));
 sg13g2_nand2b_1 _12271_ (.Y(_04081_),
    .B(_04080_),
    .A_N(_04079_));
 sg13g2_nand3_1 _12272_ (.B(_04059_),
    .C(_04069_),
    .A(_04054_),
    .Y(_04082_));
 sg13g2_nor3_1 _12273_ (.A(_04046_),
    .B(_04053_),
    .C(_04082_),
    .Y(_04083_));
 sg13g2_nand2_1 _12274_ (.Y(_04084_),
    .A(_02360_),
    .B(_04059_));
 sg13g2_nor4_1 _12275_ (.A(_04077_),
    .B(_04046_),
    .C(_04053_),
    .D(_04084_),
    .Y(_04085_));
 sg13g2_nand2b_1 _12276_ (.Y(_04086_),
    .B(_04054_),
    .A_N(_02310_));
 sg13g2_nor4_1 _12277_ (.A(_04077_),
    .B(_04046_),
    .C(_04053_),
    .D(_04086_),
    .Y(_04087_));
 sg13g2_or2_1 _12278_ (.X(_04088_),
    .B(_02310_),
    .A(_02359_));
 sg13g2_nor4_1 _12279_ (.A(_04077_),
    .B(_04046_),
    .C(_04053_),
    .D(_04088_),
    .Y(_04089_));
 sg13g2_or4_1 _12280_ (.A(_04083_),
    .B(_04085_),
    .C(_04087_),
    .D(_04089_),
    .X(_04090_));
 sg13g2_buf_1 _12281_ (.A(_04090_),
    .X(_04091_));
 sg13g2_nor2_1 _12282_ (.A(_04077_),
    .B(_04061_),
    .Y(_04092_));
 sg13g2_nor2_1 _12283_ (.A(_02359_),
    .B(_04055_),
    .Y(_04093_));
 sg13g2_nand3_1 _12284_ (.B(_04069_),
    .C(_04093_),
    .A(_04059_),
    .Y(_04094_));
 sg13g2_nand3b_1 _12285_ (.B(_04069_),
    .C(_04093_),
    .Y(_04095_),
    .A_N(_02310_));
 sg13g2_nand3b_1 _12286_ (.B(_04094_),
    .C(_04095_),
    .Y(_04096_),
    .A_N(_04092_));
 sg13g2_buf_1 _12287_ (.A(_04096_),
    .X(_04097_));
 sg13g2_nor2_1 _12288_ (.A(_04091_),
    .B(_04097_),
    .Y(_04098_));
 sg13g2_and2_1 _12289_ (.A(_04081_),
    .B(_04098_),
    .X(_04099_));
 sg13g2_buf_1 _12290_ (.A(\am_sdr0.cic1.comb1_in_del[12] ),
    .X(_04100_));
 sg13g2_xor2_1 _12291_ (.B(_04100_),
    .A(_02319_),
    .X(_04101_));
 sg13g2_xnor2_1 _12292_ (.Y(_04102_),
    .A(_04099_),
    .B(_04101_));
 sg13g2_nor2_1 _12293_ (.A(net161),
    .B(_04102_),
    .Y(_04103_));
 sg13g2_nor3_1 _12294_ (.A(_02781_),
    .B(_04074_),
    .C(_04103_),
    .Y(_00409_));
 sg13g2_buf_2 _12295_ (.A(\am_sdr0.cic1.comb1[13] ),
    .X(_04104_));
 sg13g2_nor2b_1 _12296_ (.A(_04100_),
    .B_N(_02319_),
    .Y(_04105_));
 sg13g2_nand2b_1 _12297_ (.Y(_04106_),
    .B(_04100_),
    .A_N(_02319_));
 sg13g2_o21ai_1 _12298_ (.B1(_04106_),
    .Y(_04107_),
    .A1(_04099_),
    .A2(_04105_));
 sg13g2_xor2_1 _12299_ (.B(\am_sdr0.cic1.comb1_in_del[13] ),
    .A(_02322_),
    .X(_04108_));
 sg13g2_xnor2_1 _12300_ (.Y(_04109_),
    .A(_04107_),
    .B(_04108_));
 sg13g2_nand2_1 _12301_ (.Y(_04110_),
    .A(net236),
    .B(_04109_));
 sg13g2_o21ai_1 _12302_ (.B1(_04110_),
    .Y(_04111_),
    .A1(_04104_),
    .A2(_04066_));
 sg13g2_nor2_1 _12303_ (.A(net115),
    .B(_04111_),
    .Y(_00410_));
 sg13g2_buf_1 _12304_ (.A(\am_sdr0.cic1.comb1[14] ),
    .X(_04112_));
 sg13g2_buf_1 _12305_ (.A(_04005_),
    .X(_04113_));
 sg13g2_nand2_1 _12306_ (.Y(_04114_),
    .A(_02322_),
    .B(_04106_));
 sg13g2_nor3_1 _12307_ (.A(_04091_),
    .B(_04097_),
    .C(_04114_),
    .Y(_04115_));
 sg13g2_inv_1 _12308_ (.Y(_04116_),
    .A(\am_sdr0.cic1.comb1_in_del[13] ));
 sg13g2_nand2_1 _12309_ (.Y(_04117_),
    .A(_04116_),
    .B(_04106_));
 sg13g2_nor3_1 _12310_ (.A(_04091_),
    .B(_04097_),
    .C(_04117_),
    .Y(_04118_));
 sg13g2_o21ai_1 _12311_ (.B1(_04081_),
    .Y(_04119_),
    .A1(_04115_),
    .A2(_04118_));
 sg13g2_nand2_1 _12312_ (.Y(_04120_),
    .A(_02322_),
    .B(_04116_));
 sg13g2_o21ai_1 _12313_ (.B1(_04105_),
    .Y(_04121_),
    .A1(_02322_),
    .A2(_04116_));
 sg13g2_and2_1 _12314_ (.A(_04120_),
    .B(_04121_),
    .X(_04122_));
 sg13g2_buf_1 _12315_ (.A(_04122_),
    .X(_04123_));
 sg13g2_and2_1 _12316_ (.A(_04119_),
    .B(_04123_),
    .X(_04124_));
 sg13g2_nand2b_1 _12317_ (.Y(_04125_),
    .B(\am_sdr0.cic1.comb1_in_del[14] ),
    .A_N(_02324_));
 sg13g2_buf_1 _12318_ (.A(_04125_),
    .X(_04126_));
 sg13g2_nand2b_1 _12319_ (.Y(_04127_),
    .B(_02324_),
    .A_N(\am_sdr0.cic1.comb1_in_del[14] ));
 sg13g2_buf_1 _12320_ (.A(_04127_),
    .X(_04128_));
 sg13g2_nand2_1 _12321_ (.Y(_04129_),
    .A(_04126_),
    .B(_04128_));
 sg13g2_xnor2_1 _12322_ (.Y(_04130_),
    .A(_04124_),
    .B(_04129_));
 sg13g2_nand2_1 _12323_ (.Y(_04131_),
    .A(_04113_),
    .B(_04130_));
 sg13g2_o21ai_1 _12324_ (.B1(_04131_),
    .Y(_04132_),
    .A1(_04112_),
    .A2(_04066_));
 sg13g2_nor2_1 _12325_ (.A(net115),
    .B(_04132_),
    .Y(_00411_));
 sg13g2_buf_1 _12326_ (.A(\am_sdr0.cic1.comb1[15] ),
    .X(_04133_));
 sg13g2_nand2_1 _12327_ (.Y(_04134_),
    .A(_04133_),
    .B(net113));
 sg13g2_nand2_1 _12328_ (.Y(_04135_),
    .A(_04124_),
    .B(_04128_));
 sg13g2_buf_1 _12329_ (.A(\am_sdr0.cic1.comb1_in_del[15] ),
    .X(_04136_));
 sg13g2_xnor2_1 _12330_ (.Y(_04137_),
    .A(_02325_),
    .B(_04136_));
 sg13g2_a21oi_1 _12331_ (.A1(_04126_),
    .A2(_04135_),
    .Y(_04138_),
    .B1(_04137_));
 sg13g2_nand3_1 _12332_ (.B(_04135_),
    .C(_04137_),
    .A(_04126_),
    .Y(_04139_));
 sg13g2_nand3b_1 _12333_ (.B(net236),
    .C(_04139_),
    .Y(_04140_),
    .A_N(_04138_));
 sg13g2_a21oi_1 _12334_ (.A1(_04134_),
    .A2(_04140_),
    .Y(_00412_),
    .B1(net114));
 sg13g2_buf_1 _12335_ (.A(\am_sdr0.cic1.comb1[16] ),
    .X(_04141_));
 sg13g2_nand2_1 _12336_ (.Y(_04142_),
    .A(_04141_),
    .B(net113));
 sg13g2_buf_1 _12337_ (.A(_04005_),
    .X(_04143_));
 sg13g2_and4_1 _12338_ (.A(_04136_),
    .B(_04119_),
    .C(_04123_),
    .D(_04128_),
    .X(_04144_));
 sg13g2_and4_1 _12339_ (.A(_02326_),
    .B(_04119_),
    .C(_04123_),
    .D(_04128_),
    .X(_04145_));
 sg13g2_inv_1 _12340_ (.Y(_04146_),
    .A(_04136_));
 sg13g2_a21o_1 _12341_ (.A2(_04146_),
    .A1(_02325_),
    .B1(_04126_),
    .X(_04147_));
 sg13g2_o21ai_1 _12342_ (.B1(_04147_),
    .Y(_04148_),
    .A1(_02325_),
    .A2(_04146_));
 sg13g2_or3_1 _12343_ (.A(_04144_),
    .B(_04145_),
    .C(_04148_),
    .X(_04149_));
 sg13g2_buf_1 _12344_ (.A(\am_sdr0.cic1.comb1_in_del[16] ),
    .X(_04150_));
 sg13g2_xnor2_1 _12345_ (.Y(_04151_),
    .A(_02330_),
    .B(_04150_));
 sg13g2_xnor2_1 _12346_ (.Y(_04152_),
    .A(_04149_),
    .B(_04151_));
 sg13g2_nand2_1 _12347_ (.Y(_04153_),
    .A(_04143_),
    .B(_04152_));
 sg13g2_a21oi_1 _12348_ (.A1(_04142_),
    .A2(_04153_),
    .Y(_00413_),
    .B1(net114));
 sg13g2_buf_1 _12349_ (.A(\am_sdr0.cic1.comb1[17] ),
    .X(_04154_));
 sg13g2_nor2_1 _12350_ (.A(_04154_),
    .B(net239),
    .Y(_04155_));
 sg13g2_inv_1 _12351_ (.Y(_04156_),
    .A(_04150_));
 sg13g2_nor3_1 _12352_ (.A(_04144_),
    .B(_04145_),
    .C(_04148_),
    .Y(_04157_));
 sg13g2_a21oi_1 _12353_ (.A1(_04156_),
    .A2(_04157_),
    .Y(_04158_),
    .B1(_02330_));
 sg13g2_a21oi_1 _12354_ (.A1(_04150_),
    .A2(_04149_),
    .Y(_04159_),
    .B1(_04158_));
 sg13g2_xor2_1 _12355_ (.B(\am_sdr0.cic1.comb1_in_del[17] ),
    .A(_02332_),
    .X(_04160_));
 sg13g2_xnor2_1 _12356_ (.Y(_04161_),
    .A(_04159_),
    .B(_04160_));
 sg13g2_nor2_1 _12357_ (.A(net161),
    .B(_04161_),
    .Y(_04162_));
 sg13g2_nor3_1 _12358_ (.A(_02781_),
    .B(_04155_),
    .C(_04162_),
    .Y(_00414_));
 sg13g2_inv_1 _12359_ (.Y(_04163_),
    .A(\am_sdr0.cic1.comb1_in_del[17] ));
 sg13g2_nor2_1 _12360_ (.A(_02332_),
    .B(_04163_),
    .Y(_04164_));
 sg13g2_a221oi_1 _12361_ (.B2(_04163_),
    .C1(_04157_),
    .B1(_02332_),
    .A1(_02330_),
    .Y(_04165_),
    .A2(_04156_));
 sg13g2_nand2b_1 _12362_ (.Y(_04166_),
    .B(_04150_),
    .A_N(_02330_));
 sg13g2_a21oi_1 _12363_ (.A1(_02332_),
    .A2(_04163_),
    .Y(_04167_),
    .B1(_04166_));
 sg13g2_nor3_1 _12364_ (.A(_04164_),
    .B(_04165_),
    .C(_04167_),
    .Y(_04168_));
 sg13g2_buf_1 _12365_ (.A(\am_sdr0.cic1.comb1_in_del[18] ),
    .X(_04169_));
 sg13g2_xnor2_1 _12366_ (.Y(_04170_),
    .A(_02334_),
    .B(_04169_));
 sg13g2_xnor2_1 _12367_ (.Y(_04171_),
    .A(_04168_),
    .B(_04170_));
 sg13g2_buf_1 _12368_ (.A(\am_sdr0.cic1.comb1[18] ),
    .X(_04172_));
 sg13g2_o21ai_1 _12369_ (.B1(net244),
    .Y(_04173_),
    .A1(_04172_),
    .A2(net239));
 sg13g2_a21oi_1 _12370_ (.A1(net240),
    .A2(_04171_),
    .Y(_00415_),
    .B1(_04173_));
 sg13g2_nor2b_1 _12371_ (.A(_04169_),
    .B_N(_02334_),
    .Y(_04174_));
 sg13g2_nand2b_1 _12372_ (.Y(_04175_),
    .B(_04169_),
    .A_N(_02334_));
 sg13g2_o21ai_1 _12373_ (.B1(_04175_),
    .Y(_04176_),
    .A1(_04168_),
    .A2(_04174_));
 sg13g2_xor2_1 _12374_ (.B(\am_sdr0.cic1.comb1_in_del[19] ),
    .A(\am_sdr0.cic1.integ_sample[19] ),
    .X(_04177_));
 sg13g2_xnor2_1 _12375_ (.Y(_04178_),
    .A(_04176_),
    .B(_04177_));
 sg13g2_o21ai_1 _12376_ (.B1(net244),
    .Y(_04179_),
    .A1(\am_sdr0.cic1.comb1[19] ),
    .A2(_04006_));
 sg13g2_a21oi_1 _12377_ (.A1(net240),
    .A2(_04178_),
    .Y(_00416_),
    .B1(_04179_));
 sg13g2_buf_1 _12378_ (.A(\am_sdr0.cic1.comb1[1] ),
    .X(_04180_));
 sg13g2_nand2_1 _12379_ (.Y(_04181_),
    .A(_04180_),
    .B(net113));
 sg13g2_xnor2_1 _12380_ (.Y(_04182_),
    .A(_02336_),
    .B(_04019_));
 sg13g2_xnor2_1 _12381_ (.Y(_04183_),
    .A(_04018_),
    .B(_04182_));
 sg13g2_nand2_1 _12382_ (.Y(_04184_),
    .A(net234),
    .B(_04183_));
 sg13g2_a21oi_1 _12383_ (.A1(_04181_),
    .A2(_04184_),
    .Y(_00417_),
    .B1(net114));
 sg13g2_buf_1 _12384_ (.A(\am_sdr0.cic1.comb1[2] ),
    .X(_04185_));
 sg13g2_buf_1 _12385_ (.A(net162),
    .X(_04186_));
 sg13g2_a21oi_1 _12386_ (.A1(_04018_),
    .A2(_04020_),
    .Y(_04187_),
    .B1(_04021_));
 sg13g2_xnor2_1 _12387_ (.Y(_04188_),
    .A(\am_sdr0.cic1.integ_sample[2] ),
    .B(_04016_));
 sg13g2_xnor2_1 _12388_ (.Y(_04189_),
    .A(_04187_),
    .B(_04188_));
 sg13g2_nor2_1 _12389_ (.A(net162),
    .B(_04189_),
    .Y(_04190_));
 sg13g2_a21oi_1 _12390_ (.A1(_04185_),
    .A2(net112),
    .Y(_04191_),
    .B1(_04190_));
 sg13g2_nor2_1 _12391_ (.A(net115),
    .B(_04191_),
    .Y(_00418_));
 sg13g2_buf_1 _12392_ (.A(\am_sdr0.cic1.comb1[3] ),
    .X(_04192_));
 sg13g2_nand2_1 _12393_ (.Y(_04193_),
    .A(_04192_),
    .B(net113));
 sg13g2_nor2_1 _12394_ (.A(_04017_),
    .B(_04023_),
    .Y(_04194_));
 sg13g2_xnor2_1 _12395_ (.Y(_04195_),
    .A(_02341_),
    .B(\am_sdr0.cic1.comb1_in_del[3] ));
 sg13g2_xnor2_1 _12396_ (.Y(_04196_),
    .A(_04194_),
    .B(_04195_));
 sg13g2_nand2_1 _12397_ (.Y(_04197_),
    .A(net234),
    .B(_04196_));
 sg13g2_a21oi_1 _12398_ (.A1(_04193_),
    .A2(_04197_),
    .Y(_00419_),
    .B1(_03989_));
 sg13g2_buf_1 _12399_ (.A(_01445_),
    .X(_04198_));
 sg13g2_buf_1 _12400_ (.A(\am_sdr0.cic1.comb1[4] ),
    .X(_04199_));
 sg13g2_nor2_1 _12401_ (.A(_04199_),
    .B(net239),
    .Y(_04200_));
 sg13g2_nand2_1 _12402_ (.Y(_04201_),
    .A(_04029_),
    .B(_04032_));
 sg13g2_xor2_1 _12403_ (.B(_04201_),
    .A(_04028_),
    .X(_04202_));
 sg13g2_nor2_1 _12404_ (.A(net161),
    .B(_04202_),
    .Y(_04203_));
 sg13g2_nor3_1 _12405_ (.A(net160),
    .B(_04200_),
    .C(_04203_),
    .Y(_00420_));
 sg13g2_buf_2 _12406_ (.A(\am_sdr0.cic1.comb1[5] ),
    .X(_04204_));
 sg13g2_nand2_1 _12407_ (.Y(_04205_),
    .A(_04028_),
    .B(_04029_));
 sg13g2_nand2_1 _12408_ (.Y(_04206_),
    .A(_04205_),
    .B(_04032_));
 sg13g2_xor2_1 _12409_ (.B(_04030_),
    .A(_02348_),
    .X(_04207_));
 sg13g2_xnor2_1 _12410_ (.Y(_04208_),
    .A(_04206_),
    .B(_04207_));
 sg13g2_nand2_1 _12411_ (.Y(_04209_),
    .A(net235),
    .B(_04208_));
 sg13g2_o21ai_1 _12412_ (.B1(_04209_),
    .Y(_04210_),
    .A1(_04204_),
    .A2(net237));
 sg13g2_nor2_1 _12413_ (.A(_03963_),
    .B(_04210_),
    .Y(_00421_));
 sg13g2_buf_2 _12414_ (.A(\am_sdr0.cic1.comb1[6] ),
    .X(_04211_));
 sg13g2_nor2_1 _12415_ (.A(_04030_),
    .B(_04206_),
    .Y(_04212_));
 sg13g2_nand2_1 _12416_ (.Y(_04213_),
    .A(_04030_),
    .B(_04206_));
 sg13g2_o21ai_1 _12417_ (.B1(_04213_),
    .Y(_04214_),
    .A1(_02348_),
    .A2(_04212_));
 sg13g2_buf_1 _12418_ (.A(_04214_),
    .X(_04215_));
 sg13g2_xor2_1 _12419_ (.B(_04042_),
    .A(_02351_),
    .X(_04216_));
 sg13g2_xnor2_1 _12420_ (.Y(_04217_),
    .A(_04215_),
    .B(_04216_));
 sg13g2_nand2_1 _12421_ (.Y(_04218_),
    .A(net235),
    .B(_04217_));
 sg13g2_o21ai_1 _12422_ (.B1(_04218_),
    .Y(_04219_),
    .A1(_04211_),
    .A2(net237));
 sg13g2_nor2_1 _12423_ (.A(_03963_),
    .B(_04219_),
    .Y(_00422_));
 sg13g2_buf_1 _12424_ (.A(_03962_),
    .X(_04220_));
 sg13g2_buf_2 _12425_ (.A(\am_sdr0.cic1.comb1[7] ),
    .X(_04221_));
 sg13g2_nor2_1 _12426_ (.A(_04042_),
    .B(_04215_),
    .Y(_04222_));
 sg13g2_nand2_1 _12427_ (.Y(_04223_),
    .A(_04042_),
    .B(_04215_));
 sg13g2_o21ai_1 _12428_ (.B1(_04223_),
    .Y(_04224_),
    .A1(_02351_),
    .A2(_04222_));
 sg13g2_buf_1 _12429_ (.A(_04224_),
    .X(_04225_));
 sg13g2_nand2_1 _12430_ (.Y(_04226_),
    .A(_04037_),
    .B(_04048_));
 sg13g2_xnor2_1 _12431_ (.Y(_04227_),
    .A(_04225_),
    .B(_04226_));
 sg13g2_nand2_1 _12432_ (.Y(_04228_),
    .A(net235),
    .B(_04227_));
 sg13g2_o21ai_1 _12433_ (.B1(_04228_),
    .Y(_04229_),
    .A1(_04221_),
    .A2(net237));
 sg13g2_nor2_1 _12434_ (.A(net111),
    .B(_04229_),
    .Y(_00423_));
 sg13g2_buf_2 _12435_ (.A(\am_sdr0.cic1.comb1[8] ),
    .X(_04230_));
 sg13g2_nand2_1 _12436_ (.Y(_04231_),
    .A(_04035_),
    .B(_04225_));
 sg13g2_nor2_1 _12437_ (.A(_04035_),
    .B(_04225_),
    .Y(_04232_));
 sg13g2_a21oi_1 _12438_ (.A1(_02353_),
    .A2(_04231_),
    .Y(_04233_),
    .B1(_04232_));
 sg13g2_xor2_1 _12439_ (.B(_04038_),
    .A(_02355_),
    .X(_04234_));
 sg13g2_xnor2_1 _12440_ (.Y(_04235_),
    .A(_04233_),
    .B(_04234_));
 sg13g2_nand2_1 _12441_ (.Y(_04236_),
    .A(net235),
    .B(_04235_));
 sg13g2_o21ai_1 _12442_ (.B1(_04236_),
    .Y(_04237_),
    .A1(_04230_),
    .A2(net237));
 sg13g2_nor2_1 _12443_ (.A(net111),
    .B(_04237_),
    .Y(_00424_));
 sg13g2_buf_1 _12444_ (.A(\am_sdr0.cic1.comb1[9] ),
    .X(_04238_));
 sg13g2_nand2_1 _12445_ (.Y(_04239_),
    .A(_04238_),
    .B(net113));
 sg13g2_nor2_1 _12446_ (.A(_04046_),
    .B(_04053_),
    .Y(_04240_));
 sg13g2_xnor2_1 _12447_ (.Y(_04241_),
    .A(_02359_),
    .B(_04054_));
 sg13g2_xnor2_1 _12448_ (.Y(_04242_),
    .A(_04240_),
    .B(_04241_));
 sg13g2_nand2_1 _12449_ (.Y(_04243_),
    .A(net234),
    .B(_04242_));
 sg13g2_a21oi_1 _12450_ (.A1(_04239_),
    .A2(_04243_),
    .Y(_00425_),
    .B1(_03989_));
 sg13g2_buf_1 _12451_ (.A(net291),
    .X(_04244_));
 sg13g2_nand2_1 _12452_ (.Y(_04245_),
    .A(_02298_),
    .B(_04244_));
 sg13g2_nand2_1 _12453_ (.Y(_04246_),
    .A(\am_sdr0.cic1.comb1_in_del[0] ),
    .B(net112));
 sg13g2_buf_1 _12454_ (.A(_03428_),
    .X(_04247_));
 sg13g2_a21oi_1 _12455_ (.A1(_04245_),
    .A2(_04246_),
    .Y(_00426_),
    .B1(net110));
 sg13g2_buf_1 _12456_ (.A(net291),
    .X(_04248_));
 sg13g2_nand2_1 _12457_ (.Y(_04249_),
    .A(_02310_),
    .B(net232));
 sg13g2_nand2_1 _12458_ (.Y(_04250_),
    .A(_04059_),
    .B(net112));
 sg13g2_a21oi_1 _12459_ (.A1(_04249_),
    .A2(_04250_),
    .Y(_00427_),
    .B1(net110));
 sg13g2_nand2_1 _12460_ (.Y(_04251_),
    .A(_02315_),
    .B(net232));
 sg13g2_nand2_1 _12461_ (.Y(_04252_),
    .A(_04069_),
    .B(net112));
 sg13g2_a21oi_1 _12462_ (.A1(_04251_),
    .A2(_04252_),
    .Y(_00428_),
    .B1(net110));
 sg13g2_nand2_1 _12463_ (.Y(_04253_),
    .A(_02319_),
    .B(net232));
 sg13g2_buf_1 _12464_ (.A(net162),
    .X(_04254_));
 sg13g2_nand2_1 _12465_ (.Y(_04255_),
    .A(_04100_),
    .B(_04254_));
 sg13g2_a21oi_1 _12466_ (.A1(_04253_),
    .A2(_04255_),
    .Y(_00429_),
    .B1(net110));
 sg13g2_nand2_1 _12467_ (.Y(_04256_),
    .A(_02322_),
    .B(net232));
 sg13g2_nand2_1 _12468_ (.Y(_04257_),
    .A(\am_sdr0.cic1.comb1_in_del[13] ),
    .B(net109));
 sg13g2_a21oi_1 _12469_ (.A1(_04256_),
    .A2(_04257_),
    .Y(_00430_),
    .B1(_04247_));
 sg13g2_nand2_1 _12470_ (.Y(_04258_),
    .A(_02324_),
    .B(_04248_));
 sg13g2_nand2_1 _12471_ (.Y(_04259_),
    .A(\am_sdr0.cic1.comb1_in_del[14] ),
    .B(net109));
 sg13g2_a21oi_1 _12472_ (.A1(_04258_),
    .A2(_04259_),
    .Y(_00431_),
    .B1(net110));
 sg13g2_nand2_1 _12473_ (.Y(_04260_),
    .A(_02325_),
    .B(net232));
 sg13g2_nand2_1 _12474_ (.Y(_04261_),
    .A(_04136_),
    .B(net109));
 sg13g2_a21oi_1 _12475_ (.A1(_04260_),
    .A2(_04261_),
    .Y(_00432_),
    .B1(net110));
 sg13g2_nand2_1 _12476_ (.Y(_04262_),
    .A(_02330_),
    .B(net232));
 sg13g2_nand2_1 _12477_ (.Y(_04263_),
    .A(_04150_),
    .B(net109));
 sg13g2_a21oi_1 _12478_ (.A1(_04262_),
    .A2(_04263_),
    .Y(_00433_),
    .B1(net110));
 sg13g2_nand2_1 _12479_ (.Y(_04264_),
    .A(_02332_),
    .B(net232));
 sg13g2_nand2_1 _12480_ (.Y(_04265_),
    .A(\am_sdr0.cic1.comb1_in_del[17] ),
    .B(net109));
 sg13g2_a21oi_1 _12481_ (.A1(_04264_),
    .A2(_04265_),
    .Y(_00434_),
    .B1(net110));
 sg13g2_nand2_1 _12482_ (.Y(_04266_),
    .A(_02334_),
    .B(net232));
 sg13g2_nand2_1 _12483_ (.Y(_04267_),
    .A(_04169_),
    .B(_04254_));
 sg13g2_a21oi_1 _12484_ (.A1(_04266_),
    .A2(_04267_),
    .Y(_00435_),
    .B1(_04247_));
 sg13g2_nand2_1 _12485_ (.Y(_04268_),
    .A(\am_sdr0.cic1.integ_sample[19] ),
    .B(_04248_));
 sg13g2_nand2_1 _12486_ (.Y(_04269_),
    .A(\am_sdr0.cic1.comb1_in_del[19] ),
    .B(net109));
 sg13g2_buf_1 _12487_ (.A(_03428_),
    .X(_04270_));
 sg13g2_a21oi_1 _12488_ (.A1(_04268_),
    .A2(_04269_),
    .Y(_00436_),
    .B1(_04270_));
 sg13g2_buf_1 _12489_ (.A(net291),
    .X(_04271_));
 sg13g2_nand2_1 _12490_ (.Y(_04272_),
    .A(_02336_),
    .B(_04271_));
 sg13g2_nand2_1 _12491_ (.Y(_04273_),
    .A(_04019_),
    .B(net109));
 sg13g2_a21oi_1 _12492_ (.A1(_04272_),
    .A2(_04273_),
    .Y(_00437_),
    .B1(_04270_));
 sg13g2_nand2_1 _12493_ (.Y(_04274_),
    .A(\am_sdr0.cic1.integ_sample[2] ),
    .B(_04271_));
 sg13g2_nand2_1 _12494_ (.Y(_04275_),
    .A(_04016_),
    .B(net109));
 sg13g2_a21oi_1 _12495_ (.A1(_04274_),
    .A2(_04275_),
    .Y(_00438_),
    .B1(net108));
 sg13g2_nand2_1 _12496_ (.Y(_04276_),
    .A(_02341_),
    .B(net231));
 sg13g2_buf_1 _12497_ (.A(net162),
    .X(_04277_));
 sg13g2_nand2_1 _12498_ (.Y(_04278_),
    .A(\am_sdr0.cic1.comb1_in_del[3] ),
    .B(net107));
 sg13g2_a21oi_1 _12499_ (.A1(_04276_),
    .A2(_04278_),
    .Y(_00439_),
    .B1(net108));
 sg13g2_nand2_1 _12500_ (.Y(_04279_),
    .A(_02345_),
    .B(net231));
 sg13g2_nand2_1 _12501_ (.Y(_04280_),
    .A(\am_sdr0.cic1.comb1_in_del[4] ),
    .B(net107));
 sg13g2_a21oi_1 _12502_ (.A1(_04279_),
    .A2(_04280_),
    .Y(_00440_),
    .B1(net108));
 sg13g2_nand2_1 _12503_ (.Y(_04281_),
    .A(_02348_),
    .B(net231));
 sg13g2_nand2_1 _12504_ (.Y(_04282_),
    .A(_04030_),
    .B(net107));
 sg13g2_a21oi_1 _12505_ (.A1(_04281_),
    .A2(_04282_),
    .Y(_00441_),
    .B1(net108));
 sg13g2_nand2_1 _12506_ (.Y(_04283_),
    .A(_02351_),
    .B(net231));
 sg13g2_nand2_1 _12507_ (.Y(_04284_),
    .A(_04042_),
    .B(net107));
 sg13g2_a21oi_1 _12508_ (.A1(_04283_),
    .A2(_04284_),
    .Y(_00442_),
    .B1(net108));
 sg13g2_nand2_1 _12509_ (.Y(_04285_),
    .A(_02353_),
    .B(net231));
 sg13g2_nand2_1 _12510_ (.Y(_04286_),
    .A(_04035_),
    .B(net107));
 sg13g2_a21oi_1 _12511_ (.A1(_04285_),
    .A2(_04286_),
    .Y(_00443_),
    .B1(net108));
 sg13g2_nand2_1 _12512_ (.Y(_04287_),
    .A(_02355_),
    .B(net231));
 sg13g2_nand2_1 _12513_ (.Y(_04288_),
    .A(_04038_),
    .B(net107));
 sg13g2_a21oi_1 _12514_ (.A1(_04287_),
    .A2(_04288_),
    .Y(_00444_),
    .B1(net108));
 sg13g2_nand2_1 _12515_ (.Y(_04289_),
    .A(_02359_),
    .B(net231));
 sg13g2_nand2_1 _12516_ (.Y(_04290_),
    .A(_04054_),
    .B(_04277_));
 sg13g2_a21oi_1 _12517_ (.A1(_04289_),
    .A2(_04290_),
    .Y(_00445_),
    .B1(net108));
 sg13g2_xnor2_1 _12518_ (.Y(_04291_),
    .A(_04004_),
    .B(\am_sdr0.cic1.comb2_in_del[0] ));
 sg13g2_o21ai_1 _12519_ (.B1(net244),
    .Y(_04292_),
    .A1(\am_sdr0.cic1.comb2[0] ),
    .A2(net236));
 sg13g2_a21oi_1 _12520_ (.A1(net240),
    .A2(_04291_),
    .Y(_00446_),
    .B1(_04292_));
 sg13g2_buf_1 _12521_ (.A(\am_sdr0.cic1.comb2[10] ),
    .X(_04293_));
 sg13g2_buf_1 _12522_ (.A(\am_sdr0.cic1.comb2_in_del[7] ),
    .X(_04294_));
 sg13g2_inv_1 _12523_ (.Y(_04295_),
    .A(_04294_));
 sg13g2_inv_1 _12524_ (.Y(_04296_),
    .A(\am_sdr0.cic1.comb2_in_del[8] ));
 sg13g2_buf_1 _12525_ (.A(\am_sdr0.cic1.comb2_in_del[9] ),
    .X(_04297_));
 sg13g2_nor2b_1 _12526_ (.A(_04297_),
    .B_N(_04238_),
    .Y(_04298_));
 sg13g2_nor3_1 _12527_ (.A(_04295_),
    .B(_04296_),
    .C(_04298_),
    .Y(_04299_));
 sg13g2_nor3_1 _12528_ (.A(_04221_),
    .B(_04296_),
    .C(_04298_),
    .Y(_04300_));
 sg13g2_buf_1 _12529_ (.A(\am_sdr0.cic1.comb2_in_del[6] ),
    .X(_04301_));
 sg13g2_inv_1 _12530_ (.Y(_04302_),
    .A(_04301_));
 sg13g2_nor2_1 _12531_ (.A(_04211_),
    .B(_04302_),
    .Y(_04303_));
 sg13g2_buf_1 _12532_ (.A(\am_sdr0.cic1.comb2_in_del[4] ),
    .X(_04304_));
 sg13g2_nand2b_1 _12533_ (.Y(_04305_),
    .B(_04304_),
    .A_N(_04199_));
 sg13g2_inv_1 _12534_ (.Y(_04306_),
    .A(_04192_));
 sg13g2_inv_1 _12535_ (.Y(_04307_),
    .A(\am_sdr0.cic1.comb2_in_del[3] ));
 sg13g2_inv_1 _12536_ (.Y(_04308_),
    .A(_04185_));
 sg13g2_buf_1 _12537_ (.A(\am_sdr0.cic1.comb2_in_del[2] ),
    .X(_04309_));
 sg13g2_nor2_1 _12538_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sg13g2_nor2b_1 _12539_ (.A(_04004_),
    .B_N(\am_sdr0.cic1.comb2_in_del[0] ),
    .Y(_04311_));
 sg13g2_buf_1 _12540_ (.A(\am_sdr0.cic1.comb2_in_del[1] ),
    .X(_04312_));
 sg13g2_nand2b_1 _12541_ (.Y(_04313_),
    .B(_04180_),
    .A_N(_04312_));
 sg13g2_nor2b_1 _12542_ (.A(_04180_),
    .B_N(_04312_),
    .Y(_04314_));
 sg13g2_a221oi_1 _12543_ (.B2(_04313_),
    .C1(_04314_),
    .B1(_04311_),
    .A1(_04308_),
    .Y(_04315_),
    .A2(_04309_));
 sg13g2_buf_1 _12544_ (.A(_04315_),
    .X(_04316_));
 sg13g2_nor3_1 _12545_ (.A(_04307_),
    .B(_04310_),
    .C(_04316_),
    .Y(_04317_));
 sg13g2_o21ai_1 _12546_ (.B1(_04307_),
    .Y(_04318_),
    .A1(_04310_),
    .A2(_04316_));
 sg13g2_o21ai_1 _12547_ (.B1(_04318_),
    .Y(_04319_),
    .A1(_04306_),
    .A2(_04317_));
 sg13g2_buf_2 _12548_ (.A(_04319_),
    .X(_04320_));
 sg13g2_buf_2 _12549_ (.A(\am_sdr0.cic1.comb2_in_del[5] ),
    .X(_04321_));
 sg13g2_nand2_1 _12550_ (.Y(_04322_),
    .A(_04321_),
    .B(_04301_));
 sg13g2_nand2b_1 _12551_ (.Y(_04323_),
    .B(_04301_),
    .A_N(_04204_));
 sg13g2_nor2b_1 _12552_ (.A(_04304_),
    .B_N(_04199_),
    .Y(_04324_));
 sg13g2_a221oi_1 _12553_ (.B2(_04323_),
    .C1(_04324_),
    .B1(_04322_),
    .A1(_04305_),
    .Y(_04325_),
    .A2(_04320_));
 sg13g2_nand2b_1 _12554_ (.Y(_04326_),
    .B(_04321_),
    .A_N(_04211_));
 sg13g2_or2_1 _12555_ (.X(_04327_),
    .B(_04211_),
    .A(_04204_));
 sg13g2_a221oi_1 _12556_ (.B2(_04327_),
    .C1(_04324_),
    .B1(_04326_),
    .A1(_04305_),
    .Y(_04328_),
    .A2(_04320_));
 sg13g2_nand2b_1 _12557_ (.Y(_04329_),
    .B(_04321_),
    .A_N(_04204_));
 sg13g2_a21oi_1 _12558_ (.A1(_04211_),
    .A2(_04302_),
    .Y(_04330_),
    .B1(_04329_));
 sg13g2_or4_1 _12559_ (.A(_04303_),
    .B(_04325_),
    .C(_04328_),
    .D(_04330_),
    .X(_04331_));
 sg13g2_buf_2 _12560_ (.A(_04331_),
    .X(_04332_));
 sg13g2_o21ai_1 _12561_ (.B1(_04332_),
    .Y(_04333_),
    .A1(_04299_),
    .A2(_04300_));
 sg13g2_nor3_1 _12562_ (.A(_04295_),
    .B(_04230_),
    .C(_04298_),
    .Y(_04334_));
 sg13g2_nor3_1 _12563_ (.A(_04221_),
    .B(_04230_),
    .C(_04298_),
    .Y(_04335_));
 sg13g2_o21ai_1 _12564_ (.B1(_04332_),
    .Y(_04336_),
    .A1(_04334_),
    .A2(_04335_));
 sg13g2_nand2b_1 _12565_ (.Y(_04337_),
    .B(_04238_),
    .A_N(_04297_));
 sg13g2_nor2_1 _12566_ (.A(_04230_),
    .B(_04296_),
    .Y(_04338_));
 sg13g2_nand3b_1 _12567_ (.B(_04294_),
    .C(_04337_),
    .Y(_04339_),
    .A_N(_04221_));
 sg13g2_a21oi_1 _12568_ (.A1(_04230_),
    .A2(_04296_),
    .Y(_04340_),
    .B1(_04339_));
 sg13g2_a21oi_1 _12569_ (.A1(_04337_),
    .A2(_04338_),
    .Y(_04341_),
    .B1(_04340_));
 sg13g2_nand2b_1 _12570_ (.Y(_04342_),
    .B(_04297_),
    .A_N(_04238_));
 sg13g2_buf_1 _12571_ (.A(_04342_),
    .X(_04343_));
 sg13g2_nand4_1 _12572_ (.B(_04336_),
    .C(_04341_),
    .A(_04333_),
    .Y(_04344_),
    .D(_04343_));
 sg13g2_buf_1 _12573_ (.A(_04344_),
    .X(_04345_));
 sg13g2_buf_1 _12574_ (.A(\am_sdr0.cic1.comb2_in_del[10] ),
    .X(_04346_));
 sg13g2_xor2_1 _12575_ (.B(_04346_),
    .A(_04008_),
    .X(_04347_));
 sg13g2_xnor2_1 _12576_ (.Y(_04348_),
    .A(_04345_),
    .B(_04347_));
 sg13g2_nand2_1 _12577_ (.Y(_04349_),
    .A(_04113_),
    .B(_04348_));
 sg13g2_o21ai_1 _12578_ (.B1(_04349_),
    .Y(_04350_),
    .A1(_04293_),
    .A2(net237));
 sg13g2_nor2_1 _12579_ (.A(net111),
    .B(_04350_),
    .Y(_00447_));
 sg13g2_buf_1 _12580_ (.A(\am_sdr0.cic1.comb2[11] ),
    .X(_04351_));
 sg13g2_nand2_1 _12581_ (.Y(_04352_),
    .A(_04351_),
    .B(net113));
 sg13g2_inv_1 _12582_ (.Y(_04353_),
    .A(_04346_));
 sg13g2_nand2b_1 _12583_ (.Y(_04354_),
    .B(_04353_),
    .A_N(_04345_));
 sg13g2_inv_1 _12584_ (.Y(_04355_),
    .A(_04008_));
 sg13g2_a21o_1 _12585_ (.A2(_04345_),
    .A1(_04346_),
    .B1(_04355_),
    .X(_04356_));
 sg13g2_buf_1 _12586_ (.A(_04356_),
    .X(_04357_));
 sg13g2_nand2_1 _12587_ (.Y(_04358_),
    .A(_04354_),
    .B(_04357_));
 sg13g2_buf_1 _12588_ (.A(\am_sdr0.cic1.comb2_in_del[11] ),
    .X(_04359_));
 sg13g2_xor2_1 _12589_ (.B(_04359_),
    .A(_04065_),
    .X(_04360_));
 sg13g2_xnor2_1 _12590_ (.Y(_04361_),
    .A(_04358_),
    .B(_04360_));
 sg13g2_nand2_1 _12591_ (.Y(_04362_),
    .A(net234),
    .B(_04361_));
 sg13g2_buf_1 _12592_ (.A(_03428_),
    .X(_04363_));
 sg13g2_a21oi_1 _12593_ (.A1(_04352_),
    .A2(_04362_),
    .Y(_00448_),
    .B1(_04363_));
 sg13g2_buf_1 _12594_ (.A(\am_sdr0.cic1.comb2[12] ),
    .X(_04364_));
 sg13g2_nand2_1 _12595_ (.Y(_04365_),
    .A(_04364_),
    .B(net113));
 sg13g2_nand3_1 _12596_ (.B(_04354_),
    .C(_04357_),
    .A(_04359_),
    .Y(_04366_));
 sg13g2_a21oi_1 _12597_ (.A1(_04354_),
    .A2(_04357_),
    .Y(_04367_),
    .B1(_04359_));
 sg13g2_a21oi_2 _12598_ (.B1(_04367_),
    .Y(_04368_),
    .A2(_04366_),
    .A1(_04065_));
 sg13g2_inv_1 _12599_ (.Y(_04369_),
    .A(\am_sdr0.cic1.comb1[12] ));
 sg13g2_buf_1 _12600_ (.A(\am_sdr0.cic1.comb2_in_del[12] ),
    .X(_04370_));
 sg13g2_nor2_1 _12601_ (.A(_04369_),
    .B(_04370_),
    .Y(_04371_));
 sg13g2_nand2_1 _12602_ (.Y(_04372_),
    .A(_04369_),
    .B(_04370_));
 sg13g2_nand2b_1 _12603_ (.Y(_04373_),
    .B(_04372_),
    .A_N(_04371_));
 sg13g2_xor2_1 _12604_ (.B(_04373_),
    .A(_04368_),
    .X(_04374_));
 sg13g2_nand2_1 _12605_ (.Y(_04375_),
    .A(net234),
    .B(_04374_));
 sg13g2_a21oi_1 _12606_ (.A1(_04365_),
    .A2(_04375_),
    .Y(_00449_),
    .B1(net106));
 sg13g2_and2_1 _12607_ (.A(_04370_),
    .B(_04368_),
    .X(_04376_));
 sg13g2_buf_1 _12608_ (.A(_04376_),
    .X(_04377_));
 sg13g2_o21ai_1 _12609_ (.B1(_04369_),
    .Y(_04378_),
    .A1(_04370_),
    .A2(_04368_));
 sg13g2_nand2b_1 _12610_ (.Y(_04379_),
    .B(_04378_),
    .A_N(_04377_));
 sg13g2_buf_1 _12611_ (.A(\am_sdr0.cic1.comb2_in_del[13] ),
    .X(_04380_));
 sg13g2_xor2_1 _12612_ (.B(_04380_),
    .A(_04104_),
    .X(_04381_));
 sg13g2_xnor2_1 _12613_ (.Y(_04382_),
    .A(_04379_),
    .B(_04381_));
 sg13g2_buf_1 _12614_ (.A(\am_sdr0.cic1.comb2[13] ),
    .X(_04383_));
 sg13g2_o21ai_1 _12615_ (.B1(_03002_),
    .Y(_04384_),
    .A1(_04383_),
    .A2(net236));
 sg13g2_a21oi_1 _12616_ (.A1(net240),
    .A2(_04382_),
    .Y(_00450_),
    .B1(_04384_));
 sg13g2_nand2b_1 _12617_ (.Y(_04385_),
    .B(_04104_),
    .A_N(_04380_));
 sg13g2_nor2_1 _12618_ (.A(_04380_),
    .B(_04377_),
    .Y(_04386_));
 sg13g2_nor2b_1 _12619_ (.A(_04377_),
    .B_N(_04104_),
    .Y(_04387_));
 sg13g2_o21ai_1 _12620_ (.B1(_04378_),
    .Y(_04388_),
    .A1(_04386_),
    .A2(_04387_));
 sg13g2_nand2_1 _12621_ (.Y(_04389_),
    .A(net364),
    .B(_04000_));
 sg13g2_inv_1 _12622_ (.Y(_00611_),
    .A(_04389_));
 sg13g2_buf_1 _12623_ (.A(\am_sdr0.cic1.comb2_in_del[14] ),
    .X(_04390_));
 sg13g2_xor2_1 _12624_ (.B(_04390_),
    .A(_04112_),
    .X(_04391_));
 sg13g2_nand2_1 _12625_ (.Y(_04392_),
    .A(_00611_),
    .B(_04391_));
 sg13g2_a21o_1 _12626_ (.A2(_04388_),
    .A1(_04385_),
    .B1(_04392_),
    .X(_04393_));
 sg13g2_nor2_1 _12627_ (.A(_04389_),
    .B(_04391_),
    .Y(_04394_));
 sg13g2_nand3_1 _12628_ (.B(_04388_),
    .C(_04394_),
    .A(_04385_),
    .Y(_04395_));
 sg13g2_buf_1 _12629_ (.A(\am_sdr0.cic1.comb2[14] ),
    .X(_04396_));
 sg13g2_nand3_1 _12630_ (.B(_04396_),
    .C(net162),
    .A(net253),
    .Y(_04397_));
 sg13g2_nand3_1 _12631_ (.B(_04395_),
    .C(_04397_),
    .A(_04393_),
    .Y(_00451_));
 sg13g2_buf_2 _12632_ (.A(\am_sdr0.cic1.comb2[15] ),
    .X(_04398_));
 sg13g2_nand2_1 _12633_ (.Y(_04399_),
    .A(_04398_),
    .B(_04012_));
 sg13g2_nor4_2 _12634_ (.A(_04360_),
    .B(_04373_),
    .C(_04381_),
    .Y(_04400_),
    .D(_04391_));
 sg13g2_and3_1 _12635_ (.X(_04401_),
    .A(_04353_),
    .B(_04343_),
    .C(_04400_));
 sg13g2_nand4_1 _12636_ (.B(_04336_),
    .C(_04341_),
    .A(_04333_),
    .Y(_04402_),
    .D(_04401_));
 sg13g2_and3_1 _12637_ (.X(_04403_),
    .A(_04008_),
    .B(_04343_),
    .C(_04400_));
 sg13g2_nand4_1 _12638_ (.B(_04336_),
    .C(_04341_),
    .A(_04333_),
    .Y(_04404_),
    .D(_04403_));
 sg13g2_inv_1 _12639_ (.Y(_04405_),
    .A(_04390_));
 sg13g2_nor2_1 _12640_ (.A(_04355_),
    .B(_04346_),
    .Y(_04406_));
 sg13g2_inv_1 _12641_ (.Y(_04407_),
    .A(_04112_));
 sg13g2_nor2b_1 _12642_ (.A(_04359_),
    .B_N(_04065_),
    .Y(_04408_));
 sg13g2_a21oi_1 _12643_ (.A1(_04408_),
    .A2(_04372_),
    .Y(_04409_),
    .B1(_04371_));
 sg13g2_nor2_1 _12644_ (.A(_04380_),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_nor2_1 _12645_ (.A(_04104_),
    .B(_04410_),
    .Y(_04411_));
 sg13g2_a221oi_1 _12646_ (.B2(_04380_),
    .C1(_04411_),
    .B1(_04409_),
    .A1(_04407_),
    .Y(_04412_),
    .A2(_04390_));
 sg13g2_a221oi_1 _12647_ (.B2(_04400_),
    .C1(_04412_),
    .B1(_04406_),
    .A1(_04112_),
    .Y(_04413_),
    .A2(_04405_));
 sg13g2_nand3_1 _12648_ (.B(_04404_),
    .C(_04413_),
    .A(_04402_),
    .Y(_04414_));
 sg13g2_buf_1 _12649_ (.A(_04414_),
    .X(_04415_));
 sg13g2_buf_1 _12650_ (.A(\am_sdr0.cic1.comb2_in_del[15] ),
    .X(_04416_));
 sg13g2_xor2_1 _12651_ (.B(_04416_),
    .A(_04133_),
    .X(_04417_));
 sg13g2_xnor2_1 _12652_ (.Y(_04418_),
    .A(_04415_),
    .B(_04417_));
 sg13g2_nand2_1 _12653_ (.Y(_04419_),
    .A(_04143_),
    .B(_04418_));
 sg13g2_a21oi_1 _12654_ (.A1(_04399_),
    .A2(_04419_),
    .Y(_00452_),
    .B1(_04363_));
 sg13g2_buf_1 _12655_ (.A(\am_sdr0.cic1.comb2[16] ),
    .X(_04420_));
 sg13g2_inv_1 _12656_ (.Y(_04421_),
    .A(_04420_));
 sg13g2_inv_1 _12657_ (.Y(_04422_),
    .A(_04416_));
 sg13g2_nor2_1 _12658_ (.A(_04422_),
    .B(_04415_),
    .Y(_04423_));
 sg13g2_a21oi_1 _12659_ (.A1(_04422_),
    .A2(_04415_),
    .Y(_04424_),
    .B1(_04133_));
 sg13g2_or2_1 _12660_ (.X(_04425_),
    .B(_04424_),
    .A(_04423_));
 sg13g2_xor2_1 _12661_ (.B(\am_sdr0.cic1.comb2_in_del[16] ),
    .A(_04141_),
    .X(_04426_));
 sg13g2_xnor2_1 _12662_ (.Y(_04427_),
    .A(_04425_),
    .B(_04426_));
 sg13g2_mux2_1 _12663_ (.A0(_04421_),
    .A1(_04427_),
    .S(net236),
    .X(_04428_));
 sg13g2_nor2_1 _12664_ (.A(_04220_),
    .B(_04428_),
    .Y(_00453_));
 sg13g2_buf_1 _12665_ (.A(\am_sdr0.cic1.comb2[17] ),
    .X(_04429_));
 sg13g2_inv_1 _12666_ (.Y(_04430_),
    .A(\am_sdr0.cic1.comb2_in_del[16] ));
 sg13g2_a221oi_1 _12667_ (.B2(_04430_),
    .C1(_04415_),
    .B1(_04141_),
    .A1(_04133_),
    .Y(_04431_),
    .A2(_04422_));
 sg13g2_buf_1 _12668_ (.A(_04431_),
    .X(_04432_));
 sg13g2_nand2b_1 _12669_ (.Y(_04433_),
    .B(_04416_),
    .A_N(_04133_));
 sg13g2_a21o_1 _12670_ (.A2(_04430_),
    .A1(_04141_),
    .B1(_04433_),
    .X(_04434_));
 sg13g2_o21ai_1 _12671_ (.B1(_04434_),
    .Y(_04435_),
    .A1(_04141_),
    .A2(_04430_));
 sg13g2_nor2_1 _12672_ (.A(_04432_),
    .B(_04435_),
    .Y(_04436_));
 sg13g2_buf_1 _12673_ (.A(\am_sdr0.cic1.comb2_in_del[17] ),
    .X(_04437_));
 sg13g2_xnor2_1 _12674_ (.Y(_04438_),
    .A(_04154_),
    .B(_04437_));
 sg13g2_xnor2_1 _12675_ (.Y(_04439_),
    .A(_04436_),
    .B(_04438_));
 sg13g2_nor2_1 _12676_ (.A(net162),
    .B(_04439_),
    .Y(_04440_));
 sg13g2_a21oi_1 _12677_ (.A1(_04429_),
    .A2(net112),
    .Y(_04441_),
    .B1(_04440_));
 sg13g2_nor2_1 _12678_ (.A(_04220_),
    .B(_04441_),
    .Y(_00454_));
 sg13g2_buf_1 _12679_ (.A(\am_sdr0.cic1.comb2[18] ),
    .X(_04442_));
 sg13g2_nor2_1 _12680_ (.A(_04442_),
    .B(_04006_),
    .Y(_04443_));
 sg13g2_nor3_1 _12681_ (.A(_04437_),
    .B(_04432_),
    .C(_04435_),
    .Y(_04444_));
 sg13g2_o21ai_1 _12682_ (.B1(_04437_),
    .Y(_04445_),
    .A1(_04432_),
    .A2(_04435_));
 sg13g2_o21ai_1 _12683_ (.B1(_04445_),
    .Y(_04446_),
    .A1(_04154_),
    .A2(_04444_));
 sg13g2_buf_1 _12684_ (.A(_04446_),
    .X(_04447_));
 sg13g2_buf_1 _12685_ (.A(\am_sdr0.cic1.comb2_in_del[18] ),
    .X(_04448_));
 sg13g2_xnor2_1 _12686_ (.Y(_04449_),
    .A(_04172_),
    .B(_04448_));
 sg13g2_xnor2_1 _12687_ (.Y(_04450_),
    .A(_04447_),
    .B(_04449_));
 sg13g2_nor2_1 _12688_ (.A(net161),
    .B(_04450_),
    .Y(_04451_));
 sg13g2_nor3_1 _12689_ (.A(net160),
    .B(_04443_),
    .C(_04451_),
    .Y(_00455_));
 sg13g2_xor2_1 _12690_ (.B(\am_sdr0.cic1.comb2_in_del[19] ),
    .A(\am_sdr0.cic1.comb1[19] ),
    .X(_04452_));
 sg13g2_nand2_1 _12691_ (.Y(_04453_),
    .A(_04448_),
    .B(_04447_));
 sg13g2_nor2_1 _12692_ (.A(_04448_),
    .B(_04447_),
    .Y(_04454_));
 sg13g2_a21oi_1 _12693_ (.A1(_04172_),
    .A2(_04453_),
    .Y(_04455_),
    .B1(_04454_));
 sg13g2_xnor2_1 _12694_ (.Y(_04456_),
    .A(_04452_),
    .B(_04455_));
 sg13g2_nand3_1 _12695_ (.B(\am_sdr0.cic1.comb2[19] ),
    .C(net112),
    .A(net254),
    .Y(_04457_));
 sg13g2_o21ai_1 _12696_ (.B1(_04457_),
    .Y(_00456_),
    .A1(_04389_),
    .A2(_04456_));
 sg13g2_nand2_1 _12697_ (.Y(_04458_),
    .A(\am_sdr0.cic1.comb2[1] ),
    .B(net112));
 sg13g2_xnor2_1 _12698_ (.Y(_04459_),
    .A(_04180_),
    .B(_04312_));
 sg13g2_xnor2_1 _12699_ (.Y(_04460_),
    .A(_04311_),
    .B(_04459_));
 sg13g2_nand2_1 _12700_ (.Y(_04461_),
    .A(net234),
    .B(_04460_));
 sg13g2_a21oi_1 _12701_ (.A1(_04458_),
    .A2(_04461_),
    .Y(_00457_),
    .B1(net106));
 sg13g2_buf_1 _12702_ (.A(\am_sdr0.cic1.comb2[2] ),
    .X(_04462_));
 sg13g2_nand2_1 _12703_ (.Y(_04463_),
    .A(_04462_),
    .B(net112));
 sg13g2_a21oi_1 _12704_ (.A1(_04311_),
    .A2(_04313_),
    .Y(_04464_),
    .B1(_04314_));
 sg13g2_xor2_1 _12705_ (.B(_04309_),
    .A(_04185_),
    .X(_04465_));
 sg13g2_xnor2_1 _12706_ (.Y(_04466_),
    .A(_04464_),
    .B(_04465_));
 sg13g2_nand2_1 _12707_ (.Y(_04467_),
    .A(net234),
    .B(_04466_));
 sg13g2_a21oi_1 _12708_ (.A1(_04463_),
    .A2(_04467_),
    .Y(_00458_),
    .B1(net106));
 sg13g2_nand2_1 _12709_ (.Y(_04468_),
    .A(\am_sdr0.cic1.comb2[3] ),
    .B(_04186_));
 sg13g2_nor2_1 _12710_ (.A(_04310_),
    .B(_04316_),
    .Y(_04469_));
 sg13g2_xnor2_1 _12711_ (.Y(_04470_),
    .A(_04192_),
    .B(\am_sdr0.cic1.comb2_in_del[3] ));
 sg13g2_xnor2_1 _12712_ (.Y(_04471_),
    .A(_04469_),
    .B(_04470_));
 sg13g2_nand2_1 _12713_ (.Y(_04472_),
    .A(net234),
    .B(_04471_));
 sg13g2_a21oi_1 _12714_ (.A1(_04468_),
    .A2(_04472_),
    .Y(_00459_),
    .B1(net106));
 sg13g2_buf_1 _12715_ (.A(\am_sdr0.cic1.comb2[4] ),
    .X(_04473_));
 sg13g2_nor2_1 _12716_ (.A(_04473_),
    .B(net239),
    .Y(_04474_));
 sg13g2_xor2_1 _12717_ (.B(_04304_),
    .A(_04199_),
    .X(_04475_));
 sg13g2_xnor2_1 _12718_ (.Y(_04476_),
    .A(_04320_),
    .B(_04475_));
 sg13g2_nor2_1 _12719_ (.A(net161),
    .B(_04476_),
    .Y(_04477_));
 sg13g2_nor3_1 _12720_ (.A(net160),
    .B(_04474_),
    .C(_04477_),
    .Y(_00460_));
 sg13g2_buf_1 _12721_ (.A(\am_sdr0.cic1.comb2[5] ),
    .X(_04478_));
 sg13g2_a21oi_2 _12722_ (.B1(_04324_),
    .Y(_04479_),
    .A2(_04320_),
    .A1(_04305_));
 sg13g2_xor2_1 _12723_ (.B(_04321_),
    .A(_04204_),
    .X(_04480_));
 sg13g2_xnor2_1 _12724_ (.Y(_04481_),
    .A(_04479_),
    .B(_04480_));
 sg13g2_nand2_1 _12725_ (.Y(_04482_),
    .A(net235),
    .B(_04481_));
 sg13g2_o21ai_1 _12726_ (.B1(_04482_),
    .Y(_04483_),
    .A1(_04478_),
    .A2(net239));
 sg13g2_nor2_1 _12727_ (.A(net111),
    .B(_04483_),
    .Y(_00461_));
 sg13g2_nand2_1 _12728_ (.Y(_04484_),
    .A(_04321_),
    .B(_04479_));
 sg13g2_nor2_1 _12729_ (.A(_04321_),
    .B(_04479_),
    .Y(_04485_));
 sg13g2_a21oi_1 _12730_ (.A1(_04204_),
    .A2(_04484_),
    .Y(_04486_),
    .B1(_04485_));
 sg13g2_xnor2_1 _12731_ (.Y(_04487_),
    .A(_04211_),
    .B(_04301_));
 sg13g2_xnor2_1 _12732_ (.Y(_04488_),
    .A(_04486_),
    .B(_04487_));
 sg13g2_buf_1 _12733_ (.A(\am_sdr0.cic1.comb2[6] ),
    .X(_04489_));
 sg13g2_nor2b_1 _12734_ (.A(net235),
    .B_N(_04489_),
    .Y(_04490_));
 sg13g2_a21oi_1 _12735_ (.A1(net233),
    .A2(_04488_),
    .Y(_04491_),
    .B1(_04490_));
 sg13g2_nor2_1 _12736_ (.A(net111),
    .B(_04491_),
    .Y(_00462_));
 sg13g2_xnor2_1 _12737_ (.Y(_04492_),
    .A(_04221_),
    .B(_04294_));
 sg13g2_xnor2_1 _12738_ (.Y(_04493_),
    .A(_04332_),
    .B(_04492_));
 sg13g2_buf_1 _12739_ (.A(\am_sdr0.cic1.comb2[7] ),
    .X(_04494_));
 sg13g2_nor2b_1 _12740_ (.A(net235),
    .B_N(_04494_),
    .Y(_04495_));
 sg13g2_a21oi_1 _12741_ (.A1(net233),
    .A2(_04493_),
    .Y(_04496_),
    .B1(_04495_));
 sg13g2_nor2_1 _12742_ (.A(net111),
    .B(_04496_),
    .Y(_00463_));
 sg13g2_nand2_1 _12743_ (.Y(_04497_),
    .A(_04294_),
    .B(_04332_));
 sg13g2_nor2_1 _12744_ (.A(_04294_),
    .B(_04332_),
    .Y(_04498_));
 sg13g2_a21oi_1 _12745_ (.A1(_04221_),
    .A2(_04497_),
    .Y(_04499_),
    .B1(_04498_));
 sg13g2_nand2_1 _12746_ (.Y(_04500_),
    .A(_04230_),
    .B(_04296_));
 sg13g2_nand2b_1 _12747_ (.Y(_04501_),
    .B(_04500_),
    .A_N(_04338_));
 sg13g2_xnor2_1 _12748_ (.Y(_04502_),
    .A(_04499_),
    .B(_04501_));
 sg13g2_nand2_1 _12749_ (.Y(_04503_),
    .A(net235),
    .B(_04502_));
 sg13g2_o21ai_1 _12750_ (.B1(_04503_),
    .Y(_04504_),
    .A1(\am_sdr0.cic1.comb2[8] ),
    .A2(net239));
 sg13g2_nor2_1 _12751_ (.A(net111),
    .B(_04504_),
    .Y(_00464_));
 sg13g2_buf_1 _12752_ (.A(\am_sdr0.cic1.comb2[9] ),
    .X(_04505_));
 sg13g2_nand2_1 _12753_ (.Y(_04506_),
    .A(_04505_),
    .B(_04186_));
 sg13g2_a21oi_1 _12754_ (.A1(_04499_),
    .A2(_04500_),
    .Y(_04507_),
    .B1(_04338_));
 sg13g2_nand2_1 _12755_ (.Y(_04508_),
    .A(_04337_),
    .B(_04343_));
 sg13g2_xnor2_1 _12756_ (.Y(_04509_),
    .A(_04507_),
    .B(_04508_));
 sg13g2_nand2_1 _12757_ (.Y(_04510_),
    .A(net237),
    .B(_04509_));
 sg13g2_a21oi_1 _12758_ (.A1(_04506_),
    .A2(_04510_),
    .Y(_00465_),
    .B1(net106));
 sg13g2_nand2_1 _12759_ (.Y(_04511_),
    .A(_04004_),
    .B(net231));
 sg13g2_nand2_1 _12760_ (.Y(_04512_),
    .A(\am_sdr0.cic1.comb2_in_del[0] ),
    .B(_04277_));
 sg13g2_a21oi_1 _12761_ (.A1(_04511_),
    .A2(_04512_),
    .Y(_00466_),
    .B1(net106));
 sg13g2_buf_1 _12762_ (.A(net291),
    .X(_04513_));
 sg13g2_nand2_1 _12763_ (.Y(_04514_),
    .A(_04008_),
    .B(net230));
 sg13g2_nand2_1 _12764_ (.Y(_04515_),
    .A(_04346_),
    .B(net107));
 sg13g2_a21oi_1 _12765_ (.A1(_04514_),
    .A2(_04515_),
    .Y(_00467_),
    .B1(net106));
 sg13g2_nand2_1 _12766_ (.Y(_04516_),
    .A(_04065_),
    .B(net230));
 sg13g2_nand2_1 _12767_ (.Y(_04517_),
    .A(_04359_),
    .B(net107));
 sg13g2_a21oi_1 _12768_ (.A1(_04516_),
    .A2(_04517_),
    .Y(_00468_),
    .B1(net106));
 sg13g2_nand2_1 _12769_ (.Y(_04518_),
    .A(\am_sdr0.cic1.comb1[12] ),
    .B(net230));
 sg13g2_buf_1 _12770_ (.A(_04010_),
    .X(_04519_));
 sg13g2_nand2_1 _12771_ (.Y(_04520_),
    .A(_04370_),
    .B(net159));
 sg13g2_buf_1 _12772_ (.A(_03428_),
    .X(_04521_));
 sg13g2_a21oi_1 _12773_ (.A1(_04518_),
    .A2(_04520_),
    .Y(_00469_),
    .B1(net105));
 sg13g2_nand2_1 _12774_ (.Y(_04522_),
    .A(_04104_),
    .B(net230));
 sg13g2_nand2_1 _12775_ (.Y(_04523_),
    .A(_04380_),
    .B(net159));
 sg13g2_a21oi_1 _12776_ (.A1(_04522_),
    .A2(_04523_),
    .Y(_00470_),
    .B1(net105));
 sg13g2_nand2_1 _12777_ (.Y(_04524_),
    .A(_04112_),
    .B(net230));
 sg13g2_nand2_1 _12778_ (.Y(_04525_),
    .A(_04390_),
    .B(net159));
 sg13g2_a21oi_1 _12779_ (.A1(_04524_),
    .A2(_04525_),
    .Y(_00471_),
    .B1(net105));
 sg13g2_nand2_1 _12780_ (.Y(_04526_),
    .A(_04133_),
    .B(net230));
 sg13g2_nand2_1 _12781_ (.Y(_04527_),
    .A(_04416_),
    .B(net159));
 sg13g2_a21oi_1 _12782_ (.A1(_04526_),
    .A2(_04527_),
    .Y(_00472_),
    .B1(net105));
 sg13g2_nand2_1 _12783_ (.Y(_04528_),
    .A(_04141_),
    .B(net230));
 sg13g2_nand2_1 _12784_ (.Y(_04529_),
    .A(\am_sdr0.cic1.comb2_in_del[16] ),
    .B(net159));
 sg13g2_a21oi_1 _12785_ (.A1(_04528_),
    .A2(_04529_),
    .Y(_00473_),
    .B1(net105));
 sg13g2_nand2_1 _12786_ (.Y(_04530_),
    .A(_04154_),
    .B(net230));
 sg13g2_nand2_1 _12787_ (.Y(_04531_),
    .A(_04437_),
    .B(net159));
 sg13g2_a21oi_1 _12788_ (.A1(_04530_),
    .A2(_04531_),
    .Y(_00474_),
    .B1(net105));
 sg13g2_nand2_1 _12789_ (.Y(_04532_),
    .A(_04172_),
    .B(_04513_));
 sg13g2_nand2_1 _12790_ (.Y(_04533_),
    .A(_04448_),
    .B(_04519_));
 sg13g2_a21oi_1 _12791_ (.A1(_04532_),
    .A2(_04533_),
    .Y(_00475_),
    .B1(_04521_));
 sg13g2_nand2_1 _12792_ (.Y(_04534_),
    .A(\am_sdr0.cic1.comb1[19] ),
    .B(_04513_));
 sg13g2_nand2_1 _12793_ (.Y(_04535_),
    .A(\am_sdr0.cic1.comb2_in_del[19] ),
    .B(_04519_));
 sg13g2_a21oi_1 _12794_ (.A1(_04534_),
    .A2(_04535_),
    .Y(_00476_),
    .B1(_04521_));
 sg13g2_buf_1 _12795_ (.A(net291),
    .X(_04536_));
 sg13g2_nand2_1 _12796_ (.Y(_04537_),
    .A(_04180_),
    .B(_04536_));
 sg13g2_nand2_1 _12797_ (.Y(_04538_),
    .A(_04312_),
    .B(net159));
 sg13g2_a21oi_1 _12798_ (.A1(_04537_),
    .A2(_04538_),
    .Y(_00477_),
    .B1(net105));
 sg13g2_nand2_1 _12799_ (.Y(_04539_),
    .A(_04185_),
    .B(_04536_));
 sg13g2_nand2_1 _12800_ (.Y(_04540_),
    .A(_04309_),
    .B(net159));
 sg13g2_a21oi_1 _12801_ (.A1(_04539_),
    .A2(_04540_),
    .Y(_00478_),
    .B1(net105));
 sg13g2_nand2_1 _12802_ (.Y(_04541_),
    .A(_04192_),
    .B(net229));
 sg13g2_buf_1 _12803_ (.A(_04010_),
    .X(_04542_));
 sg13g2_nand2_1 _12804_ (.Y(_04543_),
    .A(\am_sdr0.cic1.comb2_in_del[3] ),
    .B(_04542_));
 sg13g2_buf_1 _12805_ (.A(_03428_),
    .X(_04544_));
 sg13g2_a21oi_1 _12806_ (.A1(_04541_),
    .A2(_04543_),
    .Y(_00479_),
    .B1(_04544_));
 sg13g2_nand2_1 _12807_ (.Y(_04545_),
    .A(_04199_),
    .B(net229));
 sg13g2_nand2_1 _12808_ (.Y(_04546_),
    .A(_04304_),
    .B(net158));
 sg13g2_a21oi_1 _12809_ (.A1(_04545_),
    .A2(_04546_),
    .Y(_00480_),
    .B1(net104));
 sg13g2_nand2_1 _12810_ (.Y(_04547_),
    .A(_04204_),
    .B(net229));
 sg13g2_nand2_1 _12811_ (.Y(_04548_),
    .A(_04321_),
    .B(net158));
 sg13g2_a21oi_1 _12812_ (.A1(_04547_),
    .A2(_04548_),
    .Y(_00481_),
    .B1(net104));
 sg13g2_nand2_1 _12813_ (.Y(_04549_),
    .A(_04211_),
    .B(net229));
 sg13g2_nand2_1 _12814_ (.Y(_04550_),
    .A(_04301_),
    .B(net158));
 sg13g2_a21oi_1 _12815_ (.A1(_04549_),
    .A2(_04550_),
    .Y(_00482_),
    .B1(net104));
 sg13g2_nand2_1 _12816_ (.Y(_04551_),
    .A(_04221_),
    .B(net229));
 sg13g2_nand2_1 _12817_ (.Y(_04552_),
    .A(_04294_),
    .B(net158));
 sg13g2_a21oi_1 _12818_ (.A1(_04551_),
    .A2(_04552_),
    .Y(_00483_),
    .B1(net104));
 sg13g2_nand2_1 _12819_ (.Y(_04553_),
    .A(_04230_),
    .B(net229));
 sg13g2_nand2_1 _12820_ (.Y(_04554_),
    .A(\am_sdr0.cic1.comb2_in_del[8] ),
    .B(net158));
 sg13g2_a21oi_1 _12821_ (.A1(_04553_),
    .A2(_04554_),
    .Y(_00484_),
    .B1(net104));
 sg13g2_nand2_1 _12822_ (.Y(_04555_),
    .A(_04238_),
    .B(net229));
 sg13g2_nand2_1 _12823_ (.Y(_04556_),
    .A(_04297_),
    .B(net158));
 sg13g2_a21oi_1 _12824_ (.A1(_04555_),
    .A2(_04556_),
    .Y(_00485_),
    .B1(net104));
 sg13g2_nand2b_1 _12825_ (.Y(_04557_),
    .B(\am_sdr0.cic1.comb3_in_del[6] ),
    .A_N(_04489_));
 sg13g2_nand2_1 _12826_ (.Y(_04558_),
    .A(_04478_),
    .B(_04557_));
 sg13g2_nand2b_1 _12827_ (.Y(_04559_),
    .B(_04557_),
    .A_N(\am_sdr0.cic1.comb3_in_del[5] ));
 sg13g2_inv_1 _12828_ (.Y(_04560_),
    .A(\am_sdr0.cic1.comb2[3] ));
 sg13g2_nand2b_1 _12829_ (.Y(_04561_),
    .B(_04462_),
    .A_N(\am_sdr0.cic1.comb3_in_del[2] ));
 sg13g2_nand2b_1 _12830_ (.Y(_04562_),
    .B(\am_sdr0.cic1.comb3_in_del[2] ),
    .A_N(_04462_));
 sg13g2_inv_1 _12831_ (.Y(_04563_),
    .A(\am_sdr0.cic1.comb2[1] ));
 sg13g2_nor2b_1 _12832_ (.A(\am_sdr0.cic1.comb2[0] ),
    .B_N(\am_sdr0.cic1.comb3_in_del[0] ),
    .Y(_04564_));
 sg13g2_nand2_1 _12833_ (.Y(_04565_),
    .A(_04563_),
    .B(_04564_));
 sg13g2_o21ai_1 _12834_ (.B1(\am_sdr0.cic1.comb3_in_del[1] ),
    .Y(_04566_),
    .A1(_04563_),
    .A2(_04564_));
 sg13g2_nand3_1 _12835_ (.B(_04565_),
    .C(_04566_),
    .A(_04562_),
    .Y(_04567_));
 sg13g2_a22oi_1 _12836_ (.Y(_04568_),
    .B1(_04561_),
    .B2(_04567_),
    .A2(_04560_),
    .A1(\am_sdr0.cic1.comb3_in_del[3] ));
 sg13g2_nand2b_1 _12837_ (.Y(_04569_),
    .B(_04473_),
    .A_N(\am_sdr0.cic1.comb3_in_del[4] ));
 sg13g2_o21ai_1 _12838_ (.B1(_04569_),
    .Y(_04570_),
    .A1(\am_sdr0.cic1.comb3_in_del[3] ),
    .A2(_04560_));
 sg13g2_nand2b_1 _12839_ (.Y(_04571_),
    .B(\am_sdr0.cic1.comb3_in_del[4] ),
    .A_N(_04473_));
 sg13g2_o21ai_1 _12840_ (.B1(_04571_),
    .Y(_04572_),
    .A1(_04568_),
    .A2(_04570_));
 sg13g2_a21o_1 _12841_ (.A2(_04559_),
    .A1(_04558_),
    .B1(_04572_),
    .X(_04573_));
 sg13g2_nor2b_1 _12842_ (.A(\am_sdr0.cic1.comb3_in_del[5] ),
    .B_N(_04478_),
    .Y(_04574_));
 sg13g2_nor2b_1 _12843_ (.A(\am_sdr0.cic1.comb3_in_del[6] ),
    .B_N(_04489_),
    .Y(_04575_));
 sg13g2_a21oi_1 _12844_ (.A1(_04557_),
    .A2(_04574_),
    .Y(_04576_),
    .B1(_04575_));
 sg13g2_inv_1 _12845_ (.Y(_04577_),
    .A(\am_sdr0.cic1.comb2[8] ));
 sg13g2_nand2_1 _12846_ (.Y(_04578_),
    .A(\am_sdr0.cic1.comb3_in_del[8] ),
    .B(_04577_));
 sg13g2_nand2_1 _12847_ (.Y(_04579_),
    .A(_04494_),
    .B(_04578_));
 sg13g2_nand2b_1 _12848_ (.Y(_04580_),
    .B(_04578_),
    .A_N(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_a22oi_1 _12849_ (.Y(_04581_),
    .B1(_04579_),
    .B2(_04580_),
    .A2(_04576_),
    .A1(_04573_));
 sg13g2_nand3b_1 _12850_ (.B(_04494_),
    .C(_04578_),
    .Y(_04582_),
    .A_N(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_o21ai_1 _12851_ (.B1(_04582_),
    .Y(_04583_),
    .A1(\am_sdr0.cic1.comb3_in_del[8] ),
    .A2(_04577_));
 sg13g2_nor2b_1 _12852_ (.A(\am_sdr0.cic1.comb3_in_del[11] ),
    .B_N(_04351_),
    .Y(_04584_));
 sg13g2_nand2b_1 _12853_ (.Y(_04585_),
    .B(\am_sdr0.cic1.comb3_in_del[11] ),
    .A_N(_04351_));
 sg13g2_nand2b_1 _12854_ (.Y(_04586_),
    .B(_04585_),
    .A_N(_04584_));
 sg13g2_xor2_1 _12855_ (.B(_04293_),
    .A(\am_sdr0.cic1.comb3_in_del[10] ),
    .X(_04587_));
 sg13g2_nor2b_1 _12856_ (.A(\am_sdr0.cic1.comb3_in_del[9] ),
    .B_N(_04505_),
    .Y(_04588_));
 sg13g2_nor2b_1 _12857_ (.A(_04505_),
    .B_N(\am_sdr0.cic1.comb3_in_del[9] ),
    .Y(_04589_));
 sg13g2_or3_1 _12858_ (.A(_04587_),
    .B(_04588_),
    .C(_04589_),
    .X(_04590_));
 sg13g2_nor2_1 _12859_ (.A(_04586_),
    .B(_04590_),
    .Y(_04591_));
 sg13g2_o21ai_1 _12860_ (.B1(_04591_),
    .Y(_04592_),
    .A1(_04581_),
    .A2(_04583_));
 sg13g2_nor2_1 _12861_ (.A(_04293_),
    .B(_04588_),
    .Y(_04593_));
 sg13g2_nand2_1 _12862_ (.Y(_04594_),
    .A(_04293_),
    .B(_04588_));
 sg13g2_o21ai_1 _12863_ (.B1(_04594_),
    .Y(_04595_),
    .A1(\am_sdr0.cic1.comb3_in_del[10] ),
    .A2(_04593_));
 sg13g2_o21ai_1 _12864_ (.B1(_04585_),
    .Y(_04596_),
    .A1(_04584_),
    .A2(_04595_));
 sg13g2_nand2_1 _12865_ (.Y(_04597_),
    .A(_04592_),
    .B(_04596_));
 sg13g2_buf_1 _12866_ (.A(\am_sdr0.cic1.comb3_in_del[12] ),
    .X(_04598_));
 sg13g2_xor2_1 _12867_ (.B(_04598_),
    .A(_04364_),
    .X(_04599_));
 sg13g2_xnor2_1 _12868_ (.Y(_04600_),
    .A(_04597_),
    .B(_04599_));
 sg13g2_nor2b_1 _12869_ (.A(net291),
    .B_N(\am_sdr0.cic1.comb3[12] ),
    .Y(_04601_));
 sg13g2_a21oi_1 _12870_ (.A1(_04244_),
    .A2(_04600_),
    .Y(_04602_),
    .B1(_04601_));
 sg13g2_nor2_1 _12871_ (.A(net111),
    .B(_04602_),
    .Y(_00486_));
 sg13g2_nor2_1 _12872_ (.A(net236),
    .B(\am_sdr0.cic1.comb3[13] ),
    .Y(_04603_));
 sg13g2_nor3_1 _12873_ (.A(_04586_),
    .B(_04590_),
    .C(_04599_),
    .Y(_04604_));
 sg13g2_o21ai_1 _12874_ (.B1(_04604_),
    .Y(_04605_),
    .A1(_04581_),
    .A2(_04583_));
 sg13g2_buf_1 _12875_ (.A(_04605_),
    .X(_04606_));
 sg13g2_inv_1 _12876_ (.Y(_04607_),
    .A(_04598_));
 sg13g2_inv_1 _12877_ (.Y(_04608_),
    .A(_04364_));
 sg13g2_o21ai_1 _12878_ (.B1(_04596_),
    .Y(_04609_),
    .A1(_04608_),
    .A2(_04598_));
 sg13g2_o21ai_1 _12879_ (.B1(_04609_),
    .Y(_04610_),
    .A1(_04364_),
    .A2(_04607_));
 sg13g2_buf_1 _12880_ (.A(_04610_),
    .X(_04611_));
 sg13g2_nand2_2 _12881_ (.Y(_04612_),
    .A(_04606_),
    .B(_04611_));
 sg13g2_buf_2 _12882_ (.A(\am_sdr0.cic1.comb3_in_del[13] ),
    .X(_04613_));
 sg13g2_xor2_1 _12883_ (.B(_04613_),
    .A(_04383_),
    .X(_04614_));
 sg13g2_xnor2_1 _12884_ (.Y(_04615_),
    .A(_04612_),
    .B(_04614_));
 sg13g2_nor2_1 _12885_ (.A(net162),
    .B(_04615_),
    .Y(_04616_));
 sg13g2_nor3_1 _12886_ (.A(net160),
    .B(_04603_),
    .C(_04616_),
    .Y(_00487_));
 sg13g2_buf_1 _12887_ (.A(_03962_),
    .X(_04617_));
 sg13g2_inv_1 _12888_ (.Y(_04618_),
    .A(_04612_));
 sg13g2_inv_1 _12889_ (.Y(_04619_),
    .A(_04613_));
 sg13g2_a21oi_1 _12890_ (.A1(_04619_),
    .A2(_04612_),
    .Y(_04620_),
    .B1(_04383_));
 sg13g2_a21oi_1 _12891_ (.A1(_04613_),
    .A2(_04618_),
    .Y(_04621_),
    .B1(_04620_));
 sg13g2_buf_2 _12892_ (.A(\am_sdr0.cic1.comb3_in_del[14] ),
    .X(_04622_));
 sg13g2_xor2_1 _12893_ (.B(_04622_),
    .A(_04396_),
    .X(_04623_));
 sg13g2_xnor2_1 _12894_ (.Y(_04624_),
    .A(_04621_),
    .B(_04623_));
 sg13g2_nor2b_1 _12895_ (.A(net291),
    .B_N(\am_sdr0.cic1.comb3[14] ),
    .Y(_04625_));
 sg13g2_a21oi_1 _12896_ (.A1(net233),
    .A2(_04624_),
    .Y(_04626_),
    .B1(_04625_));
 sg13g2_nor2_1 _12897_ (.A(_04617_),
    .B(_04626_),
    .Y(_00488_));
 sg13g2_nand2_1 _12898_ (.Y(_04627_),
    .A(net113),
    .B(\am_sdr0.cic1.comb3[15] ));
 sg13g2_nor2_1 _12899_ (.A(_04613_),
    .B(_04622_),
    .Y(_04628_));
 sg13g2_inv_1 _12900_ (.Y(_04629_),
    .A(_04383_));
 sg13g2_nor2_1 _12901_ (.A(_04629_),
    .B(_04622_),
    .Y(_04630_));
 sg13g2_o21ai_1 _12902_ (.B1(_04612_),
    .Y(_04631_),
    .A1(_04628_),
    .A2(_04630_));
 sg13g2_buf_1 _12903_ (.A(_04631_),
    .X(_04632_));
 sg13g2_nor3_1 _12904_ (.A(_04629_),
    .B(_04613_),
    .C(_04622_),
    .Y(_04633_));
 sg13g2_nor2_1 _12905_ (.A(_04396_),
    .B(_04633_),
    .Y(_04634_));
 sg13g2_nand4_1 _12906_ (.B(_04622_),
    .C(_04606_),
    .A(_04613_),
    .Y(_04635_),
    .D(_04611_));
 sg13g2_nand4_1 _12907_ (.B(_04622_),
    .C(_04606_),
    .A(_04629_),
    .Y(_04636_),
    .D(_04611_));
 sg13g2_nand3_1 _12908_ (.B(_04613_),
    .C(_04622_),
    .A(_04629_),
    .Y(_04637_));
 sg13g2_nand3_1 _12909_ (.B(_04636_),
    .C(_04637_),
    .A(_04635_),
    .Y(_04638_));
 sg13g2_buf_1 _12910_ (.A(_04638_),
    .X(_04639_));
 sg13g2_a21oi_2 _12911_ (.B1(_04639_),
    .Y(_04640_),
    .A2(_04634_),
    .A1(_04632_));
 sg13g2_buf_1 _12912_ (.A(\am_sdr0.cic1.comb3_in_del[15] ),
    .X(_04641_));
 sg13g2_xor2_1 _12913_ (.B(_04641_),
    .A(_04398_),
    .X(_04642_));
 sg13g2_xnor2_1 _12914_ (.Y(_04643_),
    .A(_04640_),
    .B(_04642_));
 sg13g2_nand2_1 _12915_ (.Y(_04644_),
    .A(net237),
    .B(_04643_));
 sg13g2_a21oi_1 _12916_ (.A1(_04627_),
    .A2(_04644_),
    .Y(_00489_),
    .B1(net104));
 sg13g2_inv_1 _12917_ (.Y(_04645_),
    .A(_04640_));
 sg13g2_inv_1 _12918_ (.Y(_04646_),
    .A(_04641_));
 sg13g2_a21oi_1 _12919_ (.A1(_04646_),
    .A2(_04640_),
    .Y(_04647_),
    .B1(_04398_));
 sg13g2_a21oi_1 _12920_ (.A1(_04641_),
    .A2(_04645_),
    .Y(_04648_),
    .B1(_04647_));
 sg13g2_buf_1 _12921_ (.A(\am_sdr0.cic1.comb3_in_del[16] ),
    .X(_04649_));
 sg13g2_xor2_1 _12922_ (.B(_04649_),
    .A(_04420_),
    .X(_04650_));
 sg13g2_xnor2_1 _12923_ (.Y(_04651_),
    .A(_04648_),
    .B(_04650_));
 sg13g2_nor2b_1 _12924_ (.A(_04001_),
    .B_N(\am_sdr0.cic1.comb3[16] ),
    .Y(_04652_));
 sg13g2_a21oi_1 _12925_ (.A1(net233),
    .A2(_04651_),
    .Y(_04653_),
    .B1(_04652_));
 sg13g2_nor2_1 _12926_ (.A(_04617_),
    .B(_04653_),
    .Y(_00490_));
 sg13g2_nor2_1 _12927_ (.A(_04421_),
    .B(_04649_),
    .Y(_04654_));
 sg13g2_or2_1 _12928_ (.X(_04655_),
    .B(_04649_),
    .A(_04641_));
 sg13g2_nand2b_1 _12929_ (.Y(_04656_),
    .B(_04398_),
    .A_N(_04649_));
 sg13g2_a221oi_1 _12930_ (.B2(_04656_),
    .C1(_04639_),
    .B1(_04655_),
    .A1(_04632_),
    .Y(_04657_),
    .A2(_04634_));
 sg13g2_nand2_1 _12931_ (.Y(_04658_),
    .A(_04646_),
    .B(_04420_));
 sg13g2_nand2_1 _12932_ (.Y(_04659_),
    .A(_04398_),
    .B(_04420_));
 sg13g2_a221oi_1 _12933_ (.B2(_04659_),
    .C1(_04639_),
    .B1(_04658_),
    .A1(_04632_),
    .Y(_04660_),
    .A2(_04634_));
 sg13g2_nand2_1 _12934_ (.Y(_04661_),
    .A(_04398_),
    .B(_04646_));
 sg13g2_a21oi_1 _12935_ (.A1(_04421_),
    .A2(_04649_),
    .Y(_04662_),
    .B1(_04661_));
 sg13g2_nor4_2 _12936_ (.A(_04654_),
    .B(_04657_),
    .C(_04660_),
    .Y(_04663_),
    .D(_04662_));
 sg13g2_buf_1 _12937_ (.A(\am_sdr0.cic1.comb3_in_del[17] ),
    .X(_04664_));
 sg13g2_xor2_1 _12938_ (.B(_04664_),
    .A(_04429_),
    .X(_04665_));
 sg13g2_xnor2_1 _12939_ (.Y(_04666_),
    .A(_04663_),
    .B(_04665_));
 sg13g2_o21ai_1 _12940_ (.B1(_03002_),
    .Y(_04667_),
    .A1(net236),
    .A2(\am_sdr0.cic1.comb3[17] ));
 sg13g2_a21oi_1 _12941_ (.A1(net240),
    .A2(_04666_),
    .Y(_00491_),
    .B1(_04667_));
 sg13g2_nand2_1 _12942_ (.Y(_04668_),
    .A(_04011_),
    .B(\am_sdr0.cic1.comb3[18] ));
 sg13g2_inv_1 _12943_ (.Y(_04669_),
    .A(_04429_));
 sg13g2_a21o_1 _12944_ (.A2(_04663_),
    .A1(_04664_),
    .B1(_04669_),
    .X(_04670_));
 sg13g2_or2_1 _12945_ (.X(_04671_),
    .B(_04663_),
    .A(_04664_));
 sg13g2_buf_1 _12946_ (.A(\am_sdr0.cic1.comb3_in_del[18] ),
    .X(_04672_));
 sg13g2_xor2_1 _12947_ (.B(_04672_),
    .A(_04442_),
    .X(_04673_));
 sg13g2_nand2_1 _12948_ (.Y(_04674_),
    .A(_04000_),
    .B(_04673_));
 sg13g2_a21o_1 _12949_ (.A2(_04671_),
    .A1(_04670_),
    .B1(_04674_),
    .X(_04675_));
 sg13g2_nor2_1 _12950_ (.A(_04010_),
    .B(_04673_),
    .Y(_04676_));
 sg13g2_nand3_1 _12951_ (.B(_04671_),
    .C(_04676_),
    .A(_04670_),
    .Y(_04677_));
 sg13g2_nand3_1 _12952_ (.B(_04675_),
    .C(_04677_),
    .A(_04668_),
    .Y(_04678_));
 sg13g2_and2_1 _12953_ (.A(_02809_),
    .B(_04678_),
    .X(_00492_));
 sg13g2_o21ai_1 _12954_ (.B1(net301),
    .Y(_04679_),
    .A1(_04067_),
    .A2(\am_sdr0.cic1.comb3[19] ));
 sg13g2_inv_1 _12955_ (.Y(_04680_),
    .A(_04442_));
 sg13g2_nor2_1 _12956_ (.A(_04680_),
    .B(_04672_),
    .Y(_04681_));
 sg13g2_a221oi_1 _12957_ (.B2(_04672_),
    .C1(_04663_),
    .B1(_04680_),
    .A1(_04669_),
    .Y(_04682_),
    .A2(_04664_));
 sg13g2_nand2b_1 _12958_ (.Y(_04683_),
    .B(_04429_),
    .A_N(_04664_));
 sg13g2_a21oi_1 _12959_ (.A1(_04680_),
    .A2(_04672_),
    .Y(_04684_),
    .B1(_04683_));
 sg13g2_nor3_1 _12960_ (.A(_04681_),
    .B(_04682_),
    .C(_04684_),
    .Y(_04685_));
 sg13g2_xor2_1 _12961_ (.B(\am_sdr0.cic1.comb3_in_del[19] ),
    .A(\am_sdr0.cic1.comb2[19] ),
    .X(_04686_));
 sg13g2_and3_1 _12962_ (.X(_04687_),
    .A(_04067_),
    .B(_04685_),
    .C(_04686_));
 sg13g2_nor3_1 _12963_ (.A(_04011_),
    .B(_04685_),
    .C(_04686_),
    .Y(_04688_));
 sg13g2_nor3_1 _12964_ (.A(_04679_),
    .B(_04687_),
    .C(_04688_),
    .Y(_00493_));
 sg13g2_nand2_1 _12965_ (.Y(_04689_),
    .A(\am_sdr0.cic1.comb2[0] ),
    .B(net229));
 sg13g2_nand2_1 _12966_ (.Y(_04690_),
    .A(\am_sdr0.cic1.comb3_in_del[0] ),
    .B(_04542_));
 sg13g2_a21oi_1 _12967_ (.A1(_04689_),
    .A2(_04690_),
    .Y(_00494_),
    .B1(_04544_));
 sg13g2_buf_1 _12968_ (.A(_04005_),
    .X(_04691_));
 sg13g2_nand2_1 _12969_ (.Y(_04692_),
    .A(_04293_),
    .B(net228));
 sg13g2_nand2_1 _12970_ (.Y(_04693_),
    .A(\am_sdr0.cic1.comb3_in_del[10] ),
    .B(net158));
 sg13g2_a21oi_1 _12971_ (.A1(_04692_),
    .A2(_04693_),
    .Y(_00495_),
    .B1(net104));
 sg13g2_nand2_1 _12972_ (.Y(_04694_),
    .A(_04351_),
    .B(net228));
 sg13g2_nand2_1 _12973_ (.Y(_04695_),
    .A(\am_sdr0.cic1.comb3_in_del[11] ),
    .B(net158));
 sg13g2_buf_1 _12974_ (.A(_02778_),
    .X(_04696_));
 sg13g2_buf_1 _12975_ (.A(_04696_),
    .X(_04697_));
 sg13g2_a21oi_1 _12976_ (.A1(_04694_),
    .A2(_04695_),
    .Y(_00496_),
    .B1(net102));
 sg13g2_nand2_1 _12977_ (.Y(_04698_),
    .A(_04364_),
    .B(net228));
 sg13g2_buf_1 _12978_ (.A(_04010_),
    .X(_04699_));
 sg13g2_nand2_1 _12979_ (.Y(_04700_),
    .A(_04598_),
    .B(net157));
 sg13g2_a21oi_1 _12980_ (.A1(_04698_),
    .A2(_04700_),
    .Y(_00497_),
    .B1(net102));
 sg13g2_nand2_1 _12981_ (.Y(_04701_),
    .A(_04383_),
    .B(net228));
 sg13g2_nand2_1 _12982_ (.Y(_04702_),
    .A(_04613_),
    .B(net157));
 sg13g2_a21oi_1 _12983_ (.A1(_04701_),
    .A2(_04702_),
    .Y(_00498_),
    .B1(net102));
 sg13g2_nand2_1 _12984_ (.Y(_04703_),
    .A(_04396_),
    .B(net228));
 sg13g2_nand2_1 _12985_ (.Y(_04704_),
    .A(_04622_),
    .B(net157));
 sg13g2_a21oi_1 _12986_ (.A1(_04703_),
    .A2(_04704_),
    .Y(_00499_),
    .B1(net102));
 sg13g2_nand2_1 _12987_ (.Y(_04705_),
    .A(_04398_),
    .B(net228));
 sg13g2_nand2_1 _12988_ (.Y(_04706_),
    .A(_04641_),
    .B(net157));
 sg13g2_a21oi_1 _12989_ (.A1(_04705_),
    .A2(_04706_),
    .Y(_00500_),
    .B1(net102));
 sg13g2_nand2_1 _12990_ (.Y(_04707_),
    .A(_04420_),
    .B(net228));
 sg13g2_nand2_1 _12991_ (.Y(_04708_),
    .A(_04649_),
    .B(net157));
 sg13g2_a21oi_1 _12992_ (.A1(_04707_),
    .A2(_04708_),
    .Y(_00501_),
    .B1(net102));
 sg13g2_nand2_1 _12993_ (.Y(_04709_),
    .A(_04429_),
    .B(net228));
 sg13g2_nand2_1 _12994_ (.Y(_04710_),
    .A(_04664_),
    .B(net157));
 sg13g2_a21oi_1 _12995_ (.A1(_04709_),
    .A2(_04710_),
    .Y(_00502_),
    .B1(net102));
 sg13g2_nand2_1 _12996_ (.Y(_04711_),
    .A(_04442_),
    .B(_04691_));
 sg13g2_nand2_1 _12997_ (.Y(_04712_),
    .A(_04672_),
    .B(_04699_));
 sg13g2_a21oi_1 _12998_ (.A1(_04711_),
    .A2(_04712_),
    .Y(_00503_),
    .B1(_04697_));
 sg13g2_nand2_1 _12999_ (.Y(_04713_),
    .A(\am_sdr0.cic1.comb2[19] ),
    .B(_04691_));
 sg13g2_nand2_1 _13000_ (.Y(_04714_),
    .A(\am_sdr0.cic1.comb3_in_del[19] ),
    .B(_04699_));
 sg13g2_a21oi_1 _13001_ (.A1(_04713_),
    .A2(_04714_),
    .Y(_00504_),
    .B1(_04697_));
 sg13g2_nand2_1 _13002_ (.Y(_04715_),
    .A(\am_sdr0.cic1.comb2[1] ),
    .B(_04014_));
 sg13g2_nand2_1 _13003_ (.Y(_04716_),
    .A(\am_sdr0.cic1.comb3_in_del[1] ),
    .B(net157));
 sg13g2_a21oi_1 _13004_ (.A1(_04715_),
    .A2(_04716_),
    .Y(_00505_),
    .B1(net102));
 sg13g2_nand2_1 _13005_ (.Y(_04717_),
    .A(_04462_),
    .B(net238));
 sg13g2_nand2_1 _13006_ (.Y(_04718_),
    .A(\am_sdr0.cic1.comb3_in_del[2] ),
    .B(net157));
 sg13g2_buf_1 _13007_ (.A(_04696_),
    .X(_04719_));
 sg13g2_a21oi_1 _13008_ (.A1(_04717_),
    .A2(_04718_),
    .Y(_00506_),
    .B1(net101));
 sg13g2_nand2_1 _13009_ (.Y(_04720_),
    .A(\am_sdr0.cic1.comb2[3] ),
    .B(net238));
 sg13g2_buf_1 _13010_ (.A(_04010_),
    .X(_04721_));
 sg13g2_nand2_1 _13011_ (.Y(_04722_),
    .A(\am_sdr0.cic1.comb3_in_del[3] ),
    .B(net156));
 sg13g2_a21oi_1 _13012_ (.A1(_04720_),
    .A2(_04722_),
    .Y(_00507_),
    .B1(net101));
 sg13g2_nand2_1 _13013_ (.Y(_04723_),
    .A(_04473_),
    .B(net238));
 sg13g2_nand2_1 _13014_ (.Y(_04724_),
    .A(\am_sdr0.cic1.comb3_in_del[4] ),
    .B(net156));
 sg13g2_a21oi_1 _13015_ (.A1(_04723_),
    .A2(_04724_),
    .Y(_00508_),
    .B1(net101));
 sg13g2_nand2_1 _13016_ (.Y(_04725_),
    .A(_04478_),
    .B(net238));
 sg13g2_nand2_1 _13017_ (.Y(_04726_),
    .A(\am_sdr0.cic1.comb3_in_del[5] ),
    .B(net156));
 sg13g2_a21oi_1 _13018_ (.A1(_04725_),
    .A2(_04726_),
    .Y(_00509_),
    .B1(net101));
 sg13g2_nand2_1 _13019_ (.Y(_04727_),
    .A(_04489_),
    .B(net238));
 sg13g2_nand2_1 _13020_ (.Y(_04728_),
    .A(\am_sdr0.cic1.comb3_in_del[6] ),
    .B(net156));
 sg13g2_a21oi_1 _13021_ (.A1(_04727_),
    .A2(_04728_),
    .Y(_00510_),
    .B1(_04719_));
 sg13g2_nand2_1 _13022_ (.Y(_04729_),
    .A(_04494_),
    .B(net238));
 sg13g2_nand2_1 _13023_ (.Y(_04730_),
    .A(\am_sdr0.cic1.comb3_in_del[7] ),
    .B(net156));
 sg13g2_a21oi_1 _13024_ (.A1(_04729_),
    .A2(_04730_),
    .Y(_00511_),
    .B1(net101));
 sg13g2_nand2_1 _13025_ (.Y(_04731_),
    .A(\am_sdr0.cic1.comb2[8] ),
    .B(net238));
 sg13g2_nand2_1 _13026_ (.Y(_04732_),
    .A(\am_sdr0.cic1.comb3_in_del[8] ),
    .B(net156));
 sg13g2_a21oi_1 _13027_ (.A1(_04731_),
    .A2(_04732_),
    .Y(_00512_),
    .B1(net101));
 sg13g2_nand2_1 _13028_ (.Y(_04733_),
    .A(_04505_),
    .B(net238));
 sg13g2_nand2_1 _13029_ (.Y(_04734_),
    .A(\am_sdr0.cic1.comb3_in_del[9] ),
    .B(_04721_));
 sg13g2_a21oi_1 _13030_ (.A1(_04733_),
    .A2(_04734_),
    .Y(_00513_),
    .B1(net101));
 sg13g2_xnor2_1 _13031_ (.Y(_04735_),
    .A(\am_sdr0.Q_out[0] ),
    .B(\am_sdr0.cic1.integ1[0] ));
 sg13g2_nor2_1 _13032_ (.A(net103),
    .B(_04735_),
    .Y(_00522_));
 sg13g2_buf_2 _13033_ (.A(\am_sdr0.cic1.integ1[9] ),
    .X(_04736_));
 sg13g2_buf_1 _13034_ (.A(\am_sdr0.cic1.integ1[6] ),
    .X(_04737_));
 sg13g2_buf_1 _13035_ (.A(\am_sdr0.cic1.integ1[5] ),
    .X(_04738_));
 sg13g2_inv_1 _13036_ (.Y(_04739_),
    .A(_04738_));
 sg13g2_buf_2 _13037_ (.A(\am_sdr0.cic1.integ1[4] ),
    .X(_04740_));
 sg13g2_inv_1 _13038_ (.Y(_04741_),
    .A(\am_sdr0.Q_out[3] ));
 sg13g2_nor2_1 _13039_ (.A(\am_sdr0.Q_out[1] ),
    .B(\am_sdr0.cic1.integ1[1] ),
    .Y(_04742_));
 sg13g2_a22oi_1 _13040_ (.Y(_04743_),
    .B1(\am_sdr0.Q_out[1] ),
    .B2(\am_sdr0.cic1.integ1[1] ),
    .A2(\am_sdr0.cic1.integ1[0] ),
    .A1(\am_sdr0.Q_out[0] ));
 sg13g2_nand2_1 _13041_ (.Y(_04744_),
    .A(\am_sdr0.Q_out[2] ),
    .B(\am_sdr0.cic1.integ1[2] ));
 sg13g2_o21ai_1 _13042_ (.B1(_04744_),
    .Y(_04745_),
    .A1(_04742_),
    .A2(_04743_));
 sg13g2_or2_1 _13043_ (.X(_04746_),
    .B(\am_sdr0.cic1.integ1[2] ),
    .A(\am_sdr0.Q_out[2] ));
 sg13g2_buf_1 _13044_ (.A(_04746_),
    .X(_04747_));
 sg13g2_buf_2 _13045_ (.A(\am_sdr0.cic1.integ1[3] ),
    .X(_04748_));
 sg13g2_a21oi_1 _13046_ (.A1(_04745_),
    .A2(_04747_),
    .Y(_04749_),
    .B1(_04748_));
 sg13g2_nand3_1 _13047_ (.B(_04745_),
    .C(_04747_),
    .A(_04748_),
    .Y(_04750_));
 sg13g2_o21ai_1 _13048_ (.B1(_04750_),
    .Y(_04751_),
    .A1(_04741_),
    .A2(_04749_));
 sg13g2_buf_1 _13049_ (.A(_04751_),
    .X(_04752_));
 sg13g2_nand2_1 _13050_ (.Y(_04753_),
    .A(_04740_),
    .B(_04752_));
 sg13g2_o21ai_1 _13051_ (.B1(\am_sdr0.Q_out[4] ),
    .Y(_04754_),
    .A1(_04740_),
    .A2(_04752_));
 sg13g2_buf_1 _13052_ (.A(_04754_),
    .X(_04755_));
 sg13g2_nand3_1 _13053_ (.B(_04753_),
    .C(_04755_),
    .A(_04739_),
    .Y(_04756_));
 sg13g2_a21oi_1 _13054_ (.A1(_04753_),
    .A2(_04755_),
    .Y(_04757_),
    .B1(_04739_));
 sg13g2_a21o_1 _13055_ (.A2(_04756_),
    .A1(\am_sdr0.Q_out[5] ),
    .B1(_04757_),
    .X(_04758_));
 sg13g2_buf_1 _13056_ (.A(_04758_),
    .X(_04759_));
 sg13g2_nand2_1 _13057_ (.Y(_04760_),
    .A(_04737_),
    .B(_04759_));
 sg13g2_o21ai_1 _13058_ (.B1(\am_sdr0.Q_out[6] ),
    .Y(_04761_),
    .A1(_04737_),
    .A2(_04759_));
 sg13g2_buf_1 _13059_ (.A(_04761_),
    .X(_04762_));
 sg13g2_buf_2 _13060_ (.A(\am_sdr0.cic1.integ1[8] ),
    .X(_04763_));
 sg13g2_inv_1 _13061_ (.Y(_04764_),
    .A(_04763_));
 sg13g2_a21oi_1 _13062_ (.A1(_04760_),
    .A2(_04762_),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_buf_1 _13063_ (.A(\am_sdr0.Q_out[7] ),
    .X(_04766_));
 sg13g2_a21oi_1 _13064_ (.A1(_04736_),
    .A2(_04765_),
    .Y(_04767_),
    .B1(net346));
 sg13g2_inv_2 _13065_ (.Y(_04768_),
    .A(_04736_));
 sg13g2_nand4_1 _13066_ (.B(_04768_),
    .C(_04760_),
    .A(_04764_),
    .Y(_04769_),
    .D(_04762_));
 sg13g2_buf_2 _13067_ (.A(\am_sdr0.cic1.integ1[7] ),
    .X(_04770_));
 sg13g2_a21oi_1 _13068_ (.A1(net346),
    .A2(_04769_),
    .Y(_04771_),
    .B1(_04770_));
 sg13g2_nor2_2 _13069_ (.A(_04767_),
    .B(_04771_),
    .Y(_04772_));
 sg13g2_buf_1 _13070_ (.A(net346),
    .X(_04773_));
 sg13g2_buf_1 _13071_ (.A(net290),
    .X(_04774_));
 sg13g2_buf_1 _13072_ (.A(\am_sdr0.cic1.integ1[10] ),
    .X(_04775_));
 sg13g2_xor2_1 _13073_ (.B(net345),
    .A(net227),
    .X(_04776_));
 sg13g2_xnor2_1 _13074_ (.Y(_04777_),
    .A(_04772_),
    .B(_04776_));
 sg13g2_nor2_1 _13075_ (.A(net103),
    .B(_04777_),
    .Y(_00523_));
 sg13g2_inv_1 _13076_ (.Y(_04778_),
    .A(_04770_));
 sg13g2_inv_1 _13077_ (.Y(_04779_),
    .A(net345));
 sg13g2_nor2_1 _13078_ (.A(_04768_),
    .B(_04779_),
    .Y(_04780_));
 sg13g2_a21oi_1 _13079_ (.A1(_04765_),
    .A2(_04780_),
    .Y(_04781_),
    .B1(net346));
 sg13g2_o21ai_1 _13080_ (.B1(net346),
    .Y(_04782_),
    .A1(net345),
    .A2(_04769_));
 sg13g2_o21ai_1 _13081_ (.B1(_04782_),
    .Y(_04783_),
    .A1(_04778_),
    .A2(_04781_));
 sg13g2_buf_1 _13082_ (.A(_04783_),
    .X(_04784_));
 sg13g2_buf_2 _13083_ (.A(\am_sdr0.cic1.integ1[11] ),
    .X(_04785_));
 sg13g2_xor2_1 _13084_ (.B(_04785_),
    .A(net227),
    .X(_04786_));
 sg13g2_xnor2_1 _13085_ (.Y(_04787_),
    .A(_04784_),
    .B(_04786_));
 sg13g2_nor2_1 _13086_ (.A(net103),
    .B(_04787_),
    .Y(_00524_));
 sg13g2_buf_1 _13087_ (.A(\am_sdr0.cic1.integ1[12] ),
    .X(_04788_));
 sg13g2_inv_1 _13088_ (.Y(_04789_),
    .A(_04785_));
 sg13g2_nor2_1 _13089_ (.A(net346),
    .B(_04789_),
    .Y(_04790_));
 sg13g2_nand2_1 _13090_ (.Y(_04791_),
    .A(_04784_),
    .B(_04790_));
 sg13g2_nor2_1 _13091_ (.A(net345),
    .B(_04785_),
    .Y(_04792_));
 sg13g2_nand3_1 _13092_ (.B(_04771_),
    .C(_04792_),
    .A(net227),
    .Y(_04793_));
 sg13g2_buf_1 _13093_ (.A(_04793_),
    .X(_04794_));
 sg13g2_nand3_1 _13094_ (.B(_04791_),
    .C(_04794_),
    .A(_04788_),
    .Y(_04795_));
 sg13g2_a21o_1 _13095_ (.A2(_04794_),
    .A1(_04791_),
    .B1(net344),
    .X(_04796_));
 sg13g2_a21oi_1 _13096_ (.A1(_04795_),
    .A2(_04796_),
    .Y(_00525_),
    .B1(_04719_));
 sg13g2_buf_2 _13097_ (.A(\am_sdr0.cic1.integ1[13] ),
    .X(_04797_));
 sg13g2_inv_1 _13098_ (.Y(_04798_),
    .A(_04791_));
 sg13g2_nor2_1 _13099_ (.A(net344),
    .B(_04794_),
    .Y(_04799_));
 sg13g2_a21oi_1 _13100_ (.A1(net344),
    .A2(_04798_),
    .Y(_04800_),
    .B1(_04799_));
 sg13g2_xor2_1 _13101_ (.B(_04800_),
    .A(_04797_),
    .X(_04801_));
 sg13g2_nor2_1 _13102_ (.A(net103),
    .B(_04801_),
    .Y(_00526_));
 sg13g2_buf_1 _13103_ (.A(\am_sdr0.cic1.integ1[14] ),
    .X(_04802_));
 sg13g2_and2_1 _13104_ (.A(net344),
    .B(_04797_),
    .X(_04803_));
 sg13g2_buf_1 _13105_ (.A(_04803_),
    .X(_04804_));
 sg13g2_nor2_1 _13106_ (.A(_04788_),
    .B(_04797_),
    .Y(_04805_));
 sg13g2_nor2b_1 _13107_ (.A(_04794_),
    .B_N(_04805_),
    .Y(_04806_));
 sg13g2_a21oi_1 _13108_ (.A1(_04798_),
    .A2(_04804_),
    .Y(_04807_),
    .B1(_04806_));
 sg13g2_xor2_1 _13109_ (.B(_04807_),
    .A(net343),
    .X(_04808_));
 sg13g2_nor2_1 _13110_ (.A(net103),
    .B(_04808_),
    .Y(_00527_));
 sg13g2_nand2_2 _13111_ (.Y(_04809_),
    .A(_04760_),
    .B(_04762_));
 sg13g2_nand3_1 _13112_ (.B(net343),
    .C(_04804_),
    .A(_04785_),
    .Y(_04810_));
 sg13g2_nor4_1 _13113_ (.A(_04778_),
    .B(_04768_),
    .C(_04779_),
    .D(_04810_),
    .Y(_04811_));
 sg13g2_a21o_1 _13114_ (.A2(_04811_),
    .A1(_04809_),
    .B1(net346),
    .X(_04812_));
 sg13g2_nand2b_1 _13115_ (.Y(_04813_),
    .B(_04805_),
    .A_N(net343));
 sg13g2_nand3_1 _13116_ (.B(_04768_),
    .C(_04792_),
    .A(_04778_),
    .Y(_04814_));
 sg13g2_or3_1 _13117_ (.A(_04809_),
    .B(_04813_),
    .C(_04814_),
    .X(_04815_));
 sg13g2_a22oi_1 _13118_ (.Y(_04816_),
    .B1(_04815_),
    .B2(net290),
    .A2(_04812_),
    .A1(_04763_));
 sg13g2_buf_1 _13119_ (.A(_04816_),
    .X(_04817_));
 sg13g2_buf_1 _13120_ (.A(\am_sdr0.cic1.integ1[15] ),
    .X(_04818_));
 sg13g2_xnor2_1 _13121_ (.Y(_04819_),
    .A(_04774_),
    .B(net342));
 sg13g2_xnor2_1 _13122_ (.Y(_04820_),
    .A(_04817_),
    .B(_04819_));
 sg13g2_nor2_1 _13123_ (.A(net103),
    .B(_04820_),
    .Y(_00528_));
 sg13g2_inv_1 _13124_ (.Y(_04821_),
    .A(net342));
 sg13g2_nor2_1 _13125_ (.A(_04821_),
    .B(_04810_),
    .Y(_04822_));
 sg13g2_a21oi_1 _13126_ (.A1(_04772_),
    .A2(_04822_),
    .Y(_04823_),
    .B1(net290));
 sg13g2_nor2_1 _13127_ (.A(net342),
    .B(_04813_),
    .Y(_04824_));
 sg13g2_nand2_1 _13128_ (.Y(_04825_),
    .A(_04789_),
    .B(_04824_));
 sg13g2_o21ai_1 _13129_ (.B1(net290),
    .Y(_04826_),
    .A1(_04772_),
    .A2(_04825_));
 sg13g2_o21ai_1 _13130_ (.B1(_04826_),
    .Y(_04827_),
    .A1(_04779_),
    .A2(_04823_));
 sg13g2_buf_1 _13131_ (.A(_04827_),
    .X(_04828_));
 sg13g2_buf_1 _13132_ (.A(\am_sdr0.cic1.integ1[16] ),
    .X(_04829_));
 sg13g2_buf_1 _13133_ (.A(_04829_),
    .X(_04830_));
 sg13g2_xor2_1 _13134_ (.B(net289),
    .A(net227),
    .X(_04831_));
 sg13g2_xnor2_1 _13135_ (.Y(_04832_),
    .A(_04828_),
    .B(_04831_));
 sg13g2_nor2_1 _13136_ (.A(net103),
    .B(_04832_),
    .Y(_00529_));
 sg13g2_and4_1 _13137_ (.A(net343),
    .B(net342),
    .C(net289),
    .D(_04804_),
    .X(_04833_));
 sg13g2_a21oi_1 _13138_ (.A1(_04784_),
    .A2(_04833_),
    .Y(_04834_),
    .B1(net290));
 sg13g2_nand2b_1 _13139_ (.Y(_04835_),
    .B(_04824_),
    .A_N(net289));
 sg13g2_o21ai_1 _13140_ (.B1(net290),
    .Y(_04836_),
    .A1(_04784_),
    .A2(_04835_));
 sg13g2_o21ai_1 _13141_ (.B1(_04836_),
    .Y(_04837_),
    .A1(_04789_),
    .A2(_04834_));
 sg13g2_buf_1 _13142_ (.A(_04837_),
    .X(_04838_));
 sg13g2_buf_1 _13143_ (.A(\am_sdr0.cic1.integ1[17] ),
    .X(_04839_));
 sg13g2_xor2_1 _13144_ (.B(net341),
    .A(_04774_),
    .X(_04840_));
 sg13g2_xnor2_1 _13145_ (.Y(_04841_),
    .A(_04838_),
    .B(_04840_));
 sg13g2_nor2_1 _13146_ (.A(net103),
    .B(_04841_),
    .Y(_00530_));
 sg13g2_buf_1 _13147_ (.A(_03962_),
    .X(_04842_));
 sg13g2_buf_2 _13148_ (.A(\am_sdr0.cic1.integ1[18] ),
    .X(_04843_));
 sg13g2_inv_1 _13149_ (.Y(_04844_),
    .A(net346));
 sg13g2_nand3_1 _13150_ (.B(_04789_),
    .C(_04805_),
    .A(net290),
    .Y(_04845_));
 sg13g2_nand3_1 _13151_ (.B(_04790_),
    .C(_04804_),
    .A(net345),
    .Y(_04846_));
 sg13g2_o21ai_1 _13152_ (.B1(_04846_),
    .Y(_04847_),
    .A1(_04775_),
    .A2(_04845_));
 sg13g2_nand2_1 _13153_ (.Y(_04848_),
    .A(_04772_),
    .B(_04847_));
 sg13g2_nand4_1 _13154_ (.B(net342),
    .C(net289),
    .A(net343),
    .Y(_04849_),
    .D(net341));
 sg13g2_nor2_1 _13155_ (.A(_04848_),
    .B(_04849_),
    .Y(_04850_));
 sg13g2_nand2_1 _13156_ (.Y(_04851_),
    .A(_04792_),
    .B(_04824_));
 sg13g2_a21oi_1 _13157_ (.A1(_04772_),
    .A2(_04847_),
    .Y(_04852_),
    .B1(_04851_));
 sg13g2_nor2_1 _13158_ (.A(net289),
    .B(net341),
    .Y(_04853_));
 sg13g2_and2_1 _13159_ (.A(net227),
    .B(_04853_),
    .X(_04854_));
 sg13g2_a22oi_1 _13160_ (.Y(_04855_),
    .B1(_04852_),
    .B2(_04854_),
    .A2(_04850_),
    .A1(_04844_));
 sg13g2_xor2_1 _13161_ (.B(_04855_),
    .A(_04843_),
    .X(_04856_));
 sg13g2_nor2_1 _13162_ (.A(net100),
    .B(_04856_),
    .Y(_00531_));
 sg13g2_buf_1 _13163_ (.A(\am_sdr0.cic1.integ1[19] ),
    .X(_04857_));
 sg13g2_buf_1 _13164_ (.A(_04857_),
    .X(_04858_));
 sg13g2_nor2b_1 _13165_ (.A(_04766_),
    .B_N(_04843_),
    .Y(_04859_));
 sg13g2_nand4_1 _13166_ (.B(net289),
    .C(net341),
    .A(net342),
    .Y(_04860_),
    .D(_04859_));
 sg13g2_nand3b_1 _13167_ (.B(_04853_),
    .C(_04766_),
    .Y(_04861_),
    .A_N(_04843_));
 sg13g2_buf_1 _13168_ (.A(_04861_),
    .X(_04862_));
 sg13g2_nand2b_1 _13169_ (.Y(_04863_),
    .B(_04821_),
    .A_N(_04862_));
 sg13g2_mux2_1 _13170_ (.A0(_04860_),
    .A1(_04863_),
    .S(_04817_),
    .X(_04864_));
 sg13g2_xnor2_1 _13171_ (.Y(_04865_),
    .A(net288),
    .B(_04864_));
 sg13g2_and2_1 _13172_ (.A(net246),
    .B(_04865_),
    .X(_00532_));
 sg13g2_nand2_1 _13173_ (.Y(_04866_),
    .A(\am_sdr0.Q_out[0] ),
    .B(\am_sdr0.cic1.integ1[0] ));
 sg13g2_xnor2_1 _13174_ (.Y(_04867_),
    .A(\am_sdr0.Q_out[1] ),
    .B(\am_sdr0.cic1.integ1[1] ));
 sg13g2_xnor2_1 _13175_ (.Y(_04868_),
    .A(_04866_),
    .B(_04867_));
 sg13g2_nor2_1 _13176_ (.A(net100),
    .B(_04868_),
    .Y(_00533_));
 sg13g2_buf_1 _13177_ (.A(\am_sdr0.cic1.integ1[20] ),
    .X(_04869_));
 sg13g2_buf_1 _13178_ (.A(_04869_),
    .X(_04870_));
 sg13g2_nor2_1 _13179_ (.A(net288),
    .B(_04862_),
    .Y(_04871_));
 sg13g2_and4_1 _13180_ (.A(net289),
    .B(net341),
    .C(net288),
    .D(_04859_),
    .X(_04872_));
 sg13g2_mux2_1 _13181_ (.A0(_04871_),
    .A1(_04872_),
    .S(_04828_),
    .X(_04873_));
 sg13g2_xnor2_1 _13182_ (.Y(_04874_),
    .A(_04870_),
    .B(_04873_));
 sg13g2_nor2_1 _13183_ (.A(net100),
    .B(_04874_),
    .Y(_00534_));
 sg13g2_buf_2 _13184_ (.A(\am_sdr0.cic1.integ1[21] ),
    .X(_04875_));
 sg13g2_or2_1 _13185_ (.X(_04876_),
    .B(_04843_),
    .A(net341));
 sg13g2_nor4_2 _13186_ (.A(_04844_),
    .B(net288),
    .C(_04870_),
    .Y(_04877_),
    .D(_04876_));
 sg13g2_and4_1 _13187_ (.A(net341),
    .B(net288),
    .C(net287),
    .D(_04859_),
    .X(_04878_));
 sg13g2_mux2_1 _13188_ (.A0(_04877_),
    .A1(_04878_),
    .S(_04838_),
    .X(_04879_));
 sg13g2_xnor2_1 _13189_ (.Y(_04880_),
    .A(_04875_),
    .B(_04879_));
 sg13g2_nor2_1 _13190_ (.A(_04842_),
    .B(_04880_),
    .Y(_00535_));
 sg13g2_buf_2 _13191_ (.A(\am_sdr0.cic1.integ1[22] ),
    .X(_04881_));
 sg13g2_inv_1 _13192_ (.Y(_04882_),
    .A(_04881_));
 sg13g2_and4_1 _13193_ (.A(net288),
    .B(net287),
    .C(_04875_),
    .D(_04859_),
    .X(_04883_));
 sg13g2_or3_1 _13194_ (.A(net288),
    .B(net287),
    .C(_04862_),
    .X(_04884_));
 sg13g2_nor2_1 _13195_ (.A(_04875_),
    .B(_04884_),
    .Y(_04885_));
 sg13g2_a22oi_1 _13196_ (.Y(_04886_),
    .B1(_04885_),
    .B2(_04852_),
    .A2(_04883_),
    .A1(_04850_));
 sg13g2_xnor2_1 _13197_ (.Y(_04887_),
    .A(_04882_),
    .B(_04886_));
 sg13g2_nor2_1 _13198_ (.A(_04842_),
    .B(_04887_),
    .Y(_00536_));
 sg13g2_buf_2 _13199_ (.A(\am_sdr0.cic1.integ1[23] ),
    .X(_04888_));
 sg13g2_a21oi_1 _13200_ (.A1(_04860_),
    .A2(_04863_),
    .Y(_04889_),
    .B1(_04817_));
 sg13g2_inv_1 _13201_ (.Y(_04890_),
    .A(_04875_));
 sg13g2_nor3_1 _13202_ (.A(_04773_),
    .B(_04890_),
    .C(_04882_),
    .Y(_04891_));
 sg13g2_nand4_1 _13203_ (.B(net287),
    .C(_04889_),
    .A(net288),
    .Y(_04892_),
    .D(_04891_));
 sg13g2_nand3_1 _13204_ (.B(_04882_),
    .C(_04885_),
    .A(_04821_),
    .Y(_04893_));
 sg13g2_a22oi_1 _13205_ (.Y(_04894_),
    .B1(_04892_),
    .B2(_04893_),
    .A2(_04889_),
    .A1(net227));
 sg13g2_xnor2_1 _13206_ (.Y(_04895_),
    .A(_04888_),
    .B(_04894_));
 sg13g2_nor2_1 _13207_ (.A(net100),
    .B(_04895_),
    .Y(_00537_));
 sg13g2_buf_2 _13208_ (.A(\am_sdr0.cic1.integ1[24] ),
    .X(_04896_));
 sg13g2_and2_1 _13209_ (.A(net297),
    .B(_04896_),
    .X(_04897_));
 sg13g2_nor2_1 _13210_ (.A(net251),
    .B(_04896_),
    .Y(_04898_));
 sg13g2_nor3_2 _13211_ (.A(_04875_),
    .B(_04881_),
    .C(_04888_),
    .Y(_04899_));
 sg13g2_nor2b_1 _13212_ (.A(_04884_),
    .B_N(_04899_),
    .Y(_04900_));
 sg13g2_or2_1 _13213_ (.X(_04901_),
    .B(_04871_),
    .A(_04872_));
 sg13g2_nand2_1 _13214_ (.Y(_04902_),
    .A(_04888_),
    .B(_04891_));
 sg13g2_a21oi_1 _13215_ (.A1(_04773_),
    .A2(_04899_),
    .Y(_04903_),
    .B1(net287));
 sg13g2_a21oi_1 _13216_ (.A1(net287),
    .A2(_04902_),
    .Y(_04904_),
    .B1(_04903_));
 sg13g2_nand3_1 _13217_ (.B(_04901_),
    .C(_04904_),
    .A(_04828_),
    .Y(_04905_));
 sg13g2_mux2_1 _13218_ (.A0(_04844_),
    .A1(_04900_),
    .S(_04905_),
    .X(_04906_));
 sg13g2_mux2_1 _13219_ (.A0(_04897_),
    .A1(_04898_),
    .S(_04906_),
    .X(_00538_));
 sg13g2_nor2_1 _13220_ (.A(net251),
    .B(\am_sdr0.cic1.integ1[25] ),
    .Y(_04907_));
 sg13g2_and2_1 _13221_ (.A(net303),
    .B(\am_sdr0.cic1.integ1[25] ),
    .X(_04908_));
 sg13g2_nand3b_1 _13222_ (.B(_04877_),
    .C(_04899_),
    .Y(_04909_),
    .A_N(_04896_));
 sg13g2_a21o_1 _13223_ (.A2(_04899_),
    .A1(net290),
    .B1(_04896_),
    .X(_04910_));
 sg13g2_o21ai_1 _13224_ (.B1(_04910_),
    .Y(_04911_),
    .A1(_04877_),
    .A2(_04878_));
 sg13g2_a21oi_1 _13225_ (.A1(_04896_),
    .A2(_04902_),
    .Y(_04912_),
    .B1(_04911_));
 sg13g2_nand2_1 _13226_ (.Y(_04913_),
    .A(_04838_),
    .B(_04912_));
 sg13g2_mux2_1 _13227_ (.A0(net227),
    .A1(_04909_),
    .S(_04913_),
    .X(_04914_));
 sg13g2_mux2_1 _13228_ (.A0(_04907_),
    .A1(_04908_),
    .S(_04914_),
    .X(_00539_));
 sg13g2_nor2_1 _13229_ (.A(_04742_),
    .B(_04743_),
    .Y(_04915_));
 sg13g2_xor2_1 _13230_ (.B(\am_sdr0.cic1.integ1[2] ),
    .A(\am_sdr0.Q_out[2] ),
    .X(_04916_));
 sg13g2_xnor2_1 _13231_ (.Y(_04917_),
    .A(_04915_),
    .B(_04916_));
 sg13g2_nor2_1 _13232_ (.A(net100),
    .B(_04917_),
    .Y(_00540_));
 sg13g2_nand2_1 _13233_ (.Y(_04918_),
    .A(_04745_),
    .B(_04747_));
 sg13g2_xnor2_1 _13234_ (.Y(_04919_),
    .A(\am_sdr0.Q_out[3] ),
    .B(_04748_));
 sg13g2_xnor2_1 _13235_ (.Y(_04920_),
    .A(_04918_),
    .B(_04919_));
 sg13g2_nor2_1 _13236_ (.A(net100),
    .B(_04920_),
    .Y(_00541_));
 sg13g2_xor2_1 _13237_ (.B(_04740_),
    .A(\am_sdr0.Q_out[4] ),
    .X(_04921_));
 sg13g2_xnor2_1 _13238_ (.Y(_04922_),
    .A(_04752_),
    .B(_04921_));
 sg13g2_nor2_1 _13239_ (.A(net100),
    .B(_04922_),
    .Y(_00542_));
 sg13g2_xnor2_1 _13240_ (.Y(_04923_),
    .A(\am_sdr0.Q_out[5] ),
    .B(_04738_));
 sg13g2_and3_1 _13241_ (.X(_04924_),
    .A(_04753_),
    .B(_04755_),
    .C(_04923_));
 sg13g2_a21oi_1 _13242_ (.A1(_04753_),
    .A2(_04755_),
    .Y(_04925_),
    .B1(_04923_));
 sg13g2_nor3_1 _13243_ (.A(net160),
    .B(_04924_),
    .C(_04925_),
    .Y(_00543_));
 sg13g2_xor2_1 _13244_ (.B(_04737_),
    .A(\am_sdr0.Q_out[6] ),
    .X(_04926_));
 sg13g2_xnor2_1 _13245_ (.Y(_04927_),
    .A(_04759_),
    .B(_04926_));
 sg13g2_nor2_1 _13246_ (.A(net100),
    .B(_04927_),
    .Y(_00544_));
 sg13g2_buf_1 _13247_ (.A(_03962_),
    .X(_04928_));
 sg13g2_nor2_1 _13248_ (.A(net227),
    .B(_04778_),
    .Y(_04929_));
 sg13g2_nor2_1 _13249_ (.A(_04844_),
    .B(_04770_),
    .Y(_04930_));
 sg13g2_nor2_1 _13250_ (.A(_04929_),
    .B(_04930_),
    .Y(_04931_));
 sg13g2_xor2_1 _13251_ (.B(_04931_),
    .A(_04809_),
    .X(_04932_));
 sg13g2_nor2_1 _13252_ (.A(net99),
    .B(_04932_),
    .Y(_00545_));
 sg13g2_mux2_1 _13253_ (.A0(_04930_),
    .A1(_04929_),
    .S(_04809_),
    .X(_04933_));
 sg13g2_xnor2_1 _13254_ (.Y(_04934_),
    .A(_04763_),
    .B(_04933_));
 sg13g2_nor2_1 _13255_ (.A(net99),
    .B(_04934_),
    .Y(_00546_));
 sg13g2_nor2_1 _13256_ (.A(_04763_),
    .B(_04809_),
    .Y(_04935_));
 sg13g2_a22oi_1 _13257_ (.Y(_04936_),
    .B1(_04930_),
    .B2(_04935_),
    .A2(_04929_),
    .A1(_04765_));
 sg13g2_xnor2_1 _13258_ (.Y(_04937_),
    .A(_04768_),
    .B(_04936_));
 sg13g2_nor2_1 _13259_ (.A(net99),
    .B(_04937_),
    .Y(_00547_));
 sg13g2_xnor2_1 _13260_ (.Y(_04938_),
    .A(_04748_),
    .B(\am_sdr0.cic1.integ2[0] ));
 sg13g2_nor2_1 _13261_ (.A(net99),
    .B(_04938_),
    .Y(_00548_));
 sg13g2_buf_2 _13262_ (.A(\am_sdr0.cic1.integ2[10] ),
    .X(_04939_));
 sg13g2_xnor2_1 _13263_ (.Y(_04940_),
    .A(_04939_),
    .B(_04797_));
 sg13g2_buf_2 _13264_ (.A(\am_sdr0.cic1.integ2[3] ),
    .X(_04941_));
 sg13g2_or2_1 _13265_ (.X(_04942_),
    .B(\am_sdr0.cic1.integ2[1] ),
    .A(_04740_));
 sg13g2_and2_1 _13266_ (.A(_04748_),
    .B(\am_sdr0.cic1.integ2[0] ),
    .X(_04943_));
 sg13g2_buf_1 _13267_ (.A(_04943_),
    .X(_04944_));
 sg13g2_and2_1 _13268_ (.A(_04740_),
    .B(\am_sdr0.cic1.integ2[1] ),
    .X(_04945_));
 sg13g2_a221oi_1 _13269_ (.B2(_04944_),
    .C1(_04945_),
    .B1(_04942_),
    .A1(_04738_),
    .Y(_04946_),
    .A2(\am_sdr0.cic1.integ2[2] ));
 sg13g2_buf_1 _13270_ (.A(_04946_),
    .X(_04947_));
 sg13g2_nor2_1 _13271_ (.A(_04738_),
    .B(\am_sdr0.cic1.integ2[2] ),
    .Y(_04948_));
 sg13g2_inv_1 _13272_ (.Y(_04949_),
    .A(_04737_));
 sg13g2_o21ai_1 _13273_ (.B1(_04949_),
    .Y(_04950_),
    .A1(_04947_),
    .A2(_04948_));
 sg13g2_buf_2 _13274_ (.A(\am_sdr0.cic1.integ2[5] ),
    .X(_04951_));
 sg13g2_nor2_1 _13275_ (.A(_04951_),
    .B(_04763_),
    .Y(_04952_));
 sg13g2_buf_2 _13276_ (.A(\am_sdr0.cic1.integ2[4] ),
    .X(_04953_));
 sg13g2_a22oi_1 _13277_ (.Y(_04954_),
    .B1(_04763_),
    .B2(_04951_),
    .A2(_04770_),
    .A1(_04953_));
 sg13g2_buf_2 _13278_ (.A(\am_sdr0.cic1.integ2[6] ),
    .X(_04955_));
 sg13g2_nand2_1 _13279_ (.Y(_04956_),
    .A(_04955_),
    .B(_04736_));
 sg13g2_o21ai_1 _13280_ (.B1(_04956_),
    .Y(_04957_),
    .A1(_04952_),
    .A2(_04954_));
 sg13g2_buf_2 _13281_ (.A(\am_sdr0.cic1.integ2[8] ),
    .X(_04958_));
 sg13g2_nand2_1 _13282_ (.Y(_04959_),
    .A(_04958_),
    .B(_04785_));
 sg13g2_nand2_1 _13283_ (.Y(_04960_),
    .A(_04779_),
    .B(_04959_));
 sg13g2_or2_1 _13284_ (.X(_04961_),
    .B(_04960_),
    .A(_04957_));
 sg13g2_buf_2 _13285_ (.A(\am_sdr0.cic1.integ2[7] ),
    .X(_04962_));
 sg13g2_nand2b_1 _13286_ (.Y(_04963_),
    .B(_04959_),
    .A_N(_04962_));
 sg13g2_or2_1 _13287_ (.X(_04964_),
    .B(_04963_),
    .A(_04957_));
 sg13g2_nor3_1 _13288_ (.A(_04949_),
    .B(_04947_),
    .C(_04948_),
    .Y(_04965_));
 sg13g2_a221oi_1 _13289_ (.B2(_04964_),
    .C1(_04965_),
    .B1(_04961_),
    .A1(_04941_),
    .Y(_04966_),
    .A2(_04950_));
 sg13g2_buf_1 _13290_ (.A(_04966_),
    .X(_04967_));
 sg13g2_nor2_1 _13291_ (.A(_04962_),
    .B(net345),
    .Y(_04968_));
 sg13g2_inv_1 _13292_ (.Y(_04969_),
    .A(_04955_));
 sg13g2_nand2_1 _13293_ (.Y(_04970_),
    .A(_04951_),
    .B(_04763_));
 sg13g2_nor2_1 _13294_ (.A(_04953_),
    .B(_04770_),
    .Y(_04971_));
 sg13g2_a221oi_1 _13295_ (.B2(_04971_),
    .C1(_04952_),
    .B1(_04970_),
    .A1(_04969_),
    .Y(_04972_),
    .A2(_04768_));
 sg13g2_a221oi_1 _13296_ (.B2(_04963_),
    .C1(_04972_),
    .B1(_04960_),
    .A1(_04955_),
    .Y(_04973_),
    .A2(_04736_));
 sg13g2_a21o_1 _13297_ (.A2(_04968_),
    .A1(_04959_),
    .B1(_04973_),
    .X(_04974_));
 sg13g2_buf_1 _13298_ (.A(_04974_),
    .X(_04975_));
 sg13g2_nor2_1 _13299_ (.A(_04958_),
    .B(_04785_),
    .Y(_04976_));
 sg13g2_nor3_2 _13300_ (.A(_04967_),
    .B(_04975_),
    .C(_04976_),
    .Y(_04977_));
 sg13g2_buf_2 _13301_ (.A(\am_sdr0.cic1.integ2[9] ),
    .X(_04978_));
 sg13g2_a21o_1 _13302_ (.A2(_04977_),
    .A1(net344),
    .B1(_04978_),
    .X(_04979_));
 sg13g2_o21ai_1 _13303_ (.B1(_04979_),
    .Y(_04980_),
    .A1(net344),
    .A2(_04977_));
 sg13g2_xnor2_1 _13304_ (.Y(_04981_),
    .A(_04940_),
    .B(_04980_));
 sg13g2_nor2_1 _13305_ (.A(net99),
    .B(_04981_),
    .Y(_00549_));
 sg13g2_nor2_1 _13306_ (.A(_04939_),
    .B(_04797_),
    .Y(_04982_));
 sg13g2_nor2_1 _13307_ (.A(_04982_),
    .B(_04976_),
    .Y(_04983_));
 sg13g2_nand2_1 _13308_ (.Y(_04984_),
    .A(net344),
    .B(_04983_));
 sg13g2_nor3_1 _13309_ (.A(_04967_),
    .B(_04975_),
    .C(_04984_),
    .Y(_04985_));
 sg13g2_nand2_1 _13310_ (.Y(_04986_),
    .A(_04978_),
    .B(_04983_));
 sg13g2_nor3_1 _13311_ (.A(_04967_),
    .B(_04975_),
    .C(_04986_),
    .Y(_04987_));
 sg13g2_nand2_1 _13312_ (.Y(_04988_),
    .A(_04978_),
    .B(\am_sdr0.cic1.integ1[12] ));
 sg13g2_nand2_1 _13313_ (.Y(_04989_),
    .A(_04939_),
    .B(_04797_));
 sg13g2_o21ai_1 _13314_ (.B1(_04989_),
    .Y(_04990_),
    .A1(_04982_),
    .A2(_04988_));
 sg13g2_nor3_2 _13315_ (.A(_04985_),
    .B(_04987_),
    .C(_04990_),
    .Y(_04991_));
 sg13g2_buf_1 _13316_ (.A(\am_sdr0.cic1.integ2[11] ),
    .X(_04992_));
 sg13g2_xnor2_1 _13317_ (.Y(_04993_),
    .A(net340),
    .B(net343));
 sg13g2_xnor2_1 _13318_ (.Y(_04994_),
    .A(_04991_),
    .B(_04993_));
 sg13g2_nor2_1 _13319_ (.A(net99),
    .B(_04994_),
    .Y(_00550_));
 sg13g2_buf_1 _13320_ (.A(\am_sdr0.cic1.integ2[12] ),
    .X(_04995_));
 sg13g2_nand2_1 _13321_ (.Y(_04996_),
    .A(_04995_),
    .B(net342));
 sg13g2_or2_1 _13322_ (.X(_04997_),
    .B(net342),
    .A(_04995_));
 sg13g2_buf_1 _13323_ (.A(_04997_),
    .X(_04998_));
 sg13g2_nand2_1 _13324_ (.Y(_04999_),
    .A(_04996_),
    .B(_04998_));
 sg13g2_nor2_1 _13325_ (.A(net340),
    .B(net343),
    .Y(_05000_));
 sg13g2_nand2_1 _13326_ (.Y(_05001_),
    .A(net340),
    .B(net343));
 sg13g2_o21ai_1 _13327_ (.B1(_05001_),
    .Y(_05002_),
    .A1(_04991_),
    .A2(_05000_));
 sg13g2_xor2_1 _13328_ (.B(_05002_),
    .A(_04999_),
    .X(_05003_));
 sg13g2_nor2_1 _13329_ (.A(net99),
    .B(_05003_),
    .Y(_00551_));
 sg13g2_and2_1 _13330_ (.A(_04995_),
    .B(_04818_),
    .X(_05004_));
 sg13g2_buf_1 _13331_ (.A(_05004_),
    .X(_05005_));
 sg13g2_a21o_1 _13332_ (.A2(_05002_),
    .A1(_04998_),
    .B1(_05005_),
    .X(_05006_));
 sg13g2_buf_1 _13333_ (.A(_05006_),
    .X(_05007_));
 sg13g2_buf_2 _13334_ (.A(\am_sdr0.cic1.integ2[13] ),
    .X(_05008_));
 sg13g2_xor2_1 _13335_ (.B(net289),
    .A(_05008_),
    .X(_05009_));
 sg13g2_xnor2_1 _13336_ (.Y(_05010_),
    .A(_05007_),
    .B(_05009_));
 sg13g2_nor2_1 _13337_ (.A(net99),
    .B(_05010_),
    .Y(_00552_));
 sg13g2_nor3_1 _13338_ (.A(_04802_),
    .B(_04829_),
    .C(_05005_),
    .Y(_05011_));
 sg13g2_nor3_1 _13339_ (.A(net340),
    .B(_04829_),
    .C(_05005_),
    .Y(_05012_));
 sg13g2_o21ai_1 _13340_ (.B1(_04991_),
    .Y(_05013_),
    .A1(_05011_),
    .A2(_05012_));
 sg13g2_nand2_1 _13341_ (.Y(_05014_),
    .A(_04996_),
    .B(_05000_));
 sg13g2_a21o_1 _13342_ (.A2(_05014_),
    .A1(_04998_),
    .B1(_04829_),
    .X(_05015_));
 sg13g2_and3_1 _13343_ (.X(_05016_),
    .A(_05008_),
    .B(_05013_),
    .C(_05015_));
 sg13g2_a21oi_1 _13344_ (.A1(_04830_),
    .A2(_05007_),
    .Y(_05017_),
    .B1(_05016_));
 sg13g2_buf_2 _13345_ (.A(\am_sdr0.cic1.integ2[14] ),
    .X(_05018_));
 sg13g2_xnor2_1 _13346_ (.Y(_05019_),
    .A(_05018_),
    .B(net341));
 sg13g2_xnor2_1 _13347_ (.Y(_05020_),
    .A(_05017_),
    .B(_05019_));
 sg13g2_nor2_1 _13348_ (.A(_04928_),
    .B(_05020_),
    .Y(_00553_));
 sg13g2_nand2_1 _13349_ (.Y(_05021_),
    .A(_05013_),
    .B(_05015_));
 sg13g2_nand2_1 _13350_ (.Y(_05022_),
    .A(_05018_),
    .B(\am_sdr0.cic1.integ1[17] ));
 sg13g2_a21oi_1 _13351_ (.A1(_05018_),
    .A2(_04839_),
    .Y(_05023_),
    .B1(_05008_));
 sg13g2_nand2_1 _13352_ (.Y(_05024_),
    .A(_04830_),
    .B(_05007_));
 sg13g2_a22oi_1 _13353_ (.Y(_05025_),
    .B1(_05023_),
    .B2(_05024_),
    .A2(_05022_),
    .A1(_05021_));
 sg13g2_o21ai_1 _13354_ (.B1(_05025_),
    .Y(_05026_),
    .A1(_05018_),
    .A2(_04839_));
 sg13g2_buf_2 _13355_ (.A(\am_sdr0.cic1.integ2[15] ),
    .X(_05027_));
 sg13g2_xnor2_1 _13356_ (.Y(_05028_),
    .A(_05027_),
    .B(_04843_));
 sg13g2_xnor2_1 _13357_ (.Y(_05029_),
    .A(_05026_),
    .B(_05028_));
 sg13g2_nor2_1 _13358_ (.A(_04928_),
    .B(_05029_),
    .Y(_00554_));
 sg13g2_buf_2 _13359_ (.A(\am_sdr0.cic1.integ2[16] ),
    .X(_05030_));
 sg13g2_xnor2_1 _13360_ (.Y(_05031_),
    .A(_05030_),
    .B(_04857_));
 sg13g2_nor2_1 _13361_ (.A(_05027_),
    .B(_04843_),
    .Y(_05032_));
 sg13g2_nand2_1 _13362_ (.Y(_05033_),
    .A(_05027_),
    .B(_04843_));
 sg13g2_o21ai_1 _13363_ (.B1(_05033_),
    .Y(_05034_),
    .A1(_05026_),
    .A2(_05032_));
 sg13g2_xnor2_1 _13364_ (.Y(_05035_),
    .A(_05031_),
    .B(_05034_));
 sg13g2_and2_1 _13365_ (.A(net246),
    .B(_05035_),
    .X(_00555_));
 sg13g2_buf_1 _13366_ (.A(_03962_),
    .X(_05036_));
 sg13g2_a21o_1 _13367_ (.A2(_04858_),
    .A1(_05030_),
    .B1(_05034_),
    .X(_05037_));
 sg13g2_o21ai_1 _13368_ (.B1(_05037_),
    .Y(_05038_),
    .A1(_05030_),
    .A2(_04858_));
 sg13g2_buf_2 _13369_ (.A(\am_sdr0.cic1.integ2[17] ),
    .X(_05039_));
 sg13g2_xnor2_1 _13370_ (.Y(_05040_),
    .A(_05039_),
    .B(_04869_));
 sg13g2_xnor2_1 _13371_ (.Y(_05041_),
    .A(_05038_),
    .B(_05040_));
 sg13g2_nor2_1 _13372_ (.A(net98),
    .B(_05041_),
    .Y(_00556_));
 sg13g2_buf_2 _13373_ (.A(\am_sdr0.cic1.integ2[18] ),
    .X(_05042_));
 sg13g2_xor2_1 _13374_ (.B(_04875_),
    .A(_05042_),
    .X(_05043_));
 sg13g2_or4_1 _13375_ (.A(_05019_),
    .B(_05028_),
    .C(_05031_),
    .D(_05040_),
    .X(_05044_));
 sg13g2_nand2_1 _13376_ (.Y(_05045_),
    .A(_05039_),
    .B(net287));
 sg13g2_o21ai_1 _13377_ (.B1(_05033_),
    .Y(_05046_),
    .A1(_05022_),
    .A2(_05032_));
 sg13g2_nand2_1 _13378_ (.Y(_05047_),
    .A(_04857_),
    .B(_05046_));
 sg13g2_o21ai_1 _13379_ (.B1(_05030_),
    .Y(_05048_),
    .A1(_04857_),
    .A2(_05046_));
 sg13g2_nand3_1 _13380_ (.B(_05047_),
    .C(_05048_),
    .A(_05045_),
    .Y(_05049_));
 sg13g2_o21ai_1 _13381_ (.B1(_05049_),
    .Y(_05050_),
    .A1(_05039_),
    .A2(net287));
 sg13g2_o21ai_1 _13382_ (.B1(_05050_),
    .Y(_05051_),
    .A1(_05017_),
    .A2(_05044_));
 sg13g2_xnor2_1 _13383_ (.Y(_05052_),
    .A(_05043_),
    .B(_05051_));
 sg13g2_nor2_1 _13384_ (.A(net98),
    .B(_05052_),
    .Y(_00557_));
 sg13g2_inv_1 _13385_ (.Y(_05053_),
    .A(_05042_));
 sg13g2_a21oi_1 _13386_ (.A1(_05042_),
    .A2(_04875_),
    .Y(_05054_),
    .B1(_05051_));
 sg13g2_a21oi_2 _13387_ (.B1(_05054_),
    .Y(_05055_),
    .A2(_04890_),
    .A1(_05053_));
 sg13g2_buf_2 _13388_ (.A(\am_sdr0.cic1.integ2[19] ),
    .X(_05056_));
 sg13g2_xor2_1 _13389_ (.B(_04881_),
    .A(_05056_),
    .X(_05057_));
 sg13g2_xnor2_1 _13390_ (.Y(_05058_),
    .A(_05055_),
    .B(_05057_));
 sg13g2_nor2_1 _13391_ (.A(net98),
    .B(_05058_),
    .Y(_00558_));
 sg13g2_xor2_1 _13392_ (.B(\am_sdr0.cic1.integ2[1] ),
    .A(_04740_),
    .X(_05059_));
 sg13g2_xnor2_1 _13393_ (.Y(_05060_),
    .A(_04944_),
    .B(_05059_));
 sg13g2_nor2_1 _13394_ (.A(_05036_),
    .B(_05060_),
    .Y(_00559_));
 sg13g2_buf_2 _13395_ (.A(\am_sdr0.cic1.integ2[20] ),
    .X(_05061_));
 sg13g2_xor2_1 _13396_ (.B(_04888_),
    .A(_05061_),
    .X(_05062_));
 sg13g2_inv_1 _13397_ (.Y(_05063_),
    .A(_05056_));
 sg13g2_o21ai_1 _13398_ (.B1(_05055_),
    .Y(_05064_),
    .A1(_05056_),
    .A2(_04881_));
 sg13g2_o21ai_1 _13399_ (.B1(_05064_),
    .Y(_05065_),
    .A1(_05063_),
    .A2(_04882_));
 sg13g2_xnor2_1 _13400_ (.Y(_05066_),
    .A(_05062_),
    .B(_05065_));
 sg13g2_nor2_1 _13401_ (.A(net98),
    .B(_05066_),
    .Y(_00560_));
 sg13g2_o21ai_1 _13402_ (.B1(_04881_),
    .Y(_05067_),
    .A1(_05061_),
    .A2(_04888_));
 sg13g2_inv_1 _13403_ (.Y(_05068_),
    .A(_05067_));
 sg13g2_nor2_1 _13404_ (.A(_04875_),
    .B(_04881_),
    .Y(_05069_));
 sg13g2_o21ai_1 _13405_ (.B1(_05056_),
    .Y(_05070_),
    .A1(_05061_),
    .A2(_04888_));
 sg13g2_a221oi_1 _13406_ (.B2(_04882_),
    .C1(_05070_),
    .B1(_05054_),
    .A1(_05053_),
    .Y(_05071_),
    .A2(_05069_));
 sg13g2_a221oi_1 _13407_ (.B2(_05068_),
    .C1(_05071_),
    .B1(_05055_),
    .A1(_05061_),
    .Y(_05072_),
    .A2(_04888_));
 sg13g2_buf_2 _13408_ (.A(\am_sdr0.cic1.integ2[21] ),
    .X(_05073_));
 sg13g2_xnor2_1 _13409_ (.Y(_05074_),
    .A(_05073_),
    .B(_04896_));
 sg13g2_xnor2_1 _13410_ (.Y(_05075_),
    .A(_05072_),
    .B(_05074_));
 sg13g2_nor2_1 _13411_ (.A(_05036_),
    .B(_05075_),
    .Y(_00561_));
 sg13g2_xor2_1 _13412_ (.B(\am_sdr0.cic1.integ1[25] ),
    .A(\am_sdr0.cic1.integ2[22] ),
    .X(_05076_));
 sg13g2_nand2_1 _13413_ (.Y(_05077_),
    .A(_05073_),
    .B(_04896_));
 sg13g2_nor2_1 _13414_ (.A(_05073_),
    .B(_04896_),
    .Y(_05078_));
 sg13g2_a21oi_1 _13415_ (.A1(_05072_),
    .A2(_05077_),
    .Y(_05079_),
    .B1(_05078_));
 sg13g2_xnor2_1 _13416_ (.Y(_05080_),
    .A(_05076_),
    .B(_05079_));
 sg13g2_nor2_1 _13417_ (.A(net98),
    .B(_05080_),
    .Y(_00562_));
 sg13g2_a21o_1 _13418_ (.A2(_04944_),
    .A1(_04942_),
    .B1(_04945_),
    .X(_05081_));
 sg13g2_xor2_1 _13419_ (.B(\am_sdr0.cic1.integ2[2] ),
    .A(_04738_),
    .X(_05082_));
 sg13g2_xnor2_1 _13420_ (.Y(_05083_),
    .A(_05081_),
    .B(_05082_));
 sg13g2_nor2_1 _13421_ (.A(net98),
    .B(_05083_),
    .Y(_00563_));
 sg13g2_nor2_1 _13422_ (.A(_04947_),
    .B(_04948_),
    .Y(_05084_));
 sg13g2_xor2_1 _13423_ (.B(_04737_),
    .A(_04941_),
    .X(_05085_));
 sg13g2_xnor2_1 _13424_ (.Y(_05086_),
    .A(_05084_),
    .B(_05085_));
 sg13g2_nor2_1 _13425_ (.A(net98),
    .B(_05086_),
    .Y(_00564_));
 sg13g2_a21o_1 _13426_ (.A2(_04950_),
    .A1(_04941_),
    .B1(_04965_),
    .X(_05087_));
 sg13g2_buf_1 _13427_ (.A(_05087_),
    .X(_05088_));
 sg13g2_xor2_1 _13428_ (.B(_04770_),
    .A(_04953_),
    .X(_05089_));
 sg13g2_xnor2_1 _13429_ (.Y(_05090_),
    .A(_05088_),
    .B(_05089_));
 sg13g2_nor2_1 _13430_ (.A(net98),
    .B(_05090_),
    .Y(_00565_));
 sg13g2_buf_1 _13431_ (.A(_03962_),
    .X(_05091_));
 sg13g2_a21oi_1 _13432_ (.A1(_04770_),
    .A2(_05088_),
    .Y(_05092_),
    .B1(_04953_));
 sg13g2_nor2_1 _13433_ (.A(_04770_),
    .B(_05088_),
    .Y(_05093_));
 sg13g2_nor2_1 _13434_ (.A(_05092_),
    .B(_05093_),
    .Y(_05094_));
 sg13g2_xor2_1 _13435_ (.B(_04763_),
    .A(_04951_),
    .X(_05095_));
 sg13g2_xnor2_1 _13436_ (.Y(_05096_),
    .A(_05094_),
    .B(_05095_));
 sg13g2_nor2_1 _13437_ (.A(net97),
    .B(_05096_),
    .Y(_00566_));
 sg13g2_xor2_1 _13438_ (.B(_04736_),
    .A(_04955_),
    .X(_05097_));
 sg13g2_nand2b_1 _13439_ (.Y(_05098_),
    .B(_05094_),
    .A_N(_04952_));
 sg13g2_nand2_1 _13440_ (.Y(_05099_),
    .A(_04970_),
    .B(_05098_));
 sg13g2_xnor2_1 _13441_ (.Y(_05100_),
    .A(_05097_),
    .B(_05099_));
 sg13g2_nor2_1 _13442_ (.A(net97),
    .B(_05100_),
    .Y(_00567_));
 sg13g2_a21oi_1 _13443_ (.A1(_04955_),
    .A2(_04736_),
    .Y(_05101_),
    .B1(_04972_));
 sg13g2_nor2_1 _13444_ (.A(_05088_),
    .B(_04957_),
    .Y(_05102_));
 sg13g2_or2_1 _13445_ (.X(_05103_),
    .B(_05102_),
    .A(_05101_));
 sg13g2_xnor2_1 _13446_ (.Y(_05104_),
    .A(_04962_),
    .B(net345));
 sg13g2_xnor2_1 _13447_ (.Y(_05105_),
    .A(_05103_),
    .B(_05104_));
 sg13g2_nor2_1 _13448_ (.A(net97),
    .B(_05105_),
    .Y(_00568_));
 sg13g2_nor2_1 _13449_ (.A(_05103_),
    .B(_04968_),
    .Y(_05106_));
 sg13g2_a21oi_1 _13450_ (.A1(_04962_),
    .A2(net345),
    .Y(_05107_),
    .B1(_05106_));
 sg13g2_xnor2_1 _13451_ (.Y(_05108_),
    .A(_04958_),
    .B(_04785_));
 sg13g2_xnor2_1 _13452_ (.Y(_05109_),
    .A(_05107_),
    .B(_05108_));
 sg13g2_nor2_1 _13453_ (.A(net97),
    .B(_05109_),
    .Y(_00569_));
 sg13g2_xor2_1 _13454_ (.B(net344),
    .A(_04978_),
    .X(_05110_));
 sg13g2_xnor2_1 _13455_ (.Y(_05111_),
    .A(_04977_),
    .B(_05110_));
 sg13g2_nor2_1 _13456_ (.A(net97),
    .B(_05111_),
    .Y(_00570_));
 sg13g2_xnor2_1 _13457_ (.Y(_05112_),
    .A(_04941_),
    .B(_02297_));
 sg13g2_nor2_1 _13458_ (.A(net97),
    .B(_05112_),
    .Y(_00571_));
 sg13g2_nor2_1 _13459_ (.A(_04995_),
    .B(_02361_),
    .Y(_05113_));
 sg13g2_inv_1 _13460_ (.Y(_05114_),
    .A(_04939_));
 sg13g2_inv_1 _13461_ (.Y(_05115_),
    .A(_04958_));
 sg13g2_nor2_1 _13462_ (.A(_04962_),
    .B(_02343_),
    .Y(_05116_));
 sg13g2_o21ai_1 _13463_ (.B1(_05116_),
    .Y(_05117_),
    .A1(_05115_),
    .A2(_02347_));
 sg13g2_o21ai_1 _13464_ (.B1(_05117_),
    .Y(_05118_),
    .A1(_04958_),
    .A2(\am_sdr0.cic1.integ3[5] ));
 sg13g2_nand2_1 _13465_ (.Y(_05119_),
    .A(_04951_),
    .B(_02338_));
 sg13g2_nor2_1 _13466_ (.A(_04951_),
    .B(_02338_),
    .Y(_05120_));
 sg13g2_nor2_1 _13467_ (.A(_04953_),
    .B(_02335_),
    .Y(_05121_));
 sg13g2_a22oi_1 _13468_ (.Y(_05122_),
    .B1(_04953_),
    .B2(_02335_),
    .A2(_02297_),
    .A1(_04941_));
 sg13g2_or3_1 _13469_ (.A(_05120_),
    .B(_05121_),
    .C(_05122_),
    .X(_05123_));
 sg13g2_buf_1 _13470_ (.A(_05123_),
    .X(_05124_));
 sg13g2_nand3_1 _13471_ (.B(_05119_),
    .C(_05124_),
    .A(_02340_),
    .Y(_05125_));
 sg13g2_or2_1 _13472_ (.X(_05126_),
    .B(_04958_),
    .A(_04962_));
 sg13g2_nand2_1 _13473_ (.Y(_05127_),
    .A(_04962_),
    .B(_02343_));
 sg13g2_a22oi_1 _13474_ (.Y(_05128_),
    .B1(_02347_),
    .B2(_05127_),
    .A2(_05115_),
    .A1(_02344_));
 sg13g2_a21oi_1 _13475_ (.A1(_05119_),
    .A2(_05124_),
    .Y(_05129_),
    .B1(_02340_));
 sg13g2_a221oi_1 _13476_ (.B2(_05128_),
    .C1(_05129_),
    .B1(_05126_),
    .A1(_04955_),
    .Y(_05130_),
    .A2(_05125_));
 sg13g2_nor2_1 _13477_ (.A(_04978_),
    .B(_02350_),
    .Y(_05131_));
 sg13g2_or3_1 _13478_ (.A(_05118_),
    .B(_05130_),
    .C(_05131_),
    .X(_05132_));
 sg13g2_buf_1 _13479_ (.A(_05132_),
    .X(_05133_));
 sg13g2_a22oi_1 _13480_ (.Y(_05134_),
    .B1(_04939_),
    .B2(\am_sdr0.cic1.integ3[7] ),
    .A2(_02350_),
    .A1(_04978_));
 sg13g2_a22oi_1 _13481_ (.Y(_05135_),
    .B1(_05133_),
    .B2(_05134_),
    .A2(_02352_),
    .A1(_05114_));
 sg13g2_buf_1 _13482_ (.A(_05135_),
    .X(_05136_));
 sg13g2_or2_1 _13483_ (.X(_05137_),
    .B(_02357_),
    .A(net340));
 sg13g2_and2_1 _13484_ (.A(net340),
    .B(_02357_),
    .X(_05138_));
 sg13g2_a21oi_1 _13485_ (.A1(_05136_),
    .A2(_05137_),
    .Y(_05139_),
    .B1(_05138_));
 sg13g2_nand2_1 _13486_ (.Y(_05140_),
    .A(_04995_),
    .B(_02361_));
 sg13g2_o21ai_1 _13487_ (.B1(_05140_),
    .Y(_05141_),
    .A1(_05113_),
    .A2(_05139_));
 sg13g2_xor2_1 _13488_ (.B(_02308_),
    .A(_05008_),
    .X(_05142_));
 sg13g2_xnor2_1 _13489_ (.Y(_05143_),
    .A(_05141_),
    .B(_05142_));
 sg13g2_nor2_1 _13490_ (.A(_05091_),
    .B(_05143_),
    .Y(_00572_));
 sg13g2_inv_1 _13491_ (.Y(_05144_),
    .A(_05008_));
 sg13g2_or2_1 _13492_ (.X(_05145_),
    .B(_02308_),
    .A(_02357_));
 sg13g2_or2_1 _13493_ (.X(_05146_),
    .B(_02308_),
    .A(net340));
 sg13g2_a221oi_1 _13494_ (.B2(_05146_),
    .C1(_05136_),
    .B1(_05145_),
    .A1(_04995_),
    .Y(_05147_),
    .A2(_02361_));
 sg13g2_or2_1 _13495_ (.X(_05148_),
    .B(_02361_),
    .A(_04995_));
 sg13g2_buf_1 _13496_ (.A(_05148_),
    .X(_05149_));
 sg13g2_nand2b_1 _13497_ (.Y(_05150_),
    .B(_05140_),
    .A_N(_05137_));
 sg13g2_a21oi_1 _13498_ (.A1(_05149_),
    .A2(_05150_),
    .Y(_05151_),
    .B1(_02308_));
 sg13g2_nor3_1 _13499_ (.A(_05144_),
    .B(_05147_),
    .C(_05151_),
    .Y(_05152_));
 sg13g2_a21o_1 _13500_ (.A2(_05141_),
    .A1(_02308_),
    .B1(_05152_),
    .X(_05153_));
 sg13g2_xor2_1 _13501_ (.B(_02313_),
    .A(_05018_),
    .X(_05154_));
 sg13g2_xnor2_1 _13502_ (.Y(_05155_),
    .A(_05153_),
    .B(_05154_));
 sg13g2_nor2_1 _13503_ (.A(net97),
    .B(_05155_),
    .Y(_00573_));
 sg13g2_and2_1 _13504_ (.A(_05027_),
    .B(_02317_),
    .X(_05156_));
 sg13g2_or2_1 _13505_ (.X(_05157_),
    .B(_02317_),
    .A(_05027_));
 sg13g2_nand2b_1 _13506_ (.Y(_05158_),
    .B(_05157_),
    .A_N(_05156_));
 sg13g2_inv_1 _13507_ (.Y(_05159_),
    .A(_05018_));
 sg13g2_o21ai_1 _13508_ (.B1(_05153_),
    .Y(_05160_),
    .A1(_05018_),
    .A2(_02313_));
 sg13g2_o21ai_1 _13509_ (.B1(_05160_),
    .Y(_05161_),
    .A1(_05159_),
    .A2(_02314_));
 sg13g2_xnor2_1 _13510_ (.Y(_05162_),
    .A(_05158_),
    .B(_05161_));
 sg13g2_and2_1 _13511_ (.A(net246),
    .B(_05162_),
    .X(_00574_));
 sg13g2_a21oi_1 _13512_ (.A1(_05157_),
    .A2(_05161_),
    .Y(_05163_),
    .B1(_05156_));
 sg13g2_xor2_1 _13513_ (.B(_02321_),
    .A(_05030_),
    .X(_05164_));
 sg13g2_xnor2_1 _13514_ (.Y(_05165_),
    .A(_05163_),
    .B(_05164_));
 sg13g2_and2_1 _13515_ (.A(net246),
    .B(_05165_),
    .X(_00575_));
 sg13g2_xnor2_1 _13516_ (.Y(_05166_),
    .A(_05039_),
    .B(_02323_));
 sg13g2_nor2_1 _13517_ (.A(_05030_),
    .B(_02321_),
    .Y(_05167_));
 sg13g2_nand2_1 _13518_ (.Y(_05168_),
    .A(_05030_),
    .B(_02321_));
 sg13g2_o21ai_1 _13519_ (.B1(_05168_),
    .Y(_05169_),
    .A1(_05163_),
    .A2(_05167_));
 sg13g2_xnor2_1 _13520_ (.Y(_05170_),
    .A(_05166_),
    .B(_05169_));
 sg13g2_and2_1 _13521_ (.A(net246),
    .B(_05170_),
    .X(_00576_));
 sg13g2_nor2_1 _13522_ (.A(_05039_),
    .B(_02323_),
    .Y(_05171_));
 sg13g2_nand3_1 _13523_ (.B(_02308_),
    .C(_05149_),
    .A(_02357_),
    .Y(_05172_));
 sg13g2_a221oi_1 _13524_ (.B2(_05134_),
    .C1(_05172_),
    .B1(_05133_),
    .A1(_05114_),
    .Y(_05173_),
    .A2(_02352_));
 sg13g2_nand3_1 _13525_ (.B(_02308_),
    .C(_05149_),
    .A(net340),
    .Y(_05174_));
 sg13g2_a221oi_1 _13526_ (.B2(_05134_),
    .C1(_05174_),
    .B1(_05133_),
    .A1(_05114_),
    .Y(_05175_),
    .A2(_02352_));
 sg13g2_nand2_1 _13527_ (.Y(_05176_),
    .A(_05149_),
    .B(_05138_));
 sg13g2_a21oi_1 _13528_ (.A1(_05140_),
    .A2(_05176_),
    .Y(_05177_),
    .B1(_02309_));
 sg13g2_nor3_1 _13529_ (.A(_05173_),
    .B(_05175_),
    .C(_05177_),
    .Y(_05178_));
 sg13g2_o21ai_1 _13530_ (.B1(_05178_),
    .Y(_05179_),
    .A1(_02314_),
    .A2(_02318_));
 sg13g2_or2_1 _13531_ (.X(_05180_),
    .B(_05179_),
    .A(_05152_));
 sg13g2_nor2_1 _13532_ (.A(_05027_),
    .B(_02317_),
    .Y(_05181_));
 sg13g2_nor2_1 _13533_ (.A(_05159_),
    .B(_05181_),
    .Y(_05182_));
 sg13g2_a21oi_1 _13534_ (.A1(_05018_),
    .A2(_02313_),
    .Y(_05183_),
    .B1(_02317_));
 sg13g2_nand2b_1 _13535_ (.Y(_05184_),
    .B(_05027_),
    .A_N(_05183_));
 sg13g2_nand2_1 _13536_ (.Y(_05185_),
    .A(_05039_),
    .B(_02323_));
 sg13g2_nand3b_1 _13537_ (.B(_05184_),
    .C(_05185_),
    .Y(_05186_),
    .A_N(_02321_));
 sg13g2_nand3b_1 _13538_ (.B(_05184_),
    .C(_05185_),
    .Y(_05187_),
    .A_N(_05030_));
 sg13g2_nand2_1 _13539_ (.Y(_05188_),
    .A(_05008_),
    .B(_02313_));
 sg13g2_nor4_1 _13540_ (.A(_05147_),
    .B(_05151_),
    .C(_05181_),
    .D(_05188_),
    .Y(_05189_));
 sg13g2_nor3_1 _13541_ (.A(_02314_),
    .B(_05178_),
    .C(_05181_),
    .Y(_05190_));
 sg13g2_or2_1 _13542_ (.X(_05191_),
    .B(_05190_),
    .A(_05189_));
 sg13g2_a221oi_1 _13543_ (.B2(_05187_),
    .C1(_05191_),
    .B1(_05186_),
    .A1(_05180_),
    .Y(_05192_),
    .A2(_05182_));
 sg13g2_and2_1 _13544_ (.A(_05185_),
    .B(_05167_),
    .X(_05193_));
 sg13g2_nor3_1 _13545_ (.A(_05171_),
    .B(_05192_),
    .C(_05193_),
    .Y(_05194_));
 sg13g2_xor2_1 _13546_ (.B(_02327_),
    .A(_05042_),
    .X(_05195_));
 sg13g2_xnor2_1 _13547_ (.Y(_05196_),
    .A(_05194_),
    .B(_05195_));
 sg13g2_nor2_1 _13548_ (.A(_05091_),
    .B(_05196_),
    .Y(_00577_));
 sg13g2_xor2_1 _13549_ (.B(_02329_),
    .A(_05056_),
    .X(_05197_));
 sg13g2_nor2_1 _13550_ (.A(_05042_),
    .B(_02327_),
    .Y(_05198_));
 sg13g2_or4_1 _13551_ (.A(_05171_),
    .B(_05192_),
    .C(_05193_),
    .D(_05198_),
    .X(_05199_));
 sg13g2_nand2_1 _13552_ (.Y(_05200_),
    .A(_05042_),
    .B(_02327_));
 sg13g2_nand2_1 _13553_ (.Y(_05201_),
    .A(_05199_),
    .B(_05200_));
 sg13g2_xnor2_1 _13554_ (.Y(_05202_),
    .A(_05197_),
    .B(_05201_));
 sg13g2_nor2_1 _13555_ (.A(net97),
    .B(_05202_),
    .Y(_00578_));
 sg13g2_buf_1 _13556_ (.A(net259),
    .X(_05203_));
 sg13g2_buf_1 _13557_ (.A(_05203_),
    .X(_05204_));
 sg13g2_nor2_1 _13558_ (.A(_05056_),
    .B(_02329_),
    .Y(_05205_));
 sg13g2_nand2_1 _13559_ (.Y(_05206_),
    .A(_05056_),
    .B(_02329_));
 sg13g2_nand3_1 _13560_ (.B(_05199_),
    .C(_05200_),
    .A(_05206_),
    .Y(_05207_));
 sg13g2_nor2b_1 _13561_ (.A(_05205_),
    .B_N(_05207_),
    .Y(_05208_));
 sg13g2_xor2_1 _13562_ (.B(_02331_),
    .A(_05061_),
    .X(_05209_));
 sg13g2_xnor2_1 _13563_ (.Y(_05210_),
    .A(_05208_),
    .B(_05209_));
 sg13g2_nor2_1 _13564_ (.A(_05204_),
    .B(_05210_),
    .Y(_00579_));
 sg13g2_xnor2_1 _13565_ (.Y(_05211_),
    .A(_05073_),
    .B(_02333_));
 sg13g2_or2_1 _13566_ (.X(_05212_),
    .B(_02331_),
    .A(_05061_));
 sg13g2_and2_1 _13567_ (.A(_05061_),
    .B(_02331_),
    .X(_05213_));
 sg13g2_a21oi_1 _13568_ (.A1(_05208_),
    .A2(_05212_),
    .Y(_05214_),
    .B1(_05213_));
 sg13g2_xnor2_1 _13569_ (.Y(_05215_),
    .A(_05211_),
    .B(_05214_));
 sg13g2_nor2_1 _13570_ (.A(_05204_),
    .B(_05215_),
    .Y(_00580_));
 sg13g2_xor2_1 _13571_ (.B(\am_sdr0.cic1.integ3[19] ),
    .A(\am_sdr0.cic1.integ2[22] ),
    .X(_05216_));
 sg13g2_and2_1 _13572_ (.A(net297),
    .B(_05216_),
    .X(_05217_));
 sg13g2_nor2_1 _13573_ (.A(net251),
    .B(_05216_),
    .Y(_05218_));
 sg13g2_nand2_1 _13574_ (.Y(_05219_),
    .A(_05073_),
    .B(_02333_));
 sg13g2_nor2_1 _13575_ (.A(_05073_),
    .B(_02333_),
    .Y(_05220_));
 sg13g2_a21oi_1 _13576_ (.A1(_05219_),
    .A2(_05214_),
    .Y(_05221_),
    .B1(_05220_));
 sg13g2_mux2_1 _13577_ (.A0(_05217_),
    .A1(_05218_),
    .S(_05221_),
    .X(_00581_));
 sg13g2_nand2_1 _13578_ (.Y(_05222_),
    .A(_04941_),
    .B(_02297_));
 sg13g2_xnor2_1 _13579_ (.Y(_05223_),
    .A(_04953_),
    .B(_02335_));
 sg13g2_xnor2_1 _13580_ (.Y(_05224_),
    .A(_05222_),
    .B(_05223_));
 sg13g2_nor2_1 _13581_ (.A(net96),
    .B(_05224_),
    .Y(_00582_));
 sg13g2_nor2_1 _13582_ (.A(_05121_),
    .B(_05122_),
    .Y(_05225_));
 sg13g2_xor2_1 _13583_ (.B(_02338_),
    .A(_04951_),
    .X(_05226_));
 sg13g2_xnor2_1 _13584_ (.Y(_05227_),
    .A(_05225_),
    .B(_05226_));
 sg13g2_nor2_1 _13585_ (.A(net96),
    .B(_05227_),
    .Y(_00583_));
 sg13g2_nand2_1 _13586_ (.Y(_05228_),
    .A(_05119_),
    .B(_05124_));
 sg13g2_xor2_1 _13587_ (.B(\am_sdr0.cic1.integ3[3] ),
    .A(_04955_),
    .X(_05229_));
 sg13g2_xnor2_1 _13588_ (.Y(_05230_),
    .A(_05228_),
    .B(_05229_));
 sg13g2_nor2_1 _13589_ (.A(net96),
    .B(_05230_),
    .Y(_00584_));
 sg13g2_a21oi_1 _13590_ (.A1(_04955_),
    .A2(_05125_),
    .Y(_05231_),
    .B1(_05129_));
 sg13g2_xnor2_1 _13591_ (.Y(_05232_),
    .A(_04962_),
    .B(_02343_));
 sg13g2_xnor2_1 _13592_ (.Y(_05233_),
    .A(_05231_),
    .B(_05232_));
 sg13g2_nor2_1 _13593_ (.A(net96),
    .B(_05233_),
    .Y(_00585_));
 sg13g2_xor2_1 _13594_ (.B(\am_sdr0.cic1.integ3[5] ),
    .A(_04958_),
    .X(_05234_));
 sg13g2_o21ai_1 _13595_ (.B1(_05127_),
    .Y(_05235_),
    .A1(_05116_),
    .A2(_05231_));
 sg13g2_xnor2_1 _13596_ (.Y(_05236_),
    .A(_05234_),
    .B(_05235_));
 sg13g2_nor2_1 _13597_ (.A(net96),
    .B(_05236_),
    .Y(_00586_));
 sg13g2_nor2_1 _13598_ (.A(_05118_),
    .B(_05130_),
    .Y(_05237_));
 sg13g2_xor2_1 _13599_ (.B(_02350_),
    .A(_04978_),
    .X(_05238_));
 sg13g2_xnor2_1 _13600_ (.Y(_05239_),
    .A(_05237_),
    .B(_05238_));
 sg13g2_nor2_1 _13601_ (.A(net96),
    .B(_05239_),
    .Y(_00587_));
 sg13g2_nand2_1 _13602_ (.Y(_05240_),
    .A(_04978_),
    .B(_02350_));
 sg13g2_nand2_1 _13603_ (.Y(_05241_),
    .A(_05133_),
    .B(_05240_));
 sg13g2_xor2_1 _13604_ (.B(\am_sdr0.cic1.integ3[7] ),
    .A(_04939_),
    .X(_05242_));
 sg13g2_xnor2_1 _13605_ (.Y(_05243_),
    .A(_05241_),
    .B(_05242_));
 sg13g2_nor2_1 _13606_ (.A(net96),
    .B(_05243_),
    .Y(_00588_));
 sg13g2_xor2_1 _13607_ (.B(_02357_),
    .A(_04992_),
    .X(_05244_));
 sg13g2_xnor2_1 _13608_ (.Y(_05245_),
    .A(_05136_),
    .B(_05244_));
 sg13g2_nor2_1 _13609_ (.A(net96),
    .B(_05245_),
    .Y(_00589_));
 sg13g2_buf_1 _13610_ (.A(_05203_),
    .X(_05246_));
 sg13g2_nand2_1 _13611_ (.Y(_05247_),
    .A(_05149_),
    .B(_05140_));
 sg13g2_xnor2_1 _13612_ (.Y(_05248_),
    .A(_05139_),
    .B(_05247_));
 sg13g2_nor2_1 _13613_ (.A(_05246_),
    .B(_05248_),
    .Y(_00590_));
 sg13g2_nand2_1 _13614_ (.Y(_05249_),
    .A(net240),
    .B(\am_sdr0.cic1.comb3[14] ));
 sg13g2_buf_1 _13615_ (.A(\am_sdr0.cic1.x_out[10] ),
    .X(_05250_));
 sg13g2_nand2_1 _13616_ (.Y(_05251_),
    .A(_05250_),
    .B(net156));
 sg13g2_a21oi_1 _13617_ (.A1(_05249_),
    .A2(_05251_),
    .Y(_00613_),
    .B1(net101));
 sg13g2_nand2_1 _13618_ (.Y(_05252_),
    .A(net240),
    .B(\am_sdr0.cic1.comb3[15] ));
 sg13g2_nand2_1 _13619_ (.Y(_05253_),
    .A(\am_sdr0.cic1.x_out[11] ),
    .B(net156));
 sg13g2_buf_1 _13620_ (.A(_04696_),
    .X(_05254_));
 sg13g2_a21oi_1 _13621_ (.A1(_05252_),
    .A2(_05253_),
    .Y(_00614_),
    .B1(net94));
 sg13g2_nand2_1 _13622_ (.Y(_05255_),
    .A(_04002_),
    .B(\am_sdr0.cic1.comb3[16] ));
 sg13g2_nand2_1 _13623_ (.Y(_05256_),
    .A(\am_sdr0.cic1.x_out[12] ),
    .B(_04721_));
 sg13g2_a21oi_1 _13624_ (.A1(_05255_),
    .A2(_05256_),
    .Y(_00615_),
    .B1(net94));
 sg13g2_nand2_1 _13625_ (.Y(_05257_),
    .A(_04002_),
    .B(\am_sdr0.cic1.comb3[17] ));
 sg13g2_nand2_1 _13626_ (.Y(_05258_),
    .A(\am_sdr0.cic1.x_out[13] ),
    .B(net161));
 sg13g2_a21oi_1 _13627_ (.A1(_05257_),
    .A2(_05258_),
    .Y(_00616_),
    .B1(net94));
 sg13g2_nand2_1 _13628_ (.Y(_05259_),
    .A(net233),
    .B(\am_sdr0.cic1.comb3[18] ));
 sg13g2_nand2_1 _13629_ (.Y(_05260_),
    .A(\am_sdr0.cic1.x_out[14] ),
    .B(net161));
 sg13g2_a21oi_1 _13630_ (.A1(_05259_),
    .A2(_05260_),
    .Y(_00617_),
    .B1(net94));
 sg13g2_nand2_1 _13631_ (.Y(_05261_),
    .A(net233),
    .B(\am_sdr0.cic1.comb3[19] ));
 sg13g2_buf_1 _13632_ (.A(\am_sdr0.cic1.x_out[15] ),
    .X(_05262_));
 sg13g2_buf_1 _13633_ (.A(_05262_),
    .X(_05263_));
 sg13g2_buf_1 _13634_ (.A(_05263_),
    .X(_05264_));
 sg13g2_nand2_1 _13635_ (.Y(_05265_),
    .A(net226),
    .B(net161));
 sg13g2_a21oi_1 _13636_ (.A1(_05261_),
    .A2(_05265_),
    .Y(_00618_),
    .B1(net94));
 sg13g2_nand2_1 _13637_ (.Y(_05266_),
    .A(net233),
    .B(\am_sdr0.cic1.comb3[12] ));
 sg13g2_buf_1 _13638_ (.A(\am_sdr0.cic1.x_out[8] ),
    .X(_05267_));
 sg13g2_nand2_1 _13639_ (.Y(_05268_),
    .A(_05267_),
    .B(_04075_));
 sg13g2_a21oi_1 _13640_ (.A1(_05266_),
    .A2(_05268_),
    .Y(_00619_),
    .B1(_05254_));
 sg13g2_nand2_1 _13641_ (.Y(_05269_),
    .A(net233),
    .B(\am_sdr0.cic1.comb3[13] ));
 sg13g2_buf_2 _13642_ (.A(\am_sdr0.cic1.x_out[9] ),
    .X(_05270_));
 sg13g2_nand2_1 _13643_ (.Y(_05271_),
    .A(_05270_),
    .B(_04075_));
 sg13g2_a21oi_1 _13644_ (.A1(_05269_),
    .A2(_05271_),
    .Y(_00620_),
    .B1(_05254_));
 sg13g2_buf_1 _13645_ (.A(\am_sdr0.cic2.sample ),
    .X(_05272_));
 sg13g2_buf_1 _13646_ (.A(_05272_),
    .X(_05273_));
 sg13g2_buf_1 _13647_ (.A(net285),
    .X(_05274_));
 sg13g2_xnor2_1 _13648_ (.Y(_05275_),
    .A(_02363_),
    .B(\am_sdr0.cic2.comb1_in_del[0] ));
 sg13g2_buf_2 _13649_ (.A(\am_sdr0.cic2.comb1[0] ),
    .X(_05276_));
 sg13g2_buf_1 _13650_ (.A(_05272_),
    .X(_05277_));
 sg13g2_buf_1 _13651_ (.A(_05277_),
    .X(_05278_));
 sg13g2_o21ai_1 _13652_ (.B1(net244),
    .Y(_05279_),
    .A1(_05276_),
    .A2(_05278_));
 sg13g2_a21oi_1 _13653_ (.A1(_05274_),
    .A2(_05275_),
    .Y(_00621_),
    .B1(_05279_));
 sg13g2_buf_1 _13654_ (.A(_05273_),
    .X(_05280_));
 sg13g2_buf_1 _13655_ (.A(\am_sdr0.cic2.comb1_in_del[8] ),
    .X(_05281_));
 sg13g2_nor2b_1 _13656_ (.A(\am_sdr0.cic2.comb1_in_del[2] ),
    .B_N(_02398_),
    .Y(_05282_));
 sg13g2_nor2b_1 _13657_ (.A(_02363_),
    .B_N(\am_sdr0.cic2.comb1_in_del[0] ),
    .Y(_05283_));
 sg13g2_buf_1 _13658_ (.A(\am_sdr0.cic2.comb1_in_del[1] ),
    .X(_05284_));
 sg13g2_nand2b_1 _13659_ (.Y(_05285_),
    .B(_02396_),
    .A_N(_05284_));
 sg13g2_nor2b_1 _13660_ (.A(_02396_),
    .B_N(_05284_),
    .Y(_05286_));
 sg13g2_a21oi_1 _13661_ (.A1(_05283_),
    .A2(_05285_),
    .Y(_05287_),
    .B1(_05286_));
 sg13g2_nand2b_1 _13662_ (.Y(_05288_),
    .B(\am_sdr0.cic2.comb1_in_del[2] ),
    .A_N(_02398_));
 sg13g2_o21ai_1 _13663_ (.B1(_05288_),
    .Y(_05289_),
    .A1(_05282_),
    .A2(_05287_));
 sg13g2_buf_2 _13664_ (.A(_05289_),
    .X(_05290_));
 sg13g2_buf_2 _13665_ (.A(\am_sdr0.cic2.comb1_in_del[3] ),
    .X(_05291_));
 sg13g2_inv_1 _13666_ (.Y(_05292_),
    .A(_05291_));
 sg13g2_buf_2 _13667_ (.A(\am_sdr0.cic2.comb1_in_del[4] ),
    .X(_05293_));
 sg13g2_nand2b_1 _13668_ (.Y(_05294_),
    .B(_02403_),
    .A_N(_05293_));
 sg13g2_buf_1 _13669_ (.A(\am_sdr0.cic2.comb1_in_del[5] ),
    .X(_05295_));
 sg13g2_o21ai_1 _13670_ (.B1(_05295_),
    .Y(_05296_),
    .A1(_02405_),
    .A2(_05294_));
 sg13g2_nand2_1 _13671_ (.Y(_05297_),
    .A(_02405_),
    .B(_05294_));
 sg13g2_a22oi_1 _13672_ (.Y(_05298_),
    .B1(_05296_),
    .B2(_05297_),
    .A2(_05292_),
    .A1(_02400_));
 sg13g2_buf_2 _13673_ (.A(\am_sdr0.cic2.comb1_in_del[6] ),
    .X(_05299_));
 sg13g2_nand2b_1 _13674_ (.Y(_05300_),
    .B(_02410_),
    .A_N(_05299_));
 sg13g2_nand2_1 _13675_ (.Y(_05301_),
    .A(_02409_),
    .B(_02410_));
 sg13g2_inv_1 _13676_ (.Y(_05302_),
    .A(_05295_));
 sg13g2_nor2b_1 _13677_ (.A(_02400_),
    .B_N(_05291_),
    .Y(_05303_));
 sg13g2_nor2b_1 _13678_ (.A(_02403_),
    .B_N(_05293_),
    .Y(_05304_));
 sg13g2_a221oi_1 _13679_ (.B2(_05303_),
    .C1(_05304_),
    .B1(_05294_),
    .A1(_02405_),
    .Y(_05305_),
    .A2(_05295_));
 sg13g2_a21oi_1 _13680_ (.A1(_02404_),
    .A2(_05302_),
    .Y(_05306_),
    .B1(_05305_));
 sg13g2_a221oi_1 _13681_ (.B2(_05301_),
    .C1(_05306_),
    .B1(_05300_),
    .A1(_05290_),
    .Y(_05307_),
    .A2(_05298_));
 sg13g2_buf_1 _13682_ (.A(\am_sdr0.cic2.comb1_in_del[7] ),
    .X(_05308_));
 sg13g2_or2_1 _13683_ (.X(_05309_),
    .B(_05308_),
    .A(_05299_));
 sg13g2_nand2b_1 _13684_ (.Y(_05310_),
    .B(_02409_),
    .A_N(_05308_));
 sg13g2_a221oi_1 _13685_ (.B2(_05310_),
    .C1(_05306_),
    .B1(_05309_),
    .A1(_05290_),
    .Y(_05311_),
    .A2(_05298_));
 sg13g2_nor2_1 _13686_ (.A(_02411_),
    .B(_05308_),
    .Y(_05312_));
 sg13g2_nand2b_1 _13687_ (.Y(_05313_),
    .B(_02409_),
    .A_N(_05299_));
 sg13g2_a21oi_1 _13688_ (.A1(_02411_),
    .A2(_05308_),
    .Y(_05314_),
    .B1(_05313_));
 sg13g2_nor4_1 _13689_ (.A(_05307_),
    .B(_05311_),
    .C(_05312_),
    .D(_05314_),
    .Y(_05315_));
 sg13g2_buf_2 _13690_ (.A(_05315_),
    .X(_05316_));
 sg13g2_nand2_1 _13691_ (.Y(_05317_),
    .A(_05281_),
    .B(_05316_));
 sg13g2_nor2_1 _13692_ (.A(_05281_),
    .B(_05316_),
    .Y(_05318_));
 sg13g2_a21oi_1 _13693_ (.A1(_02415_),
    .A2(_05317_),
    .Y(_05319_),
    .B1(_05318_));
 sg13g2_buf_1 _13694_ (.A(\am_sdr0.cic2.comb1_in_del[9] ),
    .X(_05320_));
 sg13g2_nor2b_1 _13695_ (.A(_02416_),
    .B_N(_05320_),
    .Y(_05321_));
 sg13g2_nand2b_1 _13696_ (.Y(_05322_),
    .B(_02416_),
    .A_N(_05320_));
 sg13g2_o21ai_1 _13697_ (.B1(_05322_),
    .Y(_05323_),
    .A1(_05319_),
    .A2(_05321_));
 sg13g2_buf_1 _13698_ (.A(\am_sdr0.cic2.comb1_in_del[10] ),
    .X(_05324_));
 sg13g2_xor2_1 _13699_ (.B(_05324_),
    .A(_02376_),
    .X(_05325_));
 sg13g2_xnor2_1 _13700_ (.Y(_05326_),
    .A(_05323_),
    .B(_05325_));
 sg13g2_buf_1 _13701_ (.A(_05272_),
    .X(_05327_));
 sg13g2_buf_1 _13702_ (.A(\am_sdr0.cic2.comb1[10] ),
    .X(_05328_));
 sg13g2_nor2b_1 _13703_ (.A(net283),
    .B_N(_05328_),
    .Y(_05329_));
 sg13g2_a21oi_1 _13704_ (.A1(net223),
    .A2(_05326_),
    .Y(_05330_),
    .B1(_05329_));
 sg13g2_nor2_1 _13705_ (.A(net95),
    .B(_05330_),
    .Y(_00622_));
 sg13g2_inv_1 _13706_ (.Y(_05331_),
    .A(_05281_));
 sg13g2_inv_1 _13707_ (.Y(_05332_),
    .A(_05324_));
 sg13g2_nor2_1 _13708_ (.A(_02417_),
    .B(_05320_),
    .Y(_05333_));
 sg13g2_nor3_1 _13709_ (.A(_05331_),
    .B(_05332_),
    .C(_05333_),
    .Y(_05334_));
 sg13g2_nor3_1 _13710_ (.A(_02415_),
    .B(_05332_),
    .C(_05333_),
    .Y(_05335_));
 sg13g2_o21ai_1 _13711_ (.B1(_05316_),
    .Y(_05336_),
    .A1(_05334_),
    .A2(_05335_));
 sg13g2_nor3_1 _13712_ (.A(_02415_),
    .B(_05331_),
    .C(_05333_),
    .Y(_05337_));
 sg13g2_o21ai_1 _13713_ (.B1(_05324_),
    .Y(_05338_),
    .A1(_05321_),
    .A2(_05337_));
 sg13g2_and3_1 _13714_ (.X(_05339_),
    .A(_02376_),
    .B(_05336_),
    .C(_05338_));
 sg13g2_nand2_1 _13715_ (.Y(_05340_),
    .A(_05331_),
    .B(_05332_));
 sg13g2_nand2_1 _13716_ (.Y(_05341_),
    .A(_02415_),
    .B(_05332_));
 sg13g2_a221oi_1 _13717_ (.B2(_05341_),
    .C1(_05316_),
    .B1(_05340_),
    .A1(_02417_),
    .Y(_05342_),
    .A2(_05320_));
 sg13g2_nand3b_1 _13718_ (.B(_02415_),
    .C(_05331_),
    .Y(_05343_),
    .A_N(_05321_));
 sg13g2_a21oi_1 _13719_ (.A1(_05322_),
    .A2(_05343_),
    .Y(_05344_),
    .B1(_05324_));
 sg13g2_nor3_1 _13720_ (.A(_05339_),
    .B(_05342_),
    .C(_05344_),
    .Y(_05345_));
 sg13g2_nor2b_1 _13721_ (.A(\am_sdr0.cic2.comb1_in_del[11] ),
    .B_N(_02378_),
    .Y(_05346_));
 sg13g2_nand2b_1 _13722_ (.Y(_05347_),
    .B(\am_sdr0.cic2.comb1_in_del[11] ),
    .A_N(_02378_));
 sg13g2_nand2b_1 _13723_ (.Y(_05348_),
    .B(_05347_),
    .A_N(_05346_));
 sg13g2_xor2_1 _13724_ (.B(_05348_),
    .A(_05345_),
    .X(_05349_));
 sg13g2_buf_2 _13725_ (.A(\am_sdr0.cic2.comb1[11] ),
    .X(_05350_));
 sg13g2_nor2b_1 _13726_ (.A(net283),
    .B_N(_05350_),
    .Y(_05351_));
 sg13g2_a21oi_1 _13727_ (.A1(net223),
    .A2(_05349_),
    .Y(_05352_),
    .B1(_05351_));
 sg13g2_nor2_1 _13728_ (.A(net95),
    .B(_05352_),
    .Y(_00623_));
 sg13g2_buf_1 _13729_ (.A(\am_sdr0.cic2.comb1[12] ),
    .X(_05353_));
 sg13g2_inv_1 _13730_ (.Y(_05354_),
    .A(_05272_));
 sg13g2_buf_1 _13731_ (.A(_05354_),
    .X(_05355_));
 sg13g2_buf_1 _13732_ (.A(_05355_),
    .X(_05356_));
 sg13g2_buf_1 _13733_ (.A(net155),
    .X(_05357_));
 sg13g2_buf_1 _13734_ (.A(_05355_),
    .X(_05358_));
 sg13g2_o21ai_1 _13735_ (.B1(_05347_),
    .Y(_05359_),
    .A1(_05342_),
    .A2(_05344_));
 sg13g2_nand4_1 _13736_ (.B(_05336_),
    .C(_05338_),
    .A(_02376_),
    .Y(_05360_),
    .D(_05347_));
 sg13g2_buf_1 _13737_ (.A(_05360_),
    .X(_05361_));
 sg13g2_nand2_1 _13738_ (.Y(_05362_),
    .A(_05359_),
    .B(_05361_));
 sg13g2_nor2_1 _13739_ (.A(_05346_),
    .B(_05362_),
    .Y(_05363_));
 sg13g2_buf_1 _13740_ (.A(\am_sdr0.cic2.comb1_in_del[12] ),
    .X(_05364_));
 sg13g2_xor2_1 _13741_ (.B(_05364_),
    .A(_02380_),
    .X(_05365_));
 sg13g2_xnor2_1 _13742_ (.Y(_05366_),
    .A(_05363_),
    .B(_05365_));
 sg13g2_nor2_1 _13743_ (.A(net154),
    .B(_05366_),
    .Y(_05367_));
 sg13g2_a21oi_1 _13744_ (.A1(_05353_),
    .A2(net93),
    .Y(_05368_),
    .B1(_05367_));
 sg13g2_nor2_1 _13745_ (.A(_05246_),
    .B(_05368_),
    .Y(_00624_));
 sg13g2_buf_1 _13746_ (.A(\am_sdr0.cic2.comb1[13] ),
    .X(_05369_));
 sg13g2_buf_1 _13747_ (.A(net155),
    .X(_05370_));
 sg13g2_nand2_1 _13748_ (.Y(_05371_),
    .A(_05369_),
    .B(net92));
 sg13g2_buf_1 _13749_ (.A(net284),
    .X(_05372_));
 sg13g2_nand2b_1 _13750_ (.Y(_05373_),
    .B(_05364_),
    .A_N(_02380_));
 sg13g2_nor2b_1 _13751_ (.A(_05346_),
    .B_N(_05364_),
    .Y(_05374_));
 sg13g2_nand3_1 _13752_ (.B(_05361_),
    .C(_05374_),
    .A(_05359_),
    .Y(_05375_));
 sg13g2_nor2_1 _13753_ (.A(_02380_),
    .B(_05346_),
    .Y(_05376_));
 sg13g2_nand3_1 _13754_ (.B(_05361_),
    .C(_05376_),
    .A(_05359_),
    .Y(_05377_));
 sg13g2_nand3_1 _13755_ (.B(_05375_),
    .C(_05377_),
    .A(_05373_),
    .Y(_05378_));
 sg13g2_nor2b_1 _13756_ (.A(_02382_),
    .B_N(\am_sdr0.cic2.comb1_in_del[13] ),
    .Y(_05379_));
 sg13g2_nand2b_1 _13757_ (.Y(_05380_),
    .B(_02382_),
    .A_N(\am_sdr0.cic2.comb1_in_del[13] ));
 sg13g2_nor2b_1 _13758_ (.A(_05379_),
    .B_N(_05380_),
    .Y(_05381_));
 sg13g2_xnor2_1 _13759_ (.Y(_05382_),
    .A(_05378_),
    .B(_05381_));
 sg13g2_nand2_1 _13760_ (.Y(_05383_),
    .A(_05372_),
    .B(_05382_));
 sg13g2_a21oi_1 _13761_ (.A1(_05371_),
    .A2(_05383_),
    .Y(_00625_),
    .B1(net94));
 sg13g2_buf_1 _13762_ (.A(\am_sdr0.cic2.comb1[14] ),
    .X(_05384_));
 sg13g2_buf_1 _13763_ (.A(\am_sdr0.cic2.comb1_in_del[14] ),
    .X(_05385_));
 sg13g2_xnor2_1 _13764_ (.Y(_05386_),
    .A(_02384_),
    .B(_05385_));
 sg13g2_o21ai_1 _13765_ (.B1(_05380_),
    .Y(_05387_),
    .A1(_05378_),
    .A2(_05379_));
 sg13g2_xnor2_1 _13766_ (.Y(_05388_),
    .A(_05386_),
    .B(_05387_));
 sg13g2_nor2_1 _13767_ (.A(net154),
    .B(_05388_),
    .Y(_05389_));
 sg13g2_a21oi_1 _13768_ (.A1(_05384_),
    .A2(net93),
    .Y(_05390_),
    .B1(_05389_));
 sg13g2_nor2_1 _13769_ (.A(net95),
    .B(_05390_),
    .Y(_00626_));
 sg13g2_buf_2 _13770_ (.A(\am_sdr0.cic2.comb1[15] ),
    .X(_05391_));
 sg13g2_buf_1 _13771_ (.A(net284),
    .X(_05392_));
 sg13g2_nor2b_1 _13772_ (.A(_05385_),
    .B_N(_02384_),
    .Y(_05393_));
 sg13g2_nand2b_1 _13773_ (.Y(_05394_),
    .B(_05385_),
    .A_N(_02384_));
 sg13g2_o21ai_1 _13774_ (.B1(_05394_),
    .Y(_05395_),
    .A1(_05393_),
    .A2(_05387_));
 sg13g2_buf_1 _13775_ (.A(_05395_),
    .X(_05396_));
 sg13g2_buf_1 _13776_ (.A(\am_sdr0.cic2.comb1_in_del[15] ),
    .X(_05397_));
 sg13g2_nand2b_1 _13777_ (.Y(_05398_),
    .B(_05397_),
    .A_N(_02386_));
 sg13g2_nand2b_1 _13778_ (.Y(_05399_),
    .B(_02386_),
    .A_N(_05397_));
 sg13g2_nand2_1 _13779_ (.Y(_05400_),
    .A(_05398_),
    .B(_05399_));
 sg13g2_xnor2_1 _13780_ (.Y(_05401_),
    .A(_05396_),
    .B(_05400_));
 sg13g2_nand2_1 _13781_ (.Y(_05402_),
    .A(_05327_),
    .B(_05401_));
 sg13g2_o21ai_1 _13782_ (.B1(_05402_),
    .Y(_05403_),
    .A1(_05391_),
    .A2(_05392_));
 sg13g2_nor2_1 _13783_ (.A(net95),
    .B(_05403_),
    .Y(_00627_));
 sg13g2_buf_2 _13784_ (.A(\am_sdr0.cic2.comb1[16] ),
    .X(_05404_));
 sg13g2_nor2b_1 _13785_ (.A(_02386_),
    .B_N(_05397_),
    .Y(_05405_));
 sg13g2_o21ai_1 _13786_ (.B1(_05399_),
    .Y(_05406_),
    .A1(_05396_),
    .A2(_05405_));
 sg13g2_buf_1 _13787_ (.A(_05406_),
    .X(_05407_));
 sg13g2_xnor2_1 _13788_ (.Y(_05408_),
    .A(_02388_),
    .B(\am_sdr0.cic2.comb1_in_del[16] ));
 sg13g2_xnor2_1 _13789_ (.Y(_05409_),
    .A(_05407_),
    .B(_05408_));
 sg13g2_nor2_1 _13790_ (.A(net154),
    .B(_05409_),
    .Y(_05410_));
 sg13g2_a21oi_1 _13791_ (.A1(_05404_),
    .A2(_05357_),
    .Y(_05411_),
    .B1(_05410_));
 sg13g2_nor2_1 _13792_ (.A(net95),
    .B(_05411_),
    .Y(_00628_));
 sg13g2_buf_2 _13793_ (.A(\am_sdr0.cic2.comb1[17] ),
    .X(_05412_));
 sg13g2_nand2_1 _13794_ (.Y(_05413_),
    .A(_05412_),
    .B(net92));
 sg13g2_inv_1 _13795_ (.Y(_05414_),
    .A(\am_sdr0.cic2.comb1_in_del[16] ));
 sg13g2_nand2_1 _13796_ (.Y(_05415_),
    .A(_02388_),
    .B(_05398_));
 sg13g2_nor2b_1 _13797_ (.A(_05397_),
    .B_N(_02386_),
    .Y(_05416_));
 sg13g2_o21ai_1 _13798_ (.B1(_02388_),
    .Y(_05417_),
    .A1(_05414_),
    .A2(_05416_));
 sg13g2_o21ai_1 _13799_ (.B1(_05417_),
    .Y(_05418_),
    .A1(_05396_),
    .A2(_05415_));
 sg13g2_a21oi_1 _13800_ (.A1(_05414_),
    .A2(_05407_),
    .Y(_05419_),
    .B1(_05418_));
 sg13g2_xnor2_1 _13801_ (.Y(_05420_),
    .A(_02390_),
    .B(\am_sdr0.cic2.comb1_in_del[17] ));
 sg13g2_xnor2_1 _13802_ (.Y(_05421_),
    .A(_05419_),
    .B(_05420_));
 sg13g2_nand2_1 _13803_ (.Y(_05422_),
    .A(net222),
    .B(_05421_));
 sg13g2_a21oi_1 _13804_ (.A1(_05413_),
    .A2(_05422_),
    .Y(_00629_),
    .B1(net94));
 sg13g2_buf_1 _13805_ (.A(\am_sdr0.cic2.comb1[18] ),
    .X(_05423_));
 sg13g2_nand2_1 _13806_ (.Y(_05424_),
    .A(_05423_),
    .B(net92));
 sg13g2_inv_1 _13807_ (.Y(_05425_),
    .A(\am_sdr0.cic2.comb1_in_del[17] ));
 sg13g2_nor2_1 _13808_ (.A(_02390_),
    .B(_05425_),
    .Y(_05426_));
 sg13g2_a221oi_1 _13809_ (.B2(_05414_),
    .C1(_05418_),
    .B1(_05407_),
    .A1(_02390_),
    .Y(_05427_),
    .A2(_05425_));
 sg13g2_buf_1 _13810_ (.A(_05427_),
    .X(_05428_));
 sg13g2_nor2b_1 _13811_ (.A(\am_sdr0.cic2.comb1_in_del[18] ),
    .B_N(_02392_),
    .Y(_05429_));
 sg13g2_nor2b_1 _13812_ (.A(_02392_),
    .B_N(\am_sdr0.cic2.comb1_in_del[18] ),
    .Y(_05430_));
 sg13g2_or2_1 _13813_ (.X(_05431_),
    .B(_05430_),
    .A(_05429_));
 sg13g2_nor3_1 _13814_ (.A(_05426_),
    .B(_05428_),
    .C(_05431_),
    .Y(_05432_));
 sg13g2_o21ai_1 _13815_ (.B1(_05431_),
    .Y(_05433_),
    .A1(_05426_),
    .A2(_05428_));
 sg13g2_nand3b_1 _13816_ (.B(_05433_),
    .C(_05278_),
    .Y(_05434_),
    .A_N(_05432_));
 sg13g2_a21oi_1 _13817_ (.A1(_05424_),
    .A2(_05434_),
    .Y(_00630_),
    .B1(net94));
 sg13g2_nor3_1 _13818_ (.A(_05426_),
    .B(_05428_),
    .C(_05430_),
    .Y(_05435_));
 sg13g2_nand2_1 _13819_ (.Y(_05436_),
    .A(_01558_),
    .B(_05272_));
 sg13g2_xor2_1 _13820_ (.B(\am_sdr0.cic2.comb1_in_del[19] ),
    .A(\am_sdr0.cic2.integ_sample[19] ),
    .X(_05437_));
 sg13g2_nor2b_1 _13821_ (.A(_05436_),
    .B_N(_05437_),
    .Y(_05438_));
 sg13g2_o21ai_1 _13822_ (.B1(_05438_),
    .Y(_05439_),
    .A1(_05429_),
    .A2(_05435_));
 sg13g2_or4_1 _13823_ (.A(_05429_),
    .B(_05436_),
    .C(_05435_),
    .D(_05437_),
    .X(_05440_));
 sg13g2_nand3_1 _13824_ (.B(\am_sdr0.cic2.comb1[19] ),
    .C(_05358_),
    .A(_01718_),
    .Y(_05441_));
 sg13g2_nand3_1 _13825_ (.B(_05440_),
    .C(_05441_),
    .A(_05439_),
    .Y(_00631_));
 sg13g2_buf_1 _13826_ (.A(\am_sdr0.cic2.comb1[1] ),
    .X(_05442_));
 sg13g2_nand2_1 _13827_ (.Y(_05443_),
    .A(_05442_),
    .B(net92));
 sg13g2_xnor2_1 _13828_ (.Y(_05444_),
    .A(_02396_),
    .B(_05284_));
 sg13g2_xnor2_1 _13829_ (.Y(_05445_),
    .A(_05283_),
    .B(_05444_));
 sg13g2_nand2_1 _13830_ (.Y(_05446_),
    .A(net222),
    .B(_05445_));
 sg13g2_buf_1 _13831_ (.A(_04696_),
    .X(_05447_));
 sg13g2_a21oi_1 _13832_ (.A1(_05443_),
    .A2(_05446_),
    .Y(_00632_),
    .B1(net91));
 sg13g2_buf_2 _13833_ (.A(\am_sdr0.cic2.comb1[2] ),
    .X(_05448_));
 sg13g2_nor2b_1 _13834_ (.A(_05282_),
    .B_N(_05288_),
    .Y(_05449_));
 sg13g2_xnor2_1 _13835_ (.Y(_05450_),
    .A(_05287_),
    .B(_05449_));
 sg13g2_nor2_1 _13836_ (.A(net154),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_a21oi_1 _13837_ (.A1(_05448_),
    .A2(net93),
    .Y(_05452_),
    .B1(_05451_));
 sg13g2_nor2_1 _13838_ (.A(net95),
    .B(_05452_),
    .Y(_00633_));
 sg13g2_buf_1 _13839_ (.A(\am_sdr0.cic2.comb1[3] ),
    .X(_05453_));
 sg13g2_nand2_1 _13840_ (.Y(_05454_),
    .A(_05453_),
    .B(net92));
 sg13g2_xnor2_1 _13841_ (.Y(_05455_),
    .A(_02400_),
    .B(_05291_));
 sg13g2_xnor2_1 _13842_ (.Y(_05456_),
    .A(_05290_),
    .B(_05455_));
 sg13g2_nand2_1 _13843_ (.Y(_05457_),
    .A(net222),
    .B(_05456_));
 sg13g2_a21oi_1 _13844_ (.A1(_05454_),
    .A2(_05457_),
    .Y(_00634_),
    .B1(net91));
 sg13g2_buf_1 _13845_ (.A(\am_sdr0.cic2.comb1[4] ),
    .X(_05458_));
 sg13g2_nor2_1 _13846_ (.A(_05458_),
    .B(net221),
    .Y(_05459_));
 sg13g2_nor2_1 _13847_ (.A(_05291_),
    .B(_05290_),
    .Y(_05460_));
 sg13g2_nor2_1 _13848_ (.A(_02400_),
    .B(_05460_),
    .Y(_05461_));
 sg13g2_a21oi_2 _13849_ (.B1(_05461_),
    .Y(_05462_),
    .A2(_05290_),
    .A1(_05291_));
 sg13g2_xor2_1 _13850_ (.B(_05293_),
    .A(_02403_),
    .X(_05463_));
 sg13g2_xnor2_1 _13851_ (.Y(_05464_),
    .A(_05462_),
    .B(_05463_));
 sg13g2_nor2_1 _13852_ (.A(net154),
    .B(_05464_),
    .Y(_05465_));
 sg13g2_nor3_1 _13853_ (.A(net160),
    .B(_05459_),
    .C(_05465_),
    .Y(_00635_));
 sg13g2_buf_1 _13854_ (.A(\am_sdr0.cic2.comb1[5] ),
    .X(_05466_));
 sg13g2_buf_1 _13855_ (.A(net155),
    .X(_05467_));
 sg13g2_inv_1 _13856_ (.Y(_05468_),
    .A(_05462_));
 sg13g2_inv_1 _13857_ (.Y(_05469_),
    .A(_05293_));
 sg13g2_o21ai_1 _13858_ (.B1(_02403_),
    .Y(_05470_),
    .A1(_05469_),
    .A2(_05462_));
 sg13g2_o21ai_1 _13859_ (.B1(_05470_),
    .Y(_05471_),
    .A1(_05293_),
    .A2(_05468_));
 sg13g2_xnor2_1 _13860_ (.Y(_05472_),
    .A(_02404_),
    .B(_05295_));
 sg13g2_xnor2_1 _13861_ (.Y(_05473_),
    .A(_05471_),
    .B(_05472_));
 sg13g2_nor2_1 _13862_ (.A(net155),
    .B(_05473_),
    .Y(_05474_));
 sg13g2_a21oi_1 _13863_ (.A1(_05466_),
    .A2(net90),
    .Y(_05475_),
    .B1(_05474_));
 sg13g2_nor2_1 _13864_ (.A(net95),
    .B(_05475_),
    .Y(_00636_));
 sg13g2_buf_1 _13865_ (.A(\am_sdr0.cic2.comb1[6] ),
    .X(_05476_));
 sg13g2_a21o_1 _13866_ (.A2(_05298_),
    .A1(_05290_),
    .B1(_05306_),
    .X(_05477_));
 sg13g2_buf_1 _13867_ (.A(_05477_),
    .X(_05478_));
 sg13g2_xor2_1 _13868_ (.B(_05299_),
    .A(_02409_),
    .X(_05479_));
 sg13g2_xnor2_1 _13869_ (.Y(_05480_),
    .A(_05478_),
    .B(_05479_));
 sg13g2_nand2_1 _13870_ (.Y(_05481_),
    .A(net283),
    .B(_05480_));
 sg13g2_o21ai_1 _13871_ (.B1(_05481_),
    .Y(_05482_),
    .A1(_05476_),
    .A2(net221));
 sg13g2_nor2_1 _13872_ (.A(net95),
    .B(_05482_),
    .Y(_00637_));
 sg13g2_buf_2 _13873_ (.A(\am_sdr0.cic2.comb1[7] ),
    .X(_05483_));
 sg13g2_nand2_1 _13874_ (.Y(_05484_),
    .A(_05483_),
    .B(net92));
 sg13g2_nor2_1 _13875_ (.A(_05299_),
    .B(_05478_),
    .Y(_05485_));
 sg13g2_nand2_1 _13876_ (.Y(_05486_),
    .A(_05299_),
    .B(_05478_));
 sg13g2_o21ai_1 _13877_ (.B1(_05486_),
    .Y(_05487_),
    .A1(_02409_),
    .A2(_05485_));
 sg13g2_xnor2_1 _13878_ (.Y(_05488_),
    .A(_02410_),
    .B(_05308_));
 sg13g2_xnor2_1 _13879_ (.Y(_05489_),
    .A(_05487_),
    .B(_05488_));
 sg13g2_nand2_1 _13880_ (.Y(_05490_),
    .A(net222),
    .B(_05489_));
 sg13g2_a21oi_1 _13881_ (.A1(_05484_),
    .A2(_05490_),
    .Y(_00638_),
    .B1(net91));
 sg13g2_buf_1 _13882_ (.A(_05203_),
    .X(_05491_));
 sg13g2_buf_2 _13883_ (.A(\am_sdr0.cic2.comb1[8] ),
    .X(_05492_));
 sg13g2_xor2_1 _13884_ (.B(_05281_),
    .A(_02415_),
    .X(_05493_));
 sg13g2_xnor2_1 _13885_ (.Y(_05494_),
    .A(_05316_),
    .B(_05493_));
 sg13g2_nand2_1 _13886_ (.Y(_05495_),
    .A(net283),
    .B(_05494_));
 sg13g2_o21ai_1 _13887_ (.B1(_05495_),
    .Y(_05496_),
    .A1(_05492_),
    .A2(net221));
 sg13g2_nor2_1 _13888_ (.A(net89),
    .B(_05496_),
    .Y(_00639_));
 sg13g2_nor2_1 _13889_ (.A(_05333_),
    .B(_05321_),
    .Y(_05497_));
 sg13g2_xnor2_1 _13890_ (.Y(_05498_),
    .A(_05319_),
    .B(_05497_));
 sg13g2_buf_1 _13891_ (.A(\am_sdr0.cic2.comb1[9] ),
    .X(_05499_));
 sg13g2_nor2b_1 _13892_ (.A(net283),
    .B_N(_05499_),
    .Y(_05500_));
 sg13g2_a21oi_1 _13893_ (.A1(net223),
    .A2(_05498_),
    .Y(_05501_),
    .B1(_05500_));
 sg13g2_nor2_1 _13894_ (.A(net89),
    .B(_05501_),
    .Y(_00640_));
 sg13g2_buf_1 _13895_ (.A(net285),
    .X(_05502_));
 sg13g2_nand2_1 _13896_ (.Y(_05503_),
    .A(_02363_),
    .B(net220));
 sg13g2_nand2_1 _13897_ (.Y(_05504_),
    .A(\am_sdr0.cic2.comb1_in_del[0] ),
    .B(net90));
 sg13g2_a21oi_1 _13898_ (.A1(_05503_),
    .A2(_05504_),
    .Y(_00641_),
    .B1(net91));
 sg13g2_nand2_1 _13899_ (.Y(_05505_),
    .A(_02376_),
    .B(net220));
 sg13g2_nand2_1 _13900_ (.Y(_05506_),
    .A(_05324_),
    .B(net90));
 sg13g2_a21oi_1 _13901_ (.A1(_05505_),
    .A2(_05506_),
    .Y(_00642_),
    .B1(net91));
 sg13g2_nand2_1 _13902_ (.Y(_05507_),
    .A(_02378_),
    .B(net220));
 sg13g2_nand2_1 _13903_ (.Y(_05508_),
    .A(\am_sdr0.cic2.comb1_in_del[11] ),
    .B(net90));
 sg13g2_a21oi_1 _13904_ (.A1(_05507_),
    .A2(_05508_),
    .Y(_00643_),
    .B1(net91));
 sg13g2_nand2_1 _13905_ (.Y(_05509_),
    .A(_02380_),
    .B(net220));
 sg13g2_nand2_1 _13906_ (.Y(_05510_),
    .A(_05364_),
    .B(net90));
 sg13g2_a21oi_1 _13907_ (.A1(_05509_),
    .A2(_05510_),
    .Y(_00644_),
    .B1(net91));
 sg13g2_nand2_1 _13908_ (.Y(_05511_),
    .A(_02382_),
    .B(_05502_));
 sg13g2_nand2_1 _13909_ (.Y(_05512_),
    .A(\am_sdr0.cic2.comb1_in_del[13] ),
    .B(net90));
 sg13g2_a21oi_1 _13910_ (.A1(_05511_),
    .A2(_05512_),
    .Y(_00645_),
    .B1(net91));
 sg13g2_nand2_1 _13911_ (.Y(_05513_),
    .A(_02384_),
    .B(_05502_));
 sg13g2_nand2_1 _13912_ (.Y(_05514_),
    .A(_05385_),
    .B(net90));
 sg13g2_a21oi_1 _13913_ (.A1(_05513_),
    .A2(_05514_),
    .Y(_00646_),
    .B1(_05447_));
 sg13g2_nand2_1 _13914_ (.Y(_05515_),
    .A(_02386_),
    .B(net220));
 sg13g2_nand2_1 _13915_ (.Y(_05516_),
    .A(_05397_),
    .B(net90));
 sg13g2_a21oi_1 _13916_ (.A1(_05515_),
    .A2(_05516_),
    .Y(_00647_),
    .B1(_05447_));
 sg13g2_nand2_1 _13917_ (.Y(_05517_),
    .A(_02388_),
    .B(net220));
 sg13g2_nand2_1 _13918_ (.Y(_05518_),
    .A(\am_sdr0.cic2.comb1_in_del[16] ),
    .B(_05467_));
 sg13g2_buf_1 _13919_ (.A(_04696_),
    .X(_05519_));
 sg13g2_a21oi_1 _13920_ (.A1(_05517_),
    .A2(_05518_),
    .Y(_00648_),
    .B1(net88));
 sg13g2_nand2_1 _13921_ (.Y(_05520_),
    .A(_02390_),
    .B(net220));
 sg13g2_buf_1 _13922_ (.A(net155),
    .X(_05521_));
 sg13g2_nand2_1 _13923_ (.Y(_05522_),
    .A(\am_sdr0.cic2.comb1_in_del[17] ),
    .B(_05521_));
 sg13g2_a21oi_1 _13924_ (.A1(_05520_),
    .A2(_05522_),
    .Y(_00649_),
    .B1(net88));
 sg13g2_nand2_1 _13925_ (.Y(_05523_),
    .A(_02392_),
    .B(net220));
 sg13g2_nand2_1 _13926_ (.Y(_05524_),
    .A(\am_sdr0.cic2.comb1_in_del[18] ),
    .B(net87));
 sg13g2_a21oi_1 _13927_ (.A1(_05523_),
    .A2(_05524_),
    .Y(_00650_),
    .B1(_05519_));
 sg13g2_buf_1 _13928_ (.A(net285),
    .X(_05525_));
 sg13g2_nand2_1 _13929_ (.Y(_05526_),
    .A(\am_sdr0.cic2.integ_sample[19] ),
    .B(_05525_));
 sg13g2_nand2_1 _13930_ (.Y(_05527_),
    .A(\am_sdr0.cic2.comb1_in_del[19] ),
    .B(_05521_));
 sg13g2_a21oi_1 _13931_ (.A1(_05526_),
    .A2(_05527_),
    .Y(_00651_),
    .B1(_05519_));
 sg13g2_nand2_1 _13932_ (.Y(_05528_),
    .A(_02396_),
    .B(net219));
 sg13g2_nand2_1 _13933_ (.Y(_05529_),
    .A(_05284_),
    .B(net87));
 sg13g2_a21oi_1 _13934_ (.A1(_05528_),
    .A2(_05529_),
    .Y(_00652_),
    .B1(net88));
 sg13g2_nand2_1 _13935_ (.Y(_05530_),
    .A(_02398_),
    .B(net219));
 sg13g2_nand2_1 _13936_ (.Y(_05531_),
    .A(\am_sdr0.cic2.comb1_in_del[2] ),
    .B(net87));
 sg13g2_a21oi_1 _13937_ (.A1(_05530_),
    .A2(_05531_),
    .Y(_00653_),
    .B1(net88));
 sg13g2_nand2_1 _13938_ (.Y(_05532_),
    .A(_02400_),
    .B(net219));
 sg13g2_nand2_1 _13939_ (.Y(_05533_),
    .A(_05291_),
    .B(net87));
 sg13g2_a21oi_1 _13940_ (.A1(_05532_),
    .A2(_05533_),
    .Y(_00654_),
    .B1(net88));
 sg13g2_nand2_1 _13941_ (.Y(_05534_),
    .A(_02403_),
    .B(net219));
 sg13g2_nand2_1 _13942_ (.Y(_05535_),
    .A(_05293_),
    .B(net87));
 sg13g2_a21oi_1 _13943_ (.A1(_05534_),
    .A2(_05535_),
    .Y(_00655_),
    .B1(net88));
 sg13g2_nand2_1 _13944_ (.Y(_05536_),
    .A(_02404_),
    .B(net219));
 sg13g2_nand2_1 _13945_ (.Y(_05537_),
    .A(_05295_),
    .B(net87));
 sg13g2_a21oi_1 _13946_ (.A1(_05536_),
    .A2(_05537_),
    .Y(_00656_),
    .B1(net88));
 sg13g2_nand2_1 _13947_ (.Y(_05538_),
    .A(_02409_),
    .B(net219));
 sg13g2_nand2_1 _13948_ (.Y(_05539_),
    .A(_05299_),
    .B(net87));
 sg13g2_a21oi_1 _13949_ (.A1(_05538_),
    .A2(_05539_),
    .Y(_00657_),
    .B1(net88));
 sg13g2_nand2_1 _13950_ (.Y(_05540_),
    .A(_02410_),
    .B(net219));
 sg13g2_nand2_1 _13951_ (.Y(_05541_),
    .A(_05308_),
    .B(net87));
 sg13g2_buf_1 _13952_ (.A(_04696_),
    .X(_05542_));
 sg13g2_a21oi_1 _13953_ (.A1(_05540_),
    .A2(_05541_),
    .Y(_00658_),
    .B1(net86));
 sg13g2_nand2_1 _13954_ (.Y(_05543_),
    .A(_02415_),
    .B(_05525_));
 sg13g2_buf_1 _13955_ (.A(net155),
    .X(_05544_));
 sg13g2_nand2_1 _13956_ (.Y(_05545_),
    .A(_05281_),
    .B(net85));
 sg13g2_a21oi_1 _13957_ (.A1(_05543_),
    .A2(_05545_),
    .Y(_00659_),
    .B1(net86));
 sg13g2_nand2_1 _13958_ (.Y(_05546_),
    .A(_02416_),
    .B(net219));
 sg13g2_nand2_1 _13959_ (.Y(_05547_),
    .A(_05320_),
    .B(net85));
 sg13g2_a21oi_1 _13960_ (.A1(_05546_),
    .A2(_05547_),
    .Y(_00660_),
    .B1(net86));
 sg13g2_xnor2_1 _13961_ (.Y(_05548_),
    .A(_05276_),
    .B(\am_sdr0.cic2.comb2_in_del[0] ));
 sg13g2_buf_1 _13962_ (.A(net303),
    .X(_05549_));
 sg13g2_o21ai_1 _13963_ (.B1(net218),
    .Y(_05550_),
    .A1(\am_sdr0.cic2.comb2[0] ),
    .A2(net224));
 sg13g2_a21oi_1 _13964_ (.A1(net225),
    .A2(_05548_),
    .Y(_00661_),
    .B1(_05550_));
 sg13g2_buf_1 _13965_ (.A(\am_sdr0.cic2.comb2[10] ),
    .X(_05551_));
 sg13g2_nand2_1 _13966_ (.Y(_05552_),
    .A(_05551_),
    .B(net92));
 sg13g2_buf_1 _13967_ (.A(\am_sdr0.cic2.comb2_in_del[9] ),
    .X(_05553_));
 sg13g2_nand2b_1 _13968_ (.Y(_05554_),
    .B(_05553_),
    .A_N(_05499_));
 sg13g2_nor2b_1 _13969_ (.A(_05553_),
    .B_N(_05499_),
    .Y(_05555_));
 sg13g2_buf_1 _13970_ (.A(\am_sdr0.cic2.comb2_in_del[8] ),
    .X(_05556_));
 sg13g2_inv_1 _13971_ (.Y(_05557_),
    .A(_05556_));
 sg13g2_inv_1 _13972_ (.Y(_05558_),
    .A(\am_sdr0.cic2.comb2_in_del[7] ));
 sg13g2_nor2_1 _13973_ (.A(_05483_),
    .B(_05558_),
    .Y(_05559_));
 sg13g2_inv_1 _13974_ (.Y(_05560_),
    .A(\am_sdr0.cic2.comb2_in_del[6] ));
 sg13g2_inv_1 _13975_ (.Y(_05561_),
    .A(_05453_));
 sg13g2_inv_1 _13976_ (.Y(_05562_),
    .A(_05448_));
 sg13g2_buf_1 _13977_ (.A(\am_sdr0.cic2.comb2_in_del[2] ),
    .X(_05563_));
 sg13g2_nor2_1 _13978_ (.A(_05562_),
    .B(_05563_),
    .Y(_05564_));
 sg13g2_nor2b_1 _13979_ (.A(_05276_),
    .B_N(\am_sdr0.cic2.comb2_in_del[0] ),
    .Y(_05565_));
 sg13g2_buf_8 _13980_ (.A(\am_sdr0.cic2.comb2_in_del[1] ),
    .X(_05566_));
 sg13g2_nand2b_1 _13981_ (.Y(_05567_),
    .B(_05442_),
    .A_N(_05566_));
 sg13g2_nor2b_1 _13982_ (.A(_05442_),
    .B_N(_05566_),
    .Y(_05568_));
 sg13g2_a221oi_1 _13983_ (.B2(_05567_),
    .C1(_05568_),
    .B1(_05565_),
    .A1(_05562_),
    .Y(_05569_),
    .A2(_05563_));
 sg13g2_buf_1 _13984_ (.A(_05569_),
    .X(_05570_));
 sg13g2_inv_1 _13985_ (.Y(_05571_),
    .A(\am_sdr0.cic2.comb2_in_del[3] ));
 sg13g2_o21ai_1 _13986_ (.B1(_05571_),
    .Y(_05572_),
    .A1(_05564_),
    .A2(_05570_));
 sg13g2_nor3_1 _13987_ (.A(_05571_),
    .B(_05564_),
    .C(_05570_),
    .Y(_05573_));
 sg13g2_a21oi_1 _13988_ (.A1(_05561_),
    .A2(_05572_),
    .Y(_05574_),
    .B1(_05573_));
 sg13g2_inv_1 _13989_ (.Y(_05575_),
    .A(_05458_));
 sg13g2_buf_1 _13990_ (.A(\am_sdr0.cic2.comb2_in_del[4] ),
    .X(_05576_));
 sg13g2_buf_1 _13991_ (.A(\am_sdr0.cic2.comb2_in_del[5] ),
    .X(_05577_));
 sg13g2_a21oi_1 _13992_ (.A1(_05575_),
    .A2(_05576_),
    .Y(_05578_),
    .B1(_05577_));
 sg13g2_inv_1 _13993_ (.Y(_05579_),
    .A(_05576_));
 sg13g2_nand2_1 _13994_ (.Y(_05580_),
    .A(_05458_),
    .B(_05579_));
 sg13g2_inv_1 _13995_ (.Y(_05581_),
    .A(_05466_));
 sg13g2_o21ai_1 _13996_ (.B1(_05581_),
    .Y(_05582_),
    .A1(_05577_),
    .A2(_05580_));
 sg13g2_a221oi_1 _13997_ (.B2(_05578_),
    .C1(_05582_),
    .B1(_05574_),
    .A1(_05476_),
    .Y(_05583_),
    .A2(_05560_));
 sg13g2_buf_1 _13998_ (.A(_05583_),
    .X(_05584_));
 sg13g2_a221oi_1 _13999_ (.B2(_05561_),
    .C1(_05573_),
    .B1(_05572_),
    .A1(_05575_),
    .Y(_05585_),
    .A2(_05576_));
 sg13g2_nand2_1 _14000_ (.Y(_05586_),
    .A(_05476_),
    .B(_05560_));
 sg13g2_nand3_1 _14001_ (.B(_05580_),
    .C(_05586_),
    .A(_05577_),
    .Y(_05587_));
 sg13g2_nand2b_1 _14002_ (.Y(_05588_),
    .B(\am_sdr0.cic2.comb2_in_del[6] ),
    .A_N(_05476_));
 sg13g2_o21ai_1 _14003_ (.B1(_05588_),
    .Y(_05589_),
    .A1(_05585_),
    .A2(_05587_));
 sg13g2_or2_1 _14004_ (.X(_05590_),
    .B(_05589_),
    .A(_05584_));
 sg13g2_buf_1 _14005_ (.A(_05590_),
    .X(_05591_));
 sg13g2_nand2_1 _14006_ (.Y(_05592_),
    .A(_05483_),
    .B(_05558_));
 sg13g2_o21ai_1 _14007_ (.B1(_05592_),
    .Y(_05593_),
    .A1(_05559_),
    .A2(_05591_));
 sg13g2_buf_2 _14008_ (.A(_05593_),
    .X(_05594_));
 sg13g2_nor2_1 _14009_ (.A(_05558_),
    .B(_05557_),
    .Y(_05595_));
 sg13g2_o21ai_1 _14010_ (.B1(_05595_),
    .Y(_05596_),
    .A1(_05584_),
    .A2(_05589_));
 sg13g2_nor2_1 _14011_ (.A(_05483_),
    .B(_05557_),
    .Y(_05597_));
 sg13g2_o21ai_1 _14012_ (.B1(_05597_),
    .Y(_05598_),
    .A1(_05584_),
    .A2(_05589_));
 sg13g2_nand2_1 _14013_ (.Y(_05599_),
    .A(_05556_),
    .B(_05559_));
 sg13g2_and4_1 _14014_ (.A(_05492_),
    .B(_05596_),
    .C(_05598_),
    .D(_05599_),
    .X(_05600_));
 sg13g2_a21oi_2 _14015_ (.B1(_05600_),
    .Y(_05601_),
    .A2(_05594_),
    .A1(_05557_));
 sg13g2_nand2b_1 _14016_ (.Y(_05602_),
    .B(_05601_),
    .A_N(_05555_));
 sg13g2_nand2_1 _14017_ (.Y(_05603_),
    .A(_05554_),
    .B(_05602_));
 sg13g2_nand2b_1 _14018_ (.Y(_05604_),
    .B(_05328_),
    .A_N(\am_sdr0.cic2.comb2_in_del[10] ));
 sg13g2_nand2b_1 _14019_ (.Y(_05605_),
    .B(\am_sdr0.cic2.comb2_in_del[10] ),
    .A_N(_05328_));
 sg13g2_buf_1 _14020_ (.A(_05605_),
    .X(_05606_));
 sg13g2_nand2_1 _14021_ (.Y(_05607_),
    .A(_05604_),
    .B(_05606_));
 sg13g2_xor2_1 _14022_ (.B(_05607_),
    .A(_05603_),
    .X(_05608_));
 sg13g2_nand2_1 _14023_ (.Y(_05609_),
    .A(_05372_),
    .B(_05608_));
 sg13g2_a21oi_1 _14024_ (.A1(_05552_),
    .A2(_05609_),
    .Y(_00662_),
    .B1(_05542_));
 sg13g2_buf_1 _14025_ (.A(\am_sdr0.cic2.comb2[11] ),
    .X(_05610_));
 sg13g2_inv_1 _14026_ (.Y(_05611_),
    .A(_05553_));
 sg13g2_nor2_1 _14027_ (.A(_05556_),
    .B(_05553_),
    .Y(_05612_));
 sg13g2_nand2b_1 _14028_ (.Y(_05613_),
    .B(_05604_),
    .A_N(_05499_));
 sg13g2_a221oi_1 _14029_ (.B2(_05594_),
    .C1(_05613_),
    .B1(_05612_),
    .A1(_05611_),
    .Y(_05614_),
    .A2(_05600_));
 sg13g2_buf_2 _14030_ (.A(_05614_),
    .X(_05615_));
 sg13g2_nand2_1 _14031_ (.Y(_05616_),
    .A(_05553_),
    .B(_05604_));
 sg13g2_buf_1 _14032_ (.A(_05616_),
    .X(_05617_));
 sg13g2_nor3_1 _14033_ (.A(_05558_),
    .B(_05557_),
    .C(_05617_),
    .Y(_05618_));
 sg13g2_nor3_1 _14034_ (.A(_05483_),
    .B(_05557_),
    .C(_05617_),
    .Y(_05619_));
 sg13g2_o21ai_1 _14035_ (.B1(_05591_),
    .Y(_05620_),
    .A1(_05618_),
    .A2(_05619_));
 sg13g2_nor3_1 _14036_ (.A(_05558_),
    .B(_05492_),
    .C(_05617_),
    .Y(_05621_));
 sg13g2_nor3_1 _14037_ (.A(_05483_),
    .B(_05492_),
    .C(_05617_),
    .Y(_05622_));
 sg13g2_o21ai_1 _14038_ (.B1(_05591_),
    .Y(_05623_),
    .A1(_05621_),
    .A2(_05622_));
 sg13g2_nand2b_1 _14039_ (.Y(_05624_),
    .B(_05556_),
    .A_N(_05492_));
 sg13g2_a21oi_1 _14040_ (.A1(_05599_),
    .A2(_05624_),
    .Y(_05625_),
    .B1(_05617_));
 sg13g2_nand2b_1 _14041_ (.Y(_05626_),
    .B(\am_sdr0.cic2.comb2_in_del[7] ),
    .A_N(_05483_));
 sg13g2_nor3_1 _14042_ (.A(_05492_),
    .B(_05626_),
    .C(_05617_),
    .Y(_05627_));
 sg13g2_nor2_1 _14043_ (.A(_05625_),
    .B(_05627_),
    .Y(_05628_));
 sg13g2_nand4_1 _14044_ (.B(_05620_),
    .C(_05623_),
    .A(_05606_),
    .Y(_05629_),
    .D(_05628_));
 sg13g2_buf_1 _14045_ (.A(_05629_),
    .X(_05630_));
 sg13g2_buf_2 _14046_ (.A(\am_sdr0.cic2.comb2_in_del[11] ),
    .X(_05631_));
 sg13g2_xnor2_1 _14047_ (.Y(_05632_),
    .A(_05350_),
    .B(_05631_));
 sg13g2_o21ai_1 _14048_ (.B1(_05632_),
    .Y(_05633_),
    .A1(_05615_),
    .A2(_05630_));
 sg13g2_or3_1 _14049_ (.A(_05615_),
    .B(_05630_),
    .C(_05632_),
    .X(_05634_));
 sg13g2_a21oi_1 _14050_ (.A1(_05633_),
    .A2(_05634_),
    .Y(_05635_),
    .B1(net155));
 sg13g2_a21oi_1 _14051_ (.A1(_05610_),
    .A2(_05467_),
    .Y(_05636_),
    .B1(_05635_));
 sg13g2_nor2_1 _14052_ (.A(net89),
    .B(_05636_),
    .Y(_00663_));
 sg13g2_buf_1 _14053_ (.A(\am_sdr0.cic2.comb2[12] ),
    .X(_05637_));
 sg13g2_o21ai_1 _14054_ (.B1(_05631_),
    .Y(_05638_),
    .A1(_05615_),
    .A2(_05630_));
 sg13g2_nor3_1 _14055_ (.A(_05631_),
    .B(_05615_),
    .C(_05630_),
    .Y(_05639_));
 sg13g2_a21o_1 _14056_ (.A2(_05638_),
    .A1(_05350_),
    .B1(_05639_),
    .X(_05640_));
 sg13g2_buf_1 _14057_ (.A(\am_sdr0.cic2.comb2_in_del[12] ),
    .X(_05641_));
 sg13g2_xnor2_1 _14058_ (.Y(_05642_),
    .A(_05353_),
    .B(_05641_));
 sg13g2_xnor2_1 _14059_ (.Y(_05643_),
    .A(_05640_),
    .B(_05642_));
 sg13g2_nand2_1 _14060_ (.Y(_05644_),
    .A(net283),
    .B(_05643_));
 sg13g2_o21ai_1 _14061_ (.B1(_05644_),
    .Y(_05645_),
    .A1(_05637_),
    .A2(net221));
 sg13g2_nor2_1 _14062_ (.A(net89),
    .B(_05645_),
    .Y(_00664_));
 sg13g2_buf_1 _14063_ (.A(\am_sdr0.cic2.comb2[13] ),
    .X(_05646_));
 sg13g2_nor2_1 _14064_ (.A(_05646_),
    .B(net224),
    .Y(_05647_));
 sg13g2_inv_1 _14065_ (.Y(_05648_),
    .A(_05617_));
 sg13g2_nor2_1 _14066_ (.A(_05631_),
    .B(_05641_),
    .Y(_05649_));
 sg13g2_nand2_1 _14067_ (.Y(_05650_),
    .A(_05606_),
    .B(_05649_));
 sg13g2_nand3b_1 _14068_ (.B(_05606_),
    .C(_05350_),
    .Y(_05651_),
    .A_N(_05641_));
 sg13g2_a221oi_1 _14069_ (.B2(_05651_),
    .C1(_05615_),
    .B1(_05650_),
    .A1(_05601_),
    .Y(_05652_),
    .A2(_05648_));
 sg13g2_inv_1 _14070_ (.Y(_05653_),
    .A(_05353_));
 sg13g2_nor4_1 _14071_ (.A(_05631_),
    .B(_05653_),
    .C(_05615_),
    .D(_05630_),
    .Y(_05654_));
 sg13g2_nand2_1 _14072_ (.Y(_05655_),
    .A(_05350_),
    .B(_05353_));
 sg13g2_nor3_1 _14073_ (.A(_05615_),
    .B(_05630_),
    .C(_05655_),
    .Y(_05656_));
 sg13g2_nand2b_1 _14074_ (.Y(_05657_),
    .B(_05350_),
    .A_N(_05631_));
 sg13g2_a21o_1 _14075_ (.A2(_05641_),
    .A1(_05653_),
    .B1(_05657_),
    .X(_05658_));
 sg13g2_o21ai_1 _14076_ (.B1(_05658_),
    .Y(_05659_),
    .A1(_05653_),
    .A2(_05641_));
 sg13g2_or4_1 _14077_ (.A(_05652_),
    .B(_05654_),
    .C(_05656_),
    .D(_05659_),
    .X(_05660_));
 sg13g2_buf_8 _14078_ (.A(_05660_),
    .X(_05661_));
 sg13g2_buf_1 _14079_ (.A(\am_sdr0.cic2.comb2_in_del[13] ),
    .X(_05662_));
 sg13g2_xor2_1 _14080_ (.B(_05662_),
    .A(_05369_),
    .X(_05663_));
 sg13g2_xnor2_1 _14081_ (.Y(_05664_),
    .A(_05661_),
    .B(_05663_));
 sg13g2_nor2_1 _14082_ (.A(net154),
    .B(_05664_),
    .Y(_05665_));
 sg13g2_nor3_1 _14083_ (.A(net160),
    .B(_05647_),
    .C(_05665_),
    .Y(_00665_));
 sg13g2_inv_1 _14084_ (.Y(_05666_),
    .A(\am_sdr0.cic2.comb2[14] ));
 sg13g2_nand2b_1 _14085_ (.Y(_05667_),
    .B(_05662_),
    .A_N(_05369_));
 sg13g2_nor2b_1 _14086_ (.A(_05662_),
    .B_N(_05369_),
    .Y(_05668_));
 sg13g2_a21oi_2 _14087_ (.B1(_05668_),
    .Y(_05669_),
    .A2(_05667_),
    .A1(_05661_));
 sg13g2_buf_2 _14088_ (.A(\am_sdr0.cic2.comb2_in_del[14] ),
    .X(_05670_));
 sg13g2_xor2_1 _14089_ (.B(_05670_),
    .A(_05384_),
    .X(_05671_));
 sg13g2_xnor2_1 _14090_ (.Y(_05672_),
    .A(_05669_),
    .B(_05671_));
 sg13g2_mux2_1 _14091_ (.A0(_05666_),
    .A1(_05672_),
    .S(net283),
    .X(_05673_));
 sg13g2_nor2_1 _14092_ (.A(_05491_),
    .B(_05673_),
    .Y(_00666_));
 sg13g2_nand2_1 _14093_ (.Y(_05674_),
    .A(_05670_),
    .B(_05669_));
 sg13g2_inv_1 _14094_ (.Y(_05675_),
    .A(_05384_));
 sg13g2_o21ai_1 _14095_ (.B1(_05675_),
    .Y(_05676_),
    .A1(_05670_),
    .A2(_05669_));
 sg13g2_nand2_1 _14096_ (.Y(_05677_),
    .A(_05674_),
    .B(_05676_));
 sg13g2_buf_1 _14097_ (.A(\am_sdr0.cic2.comb2_in_del[15] ),
    .X(_05678_));
 sg13g2_xor2_1 _14098_ (.B(_05678_),
    .A(_05391_),
    .X(_05679_));
 sg13g2_xnor2_1 _14099_ (.Y(_05680_),
    .A(_05677_),
    .B(_05679_));
 sg13g2_buf_1 _14100_ (.A(\am_sdr0.cic2.comb2[15] ),
    .X(_05681_));
 sg13g2_o21ai_1 _14101_ (.B1(net218),
    .Y(_05682_),
    .A1(_05681_),
    .A2(net224));
 sg13g2_a21oi_1 _14102_ (.A1(net225),
    .A2(_05680_),
    .Y(_00667_),
    .B1(_05682_));
 sg13g2_buf_1 _14103_ (.A(\am_sdr0.cic2.comb2[16] ),
    .X(_05683_));
 sg13g2_nand2_1 _14104_ (.Y(_05684_),
    .A(_05683_),
    .B(_05357_));
 sg13g2_inv_1 _14105_ (.Y(_05685_),
    .A(_05678_));
 sg13g2_nor2_1 _14106_ (.A(_05391_),
    .B(_05685_),
    .Y(_05686_));
 sg13g2_nand2_1 _14107_ (.Y(_05687_),
    .A(_05670_),
    .B(_05678_));
 sg13g2_nand2_1 _14108_ (.Y(_05688_),
    .A(_05675_),
    .B(_05678_));
 sg13g2_a221oi_1 _14109_ (.B2(_05688_),
    .C1(_05668_),
    .B1(_05687_),
    .A1(_05661_),
    .Y(_05689_),
    .A2(_05667_));
 sg13g2_nand2b_1 _14110_ (.Y(_05690_),
    .B(_05670_),
    .A_N(_05391_));
 sg13g2_or2_1 _14111_ (.X(_05691_),
    .B(_05391_),
    .A(_05384_));
 sg13g2_a221oi_1 _14112_ (.B2(_05691_),
    .C1(_05668_),
    .B1(_05690_),
    .A1(_05661_),
    .Y(_05692_),
    .A2(_05667_));
 sg13g2_nand2_1 _14113_ (.Y(_05693_),
    .A(_05675_),
    .B(_05670_));
 sg13g2_a21oi_1 _14114_ (.A1(_05391_),
    .A2(_05685_),
    .Y(_05694_),
    .B1(_05693_));
 sg13g2_nor4_2 _14115_ (.A(_05686_),
    .B(_05689_),
    .C(_05692_),
    .Y(_05695_),
    .D(_05694_));
 sg13g2_buf_1 _14116_ (.A(\am_sdr0.cic2.comb2_in_del[16] ),
    .X(_05696_));
 sg13g2_xor2_1 _14117_ (.B(_05696_),
    .A(_05404_),
    .X(_05697_));
 sg13g2_xnor2_1 _14118_ (.Y(_05698_),
    .A(_05695_),
    .B(_05697_));
 sg13g2_nand2_1 _14119_ (.Y(_05699_),
    .A(net222),
    .B(_05698_));
 sg13g2_a21oi_1 _14120_ (.A1(_05684_),
    .A2(_05699_),
    .Y(_00668_),
    .B1(_05542_));
 sg13g2_xnor2_1 _14121_ (.Y(_05700_),
    .A(_05412_),
    .B(\am_sdr0.cic2.comb2_in_del[17] ));
 sg13g2_inv_1 _14122_ (.Y(_05701_),
    .A(_05404_));
 sg13g2_a21oi_1 _14123_ (.A1(_05674_),
    .A2(_05676_),
    .Y(_05702_),
    .B1(_05685_));
 sg13g2_inv_1 _14124_ (.Y(_05703_),
    .A(_05696_));
 sg13g2_nor2_1 _14125_ (.A(_05703_),
    .B(_05695_),
    .Y(_05704_));
 sg13g2_a21oi_1 _14126_ (.A1(_05701_),
    .A2(_05702_),
    .Y(_05705_),
    .B1(_05704_));
 sg13g2_or2_1 _14127_ (.X(_05706_),
    .B(_05705_),
    .A(_05700_));
 sg13g2_nor3_1 _14128_ (.A(_05391_),
    .B(_05404_),
    .C(_05700_),
    .Y(_05707_));
 sg13g2_a21oi_1 _14129_ (.A1(_05703_),
    .A2(_05695_),
    .Y(_05708_),
    .B1(_05404_));
 sg13g2_nor2_1 _14130_ (.A(_05704_),
    .B(_05708_),
    .Y(_05709_));
 sg13g2_inv_1 _14131_ (.Y(_00826_),
    .A(_05436_));
 sg13g2_nor2_1 _14132_ (.A(_05404_),
    .B(_05700_),
    .Y(_05710_));
 sg13g2_o21ai_1 _14133_ (.B1(_05710_),
    .Y(_05711_),
    .A1(_05696_),
    .A2(_05686_));
 sg13g2_nand2_1 _14134_ (.Y(_05712_),
    .A(_00826_),
    .B(_05711_));
 sg13g2_a221oi_1 _14135_ (.B2(_05700_),
    .C1(_05712_),
    .B1(_05709_),
    .A1(_05677_),
    .Y(_05713_),
    .A2(_05707_));
 sg13g2_buf_1 _14136_ (.A(\am_sdr0.cic2.comb2[17] ),
    .X(_05714_));
 sg13g2_and3_1 _14137_ (.X(_05715_),
    .A(net297),
    .B(_05714_),
    .C(_05358_));
 sg13g2_a21o_1 _14138_ (.A2(_05713_),
    .A1(_05706_),
    .B1(_05715_),
    .X(_00669_));
 sg13g2_buf_1 _14139_ (.A(\am_sdr0.cic2.comb2[18] ),
    .X(_05716_));
 sg13g2_nand2_1 _14140_ (.Y(_05717_),
    .A(net253),
    .B(_05716_));
 sg13g2_nand2b_1 _14141_ (.Y(_05718_),
    .B(\am_sdr0.cic2.comb2_in_del[18] ),
    .A_N(_05423_));
 sg13g2_nand2b_1 _14142_ (.Y(_05719_),
    .B(_05423_),
    .A_N(\am_sdr0.cic2.comb2_in_del[18] ));
 sg13g2_nand2_1 _14143_ (.Y(_05720_),
    .A(_05718_),
    .B(_05719_));
 sg13g2_nand2b_1 _14144_ (.Y(_05721_),
    .B(_00826_),
    .A_N(_05720_));
 sg13g2_nand2_1 _14145_ (.Y(_05722_),
    .A(_00826_),
    .B(_05720_));
 sg13g2_inv_1 _14146_ (.Y(_05723_),
    .A(\am_sdr0.cic2.comb2_in_del[17] ));
 sg13g2_nor2_1 _14147_ (.A(_05412_),
    .B(_05723_),
    .Y(_05724_));
 sg13g2_a221oi_1 _14148_ (.B2(_05723_),
    .C1(_05695_),
    .B1(_05412_),
    .A1(_05404_),
    .Y(_05725_),
    .A2(_05703_));
 sg13g2_nand2_1 _14149_ (.Y(_05726_),
    .A(_05701_),
    .B(_05696_));
 sg13g2_a21oi_1 _14150_ (.A1(_05412_),
    .A2(_05723_),
    .Y(_05727_),
    .B1(_05726_));
 sg13g2_nor3_2 _14151_ (.A(_05724_),
    .B(_05725_),
    .C(_05727_),
    .Y(_05728_));
 sg13g2_mux2_1 _14152_ (.A0(_05721_),
    .A1(_05722_),
    .S(_05728_),
    .X(_05729_));
 sg13g2_o21ai_1 _14153_ (.B1(_05729_),
    .Y(_00670_),
    .A1(_05274_),
    .A2(_05717_));
 sg13g2_xnor2_1 _14154_ (.Y(_05730_),
    .A(\am_sdr0.cic2.comb1[19] ),
    .B(\am_sdr0.cic2.comb2_in_del[19] ));
 sg13g2_mux2_1 _14155_ (.A0(_05718_),
    .A1(_05719_),
    .S(_05730_),
    .X(_05731_));
 sg13g2_nor2b_1 _14156_ (.A(net284),
    .B_N(\am_sdr0.cic2.comb2[19] ),
    .Y(_05732_));
 sg13g2_a21oi_1 _14157_ (.A1(net283),
    .A2(_05731_),
    .Y(_05733_),
    .B1(_05732_));
 sg13g2_nand2_1 _14158_ (.Y(_05734_),
    .A(net284),
    .B(_05719_));
 sg13g2_nor3_1 _14159_ (.A(_05728_),
    .B(_05730_),
    .C(_05734_),
    .Y(_05735_));
 sg13g2_and4_1 _14160_ (.A(net285),
    .B(_05728_),
    .C(_05718_),
    .D(_05730_),
    .X(_05736_));
 sg13g2_nor4_1 _14161_ (.A(net191),
    .B(_05733_),
    .C(_05735_),
    .D(_05736_),
    .Y(_00671_));
 sg13g2_nand2_1 _14162_ (.Y(_05737_),
    .A(\am_sdr0.cic2.comb2[1] ),
    .B(net93));
 sg13g2_xnor2_1 _14163_ (.Y(_05738_),
    .A(_05442_),
    .B(_05566_));
 sg13g2_xnor2_1 _14164_ (.Y(_05739_),
    .A(_05565_),
    .B(_05738_));
 sg13g2_nand2_1 _14165_ (.Y(_05740_),
    .A(net222),
    .B(_05739_));
 sg13g2_a21oi_1 _14166_ (.A1(_05737_),
    .A2(_05740_),
    .Y(_00672_),
    .B1(net86));
 sg13g2_buf_1 _14167_ (.A(\am_sdr0.cic2.comb2[2] ),
    .X(_05741_));
 sg13g2_nand2_1 _14168_ (.Y(_05742_),
    .A(_05741_),
    .B(net93));
 sg13g2_a21oi_1 _14169_ (.A1(_05565_),
    .A2(_05567_),
    .Y(_05743_),
    .B1(_05568_));
 sg13g2_xor2_1 _14170_ (.B(_05563_),
    .A(_05448_),
    .X(_05744_));
 sg13g2_xnor2_1 _14171_ (.Y(_05745_),
    .A(_05743_),
    .B(_05744_));
 sg13g2_nand2_1 _14172_ (.Y(_05746_),
    .A(net222),
    .B(_05745_));
 sg13g2_a21oi_1 _14173_ (.A1(_05742_),
    .A2(_05746_),
    .Y(_00673_),
    .B1(net86));
 sg13g2_buf_1 _14174_ (.A(\am_sdr0.cic2.comb2[3] ),
    .X(_05747_));
 sg13g2_nand2_1 _14175_ (.Y(_05748_),
    .A(_05747_),
    .B(net93));
 sg13g2_nor2_1 _14176_ (.A(_05564_),
    .B(_05570_),
    .Y(_05749_));
 sg13g2_xnor2_1 _14177_ (.Y(_05750_),
    .A(_05453_),
    .B(\am_sdr0.cic2.comb2_in_del[3] ));
 sg13g2_xnor2_1 _14178_ (.Y(_05751_),
    .A(_05749_),
    .B(_05750_));
 sg13g2_nand2_1 _14179_ (.Y(_05752_),
    .A(net222),
    .B(_05751_));
 sg13g2_a21oi_1 _14180_ (.A1(_05748_),
    .A2(_05752_),
    .Y(_00674_),
    .B1(net86));
 sg13g2_buf_1 _14181_ (.A(\am_sdr0.cic2.comb2[4] ),
    .X(_05753_));
 sg13g2_nor2_1 _14182_ (.A(_05753_),
    .B(net224),
    .Y(_05754_));
 sg13g2_nand2_1 _14183_ (.Y(_05755_),
    .A(_05575_),
    .B(_05576_));
 sg13g2_nand2_1 _14184_ (.Y(_05756_),
    .A(_05580_),
    .B(_05755_));
 sg13g2_xnor2_1 _14185_ (.Y(_05757_),
    .A(_05574_),
    .B(_05756_));
 sg13g2_nor2_1 _14186_ (.A(net154),
    .B(_05757_),
    .Y(_05758_));
 sg13g2_nor3_1 _14187_ (.A(net160),
    .B(_05754_),
    .C(_05758_),
    .Y(_00675_));
 sg13g2_buf_1 _14188_ (.A(\am_sdr0.cic2.comb2[5] ),
    .X(_05759_));
 sg13g2_nand2_1 _14189_ (.Y(_05760_),
    .A(_05759_),
    .B(net93));
 sg13g2_a21oi_1 _14190_ (.A1(_05458_),
    .A2(_05579_),
    .Y(_05761_),
    .B1(_05585_));
 sg13g2_xnor2_1 _14191_ (.Y(_05762_),
    .A(_05466_),
    .B(_05577_));
 sg13g2_xnor2_1 _14192_ (.Y(_05763_),
    .A(_05761_),
    .B(_05762_));
 sg13g2_nand2_1 _14193_ (.Y(_05764_),
    .A(net221),
    .B(_05763_));
 sg13g2_a21oi_1 _14194_ (.A1(_05760_),
    .A2(_05764_),
    .Y(_00676_),
    .B1(net86));
 sg13g2_a21oi_1 _14195_ (.A1(_05574_),
    .A2(_05578_),
    .Y(_05765_),
    .B1(_05582_));
 sg13g2_a21oi_1 _14196_ (.A1(_05577_),
    .A2(_05761_),
    .Y(_05766_),
    .B1(_05765_));
 sg13g2_nand2_1 _14197_ (.Y(_05767_),
    .A(_05586_),
    .B(_05588_));
 sg13g2_xnor2_1 _14198_ (.Y(_05768_),
    .A(_05766_),
    .B(_05767_));
 sg13g2_buf_1 _14199_ (.A(\am_sdr0.cic2.comb2[6] ),
    .X(_05769_));
 sg13g2_nor2b_1 _14200_ (.A(net285),
    .B_N(_05769_),
    .Y(_05770_));
 sg13g2_a21oi_1 _14201_ (.A1(_05280_),
    .A2(_05768_),
    .Y(_05771_),
    .B1(_05770_));
 sg13g2_nor2_1 _14202_ (.A(net89),
    .B(_05771_),
    .Y(_00677_));
 sg13g2_buf_1 _14203_ (.A(\am_sdr0.cic2.comb2[7] ),
    .X(_05772_));
 sg13g2_nand2_1 _14204_ (.Y(_05773_),
    .A(_05772_),
    .B(net93));
 sg13g2_nand2_1 _14205_ (.Y(_05774_),
    .A(_05626_),
    .B(_05592_));
 sg13g2_xor2_1 _14206_ (.B(_05774_),
    .A(_05591_),
    .X(_05775_));
 sg13g2_nand2_1 _14207_ (.Y(_05776_),
    .A(net221),
    .B(_05775_));
 sg13g2_a21oi_1 _14208_ (.A1(_05773_),
    .A2(_05776_),
    .Y(_00678_),
    .B1(net86));
 sg13g2_buf_1 _14209_ (.A(\am_sdr0.cic2.comb2[8] ),
    .X(_05777_));
 sg13g2_nor2_1 _14210_ (.A(_05777_),
    .B(net224),
    .Y(_05778_));
 sg13g2_xor2_1 _14211_ (.B(_05556_),
    .A(_05492_),
    .X(_05779_));
 sg13g2_xnor2_1 _14212_ (.Y(_05780_),
    .A(_05594_),
    .B(_05779_));
 sg13g2_nor2_1 _14213_ (.A(net154),
    .B(_05780_),
    .Y(_05781_));
 sg13g2_nor3_1 _14214_ (.A(_04198_),
    .B(_05778_),
    .C(_05781_),
    .Y(_00679_));
 sg13g2_nor2b_1 _14215_ (.A(_05555_),
    .B_N(_05554_),
    .Y(_05782_));
 sg13g2_xnor2_1 _14216_ (.Y(_05783_),
    .A(_05601_),
    .B(_05782_));
 sg13g2_buf_1 _14217_ (.A(\am_sdr0.cic2.comb2[9] ),
    .X(_05784_));
 sg13g2_nor2b_1 _14218_ (.A(net285),
    .B_N(_05784_),
    .Y(_05785_));
 sg13g2_a21oi_1 _14219_ (.A1(_05280_),
    .A2(_05783_),
    .Y(_05786_),
    .B1(_05785_));
 sg13g2_nor2_1 _14220_ (.A(net89),
    .B(_05786_),
    .Y(_00680_));
 sg13g2_buf_1 _14221_ (.A(net285),
    .X(_05787_));
 sg13g2_nand2_1 _14222_ (.Y(_05788_),
    .A(_05276_),
    .B(net217));
 sg13g2_nand2_1 _14223_ (.Y(_05789_),
    .A(\am_sdr0.cic2.comb2_in_del[0] ),
    .B(net85));
 sg13g2_buf_1 _14224_ (.A(_04696_),
    .X(_05790_));
 sg13g2_a21oi_1 _14225_ (.A1(_05788_),
    .A2(_05789_),
    .Y(_00681_),
    .B1(net84));
 sg13g2_nand2_1 _14226_ (.Y(_05791_),
    .A(_05328_),
    .B(net217));
 sg13g2_nand2_1 _14227_ (.Y(_05792_),
    .A(\am_sdr0.cic2.comb2_in_del[10] ),
    .B(net85));
 sg13g2_a21oi_1 _14228_ (.A1(_05791_),
    .A2(_05792_),
    .Y(_00682_),
    .B1(net84));
 sg13g2_nand2_1 _14229_ (.Y(_05793_),
    .A(_05350_),
    .B(net217));
 sg13g2_nand2_1 _14230_ (.Y(_05794_),
    .A(_05631_),
    .B(net85));
 sg13g2_a21oi_1 _14231_ (.A1(_05793_),
    .A2(_05794_),
    .Y(_00683_),
    .B1(net84));
 sg13g2_nand2_1 _14232_ (.Y(_05795_),
    .A(_05353_),
    .B(net217));
 sg13g2_nand2_1 _14233_ (.Y(_05796_),
    .A(_05641_),
    .B(net85));
 sg13g2_a21oi_1 _14234_ (.A1(_05795_),
    .A2(_05796_),
    .Y(_00684_),
    .B1(net84));
 sg13g2_nand2_1 _14235_ (.Y(_05797_),
    .A(_05369_),
    .B(net217));
 sg13g2_nand2_1 _14236_ (.Y(_05798_),
    .A(_05662_),
    .B(net85));
 sg13g2_a21oi_1 _14237_ (.A1(_05797_),
    .A2(_05798_),
    .Y(_00685_),
    .B1(net84));
 sg13g2_nand2_1 _14238_ (.Y(_05799_),
    .A(_05384_),
    .B(net217));
 sg13g2_nand2_1 _14239_ (.Y(_05800_),
    .A(_05670_),
    .B(net85));
 sg13g2_a21oi_1 _14240_ (.A1(_05799_),
    .A2(_05800_),
    .Y(_00686_),
    .B1(net84));
 sg13g2_nand2_1 _14241_ (.Y(_05801_),
    .A(_05391_),
    .B(_05787_));
 sg13g2_nand2_1 _14242_ (.Y(_05802_),
    .A(_05678_),
    .B(_05544_));
 sg13g2_a21oi_1 _14243_ (.A1(_05801_),
    .A2(_05802_),
    .Y(_00687_),
    .B1(_05790_));
 sg13g2_nand2_1 _14244_ (.Y(_05803_),
    .A(_05404_),
    .B(net217));
 sg13g2_nand2_1 _14245_ (.Y(_05804_),
    .A(_05696_),
    .B(_05544_));
 sg13g2_a21oi_1 _14246_ (.A1(_05803_),
    .A2(_05804_),
    .Y(_00688_),
    .B1(net84));
 sg13g2_nand2_1 _14247_ (.Y(_05805_),
    .A(_05412_),
    .B(net217));
 sg13g2_buf_1 _14248_ (.A(net155),
    .X(_05806_));
 sg13g2_nand2_1 _14249_ (.Y(_05807_),
    .A(\am_sdr0.cic2.comb2_in_del[17] ),
    .B(_05806_));
 sg13g2_a21oi_1 _14250_ (.A1(_05805_),
    .A2(_05807_),
    .Y(_00689_),
    .B1(net84));
 sg13g2_nand2_1 _14251_ (.Y(_05808_),
    .A(_05423_),
    .B(_05787_));
 sg13g2_nand2_1 _14252_ (.Y(_05809_),
    .A(\am_sdr0.cic2.comb2_in_del[18] ),
    .B(_05806_));
 sg13g2_a21oi_1 _14253_ (.A1(_05808_),
    .A2(_05809_),
    .Y(_00690_),
    .B1(_05790_));
 sg13g2_buf_1 _14254_ (.A(net284),
    .X(_05810_));
 sg13g2_nand2_1 _14255_ (.Y(_05811_),
    .A(\am_sdr0.cic2.comb1[19] ),
    .B(_05810_));
 sg13g2_nand2_1 _14256_ (.Y(_05812_),
    .A(\am_sdr0.cic2.comb2_in_del[19] ),
    .B(net83));
 sg13g2_buf_1 _14257_ (.A(_02778_),
    .X(_05813_));
 sg13g2_buf_1 _14258_ (.A(_05813_),
    .X(_05814_));
 sg13g2_a21oi_1 _14259_ (.A1(_05811_),
    .A2(_05812_),
    .Y(_00691_),
    .B1(_05814_));
 sg13g2_nand2_1 _14260_ (.Y(_05815_),
    .A(_05442_),
    .B(net216));
 sg13g2_nand2_1 _14261_ (.Y(_05816_),
    .A(_05566_),
    .B(net83));
 sg13g2_a21oi_1 _14262_ (.A1(_05815_),
    .A2(_05816_),
    .Y(_00692_),
    .B1(net82));
 sg13g2_nand2_1 _14263_ (.Y(_05817_),
    .A(_05448_),
    .B(net216));
 sg13g2_nand2_1 _14264_ (.Y(_05818_),
    .A(_05563_),
    .B(net83));
 sg13g2_a21oi_1 _14265_ (.A1(_05817_),
    .A2(_05818_),
    .Y(_00693_),
    .B1(net82));
 sg13g2_nand2_1 _14266_ (.Y(_05819_),
    .A(_05453_),
    .B(net216));
 sg13g2_nand2_1 _14267_ (.Y(_05820_),
    .A(\am_sdr0.cic2.comb2_in_del[3] ),
    .B(net83));
 sg13g2_a21oi_1 _14268_ (.A1(_05819_),
    .A2(_05820_),
    .Y(_00694_),
    .B1(net82));
 sg13g2_nand2_1 _14269_ (.Y(_05821_),
    .A(_05458_),
    .B(net216));
 sg13g2_nand2_1 _14270_ (.Y(_05822_),
    .A(_05576_),
    .B(net83));
 sg13g2_a21oi_1 _14271_ (.A1(_05821_),
    .A2(_05822_),
    .Y(_00695_),
    .B1(net82));
 sg13g2_nand2_1 _14272_ (.Y(_05823_),
    .A(_05466_),
    .B(net216));
 sg13g2_nand2_1 _14273_ (.Y(_05824_),
    .A(_05577_),
    .B(net83));
 sg13g2_a21oi_1 _14274_ (.A1(_05823_),
    .A2(_05824_),
    .Y(_00696_),
    .B1(net82));
 sg13g2_nand2_1 _14275_ (.Y(_05825_),
    .A(_05476_),
    .B(net216));
 sg13g2_nand2_1 _14276_ (.Y(_05826_),
    .A(\am_sdr0.cic2.comb2_in_del[6] ),
    .B(net83));
 sg13g2_a21oi_1 _14277_ (.A1(_05825_),
    .A2(_05826_),
    .Y(_00697_),
    .B1(net82));
 sg13g2_nand2_1 _14278_ (.Y(_05827_),
    .A(_05483_),
    .B(_05810_));
 sg13g2_nand2_1 _14279_ (.Y(_05828_),
    .A(\am_sdr0.cic2.comb2_in_del[7] ),
    .B(net83));
 sg13g2_a21oi_1 _14280_ (.A1(_05827_),
    .A2(_05828_),
    .Y(_00698_),
    .B1(_05814_));
 sg13g2_nand2_1 _14281_ (.Y(_05829_),
    .A(_05492_),
    .B(net216));
 sg13g2_buf_1 _14282_ (.A(_05355_),
    .X(_05830_));
 sg13g2_nand2_1 _14283_ (.Y(_05831_),
    .A(_05556_),
    .B(net153));
 sg13g2_a21oi_1 _14284_ (.A1(_05829_),
    .A2(_05831_),
    .Y(_00699_),
    .B1(net82));
 sg13g2_nand2_1 _14285_ (.Y(_05832_),
    .A(_05499_),
    .B(net216));
 sg13g2_nand2_1 _14286_ (.Y(_05833_),
    .A(_05553_),
    .B(net153));
 sg13g2_a21oi_1 _14287_ (.A1(_05832_),
    .A2(_05833_),
    .Y(_00700_),
    .B1(net82));
 sg13g2_nand2_1 _14288_ (.Y(_05834_),
    .A(_05370_),
    .B(\am_sdr0.cic2.comb3[12] ));
 sg13g2_inv_1 _14289_ (.Y(_05835_),
    .A(\am_sdr0.cic2.comb3_in_del[2] ));
 sg13g2_inv_1 _14290_ (.Y(_05836_),
    .A(\am_sdr0.cic2.comb2[1] ));
 sg13g2_nor2b_1 _14291_ (.A(\am_sdr0.cic2.comb2[0] ),
    .B_N(\am_sdr0.cic2.comb3_in_del[0] ),
    .Y(_05837_));
 sg13g2_nand2_1 _14292_ (.Y(_05838_),
    .A(_05836_),
    .B(_05837_));
 sg13g2_o21ai_1 _14293_ (.B1(\am_sdr0.cic2.comb3_in_del[1] ),
    .Y(_05839_),
    .A1(_05836_),
    .A2(_05837_));
 sg13g2_a22oi_1 _14294_ (.Y(_05840_),
    .B1(_05838_),
    .B2(_05839_),
    .A2(_05741_),
    .A1(_05835_));
 sg13g2_nand2b_1 _14295_ (.Y(_05841_),
    .B(\am_sdr0.cic2.comb3_in_del[3] ),
    .A_N(_05747_));
 sg13g2_o21ai_1 _14296_ (.B1(_05841_),
    .Y(_05842_),
    .A1(_05835_),
    .A2(_05741_));
 sg13g2_nand2b_1 _14297_ (.Y(_05843_),
    .B(_05747_),
    .A_N(\am_sdr0.cic2.comb3_in_del[3] ));
 sg13g2_o21ai_1 _14298_ (.B1(_05843_),
    .Y(_05844_),
    .A1(_05840_),
    .A2(_05842_));
 sg13g2_nand2_1 _14299_ (.Y(_05845_),
    .A(_05753_),
    .B(_05844_));
 sg13g2_inv_1 _14300_ (.Y(_05846_),
    .A(\am_sdr0.cic2.comb3_in_del[4] ));
 sg13g2_o21ai_1 _14301_ (.B1(_05846_),
    .Y(_05847_),
    .A1(_05753_),
    .A2(_05844_));
 sg13g2_inv_1 _14302_ (.Y(_05848_),
    .A(\am_sdr0.cic2.comb3_in_del[5] ));
 sg13g2_nor2_1 _14303_ (.A(_05848_),
    .B(_05759_),
    .Y(_05849_));
 sg13g2_a21o_1 _14304_ (.A2(_05847_),
    .A1(_05845_),
    .B1(_05849_),
    .X(_05850_));
 sg13g2_a21oi_1 _14305_ (.A1(_05848_),
    .A2(_05759_),
    .Y(_05851_),
    .B1(_05769_));
 sg13g2_o21ai_1 _14306_ (.B1(_05844_),
    .Y(_05852_),
    .A1(_05846_),
    .A2(_05753_));
 sg13g2_a22oi_1 _14307_ (.Y(_05853_),
    .B1(_05846_),
    .B2(_05753_),
    .A2(_05759_),
    .A1(_05848_));
 sg13g2_a21o_1 _14308_ (.A2(_05853_),
    .A1(_05852_),
    .B1(_05849_),
    .X(_05854_));
 sg13g2_inv_1 _14309_ (.Y(_05855_),
    .A(\am_sdr0.cic2.comb3_in_del[6] ));
 sg13g2_nand2b_1 _14310_ (.Y(_05856_),
    .B(\am_sdr0.cic2.comb3_in_del[7] ),
    .A_N(_05772_));
 sg13g2_o21ai_1 _14311_ (.B1(_05856_),
    .Y(_05857_),
    .A1(_05855_),
    .A2(_05769_));
 sg13g2_a221oi_1 _14312_ (.B2(\am_sdr0.cic2.comb3_in_del[6] ),
    .C1(_05857_),
    .B1(_05854_),
    .A1(_05850_),
    .Y(_05858_),
    .A2(_05851_));
 sg13g2_buf_1 _14313_ (.A(_05858_),
    .X(_05859_));
 sg13g2_nor2b_1 _14314_ (.A(\am_sdr0.cic2.comb3_in_del[7] ),
    .B_N(_05772_),
    .Y(_05860_));
 sg13g2_xnor2_1 _14315_ (.Y(_05861_),
    .A(\am_sdr0.cic2.comb3_in_del[10] ),
    .B(_05551_));
 sg13g2_xnor2_1 _14316_ (.Y(_05862_),
    .A(\am_sdr0.cic2.comb3_in_del[9] ),
    .B(_05784_));
 sg13g2_xnor2_1 _14317_ (.Y(_05863_),
    .A(\am_sdr0.cic2.comb3_in_del[8] ),
    .B(_05777_));
 sg13g2_nand3_1 _14318_ (.B(_05862_),
    .C(_05863_),
    .A(_05861_),
    .Y(_05864_));
 sg13g2_buf_1 _14319_ (.A(_05864_),
    .X(_05865_));
 sg13g2_inv_1 _14320_ (.Y(_05866_),
    .A(_05865_));
 sg13g2_o21ai_1 _14321_ (.B1(_05866_),
    .Y(_05867_),
    .A1(_05859_),
    .A2(_05860_));
 sg13g2_inv_1 _14322_ (.Y(_05868_),
    .A(\am_sdr0.cic2.comb3_in_del[11] ));
 sg13g2_nor2b_1 _14323_ (.A(\am_sdr0.cic2.comb3_in_del[8] ),
    .B_N(_05777_),
    .Y(_05869_));
 sg13g2_nor2_1 _14324_ (.A(_05784_),
    .B(_05869_),
    .Y(_05870_));
 sg13g2_nand2_1 _14325_ (.Y(_05871_),
    .A(_05784_),
    .B(_05869_));
 sg13g2_o21ai_1 _14326_ (.B1(_05871_),
    .Y(_05872_),
    .A1(\am_sdr0.cic2.comb3_in_del[9] ),
    .A2(_05870_));
 sg13g2_nor2_1 _14327_ (.A(_05551_),
    .B(_05872_),
    .Y(_05873_));
 sg13g2_nor2_1 _14328_ (.A(\am_sdr0.cic2.comb3_in_del[10] ),
    .B(_05873_),
    .Y(_05874_));
 sg13g2_a221oi_1 _14329_ (.B2(_05872_),
    .C1(_05874_),
    .B1(_05551_),
    .A1(_05868_),
    .Y(_05875_),
    .A2(_05610_));
 sg13g2_nor2_1 _14330_ (.A(_05868_),
    .B(_05610_),
    .Y(_05876_));
 sg13g2_a21oi_1 _14331_ (.A1(_05867_),
    .A2(_05875_),
    .Y(_05877_),
    .B1(_05876_));
 sg13g2_buf_1 _14332_ (.A(\am_sdr0.cic2.comb3_in_del[12] ),
    .X(_05878_));
 sg13g2_xor2_1 _14333_ (.B(_05878_),
    .A(_05637_),
    .X(_05879_));
 sg13g2_xnor2_1 _14334_ (.Y(_05880_),
    .A(_05877_),
    .B(_05879_));
 sg13g2_nand2_1 _14335_ (.Y(_05881_),
    .A(net221),
    .B(_05880_));
 sg13g2_buf_1 _14336_ (.A(_05813_),
    .X(_05882_));
 sg13g2_a21oi_1 _14337_ (.A1(_05834_),
    .A2(_05881_),
    .Y(_00701_),
    .B1(net81));
 sg13g2_nand2_1 _14338_ (.Y(_05883_),
    .A(net92),
    .B(\am_sdr0.cic2.comb3[13] ));
 sg13g2_nor3_1 _14339_ (.A(_05878_),
    .B(_05865_),
    .C(_05876_),
    .Y(_05884_));
 sg13g2_o21ai_1 _14340_ (.B1(_05884_),
    .Y(_05885_),
    .A1(_05859_),
    .A2(_05860_));
 sg13g2_inv_1 _14341_ (.Y(_05886_),
    .A(_05637_));
 sg13g2_nor3_1 _14342_ (.A(_05886_),
    .B(_05865_),
    .C(_05876_),
    .Y(_05887_));
 sg13g2_o21ai_1 _14343_ (.B1(_05887_),
    .Y(_05888_),
    .A1(_05859_),
    .A2(_05860_));
 sg13g2_inv_1 _14344_ (.Y(_05889_),
    .A(_05878_));
 sg13g2_inv_1 _14345_ (.Y(_05890_),
    .A(_05610_));
 sg13g2_a221oi_1 _14346_ (.B2(_05890_),
    .C1(_05875_),
    .B1(\am_sdr0.cic2.comb3_in_del[11] ),
    .A1(_05886_),
    .Y(_05891_),
    .A2(_05878_));
 sg13g2_a21oi_1 _14347_ (.A1(_05637_),
    .A2(_05889_),
    .Y(_05892_),
    .B1(_05891_));
 sg13g2_and3_1 _14348_ (.X(_05893_),
    .A(_05885_),
    .B(_05888_),
    .C(_05892_));
 sg13g2_buf_1 _14349_ (.A(_05893_),
    .X(_05894_));
 sg13g2_buf_1 _14350_ (.A(\am_sdr0.cic2.comb3_in_del[13] ),
    .X(_05895_));
 sg13g2_xnor2_1 _14351_ (.Y(_05896_),
    .A(_05646_),
    .B(_05895_));
 sg13g2_xnor2_1 _14352_ (.Y(_05897_),
    .A(_05894_),
    .B(_05896_));
 sg13g2_nand2_1 _14353_ (.Y(_05898_),
    .A(net221),
    .B(_05897_));
 sg13g2_a21oi_1 _14354_ (.A1(_05883_),
    .A2(_05898_),
    .Y(_00702_),
    .B1(net81));
 sg13g2_inv_1 _14355_ (.Y(_05899_),
    .A(_05895_));
 sg13g2_nand3_1 _14356_ (.B(_05888_),
    .C(_05892_),
    .A(_05885_),
    .Y(_05900_));
 sg13g2_a21oi_1 _14357_ (.A1(_05899_),
    .A2(_05900_),
    .Y(_05901_),
    .B1(_05646_));
 sg13g2_a21oi_1 _14358_ (.A1(_05895_),
    .A2(_05894_),
    .Y(_05902_),
    .B1(_05901_));
 sg13g2_nor2_1 _14359_ (.A(_05666_),
    .B(\am_sdr0.cic2.comb3_in_del[14] ),
    .Y(_05903_));
 sg13g2_nand2_1 _14360_ (.Y(_05904_),
    .A(_05666_),
    .B(\am_sdr0.cic2.comb3_in_del[14] ));
 sg13g2_nand2b_1 _14361_ (.Y(_05905_),
    .B(_05904_),
    .A_N(_05903_));
 sg13g2_xnor2_1 _14362_ (.Y(_05906_),
    .A(_05902_),
    .B(_05905_));
 sg13g2_nor2b_1 _14363_ (.A(net285),
    .B_N(\am_sdr0.cic2.comb3[14] ),
    .Y(_05907_));
 sg13g2_a21oi_1 _14364_ (.A1(net223),
    .A2(_05906_),
    .Y(_05908_),
    .B1(_05907_));
 sg13g2_nor2_1 _14365_ (.A(net89),
    .B(_05908_),
    .Y(_00703_));
 sg13g2_a21oi_1 _14366_ (.A1(_05646_),
    .A2(_05899_),
    .Y(_05909_),
    .B1(_05903_));
 sg13g2_nand2b_1 _14367_ (.Y(_05910_),
    .B(_05895_),
    .A_N(_05646_));
 sg13g2_o21ai_1 _14368_ (.B1(_05904_),
    .Y(_05911_),
    .A1(_05910_),
    .A2(_05903_));
 sg13g2_a21o_1 _14369_ (.A2(_05909_),
    .A1(_05894_),
    .B1(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _14370_ (.A(\am_sdr0.cic2.comb3_in_del[15] ),
    .X(_05913_));
 sg13g2_xor2_1 _14371_ (.B(_05913_),
    .A(_05681_),
    .X(_05914_));
 sg13g2_xnor2_1 _14372_ (.Y(_05915_),
    .A(_05912_),
    .B(_05914_));
 sg13g2_nand2_1 _14373_ (.Y(_05916_),
    .A(_05327_),
    .B(_05915_));
 sg13g2_o21ai_1 _14374_ (.B1(_05916_),
    .Y(_05917_),
    .A1(net224),
    .A2(\am_sdr0.cic2.comb3[15] ));
 sg13g2_nor2_1 _14375_ (.A(net89),
    .B(_05917_),
    .Y(_00704_));
 sg13g2_inv_1 _14376_ (.Y(_05918_),
    .A(_05913_));
 sg13g2_a21oi_1 _14377_ (.A1(_05894_),
    .A2(_05909_),
    .Y(_05919_),
    .B1(_05911_));
 sg13g2_inv_1 _14378_ (.Y(_05920_),
    .A(_05681_));
 sg13g2_a21oi_1 _14379_ (.A1(_05913_),
    .A2(_05912_),
    .Y(_05921_),
    .B1(_05920_));
 sg13g2_a21oi_2 _14380_ (.B1(_05921_),
    .Y(_05922_),
    .A2(_05919_),
    .A1(_05918_));
 sg13g2_buf_1 _14381_ (.A(\am_sdr0.cic2.comb3_in_del[16] ),
    .X(_05923_));
 sg13g2_xor2_1 _14382_ (.B(_05923_),
    .A(_05683_),
    .X(_05924_));
 sg13g2_xnor2_1 _14383_ (.Y(_05925_),
    .A(_05922_),
    .B(_05924_));
 sg13g2_nor2_1 _14384_ (.A(_05356_),
    .B(_05925_),
    .Y(_05926_));
 sg13g2_a21oi_1 _14385_ (.A1(_05370_),
    .A2(\am_sdr0.cic2.comb3[16] ),
    .Y(_05927_),
    .B1(_05926_));
 sg13g2_nor2_1 _14386_ (.A(_05491_),
    .B(_05927_),
    .Y(_00705_));
 sg13g2_nor2_1 _14387_ (.A(_05923_),
    .B(_05922_),
    .Y(_05928_));
 sg13g2_inv_1 _14388_ (.Y(_05929_),
    .A(_05683_));
 sg13g2_a21oi_1 _14389_ (.A1(_05923_),
    .A2(_05922_),
    .Y(_05930_),
    .B1(_05929_));
 sg13g2_or2_1 _14390_ (.X(_05931_),
    .B(_05930_),
    .A(_05928_));
 sg13g2_nor2b_1 _14391_ (.A(\am_sdr0.cic2.comb3_in_del[17] ),
    .B_N(_05714_),
    .Y(_05932_));
 sg13g2_nand2b_1 _14392_ (.Y(_05933_),
    .B(\am_sdr0.cic2.comb3_in_del[17] ),
    .A_N(_05714_));
 sg13g2_nor2b_1 _14393_ (.A(_05932_),
    .B_N(_05933_),
    .Y(_05934_));
 sg13g2_xnor2_1 _14394_ (.Y(_05935_),
    .A(_05931_),
    .B(_05934_));
 sg13g2_o21ai_1 _14395_ (.B1(net218),
    .Y(_05936_),
    .A1(net224),
    .A2(\am_sdr0.cic2.comb3[17] ));
 sg13g2_a21oi_1 _14396_ (.A1(net225),
    .A2(_05935_),
    .Y(_00706_),
    .B1(_05936_));
 sg13g2_nand2b_1 _14397_ (.Y(_05937_),
    .B(_05923_),
    .A_N(_05932_));
 sg13g2_or2_1 _14398_ (.X(_05938_),
    .B(_05932_),
    .A(_05683_));
 sg13g2_a221oi_1 _14399_ (.B2(_05938_),
    .C1(_05921_),
    .B1(_05937_),
    .A1(_05918_),
    .Y(_05939_),
    .A2(_05919_));
 sg13g2_nand2_1 _14400_ (.Y(_05940_),
    .A(_05929_),
    .B(_05923_));
 sg13g2_o21ai_1 _14401_ (.B1(_05933_),
    .Y(_05941_),
    .A1(_05940_),
    .A2(_05932_));
 sg13g2_or2_1 _14402_ (.X(_05942_),
    .B(_05941_),
    .A(_05939_));
 sg13g2_buf_1 _14403_ (.A(_05942_),
    .X(_05943_));
 sg13g2_buf_1 _14404_ (.A(\am_sdr0.cic2.comb3_in_del[18] ),
    .X(_05944_));
 sg13g2_xor2_1 _14405_ (.B(_05944_),
    .A(_05716_),
    .X(_05945_));
 sg13g2_xnor2_1 _14406_ (.Y(_05946_),
    .A(_05943_),
    .B(_05945_));
 sg13g2_o21ai_1 _14407_ (.B1(net218),
    .Y(_05947_),
    .A1(net224),
    .A2(\am_sdr0.cic2.comb3[18] ));
 sg13g2_a21oi_1 _14408_ (.A1(net225),
    .A2(_05946_),
    .Y(_00707_),
    .B1(_05947_));
 sg13g2_xnor2_1 _14409_ (.Y(_05948_),
    .A(\am_sdr0.cic2.comb2[19] ),
    .B(\am_sdr0.cic2.comb3_in_del[19] ));
 sg13g2_and3_1 _14410_ (.X(_05949_),
    .A(_05944_),
    .B(_05943_),
    .C(_05948_));
 sg13g2_inv_1 _14411_ (.Y(_05950_),
    .A(_05716_));
 sg13g2_a21oi_1 _14412_ (.A1(_05950_),
    .A2(_05944_),
    .Y(_05951_),
    .B1(_05948_));
 sg13g2_nor2b_1 _14413_ (.A(_05943_),
    .B_N(_05951_),
    .Y(_05952_));
 sg13g2_o21ai_1 _14414_ (.B1(_05392_),
    .Y(_05953_),
    .A1(_05949_),
    .A2(_05952_));
 sg13g2_and2_1 _14415_ (.A(_05950_),
    .B(_05948_),
    .X(_05954_));
 sg13g2_o21ai_1 _14416_ (.B1(_05954_),
    .Y(_05955_),
    .A1(_05944_),
    .A2(_05943_));
 sg13g2_nor3_1 _14417_ (.A(_05950_),
    .B(_05944_),
    .C(_05948_),
    .Y(_05956_));
 sg13g2_nor2_1 _14418_ (.A(_05355_),
    .B(_05956_),
    .Y(_05957_));
 sg13g2_nor2_1 _14419_ (.A(net284),
    .B(\am_sdr0.cic2.comb3[19] ),
    .Y(_05958_));
 sg13g2_a21o_1 _14420_ (.A2(_05957_),
    .A1(_05955_),
    .B1(_05958_),
    .X(_05959_));
 sg13g2_a21oi_1 _14421_ (.A1(_05953_),
    .A2(_05959_),
    .Y(_00708_),
    .B1(_05882_));
 sg13g2_buf_1 _14422_ (.A(net284),
    .X(_05960_));
 sg13g2_nand2_1 _14423_ (.Y(_05961_),
    .A(\am_sdr0.cic2.comb2[0] ),
    .B(net215));
 sg13g2_nand2_1 _14424_ (.Y(_05962_),
    .A(\am_sdr0.cic2.comb3_in_del[0] ),
    .B(net153));
 sg13g2_a21oi_1 _14425_ (.A1(_05961_),
    .A2(_05962_),
    .Y(_00709_),
    .B1(net81));
 sg13g2_nand2_1 _14426_ (.Y(_05963_),
    .A(_05551_),
    .B(net215));
 sg13g2_nand2_1 _14427_ (.Y(_05964_),
    .A(\am_sdr0.cic2.comb3_in_del[10] ),
    .B(net153));
 sg13g2_a21oi_1 _14428_ (.A1(_05963_),
    .A2(_05964_),
    .Y(_00710_),
    .B1(net81));
 sg13g2_nand2_1 _14429_ (.Y(_05965_),
    .A(_05610_),
    .B(net215));
 sg13g2_nand2_1 _14430_ (.Y(_05966_),
    .A(\am_sdr0.cic2.comb3_in_del[11] ),
    .B(net153));
 sg13g2_a21oi_1 _14431_ (.A1(_05965_),
    .A2(_05966_),
    .Y(_00711_),
    .B1(net81));
 sg13g2_nand2_1 _14432_ (.Y(_05967_),
    .A(_05637_),
    .B(net215));
 sg13g2_nand2_1 _14433_ (.Y(_05968_),
    .A(_05878_),
    .B(net153));
 sg13g2_a21oi_1 _14434_ (.A1(_05967_),
    .A2(_05968_),
    .Y(_00712_),
    .B1(net81));
 sg13g2_nand2_1 _14435_ (.Y(_05969_),
    .A(_05646_),
    .B(_05960_));
 sg13g2_nand2_1 _14436_ (.Y(_05970_),
    .A(_05895_),
    .B(net153));
 sg13g2_a21oi_1 _14437_ (.A1(_05969_),
    .A2(_05970_),
    .Y(_00713_),
    .B1(net81));
 sg13g2_nand2_1 _14438_ (.Y(_05971_),
    .A(\am_sdr0.cic2.comb2[14] ),
    .B(net215));
 sg13g2_nand2_1 _14439_ (.Y(_05972_),
    .A(\am_sdr0.cic2.comb3_in_del[14] ),
    .B(net153));
 sg13g2_a21oi_1 _14440_ (.A1(_05971_),
    .A2(_05972_),
    .Y(_00714_),
    .B1(net81));
 sg13g2_nand2_1 _14441_ (.Y(_05973_),
    .A(_05681_),
    .B(net215));
 sg13g2_nand2_1 _14442_ (.Y(_05974_),
    .A(_05913_),
    .B(_05830_));
 sg13g2_a21oi_1 _14443_ (.A1(_05973_),
    .A2(_05974_),
    .Y(_00715_),
    .B1(_05882_));
 sg13g2_nand2_1 _14444_ (.Y(_05975_),
    .A(_05683_),
    .B(net215));
 sg13g2_nand2_1 _14445_ (.Y(_05976_),
    .A(_05923_),
    .B(_05830_));
 sg13g2_buf_1 _14446_ (.A(_05813_),
    .X(_05977_));
 sg13g2_a21oi_1 _14447_ (.A1(_05975_),
    .A2(_05976_),
    .Y(_00716_),
    .B1(net80));
 sg13g2_nand2_1 _14448_ (.Y(_05978_),
    .A(_05714_),
    .B(_05960_));
 sg13g2_buf_1 _14449_ (.A(_05355_),
    .X(_05979_));
 sg13g2_nand2_1 _14450_ (.Y(_05980_),
    .A(\am_sdr0.cic2.comb3_in_del[17] ),
    .B(_05979_));
 sg13g2_a21oi_1 _14451_ (.A1(_05978_),
    .A2(_05980_),
    .Y(_00717_),
    .B1(net80));
 sg13g2_nand2_1 _14452_ (.Y(_05981_),
    .A(_05716_),
    .B(net215));
 sg13g2_nand2_1 _14453_ (.Y(_05982_),
    .A(_05944_),
    .B(_05979_));
 sg13g2_a21oi_1 _14454_ (.A1(_05981_),
    .A2(_05982_),
    .Y(_00718_),
    .B1(_05977_));
 sg13g2_buf_1 _14455_ (.A(net284),
    .X(_05983_));
 sg13g2_nand2_1 _14456_ (.Y(_05984_),
    .A(\am_sdr0.cic2.comb2[19] ),
    .B(_05983_));
 sg13g2_nand2_1 _14457_ (.Y(_05985_),
    .A(\am_sdr0.cic2.comb3_in_del[19] ),
    .B(net152));
 sg13g2_a21oi_1 _14458_ (.A1(_05984_),
    .A2(_05985_),
    .Y(_00719_),
    .B1(_05977_));
 sg13g2_nand2_1 _14459_ (.Y(_05986_),
    .A(\am_sdr0.cic2.comb2[1] ),
    .B(net214));
 sg13g2_nand2_1 _14460_ (.Y(_05987_),
    .A(\am_sdr0.cic2.comb3_in_del[1] ),
    .B(net152));
 sg13g2_a21oi_1 _14461_ (.A1(_05986_),
    .A2(_05987_),
    .Y(_00720_),
    .B1(net80));
 sg13g2_nand2_1 _14462_ (.Y(_05988_),
    .A(_05741_),
    .B(net214));
 sg13g2_nand2_1 _14463_ (.Y(_05989_),
    .A(\am_sdr0.cic2.comb3_in_del[2] ),
    .B(net152));
 sg13g2_a21oi_1 _14464_ (.A1(_05988_),
    .A2(_05989_),
    .Y(_00721_),
    .B1(net80));
 sg13g2_nand2_1 _14465_ (.Y(_05990_),
    .A(_05747_),
    .B(net214));
 sg13g2_nand2_1 _14466_ (.Y(_05991_),
    .A(\am_sdr0.cic2.comb3_in_del[3] ),
    .B(net152));
 sg13g2_a21oi_1 _14467_ (.A1(_05990_),
    .A2(_05991_),
    .Y(_00722_),
    .B1(net80));
 sg13g2_nand2_1 _14468_ (.Y(_05992_),
    .A(_05753_),
    .B(net214));
 sg13g2_nand2_1 _14469_ (.Y(_05993_),
    .A(\am_sdr0.cic2.comb3_in_del[4] ),
    .B(net152));
 sg13g2_a21oi_1 _14470_ (.A1(_05992_),
    .A2(_05993_),
    .Y(_00723_),
    .B1(net80));
 sg13g2_nand2_1 _14471_ (.Y(_05994_),
    .A(_05759_),
    .B(net214));
 sg13g2_nand2_1 _14472_ (.Y(_05995_),
    .A(\am_sdr0.cic2.comb3_in_del[5] ),
    .B(net152));
 sg13g2_a21oi_1 _14473_ (.A1(_05994_),
    .A2(_05995_),
    .Y(_00724_),
    .B1(net80));
 sg13g2_nand2_1 _14474_ (.Y(_05996_),
    .A(_05769_),
    .B(net214));
 sg13g2_nand2_1 _14475_ (.Y(_05997_),
    .A(\am_sdr0.cic2.comb3_in_del[6] ),
    .B(net152));
 sg13g2_a21oi_1 _14476_ (.A1(_05996_),
    .A2(_05997_),
    .Y(_00725_),
    .B1(net80));
 sg13g2_nand2_1 _14477_ (.Y(_05998_),
    .A(_05772_),
    .B(net214));
 sg13g2_nand2_1 _14478_ (.Y(_05999_),
    .A(\am_sdr0.cic2.comb3_in_del[7] ),
    .B(net152));
 sg13g2_buf_1 _14479_ (.A(_05813_),
    .X(_06000_));
 sg13g2_a21oi_1 _14480_ (.A1(_05998_),
    .A2(_05999_),
    .Y(_00726_),
    .B1(_06000_));
 sg13g2_nand2_1 _14481_ (.Y(_06001_),
    .A(_05777_),
    .B(net214));
 sg13g2_buf_1 _14482_ (.A(_05355_),
    .X(_06002_));
 sg13g2_nand2_1 _14483_ (.Y(_06003_),
    .A(\am_sdr0.cic2.comb3_in_del[8] ),
    .B(net151));
 sg13g2_a21oi_1 _14484_ (.A1(_06001_),
    .A2(_06003_),
    .Y(_00727_),
    .B1(net79));
 sg13g2_nand2_1 _14485_ (.Y(_06004_),
    .A(_05784_),
    .B(_05983_));
 sg13g2_nand2_1 _14486_ (.Y(_06005_),
    .A(\am_sdr0.cic2.comb3_in_del[9] ),
    .B(net151));
 sg13g2_a21oi_1 _14487_ (.A1(_06004_),
    .A2(_06005_),
    .Y(_00728_),
    .B1(_06000_));
 sg13g2_buf_1 _14488_ (.A(_05203_),
    .X(_06006_));
 sg13g2_buf_1 _14489_ (.A(\am_sdr0.cic0.out_tick ),
    .X(_06007_));
 sg13g2_buf_1 _14490_ (.A(net339),
    .X(_06008_));
 sg13g2_xnor2_1 _14491_ (.Y(_06009_),
    .A(_06008_),
    .B(\am_sdr0.cic2.count[0] ));
 sg13g2_nor2_1 _14492_ (.A(net78),
    .B(_06009_),
    .Y(_00729_));
 sg13g2_nand2_1 _14493_ (.Y(_06010_),
    .A(net282),
    .B(\am_sdr0.cic2.count[0] ));
 sg13g2_xor2_1 _14494_ (.B(_06010_),
    .A(\am_sdr0.cic2.count[1] ),
    .X(_06011_));
 sg13g2_nor2_1 _14495_ (.A(net78),
    .B(_06011_),
    .Y(_00730_));
 sg13g2_xnor2_1 _14496_ (.Y(_06012_),
    .A(_02366_),
    .B(_02367_));
 sg13g2_nor2_1 _14497_ (.A(net78),
    .B(_06012_),
    .Y(_00731_));
 sg13g2_xnor2_1 _14498_ (.Y(_06013_),
    .A(_02365_),
    .B(_02368_));
 sg13g2_nor2_1 _14499_ (.A(net78),
    .B(_06013_),
    .Y(_00732_));
 sg13g2_nand2_1 _14500_ (.Y(_06014_),
    .A(_02365_),
    .B(_02368_));
 sg13g2_xor2_1 _14501_ (.B(_06014_),
    .A(\am_sdr0.cic2.count[4] ),
    .X(_06015_));
 sg13g2_nor2_1 _14502_ (.A(net78),
    .B(_06015_),
    .Y(_00733_));
 sg13g2_nand3_1 _14503_ (.B(\am_sdr0.cic2.count[4] ),
    .C(_02368_),
    .A(_02365_),
    .Y(_06016_));
 sg13g2_xor2_1 _14504_ (.B(_06016_),
    .A(\am_sdr0.cic2.count[5] ),
    .X(_06017_));
 sg13g2_nor2_1 _14505_ (.A(net78),
    .B(_06017_),
    .Y(_00734_));
 sg13g2_inv_1 _14506_ (.Y(_06018_),
    .A(\am_sdr0.cic2.count[7] ));
 sg13g2_nor3_1 _14507_ (.A(_06018_),
    .B(_02364_),
    .C(_02370_),
    .Y(_06019_));
 sg13g2_a21oi_1 _14508_ (.A1(_02364_),
    .A2(_02370_),
    .Y(_06020_),
    .B1(_06019_));
 sg13g2_nor2_1 _14509_ (.A(_06006_),
    .B(_06020_),
    .Y(_00735_));
 sg13g2_inv_1 _14510_ (.Y(_06021_),
    .A(_02364_));
 sg13g2_nor2_1 _14511_ (.A(_06021_),
    .B(_02370_),
    .Y(_06022_));
 sg13g2_xnor2_1 _14512_ (.Y(_06023_),
    .A(\am_sdr0.cic2.count[7] ),
    .B(_06022_));
 sg13g2_nor2_1 _14513_ (.A(_06006_),
    .B(_06023_),
    .Y(_00736_));
 sg13g2_nand2_1 _14514_ (.Y(_06024_),
    .A(_06008_),
    .B(\am_sdr0.cic0.x_out[8] ));
 sg13g2_xor2_1 _14515_ (.B(_06024_),
    .A(\am_sdr0.cic2.integ1[0] ),
    .X(_06025_));
 sg13g2_nor2_1 _14516_ (.A(net78),
    .B(_06025_),
    .Y(_00737_));
 sg13g2_buf_1 _14517_ (.A(\am_sdr0.cic2.integ1[10] ),
    .X(_06026_));
 sg13g2_buf_2 _14518_ (.A(\am_sdr0.cic2.integ1[5] ),
    .X(_06027_));
 sg13g2_buf_2 _14519_ (.A(\am_sdr0.cic2.integ1[4] ),
    .X(_06028_));
 sg13g2_or2_1 _14520_ (.X(_06029_),
    .B(\am_sdr0.cic2.integ1[1] ),
    .A(_03998_));
 sg13g2_and2_1 _14521_ (.A(\am_sdr0.cic0.x_out[8] ),
    .B(\am_sdr0.cic2.integ1[0] ),
    .X(_06030_));
 sg13g2_buf_1 _14522_ (.A(_06030_),
    .X(_06031_));
 sg13g2_and2_1 _14523_ (.A(_03998_),
    .B(\am_sdr0.cic2.integ1[1] ),
    .X(_06032_));
 sg13g2_a221oi_1 _14524_ (.B2(_06031_),
    .C1(_06032_),
    .B1(_06029_),
    .A1(_03977_),
    .Y(_06033_),
    .A2(\am_sdr0.cic2.integ1[2] ));
 sg13g2_nor2_1 _14525_ (.A(_03977_),
    .B(\am_sdr0.cic2.integ1[2] ),
    .Y(_06034_));
 sg13g2_inv_1 _14526_ (.Y(_06035_),
    .A(\am_sdr0.cic0.x_out[11] ));
 sg13g2_o21ai_1 _14527_ (.B1(_06035_),
    .Y(_06036_),
    .A1(_06033_),
    .A2(_06034_));
 sg13g2_buf_2 _14528_ (.A(\am_sdr0.cic2.integ1[3] ),
    .X(_06037_));
 sg13g2_nor3_1 _14529_ (.A(_06035_),
    .B(_06033_),
    .C(_06034_),
    .Y(_06038_));
 sg13g2_a221oi_1 _14530_ (.B2(_06037_),
    .C1(_06038_),
    .B1(_06036_),
    .A1(_06028_),
    .Y(_06039_),
    .A2(_03982_));
 sg13g2_nor2_1 _14531_ (.A(_06028_),
    .B(_03982_),
    .Y(_06040_));
 sg13g2_inv_1 _14532_ (.Y(_06041_),
    .A(\am_sdr0.cic0.x_out[13] ));
 sg13g2_o21ai_1 _14533_ (.B1(_06041_),
    .Y(_06042_),
    .A1(_06039_),
    .A2(_06040_));
 sg13g2_nor3_1 _14534_ (.A(_06041_),
    .B(_06039_),
    .C(_06040_),
    .Y(_06043_));
 sg13g2_a21oi_1 _14535_ (.A1(_06027_),
    .A2(_06042_),
    .Y(_06044_),
    .B1(_06043_));
 sg13g2_buf_1 _14536_ (.A(\am_sdr0.cic2.integ1[8] ),
    .X(_06045_));
 sg13g2_buf_2 _14537_ (.A(\am_sdr0.cic2.integ1[9] ),
    .X(_06046_));
 sg13g2_and2_1 _14538_ (.A(net337),
    .B(_06046_),
    .X(_06047_));
 sg13g2_buf_1 _14539_ (.A(_06047_),
    .X(_06048_));
 sg13g2_buf_1 _14540_ (.A(\am_sdr0.cic2.integ1[7] ),
    .X(_06049_));
 sg13g2_buf_1 _14541_ (.A(_06049_),
    .X(_06050_));
 sg13g2_nor2b_1 _14542_ (.A(net347),
    .B_N(net281),
    .Y(_06051_));
 sg13g2_nor2_1 _14543_ (.A(net337),
    .B(_06046_),
    .Y(_06052_));
 sg13g2_inv_1 _14544_ (.Y(_06053_),
    .A(net347));
 sg13g2_nor2_1 _14545_ (.A(net281),
    .B(_06053_),
    .Y(_06054_));
 sg13g2_a22oi_1 _14546_ (.Y(_06055_),
    .B1(_06052_),
    .B2(_06054_),
    .A2(_06051_),
    .A1(_06048_));
 sg13g2_buf_2 _14547_ (.A(\am_sdr0.cic2.integ1[6] ),
    .X(_06056_));
 sg13g2_xnor2_1 _14548_ (.Y(_06057_),
    .A(_06056_),
    .B(_03987_));
 sg13g2_nor3_1 _14549_ (.A(_06044_),
    .B(_06055_),
    .C(_06057_),
    .Y(_06058_));
 sg13g2_a21oi_1 _14550_ (.A1(net281),
    .A2(_06048_),
    .Y(_06059_),
    .B1(net347));
 sg13g2_nand2_1 _14551_ (.Y(_06060_),
    .A(_06056_),
    .B(_03987_));
 sg13g2_nand2b_1 _14552_ (.Y(_06061_),
    .B(_06052_),
    .A_N(net281));
 sg13g2_nand2_1 _14553_ (.Y(_06062_),
    .A(net347),
    .B(_06061_));
 sg13g2_o21ai_1 _14554_ (.B1(_06062_),
    .Y(_06063_),
    .A1(_06059_),
    .A2(_06060_));
 sg13g2_nor2_2 _14555_ (.A(_06058_),
    .B(_06063_),
    .Y(_06064_));
 sg13g2_xnor2_1 _14556_ (.Y(_06065_),
    .A(net241),
    .B(_06064_));
 sg13g2_nand2_1 _14557_ (.Y(_06066_),
    .A(net282),
    .B(_06065_));
 sg13g2_xor2_1 _14558_ (.B(_06066_),
    .A(net338),
    .X(_06067_));
 sg13g2_nor2_1 _14559_ (.A(net78),
    .B(_06067_),
    .Y(_00738_));
 sg13g2_buf_1 _14560_ (.A(_05203_),
    .X(_06068_));
 sg13g2_buf_1 _14561_ (.A(\am_sdr0.cic2.integ1[11] ),
    .X(_06069_));
 sg13g2_buf_1 _14562_ (.A(net339),
    .X(_06070_));
 sg13g2_buf_1 _14563_ (.A(net280),
    .X(_06071_));
 sg13g2_nor2_1 _14564_ (.A(_06056_),
    .B(_03987_),
    .Y(_06072_));
 sg13g2_a21oi_1 _14565_ (.A1(_06044_),
    .A2(_06060_),
    .Y(_06073_),
    .B1(_06072_));
 sg13g2_buf_1 _14566_ (.A(_06073_),
    .X(_06074_));
 sg13g2_nand3_1 _14567_ (.B(_06048_),
    .C(net10),
    .A(net338),
    .Y(_06075_));
 sg13g2_buf_1 _14568_ (.A(_06075_),
    .X(_06076_));
 sg13g2_nand2_1 _14569_ (.Y(_06077_),
    .A(_06053_),
    .B(_06076_));
 sg13g2_or4_1 _14570_ (.A(net337),
    .B(_06046_),
    .C(net338),
    .D(net10),
    .X(_06078_));
 sg13g2_a22oi_1 _14571_ (.Y(_06079_),
    .B1(_06078_),
    .B2(net292),
    .A2(_06077_),
    .A1(net281));
 sg13g2_buf_1 _14572_ (.A(_06079_),
    .X(_06080_));
 sg13g2_xnor2_1 _14573_ (.Y(_06081_),
    .A(net241),
    .B(_06080_));
 sg13g2_nand2_1 _14574_ (.Y(_06082_),
    .A(net213),
    .B(_06081_));
 sg13g2_xor2_1 _14575_ (.B(_06082_),
    .A(net336),
    .X(_06083_));
 sg13g2_nor2_1 _14576_ (.A(net77),
    .B(_06083_),
    .Y(_00739_));
 sg13g2_buf_1 _14577_ (.A(\am_sdr0.cic2.integ1[12] ),
    .X(_06084_));
 sg13g2_or3_1 _14578_ (.A(_06026_),
    .B(net336),
    .C(_06061_),
    .X(_06085_));
 sg13g2_buf_1 _14579_ (.A(_06085_),
    .X(_06086_));
 sg13g2_o21ai_1 _14580_ (.B1(net347),
    .Y(_06087_),
    .A1(net10),
    .A2(_06086_));
 sg13g2_nor2_1 _14581_ (.A(net10),
    .B(_06086_),
    .Y(_06088_));
 sg13g2_nor2_1 _14582_ (.A(_06053_),
    .B(_06088_),
    .Y(_06089_));
 sg13g2_nand2_1 _14583_ (.Y(_06090_),
    .A(_06050_),
    .B(net336));
 sg13g2_nor2_1 _14584_ (.A(_06076_),
    .B(_06090_),
    .Y(_06091_));
 sg13g2_nor2_1 _14585_ (.A(_06089_),
    .B(_06091_),
    .Y(_06092_));
 sg13g2_nand2_1 _14586_ (.Y(_06093_),
    .A(_06053_),
    .B(_06092_));
 sg13g2_nand3_1 _14587_ (.B(_06087_),
    .C(_06093_),
    .A(net280),
    .Y(_06094_));
 sg13g2_xor2_1 _14588_ (.B(_06094_),
    .A(net335),
    .X(_06095_));
 sg13g2_nor2_1 _14589_ (.A(net77),
    .B(_06095_),
    .Y(_00740_));
 sg13g2_buf_1 _14590_ (.A(\am_sdr0.cic2.integ1[13] ),
    .X(_06096_));
 sg13g2_buf_1 _14591_ (.A(_06096_),
    .X(_06097_));
 sg13g2_inv_1 _14592_ (.Y(_06098_),
    .A(net339));
 sg13g2_buf_1 _14593_ (.A(_06098_),
    .X(_06099_));
 sg13g2_nor2_1 _14594_ (.A(net292),
    .B(_06092_),
    .Y(_06100_));
 sg13g2_nand2b_1 _14595_ (.Y(_06101_),
    .B(net292),
    .A_N(net335));
 sg13g2_nor3_1 _14596_ (.A(_06074_),
    .B(_06086_),
    .C(_06101_),
    .Y(_06102_));
 sg13g2_a21oi_1 _14597_ (.A1(net335),
    .A2(_06100_),
    .Y(_06103_),
    .B1(_06102_));
 sg13g2_nor2_1 _14598_ (.A(net212),
    .B(_06103_),
    .Y(_06104_));
 sg13g2_xnor2_1 _14599_ (.Y(_06105_),
    .A(net279),
    .B(_06104_));
 sg13g2_nor2_1 _14600_ (.A(net77),
    .B(_06105_),
    .Y(_00741_));
 sg13g2_buf_1 _14601_ (.A(\am_sdr0.cic2.integ1[14] ),
    .X(_06106_));
 sg13g2_and2_1 _14602_ (.A(net335),
    .B(net279),
    .X(_06107_));
 sg13g2_nor4_1 _14603_ (.A(_06026_),
    .B(net336),
    .C(net279),
    .D(_06101_),
    .Y(_06108_));
 sg13g2_a22oi_1 _14604_ (.Y(_06109_),
    .B1(_06108_),
    .B2(_06064_),
    .A2(_06107_),
    .A1(_06100_));
 sg13g2_nor2_1 _14605_ (.A(net212),
    .B(_06109_),
    .Y(_06110_));
 sg13g2_xnor2_1 _14606_ (.Y(_06111_),
    .A(net334),
    .B(_06110_));
 sg13g2_nor2_1 _14607_ (.A(net77),
    .B(_06111_),
    .Y(_00742_));
 sg13g2_buf_1 _14608_ (.A(\am_sdr0.cic2.integ1[15] ),
    .X(_06112_));
 sg13g2_buf_1 _14609_ (.A(_06112_),
    .X(_06113_));
 sg13g2_and2_1 _14610_ (.A(net334),
    .B(_06107_),
    .X(_06114_));
 sg13g2_buf_1 _14611_ (.A(_06114_),
    .X(_06115_));
 sg13g2_and2_1 _14612_ (.A(_06100_),
    .B(_06115_),
    .X(_06116_));
 sg13g2_nand2_1 _14613_ (.Y(_06117_),
    .A(net241),
    .B(_06080_));
 sg13g2_or3_1 _14614_ (.A(_06084_),
    .B(net279),
    .C(net334),
    .X(_06118_));
 sg13g2_buf_1 _14615_ (.A(_06118_),
    .X(_06119_));
 sg13g2_nor2_1 _14616_ (.A(net336),
    .B(_06119_),
    .Y(_06120_));
 sg13g2_nor2b_1 _14617_ (.A(_06117_),
    .B_N(_06120_),
    .Y(_06121_));
 sg13g2_buf_1 _14618_ (.A(net339),
    .X(_06122_));
 sg13g2_o21ai_1 _14619_ (.B1(net277),
    .Y(_06123_),
    .A1(_06116_),
    .A2(_06121_));
 sg13g2_xor2_1 _14620_ (.B(_06123_),
    .A(net278),
    .X(_06124_));
 sg13g2_nor2_1 _14621_ (.A(net77),
    .B(_06124_),
    .Y(_00743_));
 sg13g2_buf_1 _14622_ (.A(\am_sdr0.cic2.integ1[16] ),
    .X(_06125_));
 sg13g2_nor4_1 _14623_ (.A(net279),
    .B(net334),
    .C(net278),
    .D(_06101_),
    .Y(_06126_));
 sg13g2_nand2_1 _14624_ (.Y(_06127_),
    .A(_06092_),
    .B(_06126_));
 sg13g2_nand3_1 _14625_ (.B(_06100_),
    .C(_06115_),
    .A(net278),
    .Y(_06128_));
 sg13g2_a21oi_1 _14626_ (.A1(_06127_),
    .A2(_06128_),
    .Y(_06129_),
    .B1(_06098_));
 sg13g2_xnor2_1 _14627_ (.Y(_06130_),
    .A(net333),
    .B(_06129_));
 sg13g2_nor2_1 _14628_ (.A(net77),
    .B(_06130_),
    .Y(_00744_));
 sg13g2_buf_1 _14629_ (.A(\am_sdr0.cic2.integ1[17] ),
    .X(_06131_));
 sg13g2_nor4_1 _14630_ (.A(net279),
    .B(net334),
    .C(net278),
    .D(net333),
    .Y(_06132_));
 sg13g2_nand2_1 _14631_ (.Y(_06133_),
    .A(_03992_),
    .B(_06132_));
 sg13g2_and2_1 _14632_ (.A(net278),
    .B(net333),
    .X(_06134_));
 sg13g2_nand4_1 _14633_ (.B(net334),
    .C(_06053_),
    .A(net279),
    .Y(_06135_),
    .D(_06134_));
 sg13g2_a21o_1 _14634_ (.A2(_06093_),
    .A1(_06084_),
    .B1(_06089_),
    .X(_06136_));
 sg13g2_buf_1 _14635_ (.A(_06136_),
    .X(_06137_));
 sg13g2_mux2_1 _14636_ (.A0(_06133_),
    .A1(_06135_),
    .S(_06137_),
    .X(_06138_));
 sg13g2_nor2_1 _14637_ (.A(net212),
    .B(_06138_),
    .Y(_06139_));
 sg13g2_xnor2_1 _14638_ (.Y(_06140_),
    .A(net332),
    .B(_06139_));
 sg13g2_nor2_1 _14639_ (.A(net77),
    .B(_06140_),
    .Y(_00745_));
 sg13g2_buf_1 _14640_ (.A(\am_sdr0.cic2.integ1[18] ),
    .X(_06141_));
 sg13g2_and4_1 _14641_ (.A(net278),
    .B(net333),
    .C(net332),
    .D(_06115_),
    .X(_06142_));
 sg13g2_nand2_1 _14642_ (.Y(_06143_),
    .A(_06069_),
    .B(_06142_));
 sg13g2_o21ai_1 _14643_ (.B1(_06053_),
    .Y(_06144_),
    .A1(_06064_),
    .A2(_06143_));
 sg13g2_nor3_1 _14644_ (.A(net278),
    .B(net333),
    .C(net332),
    .Y(_06145_));
 sg13g2_nand3_1 _14645_ (.B(_06120_),
    .C(_06145_),
    .A(_06064_),
    .Y(_06146_));
 sg13g2_a22oi_1 _14646_ (.Y(_06147_),
    .B1(_06146_),
    .B2(net292),
    .A2(_06144_),
    .A1(net338));
 sg13g2_xnor2_1 _14647_ (.Y(_06148_),
    .A(net241),
    .B(_06147_));
 sg13g2_nand2_1 _14648_ (.Y(_06149_),
    .A(_06071_),
    .B(_06148_));
 sg13g2_xor2_1 _14649_ (.B(_06149_),
    .A(net331),
    .X(_06150_));
 sg13g2_nor2_1 _14650_ (.A(_06068_),
    .B(_06150_),
    .Y(_00746_));
 sg13g2_buf_1 _14651_ (.A(\am_sdr0.cic2.integ1[19] ),
    .X(_06151_));
 sg13g2_nand2b_1 _14652_ (.Y(_06152_),
    .B(_06145_),
    .A_N(net331));
 sg13g2_buf_1 _14653_ (.A(_06152_),
    .X(_06153_));
 sg13g2_inv_1 _14654_ (.Y(_06154_),
    .A(_06153_));
 sg13g2_nor2b_1 _14655_ (.A(net347),
    .B_N(net332),
    .Y(_06155_));
 sg13g2_and3_1 _14656_ (.X(_06156_),
    .A(net278),
    .B(net333),
    .C(_06155_));
 sg13g2_a22oi_1 _14657_ (.Y(_06157_),
    .B1(_06156_),
    .B2(net331),
    .A2(_06154_),
    .A1(net292));
 sg13g2_nor2b_1 _14658_ (.A(_06157_),
    .B_N(_06116_),
    .Y(_06158_));
 sg13g2_a21oi_1 _14659_ (.A1(_06050_),
    .A2(_06115_),
    .Y(_06159_),
    .B1(net292));
 sg13g2_a21oi_1 _14660_ (.A1(net347),
    .A2(_06119_),
    .Y(_06160_),
    .B1(_06069_));
 sg13g2_nor2_1 _14661_ (.A(_06159_),
    .B(_06160_),
    .Y(_06161_));
 sg13g2_nor3_1 _14662_ (.A(_06117_),
    .B(_06153_),
    .C(_06161_),
    .Y(_06162_));
 sg13g2_o21ai_1 _14663_ (.B1(_06070_),
    .Y(_06163_),
    .A1(_06158_),
    .A2(_06162_));
 sg13g2_xor2_1 _14664_ (.B(_06163_),
    .A(net330),
    .X(_06164_));
 sg13g2_nor2_1 _14665_ (.A(_06068_),
    .B(_06164_),
    .Y(_00747_));
 sg13g2_xnor2_1 _14666_ (.Y(_06165_),
    .A(_03998_),
    .B(_06031_));
 sg13g2_nor2_1 _14667_ (.A(net212),
    .B(_06165_),
    .Y(_06166_));
 sg13g2_xnor2_1 _14668_ (.Y(_06167_),
    .A(\am_sdr0.cic2.integ1[1] ),
    .B(_06166_));
 sg13g2_nor2_1 _14669_ (.A(net77),
    .B(_06167_),
    .Y(_00748_));
 sg13g2_buf_1 _14670_ (.A(_05203_),
    .X(_06168_));
 sg13g2_buf_1 _14671_ (.A(\am_sdr0.cic2.integ1[20] ),
    .X(_06169_));
 sg13g2_buf_1 _14672_ (.A(_06169_),
    .X(_06170_));
 sg13g2_o21ai_1 _14673_ (.B1(_06087_),
    .Y(_06171_),
    .A1(_06076_),
    .A2(_06090_));
 sg13g2_or4_1 _14674_ (.A(net330),
    .B(_06171_),
    .C(_06119_),
    .D(_06153_),
    .X(_06172_));
 sg13g2_nand4_1 _14675_ (.B(net330),
    .C(_06171_),
    .A(net331),
    .Y(_06173_),
    .D(_06142_));
 sg13g2_nor2b_1 _14676_ (.A(net292),
    .B_N(_06173_),
    .Y(_06174_));
 sg13g2_a21oi_1 _14677_ (.A1(net241),
    .A2(_06172_),
    .Y(_06175_),
    .B1(_06174_));
 sg13g2_nand2_1 _14678_ (.Y(_06176_),
    .A(_06071_),
    .B(_06175_));
 sg13g2_xor2_1 _14679_ (.B(_06176_),
    .A(net276),
    .X(_06177_));
 sg13g2_nor2_1 _14680_ (.A(net76),
    .B(_06177_),
    .Y(_00749_));
 sg13g2_buf_1 _14681_ (.A(\am_sdr0.cic2.integ1[21] ),
    .X(_06178_));
 sg13g2_buf_1 _14682_ (.A(_06178_),
    .X(_06179_));
 sg13g2_nand2_1 _14683_ (.Y(_06180_),
    .A(_06135_),
    .B(_06133_));
 sg13g2_and3_1 _14684_ (.X(_06181_),
    .A(net331),
    .B(net330),
    .C(net276));
 sg13g2_and4_1 _14685_ (.A(_06137_),
    .B(_06155_),
    .C(_06180_),
    .D(_06181_),
    .X(_06182_));
 sg13g2_nor2_1 _14686_ (.A(net332),
    .B(net331),
    .Y(_06183_));
 sg13g2_nor2_1 _14687_ (.A(net330),
    .B(_06169_),
    .Y(_06184_));
 sg13g2_nand4_1 _14688_ (.B(_06132_),
    .C(_06183_),
    .A(_03992_),
    .Y(_06185_),
    .D(_06184_));
 sg13g2_a21oi_1 _14689_ (.A1(_06137_),
    .A2(_06180_),
    .Y(_06186_),
    .B1(_06185_));
 sg13g2_o21ai_1 _14690_ (.B1(net280),
    .Y(_06187_),
    .A1(_06182_),
    .A2(_06186_));
 sg13g2_xor2_1 _14691_ (.B(_06187_),
    .A(net275),
    .X(_06188_));
 sg13g2_nor2_1 _14692_ (.A(net76),
    .B(_06188_),
    .Y(_00750_));
 sg13g2_buf_2 _14693_ (.A(\am_sdr0.cic2.integ1[22] ),
    .X(_06189_));
 sg13g2_nor2b_1 _14694_ (.A(net347),
    .B_N(net275),
    .Y(_06190_));
 sg13g2_and2_1 _14695_ (.A(_06181_),
    .B(_06190_),
    .X(_06191_));
 sg13g2_nand2_1 _14696_ (.Y(_06192_),
    .A(_03991_),
    .B(_06184_));
 sg13g2_nor3_1 _14697_ (.A(net331),
    .B(net275),
    .C(_06192_),
    .Y(_06193_));
 sg13g2_mux2_1 _14698_ (.A0(_06191_),
    .A1(_06193_),
    .S(_06147_),
    .X(_06194_));
 sg13g2_nand2_1 _14699_ (.Y(_06195_),
    .A(net213),
    .B(_06194_));
 sg13g2_xor2_1 _14700_ (.B(_06195_),
    .A(_06189_),
    .X(_06196_));
 sg13g2_nor2_1 _14701_ (.A(net76),
    .B(_06196_),
    .Y(_00751_));
 sg13g2_buf_2 _14702_ (.A(\am_sdr0.cic2.integ1[23] ),
    .X(_06197_));
 sg13g2_or3_1 _14703_ (.A(net275),
    .B(_06189_),
    .C(_06192_),
    .X(_06198_));
 sg13g2_nand4_1 _14704_ (.B(net276),
    .C(_06189_),
    .A(net330),
    .Y(_06199_),
    .D(_06190_));
 sg13g2_a21oi_1 _14705_ (.A1(_06198_),
    .A2(_06199_),
    .Y(_06200_),
    .B1(_06157_));
 sg13g2_nand3b_1 _14706_ (.B(_06161_),
    .C(_06200_),
    .Y(_06201_),
    .A_N(_06076_));
 sg13g2_nor2_1 _14707_ (.A(_03993_),
    .B(_06201_),
    .Y(_06202_));
 sg13g2_nand2b_1 _14708_ (.Y(_06203_),
    .B(_06080_),
    .A_N(_06161_));
 sg13g2_or2_1 _14709_ (.X(_06204_),
    .B(_06198_),
    .A(_06153_));
 sg13g2_a21oi_1 _14710_ (.A1(_06200_),
    .A2(_06203_),
    .Y(_06205_),
    .B1(_06204_));
 sg13g2_o21ai_1 _14711_ (.B1(net280),
    .Y(_06206_),
    .A1(_06202_),
    .A2(_06205_));
 sg13g2_xor2_1 _14712_ (.B(_06206_),
    .A(_06197_),
    .X(_06207_));
 sg13g2_nor2_1 _14713_ (.A(_06168_),
    .B(_06207_),
    .Y(_00752_));
 sg13g2_buf_2 _14714_ (.A(\am_sdr0.cic2.integ1[24] ),
    .X(_06208_));
 sg13g2_nand4_1 _14715_ (.B(_06189_),
    .C(_06197_),
    .A(net276),
    .Y(_06209_),
    .D(_06190_));
 sg13g2_nor3_1 _14716_ (.A(net275),
    .B(_06189_),
    .C(_06197_),
    .Y(_06210_));
 sg13g2_nand3b_1 _14717_ (.B(net241),
    .C(_06210_),
    .Y(_06211_),
    .A_N(net276));
 sg13g2_nand2b_1 _14718_ (.Y(_06212_),
    .B(_06172_),
    .A_N(_06174_));
 sg13g2_mux2_1 _14719_ (.A0(_06209_),
    .A1(_06211_),
    .S(_06212_),
    .X(_06213_));
 sg13g2_nor2_1 _14720_ (.A(_06099_),
    .B(_06213_),
    .Y(_06214_));
 sg13g2_xnor2_1 _14721_ (.Y(_06215_),
    .A(_06208_),
    .B(_06214_));
 sg13g2_nor2_1 _14722_ (.A(_06168_),
    .B(_06215_),
    .Y(_00753_));
 sg13g2_nor2b_1 _14723_ (.A(_06208_),
    .B_N(_06210_),
    .Y(_06216_));
 sg13g2_nand4_1 _14724_ (.B(_06197_),
    .C(_06208_),
    .A(_06189_),
    .Y(_06217_),
    .D(_06190_));
 sg13g2_nand2_1 _14725_ (.Y(_06218_),
    .A(net241),
    .B(_06216_));
 sg13g2_nand2_1 _14726_ (.Y(_06219_),
    .A(_06217_),
    .B(_06218_));
 sg13g2_a22oi_1 _14727_ (.Y(_06220_),
    .B1(_06219_),
    .B2(_06182_),
    .A2(_06216_),
    .A1(_06186_));
 sg13g2_buf_1 _14728_ (.A(\am_sdr0.cic2.integ1[25] ),
    .X(_06221_));
 sg13g2_o21ai_1 _14729_ (.B1(_06221_),
    .Y(_06222_),
    .A1(net212),
    .A2(_06220_));
 sg13g2_or3_1 _14730_ (.A(net212),
    .B(_06221_),
    .C(_06220_),
    .X(_06223_));
 sg13g2_a21oi_1 _14731_ (.A1(_06222_),
    .A2(_06223_),
    .Y(_00754_),
    .B1(net79));
 sg13g2_a21o_1 _14732_ (.A2(_06031_),
    .A1(_06029_),
    .B1(_06032_),
    .X(_06224_));
 sg13g2_xor2_1 _14733_ (.B(_06224_),
    .A(_03977_),
    .X(_06225_));
 sg13g2_nand2_1 _14734_ (.Y(_06226_),
    .A(net213),
    .B(_06225_));
 sg13g2_xor2_1 _14735_ (.B(_06226_),
    .A(\am_sdr0.cic2.integ1[2] ),
    .X(_06227_));
 sg13g2_nor2_1 _14736_ (.A(net76),
    .B(_06227_),
    .Y(_00755_));
 sg13g2_nand3b_1 _14737_ (.B(net280),
    .C(_06036_),
    .Y(_06228_),
    .A_N(_06038_));
 sg13g2_xor2_1 _14738_ (.B(_06228_),
    .A(_06037_),
    .X(_06229_));
 sg13g2_nor2_1 _14739_ (.A(net76),
    .B(_06229_),
    .Y(_00756_));
 sg13g2_a21oi_1 _14740_ (.A1(_06037_),
    .A2(_06036_),
    .Y(_06230_),
    .B1(_06038_));
 sg13g2_xnor2_1 _14741_ (.Y(_06231_),
    .A(_03982_),
    .B(_06230_));
 sg13g2_nand2_1 _14742_ (.Y(_06232_),
    .A(net213),
    .B(_06231_));
 sg13g2_xor2_1 _14743_ (.B(_06232_),
    .A(_06028_),
    .X(_06233_));
 sg13g2_nor2_1 _14744_ (.A(net76),
    .B(_06233_),
    .Y(_00757_));
 sg13g2_nand3b_1 _14745_ (.B(net280),
    .C(_06042_),
    .Y(_06234_),
    .A_N(_06043_));
 sg13g2_xor2_1 _14746_ (.B(_06234_),
    .A(_06027_),
    .X(_06235_));
 sg13g2_nor2_1 _14747_ (.A(net76),
    .B(_06235_),
    .Y(_00758_));
 sg13g2_xnor2_1 _14748_ (.Y(_06236_),
    .A(_03987_),
    .B(_06044_));
 sg13g2_nand2_1 _14749_ (.Y(_06237_),
    .A(net213),
    .B(_06236_));
 sg13g2_xor2_1 _14750_ (.B(_06237_),
    .A(_06056_),
    .X(_06238_));
 sg13g2_nor2_1 _14751_ (.A(net76),
    .B(_06238_),
    .Y(_00759_));
 sg13g2_buf_1 _14752_ (.A(_05203_),
    .X(_06239_));
 sg13g2_xor2_1 _14753_ (.B(net10),
    .A(net241),
    .X(_06240_));
 sg13g2_nand2_1 _14754_ (.Y(_06241_),
    .A(net213),
    .B(_06240_));
 sg13g2_xor2_1 _14755_ (.B(_06241_),
    .A(net281),
    .X(_06242_));
 sg13g2_nor2_1 _14756_ (.A(net75),
    .B(_06242_),
    .Y(_00760_));
 sg13g2_mux2_1 _14757_ (.A0(_06054_),
    .A1(_06051_),
    .S(net10),
    .X(_06243_));
 sg13g2_nand2_1 _14758_ (.Y(_06244_),
    .A(net213),
    .B(_06243_));
 sg13g2_xor2_1 _14759_ (.B(_06244_),
    .A(net337),
    .X(_06245_));
 sg13g2_nor2_1 _14760_ (.A(net75),
    .B(_06245_),
    .Y(_00761_));
 sg13g2_nand2b_1 _14761_ (.Y(_06246_),
    .B(_06054_),
    .A_N(_06045_));
 sg13g2_nand3_1 _14762_ (.B(_06051_),
    .C(net10),
    .A(_06045_),
    .Y(_06247_));
 sg13g2_o21ai_1 _14763_ (.B1(_06247_),
    .Y(_06248_),
    .A1(net10),
    .A2(_06246_));
 sg13g2_nand2_1 _14764_ (.Y(_06249_),
    .A(net213),
    .B(_06248_));
 sg13g2_xor2_1 _14765_ (.B(_06249_),
    .A(_06046_),
    .X(_06250_));
 sg13g2_nor2_1 _14766_ (.A(net75),
    .B(_06250_),
    .Y(_00762_));
 sg13g2_buf_1 _14767_ (.A(net280),
    .X(_06251_));
 sg13g2_nand2_1 _14768_ (.Y(_06252_),
    .A(net211),
    .B(_06037_));
 sg13g2_xor2_1 _14769_ (.B(_06252_),
    .A(\am_sdr0.cic2.integ2[0] ),
    .X(_06253_));
 sg13g2_nor2_1 _14770_ (.A(net75),
    .B(_06253_),
    .Y(_00763_));
 sg13g2_buf_2 _14771_ (.A(\am_sdr0.cic2.integ2[10] ),
    .X(_06254_));
 sg13g2_buf_1 _14772_ (.A(\am_sdr0.cic2.integ2[9] ),
    .X(_06255_));
 sg13g2_nand2_1 _14773_ (.Y(_06256_),
    .A(net335),
    .B(net329));
 sg13g2_buf_2 _14774_ (.A(\am_sdr0.cic2.integ2[8] ),
    .X(_06257_));
 sg13g2_nor2_1 _14775_ (.A(\am_sdr0.cic2.integ1[11] ),
    .B(_06257_),
    .Y(_06258_));
 sg13g2_nor2_1 _14776_ (.A(\am_sdr0.cic2.integ1[12] ),
    .B(net329),
    .Y(_06259_));
 sg13g2_a21oi_1 _14777_ (.A1(_06256_),
    .A2(_06258_),
    .Y(_06260_),
    .B1(_06259_));
 sg13g2_buf_1 _14778_ (.A(\am_sdr0.cic2.integ2[6] ),
    .X(_06261_));
 sg13g2_nand2_1 _14779_ (.Y(_06262_),
    .A(_06046_),
    .B(_06261_));
 sg13g2_buf_2 _14780_ (.A(\am_sdr0.cic2.integ2[5] ),
    .X(_06263_));
 sg13g2_buf_2 _14781_ (.A(\am_sdr0.cic2.integ2[4] ),
    .X(_06264_));
 sg13g2_or2_1 _14782_ (.X(_06265_),
    .B(_06264_),
    .A(_06049_));
 sg13g2_a21oi_1 _14783_ (.A1(_06263_),
    .A2(_06265_),
    .Y(_06266_),
    .B1(net337));
 sg13g2_a221oi_1 _14784_ (.B2(_06261_),
    .C1(net337),
    .B1(_06046_),
    .A1(net281),
    .Y(_06267_),
    .A2(_06264_));
 sg13g2_buf_2 _14785_ (.A(\am_sdr0.cic2.integ2[2] ),
    .X(_06268_));
 sg13g2_buf_2 _14786_ (.A(\am_sdr0.cic2.integ2[3] ),
    .X(_06269_));
 sg13g2_a22oi_1 _14787_ (.Y(_06270_),
    .B1(_06056_),
    .B2(_06269_),
    .A2(_06268_),
    .A1(_06027_));
 sg13g2_nor2_1 _14788_ (.A(_06028_),
    .B(\am_sdr0.cic2.integ2[1] ),
    .Y(_06271_));
 sg13g2_a22oi_1 _14789_ (.Y(_06272_),
    .B1(_06028_),
    .B2(\am_sdr0.cic2.integ2[1] ),
    .A2(\am_sdr0.cic2.integ2[0] ),
    .A1(_06037_));
 sg13g2_nor2_1 _14790_ (.A(_06027_),
    .B(_06268_),
    .Y(_06273_));
 sg13g2_or3_1 _14791_ (.A(_06271_),
    .B(_06272_),
    .C(_06273_),
    .X(_06274_));
 sg13g2_nor2_1 _14792_ (.A(_06056_),
    .B(_06269_),
    .Y(_06275_));
 sg13g2_a21o_1 _14793_ (.A2(_06274_),
    .A1(_06270_),
    .B1(_06275_),
    .X(_06276_));
 sg13g2_buf_1 _14794_ (.A(_06276_),
    .X(_06277_));
 sg13g2_nand2_1 _14795_ (.Y(_06278_),
    .A(_06049_),
    .B(_06264_));
 sg13g2_o21ai_1 _14796_ (.B1(_06278_),
    .Y(_06279_),
    .A1(_06275_),
    .A2(_06270_));
 sg13g2_nor2_1 _14797_ (.A(_06049_),
    .B(_06264_),
    .Y(_06280_));
 sg13g2_nor3_1 _14798_ (.A(_06273_),
    .B(_06275_),
    .C(_06280_),
    .Y(_06281_));
 sg13g2_nor2_1 _14799_ (.A(_06271_),
    .B(_06272_),
    .Y(_06282_));
 sg13g2_nand2b_1 _14800_ (.Y(_06283_),
    .B(_06262_),
    .A_N(_06263_));
 sg13g2_a221oi_1 _14801_ (.B2(_06282_),
    .C1(_06283_),
    .B1(_06281_),
    .A1(_06265_),
    .Y(_06284_),
    .A2(_06279_));
 sg13g2_a221oi_1 _14802_ (.B2(_06277_),
    .C1(_06284_),
    .B1(_06267_),
    .A1(_06262_),
    .Y(_06285_),
    .A2(_06266_));
 sg13g2_buf_2 _14803_ (.A(_06285_),
    .X(_06286_));
 sg13g2_buf_2 _14804_ (.A(\am_sdr0.cic2.integ2[7] ),
    .X(_06287_));
 sg13g2_inv_1 _14805_ (.Y(_06288_),
    .A(_06287_));
 sg13g2_nor2_1 _14806_ (.A(_06046_),
    .B(_06261_),
    .Y(_06289_));
 sg13g2_nor2_1 _14807_ (.A(_06288_),
    .B(_06289_),
    .Y(_06290_));
 sg13g2_a221oi_1 _14808_ (.B2(_06290_),
    .C1(_06257_),
    .B1(_06286_),
    .A1(net335),
    .Y(_06291_),
    .A2(net329));
 sg13g2_a221oi_1 _14809_ (.B2(_06290_),
    .C1(net336),
    .B1(_06286_),
    .A1(net335),
    .Y(_06292_),
    .A2(net329));
 sg13g2_nor2b_1 _14810_ (.A(_06289_),
    .B_N(net338),
    .Y(_06293_));
 sg13g2_a22oi_1 _14811_ (.Y(_06294_),
    .B1(_06286_),
    .B2(_06293_),
    .A2(_06287_),
    .A1(net338));
 sg13g2_o21ai_1 _14812_ (.B1(_06294_),
    .Y(_06295_),
    .A1(_06291_),
    .A2(_06292_));
 sg13g2_a21oi_1 _14813_ (.A1(_06260_),
    .A2(_06295_),
    .Y(_06296_),
    .B1(net279));
 sg13g2_nand3_1 _14814_ (.B(_06260_),
    .C(_06295_),
    .A(_06097_),
    .Y(_06297_));
 sg13g2_nand3b_1 _14815_ (.B(net280),
    .C(_06297_),
    .Y(_06298_),
    .A_N(_06296_));
 sg13g2_xor2_1 _14816_ (.B(_06298_),
    .A(_06254_),
    .X(_06299_));
 sg13g2_nor2_1 _14817_ (.A(net75),
    .B(_06299_),
    .Y(_00764_));
 sg13g2_buf_2 _14818_ (.A(\am_sdr0.cic2.integ2[11] ),
    .X(_06300_));
 sg13g2_nand2_1 _14819_ (.Y(_06301_),
    .A(_06096_),
    .B(_06254_));
 sg13g2_or2_1 _14820_ (.X(_06302_),
    .B(_06254_),
    .A(_06097_));
 sg13g2_nand3_1 _14821_ (.B(_06295_),
    .C(_06302_),
    .A(_06260_),
    .Y(_06303_));
 sg13g2_nand2_1 _14822_ (.Y(_06304_),
    .A(_06301_),
    .B(_06303_));
 sg13g2_xor2_1 _14823_ (.B(_06304_),
    .A(net334),
    .X(_06305_));
 sg13g2_nand2_1 _14824_ (.Y(_06306_),
    .A(net211),
    .B(_06305_));
 sg13g2_xor2_1 _14825_ (.B(_06306_),
    .A(_06300_),
    .X(_06307_));
 sg13g2_nor2_1 _14826_ (.A(net75),
    .B(_06307_),
    .Y(_00765_));
 sg13g2_buf_1 _14827_ (.A(\am_sdr0.cic2.integ2[12] ),
    .X(_06308_));
 sg13g2_inv_1 _14828_ (.Y(_06309_),
    .A(_06308_));
 sg13g2_nor2_1 _14829_ (.A(net334),
    .B(_06300_),
    .Y(_06310_));
 sg13g2_a22oi_1 _14830_ (.Y(_06311_),
    .B1(net336),
    .B2(_06257_),
    .A2(_06287_),
    .A1(net338));
 sg13g2_o21ai_1 _14831_ (.B1(_06286_),
    .Y(_06312_),
    .A1(_06290_),
    .A2(_06293_));
 sg13g2_a21oi_1 _14832_ (.A1(_06311_),
    .A2(_06312_),
    .Y(_06313_),
    .B1(_06258_));
 sg13g2_nand2_1 _14833_ (.Y(_06314_),
    .A(_06106_),
    .B(_06300_));
 sg13g2_nand3_1 _14834_ (.B(_06301_),
    .C(_06314_),
    .A(_06256_),
    .Y(_06315_));
 sg13g2_nor2_1 _14835_ (.A(_06096_),
    .B(_06254_),
    .Y(_06316_));
 sg13g2_and2_1 _14836_ (.A(_06259_),
    .B(_06301_),
    .X(_06317_));
 sg13g2_o21ai_1 _14837_ (.B1(_06314_),
    .Y(_06318_),
    .A1(_06316_),
    .A2(_06317_));
 sg13g2_o21ai_1 _14838_ (.B1(_06318_),
    .Y(_06319_),
    .A1(_06313_),
    .A2(_06315_));
 sg13g2_buf_1 _14839_ (.A(_06319_),
    .X(_06320_));
 sg13g2_nor2_1 _14840_ (.A(_06310_),
    .B(_06320_),
    .Y(_06321_));
 sg13g2_xor2_1 _14841_ (.B(_06321_),
    .A(_06113_),
    .X(_06322_));
 sg13g2_nand2_1 _14842_ (.Y(_06323_),
    .A(net282),
    .B(_06322_));
 sg13g2_xnor2_1 _14843_ (.Y(_06324_),
    .A(_06309_),
    .B(_06323_));
 sg13g2_nor2_1 _14844_ (.A(net75),
    .B(_06324_),
    .Y(_00766_));
 sg13g2_buf_1 _14845_ (.A(\am_sdr0.cic2.integ2[13] ),
    .X(_06325_));
 sg13g2_buf_1 _14846_ (.A(_06325_),
    .X(_06326_));
 sg13g2_nor2_1 _14847_ (.A(_06112_),
    .B(_06308_),
    .Y(_06327_));
 sg13g2_and2_1 _14848_ (.A(_06112_),
    .B(_06308_),
    .X(_06328_));
 sg13g2_buf_1 _14849_ (.A(_06328_),
    .X(_06329_));
 sg13g2_nor2_1 _14850_ (.A(_06321_),
    .B(_06329_),
    .Y(_06330_));
 sg13g2_or2_1 _14851_ (.X(_06331_),
    .B(_06330_),
    .A(_06327_));
 sg13g2_xnor2_1 _14852_ (.Y(_06332_),
    .A(net333),
    .B(_06331_));
 sg13g2_nand2_1 _14853_ (.Y(_06333_),
    .A(_06251_),
    .B(_06332_));
 sg13g2_xor2_1 _14854_ (.B(_06333_),
    .A(net274),
    .X(_06334_));
 sg13g2_nor2_1 _14855_ (.A(net75),
    .B(_06334_),
    .Y(_00767_));
 sg13g2_buf_2 _14856_ (.A(\am_sdr0.cic2.integ2[14] ),
    .X(_06335_));
 sg13g2_nor2_1 _14857_ (.A(net333),
    .B(net274),
    .Y(_06336_));
 sg13g2_nand2_1 _14858_ (.Y(_06337_),
    .A(_06125_),
    .B(net274));
 sg13g2_o21ai_1 _14859_ (.B1(_06337_),
    .Y(_06338_),
    .A1(_06331_),
    .A2(_06336_));
 sg13g2_xor2_1 _14860_ (.B(_06338_),
    .A(net332),
    .X(_06339_));
 sg13g2_nand2_1 _14861_ (.Y(_06340_),
    .A(net211),
    .B(_06339_));
 sg13g2_xor2_1 _14862_ (.B(_06340_),
    .A(_06335_),
    .X(_06341_));
 sg13g2_nor2_1 _14863_ (.A(_06239_),
    .B(_06341_),
    .Y(_00768_));
 sg13g2_buf_2 _14864_ (.A(\am_sdr0.cic2.integ2[15] ),
    .X(_06342_));
 sg13g2_nor2_1 _14865_ (.A(_06325_),
    .B(net332),
    .Y(_06343_));
 sg13g2_nor2b_1 _14866_ (.A(_06329_),
    .B_N(_06343_),
    .Y(_06344_));
 sg13g2_o21ai_1 _14867_ (.B1(_06344_),
    .Y(_06345_),
    .A1(_06310_),
    .A2(_06320_));
 sg13g2_buf_1 _14868_ (.A(_06345_),
    .X(_06346_));
 sg13g2_nor3_1 _14869_ (.A(net274),
    .B(_06335_),
    .C(_06329_),
    .Y(_06347_));
 sg13g2_or4_1 _14870_ (.A(_06106_),
    .B(_06300_),
    .C(net274),
    .D(_06329_),
    .X(_06348_));
 sg13g2_a21oi_1 _14871_ (.A1(net332),
    .A2(_06348_),
    .Y(_06349_),
    .B1(_06335_));
 sg13g2_a21oi_2 _14872_ (.B1(_06349_),
    .Y(_06350_),
    .A2(_06347_),
    .A1(_06320_));
 sg13g2_a21oi_1 _14873_ (.A1(_06301_),
    .A2(_06314_),
    .Y(_06351_),
    .B1(_06310_));
 sg13g2_a21o_1 _14874_ (.A2(_06325_),
    .A1(_06308_),
    .B1(_06351_),
    .X(_06352_));
 sg13g2_a21o_1 _14875_ (.A2(_06335_),
    .A1(_06131_),
    .B1(_06125_),
    .X(_06353_));
 sg13g2_a221oi_1 _14876_ (.B2(_06113_),
    .C1(_06353_),
    .B1(_06352_),
    .A1(_06308_),
    .Y(_06354_),
    .A2(_06351_));
 sg13g2_nand2b_1 _14877_ (.Y(_06355_),
    .B(_06327_),
    .A_N(_06335_));
 sg13g2_and2_1 _14878_ (.A(_06353_),
    .B(_06355_),
    .X(_06356_));
 sg13g2_o21ai_1 _14879_ (.B1(_06354_),
    .Y(_06357_),
    .A1(_06310_),
    .A2(_06327_));
 sg13g2_o21ai_1 _14880_ (.B1(_06357_),
    .Y(_06358_),
    .A1(net274),
    .A2(_06356_));
 sg13g2_a221oi_1 _14881_ (.B2(_06303_),
    .C1(_06358_),
    .B1(_06354_),
    .A1(_06327_),
    .Y(_06359_),
    .A2(_06343_));
 sg13g2_buf_1 _14882_ (.A(_06359_),
    .X(_06360_));
 sg13g2_nand3_1 _14883_ (.B(_06350_),
    .C(_06360_),
    .A(_06346_),
    .Y(_06361_));
 sg13g2_xor2_1 _14884_ (.B(_06361_),
    .A(_06141_),
    .X(_06362_));
 sg13g2_nand2b_1 _14885_ (.Y(_06363_),
    .B(_06122_),
    .A_N(_06362_));
 sg13g2_xor2_1 _14886_ (.B(_06363_),
    .A(_06342_),
    .X(_06364_));
 sg13g2_nor2_1 _14887_ (.A(_06239_),
    .B(_06364_),
    .Y(_00769_));
 sg13g2_buf_1 _14888_ (.A(_02778_),
    .X(_06365_));
 sg13g2_buf_1 _14889_ (.A(_06365_),
    .X(_06366_));
 sg13g2_buf_2 _14890_ (.A(\am_sdr0.cic2.integ2[16] ),
    .X(_06367_));
 sg13g2_or2_1 _14891_ (.X(_06368_),
    .B(_06342_),
    .A(_06141_));
 sg13g2_nand4_1 _14892_ (.B(_06350_),
    .C(_06360_),
    .A(_06346_),
    .Y(_06369_),
    .D(_06368_));
 sg13g2_nand2_1 _14893_ (.Y(_06370_),
    .A(\am_sdr0.cic2.integ1[18] ),
    .B(_06342_));
 sg13g2_nand2_1 _14894_ (.Y(_06371_),
    .A(_06369_),
    .B(_06370_));
 sg13g2_xnor2_1 _14895_ (.Y(_06372_),
    .A(net330),
    .B(_06371_));
 sg13g2_nor2_1 _14896_ (.A(net212),
    .B(_06372_),
    .Y(_06373_));
 sg13g2_xnor2_1 _14897_ (.Y(_06374_),
    .A(_06367_),
    .B(_06373_));
 sg13g2_nor2_1 _14898_ (.A(net74),
    .B(_06374_),
    .Y(_00770_));
 sg13g2_buf_1 _14899_ (.A(\am_sdr0.cic2.integ2[17] ),
    .X(_06375_));
 sg13g2_inv_1 _14900_ (.Y(_06376_),
    .A(net328));
 sg13g2_or2_1 _14901_ (.X(_06377_),
    .B(_06367_),
    .A(net330));
 sg13g2_buf_1 _14902_ (.A(_06377_),
    .X(_06378_));
 sg13g2_and2_1 _14903_ (.A(_06342_),
    .B(_06378_),
    .X(_06379_));
 sg13g2_nand4_1 _14904_ (.B(_06350_),
    .C(_06360_),
    .A(_06346_),
    .Y(_06380_),
    .D(_06379_));
 sg13g2_and2_1 _14905_ (.A(net331),
    .B(_06378_),
    .X(_06381_));
 sg13g2_nand4_1 _14906_ (.B(_06350_),
    .C(_06360_),
    .A(_06346_),
    .Y(_06382_),
    .D(_06381_));
 sg13g2_nand2_1 _14907_ (.Y(_06383_),
    .A(_06151_),
    .B(_06367_));
 sg13g2_nand2b_1 _14908_ (.Y(_06384_),
    .B(_06378_),
    .A_N(_06370_));
 sg13g2_and2_1 _14909_ (.A(_06383_),
    .B(_06384_),
    .X(_06385_));
 sg13g2_nand3_1 _14910_ (.B(_06382_),
    .C(_06385_),
    .A(_06380_),
    .Y(_06386_));
 sg13g2_xor2_1 _14911_ (.B(_06386_),
    .A(net276),
    .X(_06387_));
 sg13g2_nand2_1 _14912_ (.Y(_06388_),
    .A(net282),
    .B(_06387_));
 sg13g2_xnor2_1 _14913_ (.Y(_06389_),
    .A(_06376_),
    .B(_06388_));
 sg13g2_nor2_1 _14914_ (.A(net74),
    .B(_06389_),
    .Y(_00771_));
 sg13g2_buf_1 _14915_ (.A(\am_sdr0.cic2.integ2[18] ),
    .X(_06390_));
 sg13g2_nand4_1 _14916_ (.B(_06380_),
    .C(_06382_),
    .A(_06376_),
    .Y(_06391_),
    .D(_06385_));
 sg13g2_and2_1 _14917_ (.A(net328),
    .B(_06378_),
    .X(_06392_));
 sg13g2_nand3_1 _14918_ (.B(_06370_),
    .C(_06383_),
    .A(_06369_),
    .Y(_06393_));
 sg13g2_buf_1 _14919_ (.A(_06393_),
    .X(_06394_));
 sg13g2_a22oi_1 _14920_ (.Y(_06395_),
    .B1(_06392_),
    .B2(_06394_),
    .A2(_06391_),
    .A1(net276));
 sg13g2_xor2_1 _14921_ (.B(_06395_),
    .A(net275),
    .X(_06396_));
 sg13g2_nor2_1 _14922_ (.A(_06099_),
    .B(_06396_),
    .Y(_06397_));
 sg13g2_xnor2_1 _14923_ (.Y(_06398_),
    .A(net327),
    .B(_06397_));
 sg13g2_nor2_1 _14924_ (.A(net74),
    .B(_06398_),
    .Y(_00772_));
 sg13g2_buf_1 _14925_ (.A(\am_sdr0.cic2.integ2[19] ),
    .X(_06399_));
 sg13g2_buf_2 _14926_ (.A(_06399_),
    .X(_06400_));
 sg13g2_nand2_1 _14927_ (.Y(_06401_),
    .A(net275),
    .B(net327));
 sg13g2_nor2_1 _14928_ (.A(_06178_),
    .B(net327),
    .Y(_06402_));
 sg13g2_a21oi_1 _14929_ (.A1(_06395_),
    .A2(_06401_),
    .Y(_06403_),
    .B1(_06402_));
 sg13g2_xor2_1 _14930_ (.B(_06403_),
    .A(_06189_),
    .X(_06404_));
 sg13g2_nand2_1 _14931_ (.Y(_06405_),
    .A(_06251_),
    .B(_06404_));
 sg13g2_xor2_1 _14932_ (.B(_06405_),
    .A(_06400_),
    .X(_06406_));
 sg13g2_nor2_1 _14933_ (.A(_06366_),
    .B(_06406_),
    .Y(_00773_));
 sg13g2_nand2_1 _14934_ (.Y(_06407_),
    .A(_06037_),
    .B(\am_sdr0.cic2.integ2[0] ));
 sg13g2_xnor2_1 _14935_ (.Y(_06408_),
    .A(_06028_),
    .B(_06407_));
 sg13g2_nand2_1 _14936_ (.Y(_06409_),
    .A(net211),
    .B(_06408_));
 sg13g2_xor2_1 _14937_ (.B(_06409_),
    .A(\am_sdr0.cic2.integ2[1] ),
    .X(_06410_));
 sg13g2_nor2_1 _14938_ (.A(net74),
    .B(_06410_),
    .Y(_00774_));
 sg13g2_buf_2 _14939_ (.A(\am_sdr0.cic2.integ2[20] ),
    .X(_06411_));
 sg13g2_and2_1 _14940_ (.A(net297),
    .B(_06411_),
    .X(_06412_));
 sg13g2_nor2_1 _14941_ (.A(net251),
    .B(_06411_),
    .Y(_06413_));
 sg13g2_nand2_1 _14942_ (.Y(_06414_),
    .A(net273),
    .B(_06386_));
 sg13g2_or2_1 _14943_ (.X(_06415_),
    .B(net327),
    .A(_06178_));
 sg13g2_o21ai_1 _14944_ (.B1(_06415_),
    .Y(_06416_),
    .A1(net276),
    .A2(net328));
 sg13g2_nand2_1 _14945_ (.Y(_06417_),
    .A(_06169_),
    .B(net328));
 sg13g2_o21ai_1 _14946_ (.B1(_06401_),
    .Y(_06418_),
    .A1(_06402_),
    .A2(_06417_));
 sg13g2_a21oi_1 _14947_ (.A1(net273),
    .A2(_06418_),
    .Y(_06419_),
    .B1(_06189_));
 sg13g2_o21ai_1 _14948_ (.B1(_06419_),
    .Y(_06420_),
    .A1(_06414_),
    .A2(_06416_));
 sg13g2_o21ai_1 _14949_ (.B1(_06420_),
    .Y(_06421_),
    .A1(net273),
    .A2(_06403_));
 sg13g2_xor2_1 _14950_ (.B(_06421_),
    .A(_06197_),
    .X(_06422_));
 sg13g2_nor2_1 _14951_ (.A(net212),
    .B(_06422_),
    .Y(_06423_));
 sg13g2_mux2_1 _14952_ (.A0(_06412_),
    .A1(_06413_),
    .S(_06423_),
    .X(_00775_));
 sg13g2_buf_2 _14953_ (.A(\am_sdr0.cic2.integ2[21] ),
    .X(_06424_));
 sg13g2_nor2_1 _14954_ (.A(_06197_),
    .B(_06411_),
    .Y(_06425_));
 sg13g2_nor2_1 _14955_ (.A(_06098_),
    .B(_06208_),
    .Y(_06426_));
 sg13g2_nand2b_1 _14956_ (.Y(_06427_),
    .B(_06426_),
    .A_N(_06425_));
 sg13g2_nand2_1 _14957_ (.Y(_06428_),
    .A(_06197_),
    .B(_06411_));
 sg13g2_nand3_1 _14958_ (.B(_06208_),
    .C(_06428_),
    .A(net339),
    .Y(_06429_));
 sg13g2_mux2_1 _14959_ (.A0(_06427_),
    .A1(_06429_),
    .S(_06421_),
    .X(_06430_));
 sg13g2_nand2b_1 _14960_ (.Y(_06431_),
    .B(_06426_),
    .A_N(_06428_));
 sg13g2_nand3_1 _14961_ (.B(_06208_),
    .C(_06425_),
    .A(net339),
    .Y(_06432_));
 sg13g2_and2_1 _14962_ (.A(_06431_),
    .B(_06432_),
    .X(_06433_));
 sg13g2_nand3_1 _14963_ (.B(_06430_),
    .C(_06433_),
    .A(_06424_),
    .Y(_06434_));
 sg13g2_a21o_1 _14964_ (.A2(_06433_),
    .A1(_06430_),
    .B1(_06424_),
    .X(_06435_));
 sg13g2_a21oi_1 _14965_ (.A1(_06434_),
    .A2(_06435_),
    .Y(_00776_),
    .B1(net79));
 sg13g2_nand2b_1 _14966_ (.Y(_06436_),
    .B(net339),
    .A_N(_06221_));
 sg13g2_nand2_1 _14967_ (.Y(_06437_),
    .A(_06007_),
    .B(_06221_));
 sg13g2_or2_1 _14968_ (.X(_06438_),
    .B(\am_sdr0.cic2.integ2[18] ),
    .A(\am_sdr0.cic2.integ2[17] ));
 sg13g2_buf_1 _14969_ (.A(_06438_),
    .X(_06439_));
 sg13g2_or2_1 _14970_ (.X(_06440_),
    .B(net327),
    .A(_06169_));
 sg13g2_a221oi_1 _14971_ (.B2(_06440_),
    .C1(net273),
    .B1(_06439_),
    .A1(_06378_),
    .Y(_06441_),
    .A2(_06394_));
 sg13g2_or2_1 _14972_ (.X(_06442_),
    .B(net275),
    .A(net328));
 sg13g2_or2_1 _14973_ (.X(_06443_),
    .B(_06179_),
    .A(_06170_));
 sg13g2_a221oi_1 _14974_ (.B2(_06443_),
    .C1(net273),
    .B1(_06442_),
    .A1(_06378_),
    .Y(_06444_),
    .A2(_06394_));
 sg13g2_nor2_1 _14975_ (.A(net273),
    .B(_06415_),
    .Y(_06445_));
 sg13g2_nor4_1 _14976_ (.A(_06169_),
    .B(net328),
    .C(net327),
    .D(net273),
    .Y(_06446_));
 sg13g2_nor4_1 _14977_ (.A(_06170_),
    .B(net328),
    .C(_06179_),
    .D(net273),
    .Y(_06447_));
 sg13g2_or3_1 _14978_ (.A(_06445_),
    .B(_06446_),
    .C(_06447_),
    .X(_06448_));
 sg13g2_nor2_1 _14979_ (.A(_06208_),
    .B(_06424_),
    .Y(_06449_));
 sg13g2_or2_1 _14980_ (.X(_06450_),
    .B(_06449_),
    .A(_06425_));
 sg13g2_nor4_1 _14981_ (.A(_06441_),
    .B(_06444_),
    .C(_06448_),
    .D(_06450_),
    .Y(_06451_));
 sg13g2_nor2_1 _14982_ (.A(_06428_),
    .B(_06449_),
    .Y(_06452_));
 sg13g2_a221oi_1 _14983_ (.B2(_06451_),
    .C1(_06452_),
    .B1(_06420_),
    .A1(_06208_),
    .Y(_06453_),
    .A2(_06424_));
 sg13g2_mux2_1 _14984_ (.A0(_06436_),
    .A1(_06437_),
    .S(_06453_),
    .X(_06454_));
 sg13g2_xor2_1 _14985_ (.B(_06454_),
    .A(\am_sdr0.cic2.integ2[22] ),
    .X(_06455_));
 sg13g2_nor2_1 _14986_ (.A(_06366_),
    .B(_06455_),
    .Y(_00777_));
 sg13g2_xor2_1 _14987_ (.B(_06282_),
    .A(_06027_),
    .X(_06456_));
 sg13g2_nand2_1 _14988_ (.Y(_06457_),
    .A(net211),
    .B(_06456_));
 sg13g2_xor2_1 _14989_ (.B(_06457_),
    .A(_06268_),
    .X(_06458_));
 sg13g2_nor2_1 _14990_ (.A(net74),
    .B(_06458_),
    .Y(_00778_));
 sg13g2_nand2_1 _14991_ (.Y(_06459_),
    .A(_06027_),
    .B(_06268_));
 sg13g2_inv_1 _14992_ (.Y(_06460_),
    .A(_06282_));
 sg13g2_a21oi_1 _14993_ (.A1(_06459_),
    .A2(_06460_),
    .Y(_06461_),
    .B1(_06273_));
 sg13g2_xor2_1 _14994_ (.B(_06461_),
    .A(_06056_),
    .X(_06462_));
 sg13g2_nand2_1 _14995_ (.Y(_06463_),
    .A(net211),
    .B(_06462_));
 sg13g2_xor2_1 _14996_ (.B(_06463_),
    .A(_06269_),
    .X(_06464_));
 sg13g2_nor2_1 _14997_ (.A(net74),
    .B(_06464_),
    .Y(_00779_));
 sg13g2_xnor2_1 _14998_ (.Y(_06465_),
    .A(net281),
    .B(_06277_));
 sg13g2_nand2_1 _14999_ (.Y(_06466_),
    .A(net211),
    .B(_06465_));
 sg13g2_xor2_1 _15000_ (.B(_06466_),
    .A(_06264_),
    .X(_06467_));
 sg13g2_nor2_1 _15001_ (.A(net74),
    .B(_06467_),
    .Y(_00780_));
 sg13g2_a21oi_1 _15002_ (.A1(_06277_),
    .A2(_06278_),
    .Y(_06468_),
    .B1(_06280_));
 sg13g2_xor2_1 _15003_ (.B(_06468_),
    .A(net337),
    .X(_06469_));
 sg13g2_nand2_1 _15004_ (.Y(_06470_),
    .A(net211),
    .B(_06469_));
 sg13g2_xor2_1 _15005_ (.B(_06470_),
    .A(_06263_),
    .X(_06471_));
 sg13g2_nor2_1 _15006_ (.A(net74),
    .B(_06471_),
    .Y(_00781_));
 sg13g2_buf_1 _15007_ (.A(_06365_),
    .X(_06472_));
 sg13g2_inv_1 _15008_ (.Y(_06473_),
    .A(_06261_));
 sg13g2_nand3b_1 _15009_ (.B(_06277_),
    .C(_06278_),
    .Y(_06474_),
    .A_N(net337));
 sg13g2_nor2_1 _15010_ (.A(_06263_),
    .B(_06468_),
    .Y(_06475_));
 sg13g2_nor2_1 _15011_ (.A(_06266_),
    .B(_06475_),
    .Y(_06476_));
 sg13g2_nand2_1 _15012_ (.Y(_06477_),
    .A(_06474_),
    .B(_06476_));
 sg13g2_xnor2_1 _15013_ (.Y(_06478_),
    .A(_06046_),
    .B(_06477_));
 sg13g2_nand2_1 _15014_ (.Y(_06479_),
    .A(net282),
    .B(_06478_));
 sg13g2_xnor2_1 _15015_ (.Y(_06480_),
    .A(_06473_),
    .B(_06479_));
 sg13g2_nor2_1 _15016_ (.A(net73),
    .B(_06480_),
    .Y(_00782_));
 sg13g2_buf_1 _15017_ (.A(net339),
    .X(_06481_));
 sg13g2_nand2b_1 _15018_ (.Y(_06482_),
    .B(_06286_),
    .A_N(_06289_));
 sg13g2_xnor2_1 _15019_ (.Y(_06483_),
    .A(net338),
    .B(_06482_));
 sg13g2_nand2_1 _15020_ (.Y(_06484_),
    .A(net272),
    .B(_06483_));
 sg13g2_xor2_1 _15021_ (.B(_06484_),
    .A(_06287_),
    .X(_06485_));
 sg13g2_nor2_1 _15022_ (.A(net73),
    .B(_06485_),
    .Y(_00783_));
 sg13g2_o21ai_1 _15023_ (.B1(_06294_),
    .Y(_06486_),
    .A1(_06288_),
    .A2(_06482_));
 sg13g2_xor2_1 _15024_ (.B(_06486_),
    .A(net336),
    .X(_06487_));
 sg13g2_nand2_1 _15025_ (.Y(_06488_),
    .A(net272),
    .B(_06487_));
 sg13g2_xor2_1 _15026_ (.B(_06488_),
    .A(_06257_),
    .X(_06489_));
 sg13g2_nor2_1 _15027_ (.A(net73),
    .B(_06489_),
    .Y(_00784_));
 sg13g2_xor2_1 _15028_ (.B(_06313_),
    .A(net335),
    .X(_06490_));
 sg13g2_nand2_1 _15029_ (.Y(_06491_),
    .A(net272),
    .B(_06490_));
 sg13g2_xor2_1 _15030_ (.B(_06491_),
    .A(net329),
    .X(_06492_));
 sg13g2_nor2_1 _15031_ (.A(net73),
    .B(_06492_),
    .Y(_00785_));
 sg13g2_nand2_1 _15032_ (.Y(_06493_),
    .A(net272),
    .B(_06269_));
 sg13g2_xor2_1 _15033_ (.B(_06493_),
    .A(\am_sdr0.cic2.integ3[0] ),
    .X(_06494_));
 sg13g2_nor2_1 _15034_ (.A(net73),
    .B(_06494_),
    .Y(_00786_));
 sg13g2_nor2_1 _15035_ (.A(_06254_),
    .B(_02412_),
    .Y(_06495_));
 sg13g2_nand2_1 _15036_ (.Y(_06496_),
    .A(_06300_),
    .B(_02414_));
 sg13g2_nor2_1 _15037_ (.A(_06300_),
    .B(_02414_),
    .Y(_06497_));
 sg13g2_a21oi_1 _15038_ (.A1(_06495_),
    .A2(_06496_),
    .Y(_06498_),
    .B1(_06497_));
 sg13g2_nand2_1 _15039_ (.Y(_06499_),
    .A(_06257_),
    .B(_02406_));
 sg13g2_nor2_1 _15040_ (.A(_06287_),
    .B(_02402_),
    .Y(_06500_));
 sg13g2_nor2_1 _15041_ (.A(_06257_),
    .B(_02406_),
    .Y(_06501_));
 sg13g2_a21oi_1 _15042_ (.A1(_06499_),
    .A2(_06500_),
    .Y(_06502_),
    .B1(_06501_));
 sg13g2_a21o_1 _15043_ (.A2(_02408_),
    .A1(net329),
    .B1(_06502_),
    .X(_06503_));
 sg13g2_o21ai_1 _15044_ (.B1(_06503_),
    .Y(_06504_),
    .A1(net329),
    .A2(_02408_));
 sg13g2_nor2_1 _15045_ (.A(_06263_),
    .B(_02397_),
    .Y(_06505_));
 sg13g2_or2_1 _15046_ (.X(_06506_),
    .B(_02395_),
    .A(_06264_));
 sg13g2_and2_1 _15047_ (.A(_06269_),
    .B(\am_sdr0.cic2.integ3[0] ),
    .X(_06507_));
 sg13g2_buf_1 _15048_ (.A(_06507_),
    .X(_06508_));
 sg13g2_and2_1 _15049_ (.A(_06264_),
    .B(_02395_),
    .X(_06509_));
 sg13g2_a221oi_1 _15050_ (.B2(_06508_),
    .C1(_06509_),
    .B1(_06506_),
    .A1(_06263_),
    .Y(_06510_),
    .A2(_02397_));
 sg13g2_buf_1 _15051_ (.A(_06510_),
    .X(_06511_));
 sg13g2_o21ai_1 _15052_ (.B1(_02399_),
    .Y(_06512_),
    .A1(_06505_),
    .A2(_06511_));
 sg13g2_o21ai_1 _15053_ (.B1(\am_sdr0.cic2.integ3[3] ),
    .Y(_06513_),
    .A1(_06263_),
    .A2(_02397_));
 sg13g2_o21ai_1 _15054_ (.B1(_06473_),
    .Y(_06514_),
    .A1(_06511_),
    .A2(_06513_));
 sg13g2_nand2_1 _15055_ (.Y(_06515_),
    .A(_06287_),
    .B(_02402_));
 sg13g2_nand2_1 _15056_ (.Y(_06516_),
    .A(_06499_),
    .B(_06515_));
 sg13g2_a221oi_1 _15057_ (.B2(_06514_),
    .C1(_06516_),
    .B1(_06512_),
    .A1(net329),
    .Y(_06517_),
    .A2(_02408_));
 sg13g2_and2_1 _15058_ (.A(_06254_),
    .B(_02412_),
    .X(_06518_));
 sg13g2_nor2b_1 _15059_ (.A(_06518_),
    .B_N(_06496_),
    .Y(_06519_));
 sg13g2_o21ai_1 _15060_ (.B1(_06519_),
    .Y(_06520_),
    .A1(_06504_),
    .A2(_06517_));
 sg13g2_nand3_1 _15061_ (.B(_06498_),
    .C(_06520_),
    .A(_02418_),
    .Y(_06521_));
 sg13g2_a21oi_1 _15062_ (.A1(_06498_),
    .A2(_06520_),
    .Y(_06522_),
    .B1(_02418_));
 sg13g2_a21oi_1 _15063_ (.A1(_06309_),
    .A2(_06521_),
    .Y(_06523_),
    .B1(_06522_));
 sg13g2_xor2_1 _15064_ (.B(_06523_),
    .A(net274),
    .X(_06524_));
 sg13g2_nand2_1 _15065_ (.Y(_06525_),
    .A(net272),
    .B(_06524_));
 sg13g2_xor2_1 _15066_ (.B(_06525_),
    .A(_02375_),
    .X(_06526_));
 sg13g2_nor2_1 _15067_ (.A(net73),
    .B(_06526_),
    .Y(_00787_));
 sg13g2_or2_1 _15068_ (.X(_06527_),
    .B(_02375_),
    .A(net274));
 sg13g2_and2_1 _15069_ (.A(_06326_),
    .B(_02375_),
    .X(_06528_));
 sg13g2_a21oi_1 _15070_ (.A1(_06523_),
    .A2(_06527_),
    .Y(_06529_),
    .B1(_06528_));
 sg13g2_xnor2_1 _15071_ (.Y(_06530_),
    .A(_06335_),
    .B(_06529_));
 sg13g2_nand2_1 _15072_ (.Y(_06531_),
    .A(net272),
    .B(_06530_));
 sg13g2_xor2_1 _15073_ (.B(_06531_),
    .A(_02377_),
    .X(_06532_));
 sg13g2_nor2_1 _15074_ (.A(net73),
    .B(_06532_),
    .Y(_00788_));
 sg13g2_or2_1 _15075_ (.X(_06533_),
    .B(_02377_),
    .A(_06335_));
 sg13g2_buf_1 _15076_ (.A(_06533_),
    .X(_06534_));
 sg13g2_nand2_1 _15077_ (.Y(_06535_),
    .A(_02375_),
    .B(_06534_));
 sg13g2_nand2_1 _15078_ (.Y(_06536_),
    .A(_06326_),
    .B(_06534_));
 sg13g2_a221oi_1 _15079_ (.B2(_06536_),
    .C1(_06522_),
    .B1(_06535_),
    .A1(_06309_),
    .Y(_06537_),
    .A2(_06521_));
 sg13g2_buf_1 _15080_ (.A(_06537_),
    .X(_06538_));
 sg13g2_and2_1 _15081_ (.A(_06335_),
    .B(_02377_),
    .X(_06539_));
 sg13g2_a21o_1 _15082_ (.A2(_06534_),
    .A1(_06528_),
    .B1(_06539_),
    .X(_06540_));
 sg13g2_buf_1 _15083_ (.A(_06540_),
    .X(_06541_));
 sg13g2_nor2_1 _15084_ (.A(_06538_),
    .B(_06541_),
    .Y(_06542_));
 sg13g2_xnor2_1 _15085_ (.Y(_06543_),
    .A(_06342_),
    .B(_06542_));
 sg13g2_nand2_1 _15086_ (.Y(_06544_),
    .A(net272),
    .B(_06543_));
 sg13g2_xor2_1 _15087_ (.B(_06544_),
    .A(_02379_),
    .X(_06545_));
 sg13g2_nor2_1 _15088_ (.A(_06472_),
    .B(_06545_),
    .Y(_00789_));
 sg13g2_nor2_1 _15089_ (.A(_06342_),
    .B(_02379_),
    .Y(_06546_));
 sg13g2_nand2_1 _15090_ (.Y(_06547_),
    .A(_06342_),
    .B(_02379_));
 sg13g2_o21ai_1 _15091_ (.B1(_06547_),
    .Y(_06548_),
    .A1(_06542_),
    .A2(_06546_));
 sg13g2_xor2_1 _15092_ (.B(_06548_),
    .A(_06367_),
    .X(_06549_));
 sg13g2_nand2_1 _15093_ (.Y(_06550_),
    .A(net272),
    .B(_06549_));
 sg13g2_xor2_1 _15094_ (.B(_06550_),
    .A(_02381_),
    .X(_06551_));
 sg13g2_nor2_1 _15095_ (.A(net73),
    .B(_06551_),
    .Y(_00790_));
 sg13g2_buf_1 _15096_ (.A(net301),
    .X(_06552_));
 sg13g2_nor2_1 _15097_ (.A(_06367_),
    .B(_02381_),
    .Y(_06553_));
 sg13g2_nor2b_1 _15098_ (.A(_06553_),
    .B_N(_02379_),
    .Y(_06554_));
 sg13g2_o21ai_1 _15099_ (.B1(_06554_),
    .Y(_06555_),
    .A1(_06538_),
    .A2(_06541_));
 sg13g2_nor2b_1 _15100_ (.A(_06553_),
    .B_N(_06342_),
    .Y(_06556_));
 sg13g2_o21ai_1 _15101_ (.B1(_06556_),
    .Y(_06557_),
    .A1(_06538_),
    .A2(_06541_));
 sg13g2_nor2_1 _15102_ (.A(_06547_),
    .B(_06553_),
    .Y(_06558_));
 sg13g2_a21oi_1 _15103_ (.A1(_06367_),
    .A2(_02381_),
    .Y(_06559_),
    .B1(_06558_));
 sg13g2_nand3_1 _15104_ (.B(_06557_),
    .C(_06559_),
    .A(_06555_),
    .Y(_06560_));
 sg13g2_buf_2 _15105_ (.A(_06560_),
    .X(_06561_));
 sg13g2_xnor2_1 _15106_ (.Y(_06562_),
    .A(_06376_),
    .B(_06561_));
 sg13g2_nand2_1 _15107_ (.Y(_06563_),
    .A(_06070_),
    .B(_06562_));
 sg13g2_xnor2_1 _15108_ (.Y(_06564_),
    .A(_02383_),
    .B(_06563_));
 sg13g2_and2_1 _15109_ (.A(net210),
    .B(_06564_),
    .X(_00791_));
 sg13g2_a21oi_1 _15110_ (.A1(_02383_),
    .A2(_06561_),
    .Y(_06565_),
    .B1(_06375_));
 sg13g2_nor2_1 _15111_ (.A(_02383_),
    .B(_06561_),
    .Y(_06566_));
 sg13g2_nor2_1 _15112_ (.A(_06565_),
    .B(_06566_),
    .Y(_06567_));
 sg13g2_xor2_1 _15113_ (.B(_06567_),
    .A(net327),
    .X(_06568_));
 sg13g2_nand2_1 _15114_ (.Y(_06569_),
    .A(_06481_),
    .B(_06568_));
 sg13g2_xor2_1 _15115_ (.B(_06569_),
    .A(_02385_),
    .X(_06570_));
 sg13g2_nor2_1 _15116_ (.A(_06472_),
    .B(_06570_),
    .Y(_00792_));
 sg13g2_buf_1 _15117_ (.A(_06365_),
    .X(_06571_));
 sg13g2_and2_1 _15118_ (.A(net327),
    .B(_02385_),
    .X(_06572_));
 sg13g2_or2_1 _15119_ (.X(_06573_),
    .B(_02385_),
    .A(_06390_));
 sg13g2_o21ai_1 _15120_ (.B1(_06573_),
    .Y(_06574_),
    .A1(_06567_),
    .A2(_06572_));
 sg13g2_xnor2_1 _15121_ (.Y(_06575_),
    .A(_06400_),
    .B(_06574_));
 sg13g2_nand2_1 _15122_ (.Y(_06576_),
    .A(_06481_),
    .B(_06575_));
 sg13g2_xor2_1 _15123_ (.B(_06576_),
    .A(_02387_),
    .X(_06577_));
 sg13g2_nor2_1 _15124_ (.A(_06571_),
    .B(_06577_),
    .Y(_00793_));
 sg13g2_or2_1 _15125_ (.X(_06578_),
    .B(_02385_),
    .A(_02383_));
 sg13g2_or2_1 _15126_ (.X(_06579_),
    .B(_02385_),
    .A(_06375_));
 sg13g2_a221oi_1 _15127_ (.B2(_06579_),
    .C1(_06561_),
    .B1(_06578_),
    .A1(_06399_),
    .Y(_06580_),
    .A2(_02387_));
 sg13g2_or2_1 _15128_ (.X(_06581_),
    .B(_02383_),
    .A(_06390_));
 sg13g2_a221oi_1 _15129_ (.B2(_06581_),
    .C1(_06561_),
    .B1(_06439_),
    .A1(_06399_),
    .Y(_06582_),
    .A2(_02387_));
 sg13g2_and2_1 _15130_ (.A(_06399_),
    .B(_02387_),
    .X(_06583_));
 sg13g2_buf_1 _15131_ (.A(_06583_),
    .X(_06584_));
 sg13g2_nor4_1 _15132_ (.A(net328),
    .B(_02383_),
    .C(_02385_),
    .D(_06584_),
    .Y(_06585_));
 sg13g2_nor3_1 _15133_ (.A(_02383_),
    .B(_06439_),
    .C(_06584_),
    .Y(_06586_));
 sg13g2_nor2_1 _15134_ (.A(_06585_),
    .B(_06586_),
    .Y(_06587_));
 sg13g2_o21ai_1 _15135_ (.B1(_06587_),
    .Y(_06588_),
    .A1(_06573_),
    .A2(_06584_));
 sg13g2_nor2_1 _15136_ (.A(_06399_),
    .B(_02387_),
    .Y(_06589_));
 sg13g2_nor4_2 _15137_ (.A(_06580_),
    .B(_06582_),
    .C(_06588_),
    .Y(_06590_),
    .D(_06589_));
 sg13g2_xor2_1 _15138_ (.B(_06590_),
    .A(_06411_),
    .X(_06591_));
 sg13g2_nand2_1 _15139_ (.Y(_06592_),
    .A(_06122_),
    .B(_06591_));
 sg13g2_xor2_1 _15140_ (.B(_06592_),
    .A(_02389_),
    .X(_06593_));
 sg13g2_nor2_1 _15141_ (.A(net72),
    .B(_06593_),
    .Y(_00794_));
 sg13g2_or2_1 _15142_ (.X(_06594_),
    .B(_02389_),
    .A(_06411_));
 sg13g2_and2_1 _15143_ (.A(_06411_),
    .B(_02389_),
    .X(_06595_));
 sg13g2_a21oi_1 _15144_ (.A1(_06590_),
    .A2(_06594_),
    .Y(_06596_),
    .B1(_06595_));
 sg13g2_xor2_1 _15145_ (.B(_06596_),
    .A(_06424_),
    .X(_06597_));
 sg13g2_nor2_1 _15146_ (.A(_06098_),
    .B(_06597_),
    .Y(_06598_));
 sg13g2_xnor2_1 _15147_ (.Y(_06599_),
    .A(_02391_),
    .B(_06598_));
 sg13g2_nor2_1 _15148_ (.A(_06571_),
    .B(_06599_),
    .Y(_00795_));
 sg13g2_nand2_1 _15149_ (.Y(_06600_),
    .A(_06424_),
    .B(_02391_));
 sg13g2_nor2_1 _15150_ (.A(_06424_),
    .B(_02391_),
    .Y(_06601_));
 sg13g2_a21oi_1 _15151_ (.A1(_06596_),
    .A2(_06600_),
    .Y(_06602_),
    .B1(_06601_));
 sg13g2_xor2_1 _15152_ (.B(_06602_),
    .A(\am_sdr0.cic2.integ2[22] ),
    .X(_06603_));
 sg13g2_nand2_1 _15153_ (.Y(_06604_),
    .A(net303),
    .B(\am_sdr0.cic2.integ3[19] ));
 sg13g2_a21oi_1 _15154_ (.A1(net282),
    .A2(_06603_),
    .Y(_06605_),
    .B1(_06604_));
 sg13g2_nand4_1 _15155_ (.B(net282),
    .C(_02393_),
    .A(net254),
    .Y(_06606_),
    .D(_06603_));
 sg13g2_nand2b_1 _15156_ (.Y(_00796_),
    .B(_06606_),
    .A_N(_06605_));
 sg13g2_xnor2_1 _15157_ (.Y(_06607_),
    .A(_06264_),
    .B(_06508_));
 sg13g2_nor2_1 _15158_ (.A(_06098_),
    .B(_06607_),
    .Y(_06608_));
 sg13g2_xnor2_1 _15159_ (.Y(_06609_),
    .A(_02395_),
    .B(_06608_));
 sg13g2_nor2_1 _15160_ (.A(net72),
    .B(_06609_),
    .Y(_00797_));
 sg13g2_a21o_1 _15161_ (.A2(_06508_),
    .A1(_06506_),
    .B1(_06509_),
    .X(_06610_));
 sg13g2_xor2_1 _15162_ (.B(_06610_),
    .A(_06263_),
    .X(_06611_));
 sg13g2_nand2_1 _15163_ (.Y(_06612_),
    .A(net277),
    .B(_06611_));
 sg13g2_xor2_1 _15164_ (.B(_06612_),
    .A(_02397_),
    .X(_06613_));
 sg13g2_nor2_1 _15165_ (.A(net72),
    .B(_06613_),
    .Y(_00798_));
 sg13g2_nor2_1 _15166_ (.A(_06505_),
    .B(_06511_),
    .Y(_06614_));
 sg13g2_xnor2_1 _15167_ (.Y(_06615_),
    .A(_06473_),
    .B(_06614_));
 sg13g2_nand2_1 _15168_ (.Y(_06616_),
    .A(net282),
    .B(_06615_));
 sg13g2_xnor2_1 _15169_ (.Y(_06617_),
    .A(_02399_),
    .B(_06616_));
 sg13g2_nor2_1 _15170_ (.A(net72),
    .B(_06617_),
    .Y(_00799_));
 sg13g2_nand2_1 _15171_ (.Y(_06618_),
    .A(_06512_),
    .B(_06514_));
 sg13g2_xnor2_1 _15172_ (.Y(_06619_),
    .A(_06287_),
    .B(_06618_));
 sg13g2_nand2_1 _15173_ (.Y(_06620_),
    .A(net277),
    .B(_06619_));
 sg13g2_xor2_1 _15174_ (.B(_06620_),
    .A(_02402_),
    .X(_06621_));
 sg13g2_nor2_1 _15175_ (.A(net72),
    .B(_06621_),
    .Y(_00800_));
 sg13g2_o21ai_1 _15176_ (.B1(_06515_),
    .Y(_06622_),
    .A1(_06618_),
    .A2(_06500_));
 sg13g2_xor2_1 _15177_ (.B(_06622_),
    .A(_06257_),
    .X(_06623_));
 sg13g2_nand2_1 _15178_ (.Y(_06624_),
    .A(net277),
    .B(_06623_));
 sg13g2_xor2_1 _15179_ (.B(_06624_),
    .A(_02406_),
    .X(_06625_));
 sg13g2_nor2_1 _15180_ (.A(net72),
    .B(_06625_),
    .Y(_00801_));
 sg13g2_a21oi_1 _15181_ (.A1(_06512_),
    .A2(_06514_),
    .Y(_06626_),
    .B1(_06516_));
 sg13g2_nand2b_1 _15182_ (.Y(_06627_),
    .B(_06502_),
    .A_N(_06626_));
 sg13g2_xnor2_1 _15183_ (.Y(_06628_),
    .A(_06255_),
    .B(_06627_));
 sg13g2_nand2_1 _15184_ (.Y(_06629_),
    .A(net277),
    .B(_06628_));
 sg13g2_xor2_1 _15185_ (.B(_06629_),
    .A(_02408_),
    .X(_06630_));
 sg13g2_nor2_1 _15186_ (.A(net72),
    .B(_06630_),
    .Y(_00802_));
 sg13g2_nor2_1 _15187_ (.A(_06504_),
    .B(_06517_),
    .Y(_06631_));
 sg13g2_xor2_1 _15188_ (.B(_06631_),
    .A(_06254_),
    .X(_06632_));
 sg13g2_nand2_1 _15189_ (.Y(_06633_),
    .A(net277),
    .B(_06632_));
 sg13g2_xor2_1 _15190_ (.B(_06633_),
    .A(_02412_),
    .X(_06634_));
 sg13g2_nor2_1 _15191_ (.A(net72),
    .B(_06634_),
    .Y(_00803_));
 sg13g2_buf_1 _15192_ (.A(_06365_),
    .X(_06635_));
 sg13g2_nor2_1 _15193_ (.A(_06518_),
    .B(_06631_),
    .Y(_06636_));
 sg13g2_nor2_1 _15194_ (.A(_06495_),
    .B(_06636_),
    .Y(_06637_));
 sg13g2_xor2_1 _15195_ (.B(_06637_),
    .A(_06300_),
    .X(_06638_));
 sg13g2_nand2_1 _15196_ (.Y(_06639_),
    .A(net277),
    .B(_06638_));
 sg13g2_xor2_1 _15197_ (.B(_06639_),
    .A(_02414_),
    .X(_06640_));
 sg13g2_nor2_1 _15198_ (.A(net71),
    .B(_06640_),
    .Y(_00804_));
 sg13g2_and2_1 _15199_ (.A(_06498_),
    .B(_06520_),
    .X(_06641_));
 sg13g2_xnor2_1 _15200_ (.Y(_06642_),
    .A(_06309_),
    .B(_06641_));
 sg13g2_nand2_1 _15201_ (.Y(_06643_),
    .A(net277),
    .B(_06642_));
 sg13g2_xor2_1 _15202_ (.B(_06643_),
    .A(_02418_),
    .X(_06644_));
 sg13g2_nor2_1 _15203_ (.A(net71),
    .B(_06644_),
    .Y(_00805_));
 sg13g2_nand2_1 _15204_ (.Y(_06645_),
    .A(net225),
    .B(\am_sdr0.cic2.comb3[14] ));
 sg13g2_nand2_1 _15205_ (.Y(_06646_),
    .A(\am_sdr0.am0.I_in[2] ),
    .B(net151));
 sg13g2_a21oi_1 _15206_ (.A1(_06645_),
    .A2(_06646_),
    .Y(_00828_),
    .B1(net79));
 sg13g2_nand2_1 _15207_ (.Y(_06647_),
    .A(net225),
    .B(\am_sdr0.cic2.comb3[15] ));
 sg13g2_nand2_1 _15208_ (.Y(_06648_),
    .A(\am_sdr0.am0.I_in[3] ),
    .B(net151));
 sg13g2_a21oi_1 _15209_ (.A1(_06647_),
    .A2(_06648_),
    .Y(_00829_),
    .B1(net79));
 sg13g2_nand2_1 _15210_ (.Y(_06649_),
    .A(net225),
    .B(\am_sdr0.cic2.comb3[16] ));
 sg13g2_nand2_1 _15211_ (.Y(_06650_),
    .A(\am_sdr0.am0.I_in[4] ),
    .B(net151));
 sg13g2_a21oi_1 _15212_ (.A1(_06649_),
    .A2(_06650_),
    .Y(_00830_),
    .B1(net79));
 sg13g2_nand2_1 _15213_ (.Y(_06651_),
    .A(net225),
    .B(\am_sdr0.cic2.comb3[17] ));
 sg13g2_nand2_1 _15214_ (.Y(_06652_),
    .A(\am_sdr0.am0.I_in[5] ),
    .B(net151));
 sg13g2_a21oi_1 _15215_ (.A1(_06651_),
    .A2(_06652_),
    .Y(_00831_),
    .B1(net79));
 sg13g2_nand2_1 _15216_ (.Y(_06653_),
    .A(net223),
    .B(\am_sdr0.cic2.comb3[18] ));
 sg13g2_nand2_1 _15217_ (.Y(_06654_),
    .A(\am_sdr0.am0.I_in[6] ),
    .B(net151));
 sg13g2_a21oi_1 _15218_ (.A1(_06653_),
    .A2(_06654_),
    .Y(_00832_),
    .B1(net79));
 sg13g2_nand2_1 _15219_ (.Y(_06655_),
    .A(net223),
    .B(\am_sdr0.cic2.comb3[19] ));
 sg13g2_nand2_1 _15220_ (.Y(_06656_),
    .A(\am_sdr0.am0.I_in[7] ),
    .B(net151));
 sg13g2_buf_1 _15221_ (.A(_05813_),
    .X(_06657_));
 sg13g2_a21oi_1 _15222_ (.A1(_06655_),
    .A2(_06656_),
    .Y(_00833_),
    .B1(net70));
 sg13g2_nand2_1 _15223_ (.Y(_06658_),
    .A(net223),
    .B(\am_sdr0.cic2.comb3[12] ));
 sg13g2_nand2_1 _15224_ (.Y(_06659_),
    .A(\am_sdr0.am0.I_in[0] ),
    .B(_06002_));
 sg13g2_a21oi_1 _15225_ (.A1(_06658_),
    .A2(_06659_),
    .Y(_00834_),
    .B1(net70));
 sg13g2_nand2_1 _15226_ (.Y(_06660_),
    .A(net223),
    .B(\am_sdr0.cic2.comb3[13] ));
 sg13g2_nand2_1 _15227_ (.Y(_06661_),
    .A(\am_sdr0.am0.I_in[1] ),
    .B(_06002_));
 sg13g2_a21oi_1 _15228_ (.A1(_06660_),
    .A2(_06661_),
    .Y(_00835_),
    .B1(net70));
 sg13g2_buf_1 _15229_ (.A(\am_sdr0.cic3.sample ),
    .X(_06662_));
 sg13g2_buf_1 _15230_ (.A(_06662_),
    .X(_06663_));
 sg13g2_buf_1 _15231_ (.A(net271),
    .X(_06664_));
 sg13g2_xnor2_1 _15232_ (.Y(_06665_),
    .A(_02421_),
    .B(\am_sdr0.cic3.comb1_in_del[0] ));
 sg13g2_buf_2 _15233_ (.A(\am_sdr0.cic3.comb1[0] ),
    .X(_06666_));
 sg13g2_buf_1 _15234_ (.A(_06662_),
    .X(_06667_));
 sg13g2_o21ai_1 _15235_ (.B1(net218),
    .Y(_06668_),
    .A1(_06666_),
    .A2(net270));
 sg13g2_a21oi_1 _15236_ (.A1(net209),
    .A2(_06665_),
    .Y(_00836_),
    .B1(_06668_));
 sg13g2_buf_1 _15237_ (.A(\am_sdr0.cic3.comb1[10] ),
    .X(_06669_));
 sg13g2_inv_1 _15238_ (.Y(_06670_),
    .A(_06662_));
 sg13g2_buf_1 _15239_ (.A(_06670_),
    .X(_06671_));
 sg13g2_buf_1 _15240_ (.A(_06671_),
    .X(_06672_));
 sg13g2_buf_1 _15241_ (.A(net150),
    .X(_06673_));
 sg13g2_nand2_1 _15242_ (.Y(_06674_),
    .A(_06669_),
    .B(net69));
 sg13g2_buf_1 _15243_ (.A(_06662_),
    .X(_06675_));
 sg13g2_buf_1 _15244_ (.A(_06675_),
    .X(_06676_));
 sg13g2_inv_1 _15245_ (.Y(_06677_),
    .A(_02468_));
 sg13g2_buf_1 _15246_ (.A(\am_sdr0.cic3.comb1_in_del[2] ),
    .X(_06678_));
 sg13g2_nor2_1 _15247_ (.A(_02464_),
    .B(_06678_),
    .Y(_06679_));
 sg13g2_nor2b_1 _15248_ (.A(_02421_),
    .B_N(\am_sdr0.cic3.comb1_in_del[0] ),
    .Y(_06680_));
 sg13g2_buf_1 _15249_ (.A(\am_sdr0.cic3.comb1_in_del[1] ),
    .X(_06681_));
 sg13g2_nand2b_1 _15250_ (.Y(_06682_),
    .B(_02463_),
    .A_N(_06681_));
 sg13g2_nor2b_1 _15251_ (.A(_02463_),
    .B_N(_06681_),
    .Y(_06683_));
 sg13g2_a221oi_1 _15252_ (.B2(_06682_),
    .C1(_06683_),
    .B1(_06680_),
    .A1(_02464_),
    .Y(_06684_),
    .A2(_06678_));
 sg13g2_buf_1 _15253_ (.A(_06684_),
    .X(_06685_));
 sg13g2_inv_1 _15254_ (.Y(_06686_),
    .A(\am_sdr0.cic3.comb1_in_del[3] ));
 sg13g2_o21ai_1 _15255_ (.B1(_06686_),
    .Y(_06687_),
    .A1(_06679_),
    .A2(_06685_));
 sg13g2_nor3_1 _15256_ (.A(_06686_),
    .B(_06679_),
    .C(_06685_),
    .Y(_06688_));
 sg13g2_a21o_1 _15257_ (.A2(_06687_),
    .A1(_06677_),
    .B1(_06688_),
    .X(_06689_));
 sg13g2_buf_1 _15258_ (.A(_06689_),
    .X(_06690_));
 sg13g2_nand2b_1 _15259_ (.Y(_06691_),
    .B(_02471_),
    .A_N(\am_sdr0.cic3.comb1_in_del[4] ));
 sg13g2_buf_1 _15260_ (.A(\am_sdr0.cic3.comb1_in_del[5] ),
    .X(_06692_));
 sg13g2_nand2b_1 _15261_ (.Y(_06693_),
    .B(\am_sdr0.cic3.comb1_in_del[4] ),
    .A_N(_02471_));
 sg13g2_buf_1 _15262_ (.A(_06693_),
    .X(_06694_));
 sg13g2_nand2b_1 _15263_ (.Y(_06695_),
    .B(_06694_),
    .A_N(_06692_));
 sg13g2_nand2_1 _15264_ (.Y(_06696_),
    .A(_02473_),
    .B(_06694_));
 sg13g2_buf_1 _15265_ (.A(\am_sdr0.cic3.comb1_in_del[7] ),
    .X(_06697_));
 sg13g2_nand2b_1 _15266_ (.Y(_06698_),
    .B(_06697_),
    .A_N(_02478_));
 sg13g2_buf_1 _15267_ (.A(_06698_),
    .X(_06699_));
 sg13g2_buf_1 _15268_ (.A(\am_sdr0.cic3.comb1_in_del[8] ),
    .X(_06700_));
 sg13g2_inv_1 _15269_ (.Y(_06701_),
    .A(_06700_));
 sg13g2_o21ai_1 _15270_ (.B1(_06701_),
    .Y(_06702_),
    .A1(_02479_),
    .A2(_06699_));
 sg13g2_nand2_1 _15271_ (.Y(_06703_),
    .A(_02479_),
    .B(_06699_));
 sg13g2_buf_1 _15272_ (.A(\am_sdr0.cic3.comb1_in_del[6] ),
    .X(_06704_));
 sg13g2_nor2b_1 _15273_ (.A(_02476_),
    .B_N(_06704_),
    .Y(_06705_));
 sg13g2_a21o_1 _15274_ (.A2(_06703_),
    .A1(_06702_),
    .B1(_06705_),
    .X(_06706_));
 sg13g2_a221oi_1 _15275_ (.B2(_06696_),
    .C1(_06706_),
    .B1(_06695_),
    .A1(_06690_),
    .Y(_06707_),
    .A2(_06691_));
 sg13g2_buf_2 _15276_ (.A(_06707_),
    .X(_06708_));
 sg13g2_nand2b_1 _15277_ (.Y(_06709_),
    .B(_02473_),
    .A_N(_06692_));
 sg13g2_nand2b_1 _15278_ (.Y(_06710_),
    .B(_02478_),
    .A_N(_06697_));
 sg13g2_nand3b_1 _15279_ (.B(_06699_),
    .C(_02476_),
    .Y(_06711_),
    .A_N(_06704_));
 sg13g2_a22oi_1 _15280_ (.Y(_06712_),
    .B1(_06710_),
    .B2(_06711_),
    .A2(_06700_),
    .A1(_02480_));
 sg13g2_a21oi_1 _15281_ (.A1(_02479_),
    .A2(_06701_),
    .Y(_06713_),
    .B1(_06712_));
 sg13g2_o21ai_1 _15282_ (.B1(_06713_),
    .Y(_06714_),
    .A1(_06706_),
    .A2(_06709_));
 sg13g2_buf_2 _15283_ (.A(_06714_),
    .X(_06715_));
 sg13g2_buf_1 _15284_ (.A(\am_sdr0.cic3.comb1_in_del[9] ),
    .X(_06716_));
 sg13g2_inv_1 _15285_ (.Y(_06717_),
    .A(_06716_));
 sg13g2_o21ai_1 _15286_ (.B1(_06717_),
    .Y(_06718_),
    .A1(_06708_),
    .A2(_06715_));
 sg13g2_nor3_1 _15287_ (.A(_06717_),
    .B(_06708_),
    .C(_06715_),
    .Y(_06719_));
 sg13g2_a21oi_1 _15288_ (.A1(_02484_),
    .A2(_06718_),
    .Y(_06720_),
    .B1(_06719_));
 sg13g2_buf_2 _15289_ (.A(\am_sdr0.cic3.comb1_in_del[10] ),
    .X(_06721_));
 sg13g2_nor2_1 _15290_ (.A(_02434_),
    .B(_06721_),
    .Y(_06722_));
 sg13g2_nand2_1 _15291_ (.Y(_06723_),
    .A(_02434_),
    .B(_06721_));
 sg13g2_nand2b_1 _15292_ (.Y(_06724_),
    .B(_06723_),
    .A_N(_06722_));
 sg13g2_xnor2_1 _15293_ (.Y(_06725_),
    .A(_06720_),
    .B(_06724_));
 sg13g2_nand2_1 _15294_ (.Y(_06726_),
    .A(net208),
    .B(_06725_));
 sg13g2_a21oi_1 _15295_ (.A1(_06674_),
    .A2(_06726_),
    .Y(_00837_),
    .B1(net70));
 sg13g2_buf_1 _15296_ (.A(\am_sdr0.cic3.comb1[11] ),
    .X(_06727_));
 sg13g2_buf_1 _15297_ (.A(_06675_),
    .X(_06728_));
 sg13g2_buf_1 _15298_ (.A(_06662_),
    .X(_06729_));
 sg13g2_o21ai_1 _15299_ (.B1(_06723_),
    .Y(_06730_),
    .A1(_06720_),
    .A2(_06722_));
 sg13g2_buf_1 _15300_ (.A(\am_sdr0.cic3.comb1_in_del[11] ),
    .X(_06731_));
 sg13g2_xor2_1 _15301_ (.B(_06731_),
    .A(_02439_),
    .X(_06732_));
 sg13g2_xnor2_1 _15302_ (.Y(_06733_),
    .A(_06730_),
    .B(_06732_));
 sg13g2_nand2_1 _15303_ (.Y(_06734_),
    .A(net269),
    .B(_06733_));
 sg13g2_o21ai_1 _15304_ (.B1(_06734_),
    .Y(_06735_),
    .A1(_06727_),
    .A2(net207));
 sg13g2_nor2_1 _15305_ (.A(net71),
    .B(_06735_),
    .Y(_00838_));
 sg13g2_nor2_1 _15306_ (.A(\am_sdr0.cic3.comb1[12] ),
    .B(net270),
    .Y(_06736_));
 sg13g2_buf_1 _15307_ (.A(_06671_),
    .X(_06737_));
 sg13g2_or2_1 _15308_ (.X(_06738_),
    .B(net326),
    .A(_06721_));
 sg13g2_inv_1 _15309_ (.Y(_06739_),
    .A(net326));
 sg13g2_nand2_1 _15310_ (.Y(_06740_),
    .A(_02433_),
    .B(_06739_));
 sg13g2_a221oi_1 _15311_ (.B2(_06740_),
    .C1(_06719_),
    .B1(_06738_),
    .A1(_02484_),
    .Y(_06741_),
    .A2(_06718_));
 sg13g2_a21oi_1 _15312_ (.A1(_06739_),
    .A2(_06722_),
    .Y(_06742_),
    .B1(_02439_));
 sg13g2_nor2b_1 _15313_ (.A(_06741_),
    .B_N(_06742_),
    .Y(_06743_));
 sg13g2_a21oi_1 _15314_ (.A1(net326),
    .A2(_06730_),
    .Y(_06744_),
    .B1(_06743_));
 sg13g2_buf_1 _15315_ (.A(\am_sdr0.cic3.comb1_in_del[12] ),
    .X(_06745_));
 sg13g2_xor2_1 _15316_ (.B(_06745_),
    .A(_02441_),
    .X(_06746_));
 sg13g2_xnor2_1 _15317_ (.Y(_06747_),
    .A(_06744_),
    .B(_06746_));
 sg13g2_nor2_1 _15318_ (.A(net149),
    .B(_06747_),
    .Y(_06748_));
 sg13g2_nor3_1 _15319_ (.A(_04198_),
    .B(_06736_),
    .C(_06748_),
    .Y(_00839_));
 sg13g2_buf_1 _15320_ (.A(\am_sdr0.cic3.comb1[13] ),
    .X(_06749_));
 sg13g2_nor2b_1 _15321_ (.A(_06745_),
    .B_N(_02441_),
    .Y(_06750_));
 sg13g2_nand2b_1 _15322_ (.Y(_06751_),
    .B(_06745_),
    .A_N(_02441_));
 sg13g2_o21ai_1 _15323_ (.B1(_06751_),
    .Y(_06752_),
    .A1(_06744_),
    .A2(_06750_));
 sg13g2_buf_1 _15324_ (.A(\am_sdr0.cic3.comb1_in_del[13] ),
    .X(_06753_));
 sg13g2_xor2_1 _15325_ (.B(_06753_),
    .A(_02442_),
    .X(_06754_));
 sg13g2_xnor2_1 _15326_ (.Y(_06755_),
    .A(_06752_),
    .B(_06754_));
 sg13g2_nand2_1 _15327_ (.Y(_06756_),
    .A(net269),
    .B(_06755_));
 sg13g2_o21ai_1 _15328_ (.B1(_06756_),
    .Y(_06757_),
    .A1(_06749_),
    .A2(net207));
 sg13g2_nor2_1 _15329_ (.A(net71),
    .B(_06757_),
    .Y(_00840_));
 sg13g2_buf_1 _15330_ (.A(\am_sdr0.cic3.comb1[14] ),
    .X(_06758_));
 sg13g2_nand3_1 _15331_ (.B(_06721_),
    .C(\am_sdr0.cic3.comb1_in_del[11] ),
    .A(_06716_),
    .Y(_06759_));
 sg13g2_nor3_1 _15332_ (.A(_06708_),
    .B(_06715_),
    .C(_06759_),
    .Y(_06760_));
 sg13g2_nand3_1 _15333_ (.B(_06721_),
    .C(net326),
    .A(_02484_),
    .Y(_06761_));
 sg13g2_nor3_1 _15334_ (.A(_06708_),
    .B(_06715_),
    .C(_06761_),
    .Y(_06762_));
 sg13g2_nand3_1 _15335_ (.B(_02434_),
    .C(_06731_),
    .A(_06716_),
    .Y(_06763_));
 sg13g2_nor3_1 _15336_ (.A(_06708_),
    .B(_06715_),
    .C(_06763_),
    .Y(_06764_));
 sg13g2_nand3_1 _15337_ (.B(_02434_),
    .C(net326),
    .A(_02484_),
    .Y(_06765_));
 sg13g2_nor3_1 _15338_ (.A(_06708_),
    .B(_06715_),
    .C(_06765_),
    .Y(_06766_));
 sg13g2_nor4_1 _15339_ (.A(_06760_),
    .B(_06762_),
    .C(_06764_),
    .D(_06766_),
    .Y(_06767_));
 sg13g2_nor2b_1 _15340_ (.A(_02433_),
    .B_N(_06721_),
    .Y(_06768_));
 sg13g2_nor2_1 _15341_ (.A(_02483_),
    .B(_06717_),
    .Y(_06769_));
 sg13g2_and2_1 _15342_ (.A(_06721_),
    .B(net326),
    .X(_06770_));
 sg13g2_nor4_1 _15343_ (.A(_02483_),
    .B(_06717_),
    .C(_02433_),
    .D(_06739_),
    .Y(_06771_));
 sg13g2_a221oi_1 _15344_ (.B2(_06770_),
    .C1(_06771_),
    .B1(_06769_),
    .A1(net326),
    .Y(_06772_),
    .A2(_06768_));
 sg13g2_nand4_1 _15345_ (.B(_06767_),
    .C(_06772_),
    .A(_02442_),
    .Y(_06773_),
    .D(_06751_));
 sg13g2_inv_1 _15346_ (.Y(_06774_),
    .A(_06753_));
 sg13g2_nand4_1 _15347_ (.B(_06767_),
    .C(_06772_),
    .A(_06774_),
    .Y(_06775_),
    .D(_06751_));
 sg13g2_a21oi_2 _15348_ (.B1(_06743_),
    .Y(_06776_),
    .A2(_06775_),
    .A1(_06773_));
 sg13g2_o21ai_1 _15349_ (.B1(_06750_),
    .Y(_06777_),
    .A1(_02442_),
    .A2(_06774_));
 sg13g2_o21ai_1 _15350_ (.B1(_06777_),
    .Y(_06778_),
    .A1(_02443_),
    .A2(_06753_));
 sg13g2_or2_1 _15351_ (.X(_06779_),
    .B(_06778_),
    .A(_06776_));
 sg13g2_nor2b_1 _15352_ (.A(_02448_),
    .B_N(\am_sdr0.cic3.comb1_in_del[14] ),
    .Y(_06780_));
 sg13g2_nor2b_2 _15353_ (.A(\am_sdr0.cic3.comb1_in_del[14] ),
    .B_N(_02448_),
    .Y(_06781_));
 sg13g2_nor2_1 _15354_ (.A(_06780_),
    .B(_06781_),
    .Y(_06782_));
 sg13g2_xnor2_1 _15355_ (.Y(_06783_),
    .A(_06779_),
    .B(_06782_));
 sg13g2_nand2_1 _15356_ (.Y(_06784_),
    .A(_06729_),
    .B(_06783_));
 sg13g2_o21ai_1 _15357_ (.B1(_06784_),
    .Y(_06785_),
    .A1(_06758_),
    .A2(_06728_));
 sg13g2_nor2_1 _15358_ (.A(net71),
    .B(_06785_),
    .Y(_00841_));
 sg13g2_buf_1 _15359_ (.A(_06663_),
    .X(_06786_));
 sg13g2_inv_1 _15360_ (.Y(_06787_),
    .A(_06780_));
 sg13g2_o21ai_1 _15361_ (.B1(_06787_),
    .Y(_06788_),
    .A1(_06779_),
    .A2(_06781_));
 sg13g2_xnor2_1 _15362_ (.Y(_06789_),
    .A(_02452_),
    .B(\am_sdr0.cic3.comb1_in_del[15] ));
 sg13g2_xnor2_1 _15363_ (.Y(_06790_),
    .A(_06788_),
    .B(_06789_));
 sg13g2_buf_2 _15364_ (.A(\am_sdr0.cic3.comb1[15] ),
    .X(_06791_));
 sg13g2_nor2b_1 _15365_ (.A(net271),
    .B_N(_06791_),
    .Y(_06792_));
 sg13g2_a21oi_1 _15366_ (.A1(net206),
    .A2(_06790_),
    .Y(_06793_),
    .B1(_06792_));
 sg13g2_nor2_1 _15367_ (.A(net71),
    .B(_06793_),
    .Y(_00842_));
 sg13g2_buf_1 _15368_ (.A(\am_sdr0.cic3.comb1[16] ),
    .X(_06794_));
 sg13g2_inv_1 _15369_ (.Y(_06795_),
    .A(_06794_));
 sg13g2_inv_1 _15370_ (.Y(_06796_),
    .A(\am_sdr0.cic3.comb1_in_del[15] ));
 sg13g2_nor4_2 _15371_ (.A(_06796_),
    .B(_06776_),
    .C(_06778_),
    .Y(_06797_),
    .D(_06781_));
 sg13g2_nor4_2 _15372_ (.A(_02452_),
    .B(_06776_),
    .C(_06778_),
    .Y(_06798_),
    .D(_06781_));
 sg13g2_a21o_1 _15373_ (.A2(_06796_),
    .A1(_02452_),
    .B1(_06787_),
    .X(_06799_));
 sg13g2_o21ai_1 _15374_ (.B1(_06799_),
    .Y(_06800_),
    .A1(_02452_),
    .A2(_06796_));
 sg13g2_nor3_2 _15375_ (.A(_06797_),
    .B(_06798_),
    .C(_06800_),
    .Y(_06801_));
 sg13g2_buf_1 _15376_ (.A(\am_sdr0.cic3.comb1_in_del[16] ),
    .X(_06802_));
 sg13g2_xnor2_1 _15377_ (.Y(_06803_),
    .A(_02454_),
    .B(_06802_));
 sg13g2_xnor2_1 _15378_ (.Y(_06804_),
    .A(_06801_),
    .B(_06803_));
 sg13g2_buf_1 _15379_ (.A(_06662_),
    .X(_06805_));
 sg13g2_mux2_1 _15380_ (.A0(_06795_),
    .A1(_06804_),
    .S(net268),
    .X(_06806_));
 sg13g2_nor2_1 _15381_ (.A(net71),
    .B(_06806_),
    .Y(_00843_));
 sg13g2_buf_1 _15382_ (.A(\am_sdr0.cic3.comb1[17] ),
    .X(_06807_));
 sg13g2_nor2_1 _15383_ (.A(_06807_),
    .B(net270),
    .Y(_06808_));
 sg13g2_or3_1 _15384_ (.A(_06797_),
    .B(_06798_),
    .C(_06800_),
    .X(_06809_));
 sg13g2_inv_1 _15385_ (.Y(_06810_),
    .A(_06802_));
 sg13g2_a21oi_1 _15386_ (.A1(_06810_),
    .A2(_06801_),
    .Y(_06811_),
    .B1(_02454_));
 sg13g2_a21oi_1 _15387_ (.A1(_06802_),
    .A2(_06809_),
    .Y(_06812_),
    .B1(_06811_));
 sg13g2_xor2_1 _15388_ (.B(\am_sdr0.cic3.comb1_in_del[17] ),
    .A(_02458_),
    .X(_06813_));
 sg13g2_xnor2_1 _15389_ (.Y(_06814_),
    .A(_06812_),
    .B(_06813_));
 sg13g2_nor2_1 _15390_ (.A(net149),
    .B(_06814_),
    .Y(_06815_));
 sg13g2_nor3_1 _15391_ (.A(net191),
    .B(_06808_),
    .C(_06815_),
    .Y(_00844_));
 sg13g2_inv_1 _15392_ (.Y(_06816_),
    .A(\am_sdr0.cic3.comb1_in_del[17] ));
 sg13g2_nor2_1 _15393_ (.A(_02458_),
    .B(_06816_),
    .Y(_06817_));
 sg13g2_a221oi_1 _15394_ (.B2(_06816_),
    .C1(_06801_),
    .B1(_02458_),
    .A1(_02454_),
    .Y(_06818_),
    .A2(_06810_));
 sg13g2_nand2b_1 _15395_ (.Y(_06819_),
    .B(_06802_),
    .A_N(_02454_));
 sg13g2_a21oi_1 _15396_ (.A1(_02458_),
    .A2(_06816_),
    .Y(_06820_),
    .B1(_06819_));
 sg13g2_nor3_1 _15397_ (.A(_06817_),
    .B(_06818_),
    .C(_06820_),
    .Y(_06821_));
 sg13g2_buf_1 _15398_ (.A(\am_sdr0.cic3.comb1_in_del[18] ),
    .X(_06822_));
 sg13g2_xnor2_1 _15399_ (.Y(_06823_),
    .A(_02461_),
    .B(_06822_));
 sg13g2_xnor2_1 _15400_ (.Y(_06824_),
    .A(_06821_),
    .B(_06823_));
 sg13g2_buf_1 _15401_ (.A(\am_sdr0.cic3.comb1[18] ),
    .X(_06825_));
 sg13g2_o21ai_1 _15402_ (.B1(net218),
    .Y(_06826_),
    .A1(_06825_),
    .A2(net270));
 sg13g2_a21oi_1 _15403_ (.A1(net209),
    .A2(_06824_),
    .Y(_00845_),
    .B1(_06826_));
 sg13g2_nor2b_1 _15404_ (.A(_06822_),
    .B_N(_02461_),
    .Y(_06827_));
 sg13g2_nand2b_1 _15405_ (.Y(_06828_),
    .B(_06822_),
    .A_N(_02461_));
 sg13g2_o21ai_1 _15406_ (.B1(_06828_),
    .Y(_06829_),
    .A1(_06821_),
    .A2(_06827_));
 sg13g2_xor2_1 _15407_ (.B(\am_sdr0.cic3.comb1_in_del[19] ),
    .A(\am_sdr0.cic3.integ_sample[19] ),
    .X(_06830_));
 sg13g2_xnor2_1 _15408_ (.Y(_06831_),
    .A(_06829_),
    .B(_06830_));
 sg13g2_o21ai_1 _15409_ (.B1(net218),
    .Y(_06832_),
    .A1(\am_sdr0.cic3.comb1[19] ),
    .A2(net270));
 sg13g2_a21oi_1 _15410_ (.A1(net209),
    .A2(_06831_),
    .Y(_00846_),
    .B1(_06832_));
 sg13g2_buf_2 _15411_ (.A(\am_sdr0.cic3.comb1[1] ),
    .X(_06833_));
 sg13g2_nand2_1 _15412_ (.Y(_06834_),
    .A(_06833_),
    .B(net69));
 sg13g2_xnor2_1 _15413_ (.Y(_06835_),
    .A(_02463_),
    .B(_06681_));
 sg13g2_xnor2_1 _15414_ (.Y(_06836_),
    .A(_06680_),
    .B(_06835_));
 sg13g2_nand2_1 _15415_ (.Y(_06837_),
    .A(net208),
    .B(_06836_));
 sg13g2_a21oi_1 _15416_ (.A1(_06834_),
    .A2(_06837_),
    .Y(_00847_),
    .B1(net70));
 sg13g2_buf_1 _15417_ (.A(\am_sdr0.cic3.comb1[2] ),
    .X(_06838_));
 sg13g2_buf_1 _15418_ (.A(_06672_),
    .X(_06839_));
 sg13g2_a21oi_1 _15419_ (.A1(_06680_),
    .A2(_06682_),
    .Y(_06840_),
    .B1(_06683_));
 sg13g2_xnor2_1 _15420_ (.Y(_06841_),
    .A(\am_sdr0.cic3.integ_sample[2] ),
    .B(_06678_));
 sg13g2_xnor2_1 _15421_ (.Y(_06842_),
    .A(_06840_),
    .B(_06841_));
 sg13g2_nor2_1 _15422_ (.A(net150),
    .B(_06842_),
    .Y(_06843_));
 sg13g2_a21oi_1 _15423_ (.A1(_06838_),
    .A2(net68),
    .Y(_06844_),
    .B1(_06843_));
 sg13g2_nor2_1 _15424_ (.A(net71),
    .B(_06844_),
    .Y(_00848_));
 sg13g2_buf_1 _15425_ (.A(\am_sdr0.cic3.comb1[3] ),
    .X(_06845_));
 sg13g2_nand2_1 _15426_ (.Y(_06846_),
    .A(_06845_),
    .B(net69));
 sg13g2_nor2_1 _15427_ (.A(_06679_),
    .B(_06685_),
    .Y(_06847_));
 sg13g2_xnor2_1 _15428_ (.Y(_06848_),
    .A(_02468_),
    .B(\am_sdr0.cic3.comb1_in_del[3] ));
 sg13g2_xnor2_1 _15429_ (.Y(_06849_),
    .A(_06847_),
    .B(_06848_));
 sg13g2_nand2_1 _15430_ (.Y(_06850_),
    .A(net208),
    .B(_06849_));
 sg13g2_a21oi_1 _15431_ (.A1(_06846_),
    .A2(_06850_),
    .Y(_00849_),
    .B1(_06657_));
 sg13g2_buf_1 _15432_ (.A(\am_sdr0.cic3.comb1[4] ),
    .X(_06851_));
 sg13g2_nor2_1 _15433_ (.A(_06851_),
    .B(net270),
    .Y(_06852_));
 sg13g2_nand2_1 _15434_ (.Y(_06853_),
    .A(_06691_),
    .B(_06694_));
 sg13g2_xor2_1 _15435_ (.B(_06853_),
    .A(_06690_),
    .X(_06854_));
 sg13g2_nor2_1 _15436_ (.A(net149),
    .B(_06854_),
    .Y(_06855_));
 sg13g2_nor3_1 _15437_ (.A(net191),
    .B(_06852_),
    .C(_06855_),
    .Y(_00850_));
 sg13g2_buf_2 _15438_ (.A(\am_sdr0.cic3.comb1[5] ),
    .X(_06856_));
 sg13g2_nand2_1 _15439_ (.Y(_06857_),
    .A(_06690_),
    .B(_06691_));
 sg13g2_nand2_1 _15440_ (.Y(_06858_),
    .A(_06857_),
    .B(_06694_));
 sg13g2_xor2_1 _15441_ (.B(_06692_),
    .A(_02473_),
    .X(_06859_));
 sg13g2_xnor2_1 _15442_ (.Y(_06860_),
    .A(_06858_),
    .B(_06859_));
 sg13g2_nand2_1 _15443_ (.Y(_06861_),
    .A(net269),
    .B(_06860_));
 sg13g2_o21ai_1 _15444_ (.B1(_06861_),
    .Y(_06862_),
    .A1(_06856_),
    .A2(net207));
 sg13g2_nor2_1 _15445_ (.A(_06635_),
    .B(_06862_),
    .Y(_00851_));
 sg13g2_buf_1 _15446_ (.A(\am_sdr0.cic3.comb1[6] ),
    .X(_06863_));
 sg13g2_nor2_1 _15447_ (.A(_06692_),
    .B(_06858_),
    .Y(_06864_));
 sg13g2_nand2_1 _15448_ (.Y(_06865_),
    .A(_06692_),
    .B(_06858_));
 sg13g2_o21ai_1 _15449_ (.B1(_06865_),
    .Y(_06866_),
    .A1(_02473_),
    .A2(_06864_));
 sg13g2_buf_1 _15450_ (.A(_06866_),
    .X(_06867_));
 sg13g2_xor2_1 _15451_ (.B(_06704_),
    .A(_02476_),
    .X(_06868_));
 sg13g2_xnor2_1 _15452_ (.Y(_06869_),
    .A(_06867_),
    .B(_06868_));
 sg13g2_nand2_1 _15453_ (.Y(_06870_),
    .A(net269),
    .B(_06869_));
 sg13g2_o21ai_1 _15454_ (.B1(_06870_),
    .Y(_06871_),
    .A1(_06863_),
    .A2(net207));
 sg13g2_nor2_1 _15455_ (.A(_06635_),
    .B(_06871_),
    .Y(_00852_));
 sg13g2_buf_1 _15456_ (.A(_06365_),
    .X(_06872_));
 sg13g2_buf_1 _15457_ (.A(\am_sdr0.cic3.comb1[7] ),
    .X(_06873_));
 sg13g2_nor2_1 _15458_ (.A(_06704_),
    .B(_06867_),
    .Y(_06874_));
 sg13g2_nand2_1 _15459_ (.Y(_06875_),
    .A(_06704_),
    .B(_06867_));
 sg13g2_o21ai_1 _15460_ (.B1(_06875_),
    .Y(_06876_),
    .A1(_02476_),
    .A2(_06874_));
 sg13g2_buf_1 _15461_ (.A(_06876_),
    .X(_06877_));
 sg13g2_nand2_1 _15462_ (.Y(_06878_),
    .A(_06699_),
    .B(_06710_));
 sg13g2_xnor2_1 _15463_ (.Y(_06879_),
    .A(_06877_),
    .B(_06878_));
 sg13g2_nand2_1 _15464_ (.Y(_06880_),
    .A(net269),
    .B(_06879_));
 sg13g2_o21ai_1 _15465_ (.B1(_06880_),
    .Y(_06881_),
    .A1(_06873_),
    .A2(net207));
 sg13g2_nor2_1 _15466_ (.A(net67),
    .B(_06881_),
    .Y(_00853_));
 sg13g2_buf_1 _15467_ (.A(\am_sdr0.cic3.comb1[8] ),
    .X(_06882_));
 sg13g2_nand2_1 _15468_ (.Y(_06883_),
    .A(_06697_),
    .B(_06877_));
 sg13g2_nor2_1 _15469_ (.A(_06697_),
    .B(_06877_),
    .Y(_06884_));
 sg13g2_a21oi_1 _15470_ (.A1(_02478_),
    .A2(_06883_),
    .Y(_06885_),
    .B1(_06884_));
 sg13g2_xor2_1 _15471_ (.B(_06700_),
    .A(_02479_),
    .X(_06886_));
 sg13g2_xnor2_1 _15472_ (.Y(_06887_),
    .A(_06885_),
    .B(_06886_));
 sg13g2_nand2_1 _15473_ (.Y(_06888_),
    .A(net269),
    .B(_06887_));
 sg13g2_o21ai_1 _15474_ (.B1(_06888_),
    .Y(_06889_),
    .A1(_06882_),
    .A2(net207));
 sg13g2_nor2_1 _15475_ (.A(net67),
    .B(_06889_),
    .Y(_00854_));
 sg13g2_buf_1 _15476_ (.A(\am_sdr0.cic3.comb1[9] ),
    .X(_06890_));
 sg13g2_nand2_1 _15477_ (.Y(_06891_),
    .A(_06890_),
    .B(net69));
 sg13g2_nor2_1 _15478_ (.A(_06708_),
    .B(_06715_),
    .Y(_06892_));
 sg13g2_xnor2_1 _15479_ (.Y(_06893_),
    .A(_02483_),
    .B(_06716_));
 sg13g2_xnor2_1 _15480_ (.Y(_06894_),
    .A(_06892_),
    .B(_06893_));
 sg13g2_nand2_1 _15481_ (.Y(_06895_),
    .A(net208),
    .B(_06894_));
 sg13g2_a21oi_1 _15482_ (.A1(_06891_),
    .A2(_06895_),
    .Y(_00855_),
    .B1(_06657_));
 sg13g2_buf_1 _15483_ (.A(net271),
    .X(_06896_));
 sg13g2_nand2_1 _15484_ (.Y(_06897_),
    .A(_02421_),
    .B(net205));
 sg13g2_nand2_1 _15485_ (.Y(_06898_),
    .A(\am_sdr0.cic3.comb1_in_del[0] ),
    .B(net68));
 sg13g2_a21oi_1 _15486_ (.A1(_06897_),
    .A2(_06898_),
    .Y(_00856_),
    .B1(net70));
 sg13g2_nand2_1 _15487_ (.Y(_06899_),
    .A(_02433_),
    .B(net205));
 sg13g2_nand2_1 _15488_ (.Y(_06900_),
    .A(_06721_),
    .B(net68));
 sg13g2_a21oi_1 _15489_ (.A1(_06899_),
    .A2(_06900_),
    .Y(_00857_),
    .B1(net70));
 sg13g2_nand2_1 _15490_ (.Y(_06901_),
    .A(_02439_),
    .B(net205));
 sg13g2_nand2_1 _15491_ (.Y(_06902_),
    .A(net326),
    .B(net68));
 sg13g2_a21oi_1 _15492_ (.A1(_06901_),
    .A2(_06902_),
    .Y(_00858_),
    .B1(net70));
 sg13g2_nand2_1 _15493_ (.Y(_06903_),
    .A(_02441_),
    .B(net205));
 sg13g2_nand2_1 _15494_ (.Y(_06904_),
    .A(_06745_),
    .B(net68));
 sg13g2_buf_1 _15495_ (.A(_05813_),
    .X(_06905_));
 sg13g2_a21oi_1 _15496_ (.A1(_06903_),
    .A2(_06904_),
    .Y(_00859_),
    .B1(net66));
 sg13g2_nand2_1 _15497_ (.Y(_06906_),
    .A(_02442_),
    .B(net205));
 sg13g2_nand2_1 _15498_ (.Y(_06907_),
    .A(_06753_),
    .B(net68));
 sg13g2_a21oi_1 _15499_ (.A1(_06906_),
    .A2(_06907_),
    .Y(_00860_),
    .B1(net66));
 sg13g2_nand2_1 _15500_ (.Y(_06908_),
    .A(_02448_),
    .B(net205));
 sg13g2_nand2_1 _15501_ (.Y(_06909_),
    .A(\am_sdr0.cic3.comb1_in_del[14] ),
    .B(net68));
 sg13g2_a21oi_1 _15502_ (.A1(_06908_),
    .A2(_06909_),
    .Y(_00861_),
    .B1(net66));
 sg13g2_nand2_1 _15503_ (.Y(_06910_),
    .A(_02452_),
    .B(net205));
 sg13g2_buf_1 _15504_ (.A(net150),
    .X(_06911_));
 sg13g2_nand2_1 _15505_ (.Y(_06912_),
    .A(\am_sdr0.cic3.comb1_in_del[15] ),
    .B(net65));
 sg13g2_a21oi_1 _15506_ (.A1(_06910_),
    .A2(_06912_),
    .Y(_00862_),
    .B1(net66));
 sg13g2_nand2_1 _15507_ (.Y(_06913_),
    .A(_02454_),
    .B(net205));
 sg13g2_nand2_1 _15508_ (.Y(_06914_),
    .A(_06802_),
    .B(net65));
 sg13g2_a21oi_1 _15509_ (.A1(_06913_),
    .A2(_06914_),
    .Y(_00863_),
    .B1(net66));
 sg13g2_nand2_1 _15510_ (.Y(_06915_),
    .A(_02458_),
    .B(_06896_));
 sg13g2_nand2_1 _15511_ (.Y(_06916_),
    .A(\am_sdr0.cic3.comb1_in_del[17] ),
    .B(net65));
 sg13g2_a21oi_1 _15512_ (.A1(_06915_),
    .A2(_06916_),
    .Y(_00864_),
    .B1(_06905_));
 sg13g2_nand2_1 _15513_ (.Y(_06917_),
    .A(_02461_),
    .B(_06896_));
 sg13g2_nand2_1 _15514_ (.Y(_06918_),
    .A(_06822_),
    .B(_06911_));
 sg13g2_a21oi_1 _15515_ (.A1(_06917_),
    .A2(_06918_),
    .Y(_00865_),
    .B1(_06905_));
 sg13g2_buf_1 _15516_ (.A(_06675_),
    .X(_06919_));
 sg13g2_nand2_1 _15517_ (.Y(_06920_),
    .A(\am_sdr0.cic3.integ_sample[19] ),
    .B(_06919_));
 sg13g2_nand2_1 _15518_ (.Y(_06921_),
    .A(\am_sdr0.cic3.comb1_in_del[19] ),
    .B(_06911_));
 sg13g2_a21oi_1 _15519_ (.A1(_06920_),
    .A2(_06921_),
    .Y(_00866_),
    .B1(net66));
 sg13g2_nand2_1 _15520_ (.Y(_06922_),
    .A(_02463_),
    .B(net204));
 sg13g2_nand2_1 _15521_ (.Y(_06923_),
    .A(_06681_),
    .B(net65));
 sg13g2_a21oi_1 _15522_ (.A1(_06922_),
    .A2(_06923_),
    .Y(_00867_),
    .B1(net66));
 sg13g2_nand2_1 _15523_ (.Y(_06924_),
    .A(\am_sdr0.cic3.integ_sample[2] ),
    .B(net204));
 sg13g2_nand2_1 _15524_ (.Y(_06925_),
    .A(_06678_),
    .B(net65));
 sg13g2_a21oi_1 _15525_ (.A1(_06924_),
    .A2(_06925_),
    .Y(_00868_),
    .B1(net66));
 sg13g2_nand2_1 _15526_ (.Y(_06926_),
    .A(_02468_),
    .B(net204));
 sg13g2_nand2_1 _15527_ (.Y(_06927_),
    .A(\am_sdr0.cic3.comb1_in_del[3] ),
    .B(net65));
 sg13g2_buf_1 _15528_ (.A(_05813_),
    .X(_06928_));
 sg13g2_a21oi_1 _15529_ (.A1(_06926_),
    .A2(_06927_),
    .Y(_00869_),
    .B1(net64));
 sg13g2_nand2_1 _15530_ (.Y(_06929_),
    .A(_02471_),
    .B(net204));
 sg13g2_nand2_1 _15531_ (.Y(_06930_),
    .A(\am_sdr0.cic3.comb1_in_del[4] ),
    .B(net65));
 sg13g2_a21oi_1 _15532_ (.A1(_06929_),
    .A2(_06930_),
    .Y(_00870_),
    .B1(net64));
 sg13g2_nand2_1 _15533_ (.Y(_06931_),
    .A(_02473_),
    .B(net204));
 sg13g2_nand2_1 _15534_ (.Y(_06932_),
    .A(_06692_),
    .B(net65));
 sg13g2_a21oi_1 _15535_ (.A1(_06931_),
    .A2(_06932_),
    .Y(_00871_),
    .B1(net64));
 sg13g2_nand2_1 _15536_ (.Y(_06933_),
    .A(_02476_),
    .B(net204));
 sg13g2_buf_1 _15537_ (.A(net150),
    .X(_06934_));
 sg13g2_nand2_1 _15538_ (.Y(_06935_),
    .A(_06704_),
    .B(net63));
 sg13g2_a21oi_1 _15539_ (.A1(_06933_),
    .A2(_06935_),
    .Y(_00872_),
    .B1(net64));
 sg13g2_nand2_1 _15540_ (.Y(_06936_),
    .A(_02478_),
    .B(net204));
 sg13g2_nand2_1 _15541_ (.Y(_06937_),
    .A(_06697_),
    .B(net63));
 sg13g2_a21oi_1 _15542_ (.A1(_06936_),
    .A2(_06937_),
    .Y(_00873_),
    .B1(net64));
 sg13g2_nand2_1 _15543_ (.Y(_06938_),
    .A(_02479_),
    .B(net204));
 sg13g2_nand2_1 _15544_ (.Y(_06939_),
    .A(_06700_),
    .B(net63));
 sg13g2_a21oi_1 _15545_ (.A1(_06938_),
    .A2(_06939_),
    .Y(_00874_),
    .B1(net64));
 sg13g2_nand2_1 _15546_ (.Y(_06940_),
    .A(_02483_),
    .B(_06919_));
 sg13g2_nand2_1 _15547_ (.Y(_06941_),
    .A(_06716_),
    .B(net63));
 sg13g2_a21oi_1 _15548_ (.A1(_06940_),
    .A2(_06941_),
    .Y(_00875_),
    .B1(net64));
 sg13g2_xnor2_1 _15549_ (.Y(_06942_),
    .A(_06666_),
    .B(\am_sdr0.cic3.comb2_in_del[0] ));
 sg13g2_o21ai_1 _15550_ (.B1(net218),
    .Y(_06943_),
    .A1(\am_sdr0.cic3.comb2[0] ),
    .A2(_06805_));
 sg13g2_a21oi_1 _15551_ (.A1(net209),
    .A2(_06942_),
    .Y(_00876_),
    .B1(_06943_));
 sg13g2_buf_1 _15552_ (.A(\am_sdr0.cic3.comb2[10] ),
    .X(_06944_));
 sg13g2_nand2_1 _15553_ (.Y(_06945_),
    .A(_06944_),
    .B(_06673_));
 sg13g2_buf_1 _15554_ (.A(\am_sdr0.cic3.comb2_in_del[8] ),
    .X(_06946_));
 sg13g2_buf_1 _15555_ (.A(\am_sdr0.cic3.comb2_in_del[9] ),
    .X(_06947_));
 sg13g2_nor2_1 _15556_ (.A(_06946_),
    .B(_06947_),
    .Y(_06948_));
 sg13g2_nor2b_1 _15557_ (.A(_06947_),
    .B_N(_06882_),
    .Y(_06949_));
 sg13g2_buf_1 _15558_ (.A(\am_sdr0.cic3.comb2_in_del[5] ),
    .X(_06950_));
 sg13g2_inv_1 _15559_ (.Y(_06951_),
    .A(_06950_));
 sg13g2_buf_1 _15560_ (.A(\am_sdr0.cic3.comb2_in_del[4] ),
    .X(_06952_));
 sg13g2_nand2b_1 _15561_ (.Y(_06953_),
    .B(_06952_),
    .A_N(_06851_));
 sg13g2_inv_1 _15562_ (.Y(_06954_),
    .A(_06845_));
 sg13g2_inv_1 _15563_ (.Y(_06955_),
    .A(\am_sdr0.cic3.comb2_in_del[3] ));
 sg13g2_inv_1 _15564_ (.Y(_06956_),
    .A(_06838_));
 sg13g2_buf_1 _15565_ (.A(\am_sdr0.cic3.comb2_in_del[2] ),
    .X(_06957_));
 sg13g2_nor2_1 _15566_ (.A(_06956_),
    .B(_06957_),
    .Y(_06958_));
 sg13g2_nor2b_1 _15567_ (.A(_06666_),
    .B_N(\am_sdr0.cic3.comb2_in_del[0] ),
    .Y(_06959_));
 sg13g2_buf_1 _15568_ (.A(\am_sdr0.cic3.comb2_in_del[1] ),
    .X(_06960_));
 sg13g2_nand2b_1 _15569_ (.Y(_06961_),
    .B(_06833_),
    .A_N(_06960_));
 sg13g2_nor2b_1 _15570_ (.A(_06833_),
    .B_N(_06960_),
    .Y(_06962_));
 sg13g2_a221oi_1 _15571_ (.B2(_06961_),
    .C1(_06962_),
    .B1(_06959_),
    .A1(_06956_),
    .Y(_06963_),
    .A2(_06957_));
 sg13g2_buf_1 _15572_ (.A(_06963_),
    .X(_06964_));
 sg13g2_nor3_1 _15573_ (.A(_06955_),
    .B(_06958_),
    .C(_06964_),
    .Y(_06965_));
 sg13g2_o21ai_1 _15574_ (.B1(_06955_),
    .Y(_06966_),
    .A1(_06958_),
    .A2(_06964_));
 sg13g2_o21ai_1 _15575_ (.B1(_06966_),
    .Y(_06967_),
    .A1(_06954_),
    .A2(_06965_));
 sg13g2_buf_2 _15576_ (.A(_06967_),
    .X(_06968_));
 sg13g2_nor2b_1 _15577_ (.A(\am_sdr0.cic3.comb2_in_del[6] ),
    .B_N(_06863_),
    .Y(_06969_));
 sg13g2_nor2b_1 _15578_ (.A(_06952_),
    .B_N(_06851_),
    .Y(_06970_));
 sg13g2_or2_1 _15579_ (.X(_06971_),
    .B(_06970_),
    .A(_06969_));
 sg13g2_a221oi_1 _15580_ (.B2(_06968_),
    .C1(_06971_),
    .B1(_06953_),
    .A1(_06856_),
    .Y(_06972_),
    .A2(_06951_));
 sg13g2_buf_1 _15581_ (.A(_06972_),
    .X(_06973_));
 sg13g2_nand2b_1 _15582_ (.Y(_06974_),
    .B(_06950_),
    .A_N(_06856_));
 sg13g2_nand2b_1 _15583_ (.Y(_06975_),
    .B(\am_sdr0.cic3.comb2_in_del[6] ),
    .A_N(_06863_));
 sg13g2_o21ai_1 _15584_ (.B1(_06975_),
    .Y(_06976_),
    .A1(_06969_),
    .A2(_06974_));
 sg13g2_buf_1 _15585_ (.A(\am_sdr0.cic3.comb2_in_del[7] ),
    .X(_06977_));
 sg13g2_o21ai_1 _15586_ (.B1(_06977_),
    .Y(_06978_),
    .A1(_06973_),
    .A2(_06976_));
 sg13g2_nor3_1 _15587_ (.A(_06977_),
    .B(_06973_),
    .C(_06976_),
    .Y(_06979_));
 sg13g2_a21o_1 _15588_ (.A2(_06978_),
    .A1(_06873_),
    .B1(_06979_),
    .X(_06980_));
 sg13g2_buf_2 _15589_ (.A(_06980_),
    .X(_06981_));
 sg13g2_o21ai_1 _15590_ (.B1(_06981_),
    .Y(_06982_),
    .A1(_06948_),
    .A2(_06949_));
 sg13g2_inv_1 _15591_ (.Y(_06983_),
    .A(_06947_));
 sg13g2_nor2b_1 _15592_ (.A(_06946_),
    .B_N(_06882_),
    .Y(_06984_));
 sg13g2_a21oi_1 _15593_ (.A1(_06983_),
    .A2(_06984_),
    .Y(_06985_),
    .B1(_06890_));
 sg13g2_inv_1 _15594_ (.Y(_06986_),
    .A(_06946_));
 sg13g2_a21oi_1 _15595_ (.A1(_06986_),
    .A2(_06981_),
    .Y(_06987_),
    .B1(_06983_));
 sg13g2_o21ai_1 _15596_ (.B1(_06882_),
    .Y(_06988_),
    .A1(_06986_),
    .A2(_06981_));
 sg13g2_buf_1 _15597_ (.A(_06988_),
    .X(_06989_));
 sg13g2_a22oi_1 _15598_ (.Y(_06990_),
    .B1(_06987_),
    .B2(_06989_),
    .A2(_06985_),
    .A1(_06982_));
 sg13g2_buf_1 _15599_ (.A(_06990_),
    .X(_06991_));
 sg13g2_buf_1 _15600_ (.A(\am_sdr0.cic3.comb2_in_del[10] ),
    .X(_06992_));
 sg13g2_xor2_1 _15601_ (.B(_06992_),
    .A(_06669_),
    .X(_06993_));
 sg13g2_xnor2_1 _15602_ (.Y(_06994_),
    .A(_06991_),
    .B(_06993_));
 sg13g2_nand2_1 _15603_ (.Y(_06995_),
    .A(_06676_),
    .B(_06994_));
 sg13g2_a21oi_1 _15604_ (.A1(_06945_),
    .A2(_06995_),
    .Y(_00877_),
    .B1(net64));
 sg13g2_buf_1 _15605_ (.A(\am_sdr0.cic3.comb2[11] ),
    .X(_06996_));
 sg13g2_nor2_1 _15606_ (.A(_06996_),
    .B(net270),
    .Y(_06997_));
 sg13g2_inv_1 _15607_ (.Y(_06998_),
    .A(_06992_));
 sg13g2_a21oi_1 _15608_ (.A1(_06998_),
    .A2(_06991_),
    .Y(_06999_),
    .B1(_06669_));
 sg13g2_nor2_1 _15609_ (.A(_06998_),
    .B(_06991_),
    .Y(_07000_));
 sg13g2_nor2_1 _15610_ (.A(_06999_),
    .B(_07000_),
    .Y(_07001_));
 sg13g2_buf_1 _15611_ (.A(\am_sdr0.cic3.comb2_in_del[11] ),
    .X(_07002_));
 sg13g2_nor2b_1 _15612_ (.A(_07002_),
    .B_N(_06727_),
    .Y(_07003_));
 sg13g2_nand2b_1 _15613_ (.Y(_07004_),
    .B(_07002_),
    .A_N(_06727_));
 sg13g2_nor2b_1 _15614_ (.A(_07003_),
    .B_N(_07004_),
    .Y(_07005_));
 sg13g2_xor2_1 _15615_ (.B(_07005_),
    .A(_07001_),
    .X(_07006_));
 sg13g2_nor2_1 _15616_ (.A(net149),
    .B(_07006_),
    .Y(_07007_));
 sg13g2_nor3_1 _15617_ (.A(net191),
    .B(_06997_),
    .C(_07007_),
    .Y(_00878_));
 sg13g2_buf_1 _15618_ (.A(\am_sdr0.cic3.comb2[12] ),
    .X(_07008_));
 sg13g2_nor2_1 _15619_ (.A(_07008_),
    .B(_06667_),
    .Y(_07009_));
 sg13g2_o21ai_1 _15620_ (.B1(_07002_),
    .Y(_07010_),
    .A1(_06999_),
    .A2(_07000_));
 sg13g2_nor3_1 _15621_ (.A(_07002_),
    .B(_06999_),
    .C(_07000_),
    .Y(_07011_));
 sg13g2_a21oi_2 _15622_ (.B1(_07011_),
    .Y(_07012_),
    .A2(_07010_),
    .A1(_06727_));
 sg13g2_inv_1 _15623_ (.Y(_07013_),
    .A(\am_sdr0.cic3.comb1[12] ));
 sg13g2_buf_2 _15624_ (.A(\am_sdr0.cic3.comb2_in_del[12] ),
    .X(_07014_));
 sg13g2_nor2_1 _15625_ (.A(_07013_),
    .B(_07014_),
    .Y(_07015_));
 sg13g2_nand2_1 _15626_ (.Y(_07016_),
    .A(_07013_),
    .B(_07014_));
 sg13g2_nor2b_1 _15627_ (.A(_07015_),
    .B_N(_07016_),
    .Y(_07017_));
 sg13g2_xnor2_1 _15628_ (.Y(_07018_),
    .A(_07012_),
    .B(_07017_));
 sg13g2_nor2_1 _15629_ (.A(_06737_),
    .B(_07018_),
    .Y(_07019_));
 sg13g2_nor3_1 _15630_ (.A(net191),
    .B(_07009_),
    .C(_07019_),
    .Y(_00879_));
 sg13g2_buf_1 _15631_ (.A(\am_sdr0.cic3.comb2[13] ),
    .X(_07020_));
 sg13g2_nand2_1 _15632_ (.Y(_07021_),
    .A(_07020_),
    .B(net150));
 sg13g2_nand2_1 _15633_ (.Y(_07022_),
    .A(_07014_),
    .B(_07012_));
 sg13g2_o21ai_1 _15634_ (.B1(_07013_),
    .Y(_07023_),
    .A1(_07014_),
    .A2(_07012_));
 sg13g2_nand2b_1 _15635_ (.Y(_07024_),
    .B(_06749_),
    .A_N(\am_sdr0.cic3.comb2_in_del[13] ));
 sg13g2_buf_1 _15636_ (.A(_07024_),
    .X(_07025_));
 sg13g2_nand2b_1 _15637_ (.Y(_07026_),
    .B(\am_sdr0.cic3.comb2_in_del[13] ),
    .A_N(_06749_));
 sg13g2_buf_1 _15638_ (.A(_07026_),
    .X(_07027_));
 sg13g2_a21oi_1 _15639_ (.A1(_07025_),
    .A2(_07027_),
    .Y(_07028_),
    .B1(_06671_));
 sg13g2_nand3_1 _15640_ (.B(_07023_),
    .C(_07028_),
    .A(_07022_),
    .Y(_07029_));
 sg13g2_nand3_1 _15641_ (.B(_07025_),
    .C(_07027_),
    .A(_06662_),
    .Y(_07030_));
 sg13g2_a21o_1 _15642_ (.A2(_07023_),
    .A1(_07022_),
    .B1(_07030_),
    .X(_07031_));
 sg13g2_nand3_1 _15643_ (.B(_07029_),
    .C(_07031_),
    .A(_07021_),
    .Y(_07032_));
 sg13g2_and2_1 _15644_ (.A(net210),
    .B(_07032_),
    .X(_00880_));
 sg13g2_buf_1 _15645_ (.A(\am_sdr0.cic3.comb2[14] ),
    .X(_07033_));
 sg13g2_nand2_1 _15646_ (.Y(_07034_),
    .A(_07033_),
    .B(net69));
 sg13g2_and4_1 _15647_ (.A(_07005_),
    .B(_07017_),
    .C(_07025_),
    .D(_07027_),
    .X(_07035_));
 sg13g2_buf_1 _15648_ (.A(_07035_),
    .X(_07036_));
 sg13g2_nor2b_1 _15649_ (.A(_06993_),
    .B_N(_07036_),
    .Y(_07037_));
 sg13g2_nor2b_1 _15650_ (.A(_06992_),
    .B_N(_06669_),
    .Y(_07038_));
 sg13g2_a21oi_1 _15651_ (.A1(_07038_),
    .A2(_07004_),
    .Y(_07039_),
    .B1(_07003_));
 sg13g2_nand2_1 _15652_ (.Y(_07040_),
    .A(_07014_),
    .B(_07039_));
 sg13g2_o21ai_1 _15653_ (.B1(_07013_),
    .Y(_07041_),
    .A1(_07014_),
    .A2(_07039_));
 sg13g2_nand3_1 _15654_ (.B(_07040_),
    .C(_07041_),
    .A(_07027_),
    .Y(_07042_));
 sg13g2_nand2_1 _15655_ (.Y(_07043_),
    .A(_07025_),
    .B(_07042_));
 sg13g2_a21oi_1 _15656_ (.A1(_06991_),
    .A2(_07037_),
    .Y(_07044_),
    .B1(_07043_));
 sg13g2_buf_1 _15657_ (.A(\am_sdr0.cic3.comb2_in_del[14] ),
    .X(_07045_));
 sg13g2_xnor2_1 _15658_ (.Y(_07046_),
    .A(_06758_),
    .B(_07045_));
 sg13g2_xnor2_1 _15659_ (.Y(_07047_),
    .A(_07044_),
    .B(_07046_));
 sg13g2_nand2_1 _15660_ (.Y(_07048_),
    .A(net208),
    .B(_07047_));
 sg13g2_a21oi_1 _15661_ (.A1(_07034_),
    .A2(_07048_),
    .Y(_00881_),
    .B1(_06928_));
 sg13g2_buf_1 _15662_ (.A(\am_sdr0.cic3.comb2[15] ),
    .X(_07049_));
 sg13g2_nand2_1 _15663_ (.Y(_07050_),
    .A(_07049_),
    .B(_06673_));
 sg13g2_inv_1 _15664_ (.Y(_07051_),
    .A(_07045_));
 sg13g2_a21oi_1 _15665_ (.A1(_07051_),
    .A2(_07043_),
    .Y(_07052_),
    .B1(_06758_));
 sg13g2_nand3_1 _15666_ (.B(_06991_),
    .C(_07037_),
    .A(_07051_),
    .Y(_07053_));
 sg13g2_buf_1 _15667_ (.A(_07053_),
    .X(_07054_));
 sg13g2_nand2_1 _15668_ (.Y(_07055_),
    .A(_07038_),
    .B(_07036_));
 sg13g2_a21oi_1 _15669_ (.A1(_07003_),
    .A2(_07016_),
    .Y(_07056_),
    .B1(_07015_));
 sg13g2_nand2b_1 _15670_ (.Y(_07057_),
    .B(_07027_),
    .A_N(_07056_));
 sg13g2_nand4_1 _15671_ (.B(_07025_),
    .C(_07055_),
    .A(_07045_),
    .Y(_07058_),
    .D(_07057_));
 sg13g2_nand2_1 _15672_ (.Y(_07059_),
    .A(_06998_),
    .B(_07036_));
 sg13g2_a221oi_1 _15673_ (.B2(_06989_),
    .C1(_07059_),
    .B1(_06987_),
    .A1(_06982_),
    .Y(_07060_),
    .A2(_06985_));
 sg13g2_nand2_1 _15674_ (.Y(_07061_),
    .A(_06669_),
    .B(_07036_));
 sg13g2_a221oi_1 _15675_ (.B2(_06989_),
    .C1(_07061_),
    .B1(_06987_),
    .A1(_06982_),
    .Y(_07062_),
    .A2(_06985_));
 sg13g2_nor3_1 _15676_ (.A(_07058_),
    .B(_07060_),
    .C(_07062_),
    .Y(_07063_));
 sg13g2_a21o_1 _15677_ (.A2(_07054_),
    .A1(_07052_),
    .B1(_07063_),
    .X(_07064_));
 sg13g2_buf_1 _15678_ (.A(_07064_),
    .X(_07065_));
 sg13g2_buf_2 _15679_ (.A(\am_sdr0.cic3.comb2_in_del[15] ),
    .X(_07066_));
 sg13g2_xnor2_1 _15680_ (.Y(_07067_),
    .A(_06791_),
    .B(_07066_));
 sg13g2_xnor2_1 _15681_ (.Y(_07068_),
    .A(_07065_),
    .B(_07067_));
 sg13g2_nand2_1 _15682_ (.Y(_07069_),
    .A(_06676_),
    .B(_07068_));
 sg13g2_a21oi_1 _15683_ (.A1(_07050_),
    .A2(_07069_),
    .Y(_00882_),
    .B1(_06928_));
 sg13g2_nor2_1 _15684_ (.A(_07066_),
    .B(_07065_),
    .Y(_07070_));
 sg13g2_nand2_1 _15685_ (.Y(_07071_),
    .A(_07066_),
    .B(_07065_));
 sg13g2_o21ai_1 _15686_ (.B1(_07071_),
    .Y(_07072_),
    .A1(_06791_),
    .A2(_07070_));
 sg13g2_buf_1 _15687_ (.A(\am_sdr0.cic3.comb2_in_del[16] ),
    .X(_07073_));
 sg13g2_xor2_1 _15688_ (.B(_07073_),
    .A(_06794_),
    .X(_07074_));
 sg13g2_xnor2_1 _15689_ (.Y(_07075_),
    .A(_07072_),
    .B(_07074_));
 sg13g2_buf_1 _15690_ (.A(\am_sdr0.cic3.comb2[16] ),
    .X(_07076_));
 sg13g2_o21ai_1 _15691_ (.B1(_05549_),
    .Y(_07077_),
    .A1(_07076_),
    .A2(_06805_));
 sg13g2_a21oi_1 _15692_ (.A1(net209),
    .A2(_07075_),
    .Y(_00883_),
    .B1(_07077_));
 sg13g2_buf_1 _15693_ (.A(\am_sdr0.cic3.comb2[17] ),
    .X(_07078_));
 sg13g2_nor2_1 _15694_ (.A(_06795_),
    .B(_07073_),
    .Y(_07079_));
 sg13g2_or2_1 _15695_ (.X(_07080_),
    .B(_07073_),
    .A(_07066_));
 sg13g2_nand2b_1 _15696_ (.Y(_07081_),
    .B(_06791_),
    .A_N(_07073_));
 sg13g2_a221oi_1 _15697_ (.B2(_07081_),
    .C1(_07063_),
    .B1(_07080_),
    .A1(_07052_),
    .Y(_07082_),
    .A2(_07054_));
 sg13g2_nand2b_1 _15698_ (.Y(_07083_),
    .B(_06794_),
    .A_N(_07066_));
 sg13g2_nand2_1 _15699_ (.Y(_07084_),
    .A(_06791_),
    .B(_06794_));
 sg13g2_a221oi_1 _15700_ (.B2(_07084_),
    .C1(_07063_),
    .B1(_07083_),
    .A1(_07052_),
    .Y(_07085_),
    .A2(_07054_));
 sg13g2_nand2b_1 _15701_ (.Y(_07086_),
    .B(_06791_),
    .A_N(_07066_));
 sg13g2_a21oi_1 _15702_ (.A1(_06795_),
    .A2(_07073_),
    .Y(_07087_),
    .B1(_07086_));
 sg13g2_nor4_2 _15703_ (.A(_07079_),
    .B(_07082_),
    .C(_07085_),
    .Y(_07088_),
    .D(_07087_));
 sg13g2_nor2b_1 _15704_ (.A(_06807_),
    .B_N(\am_sdr0.cic3.comb2_in_del[17] ),
    .Y(_07089_));
 sg13g2_nand2b_1 _15705_ (.Y(_07090_),
    .B(_06807_),
    .A_N(\am_sdr0.cic3.comb2_in_del[17] ));
 sg13g2_nand2b_1 _15706_ (.Y(_07091_),
    .B(_07090_),
    .A_N(_07089_));
 sg13g2_xnor2_1 _15707_ (.Y(_07092_),
    .A(_07088_),
    .B(_07091_));
 sg13g2_nand2_1 _15708_ (.Y(_07093_),
    .A(_06729_),
    .B(_07092_));
 sg13g2_o21ai_1 _15709_ (.B1(_07093_),
    .Y(_07094_),
    .A1(_07078_),
    .A2(net207));
 sg13g2_nor2_1 _15710_ (.A(net67),
    .B(_07094_),
    .Y(_00884_));
 sg13g2_buf_1 _15711_ (.A(\am_sdr0.cic3.comb2[18] ),
    .X(_07095_));
 sg13g2_nor2_1 _15712_ (.A(_07095_),
    .B(net270),
    .Y(_07096_));
 sg13g2_buf_1 _15713_ (.A(\am_sdr0.cic3.comb2_in_del[18] ),
    .X(_07097_));
 sg13g2_xor2_1 _15714_ (.B(_07097_),
    .A(_06825_),
    .X(_07098_));
 sg13g2_a21oi_1 _15715_ (.A1(_07088_),
    .A2(_07090_),
    .Y(_07099_),
    .B1(_07089_));
 sg13g2_xnor2_1 _15716_ (.Y(_07100_),
    .A(_07098_),
    .B(_07099_));
 sg13g2_nor2_1 _15717_ (.A(net149),
    .B(_07100_),
    .Y(_07101_));
 sg13g2_nor3_1 _15718_ (.A(_01446_),
    .B(_07096_),
    .C(_07101_),
    .Y(_00885_));
 sg13g2_nand2b_1 _15719_ (.Y(_07102_),
    .B(_07097_),
    .A_N(_06825_));
 sg13g2_nor2b_1 _15720_ (.A(_07097_),
    .B_N(_06825_),
    .Y(_07103_));
 sg13g2_a21oi_1 _15721_ (.A1(_07102_),
    .A2(_07099_),
    .Y(_07104_),
    .B1(_07103_));
 sg13g2_xor2_1 _15722_ (.B(\am_sdr0.cic3.comb2_in_del[19] ),
    .A(\am_sdr0.cic3.comb1[19] ),
    .X(_07105_));
 sg13g2_and3_1 _15723_ (.X(_07106_),
    .A(net268),
    .B(_07104_),
    .C(_07105_));
 sg13g2_nor3_1 _15724_ (.A(net149),
    .B(_07104_),
    .C(_07105_),
    .Y(_07107_));
 sg13g2_o21ai_1 _15725_ (.B1(net253),
    .Y(_07108_),
    .A1(\am_sdr0.cic3.comb2[19] ),
    .A2(net268));
 sg13g2_nor3_1 _15726_ (.A(_07106_),
    .B(_07107_),
    .C(_07108_),
    .Y(_00886_));
 sg13g2_nand2_1 _15727_ (.Y(_07109_),
    .A(\am_sdr0.cic3.comb2[1] ),
    .B(net69));
 sg13g2_xnor2_1 _15728_ (.Y(_07110_),
    .A(_06833_),
    .B(_06960_));
 sg13g2_xnor2_1 _15729_ (.Y(_07111_),
    .A(_06959_),
    .B(_07110_));
 sg13g2_nand2_1 _15730_ (.Y(_07112_),
    .A(net208),
    .B(_07111_));
 sg13g2_buf_2 _15731_ (.A(_02778_),
    .X(_07113_));
 sg13g2_buf_1 _15732_ (.A(_07113_),
    .X(_07114_));
 sg13g2_a21oi_1 _15733_ (.A1(_07109_),
    .A2(_07112_),
    .Y(_00887_),
    .B1(net62));
 sg13g2_buf_1 _15734_ (.A(\am_sdr0.cic3.comb2[2] ),
    .X(_07115_));
 sg13g2_nand2_1 _15735_ (.Y(_07116_),
    .A(_07115_),
    .B(net69));
 sg13g2_a21oi_1 _15736_ (.A1(_06959_),
    .A2(_06961_),
    .Y(_07117_),
    .B1(_06962_));
 sg13g2_xor2_1 _15737_ (.B(_06957_),
    .A(_06838_),
    .X(_07118_));
 sg13g2_xnor2_1 _15738_ (.Y(_07119_),
    .A(_07117_),
    .B(_07118_));
 sg13g2_nand2_1 _15739_ (.Y(_07120_),
    .A(net208),
    .B(_07119_));
 sg13g2_a21oi_1 _15740_ (.A1(_07116_),
    .A2(_07120_),
    .Y(_00888_),
    .B1(net62));
 sg13g2_nand2_1 _15741_ (.Y(_07121_),
    .A(\am_sdr0.cic3.comb2[3] ),
    .B(net69));
 sg13g2_nor2_1 _15742_ (.A(_06958_),
    .B(_06964_),
    .Y(_07122_));
 sg13g2_xnor2_1 _15743_ (.Y(_07123_),
    .A(_06845_),
    .B(\am_sdr0.cic3.comb2_in_del[3] ));
 sg13g2_xnor2_1 _15744_ (.Y(_07124_),
    .A(_07122_),
    .B(_07123_));
 sg13g2_nand2_1 _15745_ (.Y(_07125_),
    .A(net208),
    .B(_07124_));
 sg13g2_a21oi_1 _15746_ (.A1(_07121_),
    .A2(_07125_),
    .Y(_00889_),
    .B1(_07114_));
 sg13g2_buf_1 _15747_ (.A(\am_sdr0.cic3.comb2[4] ),
    .X(_07126_));
 sg13g2_nor2_1 _15748_ (.A(_07126_),
    .B(_06667_),
    .Y(_07127_));
 sg13g2_xor2_1 _15749_ (.B(_06952_),
    .A(_06851_),
    .X(_07128_));
 sg13g2_xnor2_1 _15750_ (.Y(_07129_),
    .A(_06968_),
    .B(_07128_));
 sg13g2_nor2_1 _15751_ (.A(_06737_),
    .B(_07129_),
    .Y(_07130_));
 sg13g2_nor3_1 _15752_ (.A(_01446_),
    .B(_07127_),
    .C(_07130_),
    .Y(_00890_));
 sg13g2_a21oi_2 _15753_ (.B1(_06970_),
    .Y(_07131_),
    .A2(_06968_),
    .A1(_06953_));
 sg13g2_xor2_1 _15754_ (.B(_06950_),
    .A(_06856_),
    .X(_07132_));
 sg13g2_xnor2_1 _15755_ (.Y(_07133_),
    .A(_07131_),
    .B(_07132_));
 sg13g2_nor2_1 _15756_ (.A(net150),
    .B(_07133_),
    .Y(_07134_));
 sg13g2_a21oi_1 _15757_ (.A1(\am_sdr0.cic3.comb2[5] ),
    .A2(_06839_),
    .Y(_07135_),
    .B1(_07134_));
 sg13g2_nor2_1 _15758_ (.A(net67),
    .B(_07135_),
    .Y(_00891_));
 sg13g2_nand2_1 _15759_ (.Y(_07136_),
    .A(\am_sdr0.cic3.comb2[6] ),
    .B(_06839_));
 sg13g2_nand2_1 _15760_ (.Y(_07137_),
    .A(_06950_),
    .B(_07131_));
 sg13g2_nor2_1 _15761_ (.A(_06950_),
    .B(_07131_),
    .Y(_07138_));
 sg13g2_a21oi_1 _15762_ (.A1(_06856_),
    .A2(_07137_),
    .Y(_07139_),
    .B1(_07138_));
 sg13g2_nor2b_1 _15763_ (.A(_06969_),
    .B_N(_06975_),
    .Y(_07140_));
 sg13g2_xnor2_1 _15764_ (.Y(_07141_),
    .A(_07139_),
    .B(_07140_));
 sg13g2_nand2_1 _15765_ (.Y(_07142_),
    .A(net207),
    .B(_07141_));
 sg13g2_a21oi_1 _15766_ (.A1(_07136_),
    .A2(_07142_),
    .Y(_00892_),
    .B1(_07114_));
 sg13g2_buf_1 _15767_ (.A(\am_sdr0.cic3.comb2[7] ),
    .X(_07143_));
 sg13g2_nor2_1 _15768_ (.A(_06973_),
    .B(_06976_),
    .Y(_07144_));
 sg13g2_xnor2_1 _15769_ (.Y(_07145_),
    .A(_06873_),
    .B(_06977_));
 sg13g2_xnor2_1 _15770_ (.Y(_07146_),
    .A(_07144_),
    .B(_07145_));
 sg13g2_nor2_1 _15771_ (.A(net150),
    .B(_07146_),
    .Y(_07147_));
 sg13g2_a21oi_1 _15772_ (.A1(_07143_),
    .A2(net68),
    .Y(_07148_),
    .B1(_07147_));
 sg13g2_nor2_1 _15773_ (.A(_06872_),
    .B(_07148_),
    .Y(_00893_));
 sg13g2_buf_1 _15774_ (.A(\am_sdr0.cic3.comb2[8] ),
    .X(_07149_));
 sg13g2_xnor2_1 _15775_ (.Y(_07150_),
    .A(_06882_),
    .B(_06946_));
 sg13g2_xnor2_1 _15776_ (.Y(_07151_),
    .A(_06981_),
    .B(_07150_));
 sg13g2_nand2_1 _15777_ (.Y(_07152_),
    .A(net269),
    .B(_07151_));
 sg13g2_o21ai_1 _15778_ (.B1(_07152_),
    .Y(_07153_),
    .A1(_07149_),
    .A2(_06728_));
 sg13g2_nor2_1 _15779_ (.A(_06872_),
    .B(_07153_),
    .Y(_00894_));
 sg13g2_inv_1 _15780_ (.Y(_07154_),
    .A(_06981_));
 sg13g2_o21ai_1 _15781_ (.B1(_06989_),
    .Y(_07155_),
    .A1(_06946_),
    .A2(_07154_));
 sg13g2_xor2_1 _15782_ (.B(_06947_),
    .A(_06890_),
    .X(_07156_));
 sg13g2_xnor2_1 _15783_ (.Y(_07157_),
    .A(_07155_),
    .B(_07156_));
 sg13g2_buf_1 _15784_ (.A(\am_sdr0.cic3.comb2[9] ),
    .X(_07158_));
 sg13g2_nor2b_1 _15785_ (.A(net271),
    .B_N(_07158_),
    .Y(_07159_));
 sg13g2_a21oi_1 _15786_ (.A1(_06786_),
    .A2(_07157_),
    .Y(_07160_),
    .B1(_07159_));
 sg13g2_nor2_1 _15787_ (.A(net67),
    .B(_07160_),
    .Y(_00895_));
 sg13g2_buf_1 _15788_ (.A(_06675_),
    .X(_07161_));
 sg13g2_nand2_1 _15789_ (.Y(_07162_),
    .A(_06666_),
    .B(_07161_));
 sg13g2_nand2_1 _15790_ (.Y(_07163_),
    .A(\am_sdr0.cic3.comb2_in_del[0] ),
    .B(net63));
 sg13g2_a21oi_1 _15791_ (.A1(_07162_),
    .A2(_07163_),
    .Y(_00896_),
    .B1(net62));
 sg13g2_nand2_1 _15792_ (.Y(_07164_),
    .A(_06669_),
    .B(net203));
 sg13g2_nand2_1 _15793_ (.Y(_07165_),
    .A(_06992_),
    .B(net63));
 sg13g2_a21oi_1 _15794_ (.A1(_07164_),
    .A2(_07165_),
    .Y(_00897_),
    .B1(net62));
 sg13g2_nand2_1 _15795_ (.Y(_07166_),
    .A(_06727_),
    .B(net203));
 sg13g2_nand2_1 _15796_ (.Y(_07167_),
    .A(_07002_),
    .B(net63));
 sg13g2_a21oi_1 _15797_ (.A1(_07166_),
    .A2(_07167_),
    .Y(_00898_),
    .B1(net62));
 sg13g2_nand2_1 _15798_ (.Y(_07168_),
    .A(\am_sdr0.cic3.comb1[12] ),
    .B(net203));
 sg13g2_nand2_1 _15799_ (.Y(_07169_),
    .A(_07014_),
    .B(net63));
 sg13g2_a21oi_1 _15800_ (.A1(_07168_),
    .A2(_07169_),
    .Y(_00899_),
    .B1(net62));
 sg13g2_nand2_1 _15801_ (.Y(_07170_),
    .A(_06749_),
    .B(net203));
 sg13g2_nand2_1 _15802_ (.Y(_07171_),
    .A(\am_sdr0.cic3.comb2_in_del[13] ),
    .B(_06934_));
 sg13g2_a21oi_1 _15803_ (.A1(_07170_),
    .A2(_07171_),
    .Y(_00900_),
    .B1(net62));
 sg13g2_nand2_1 _15804_ (.Y(_07172_),
    .A(_06758_),
    .B(_07161_));
 sg13g2_nand2_1 _15805_ (.Y(_07173_),
    .A(_07045_),
    .B(_06934_));
 sg13g2_a21oi_1 _15806_ (.A1(_07172_),
    .A2(_07173_),
    .Y(_00901_),
    .B1(net62));
 sg13g2_nand2_1 _15807_ (.Y(_07174_),
    .A(_06791_),
    .B(net203));
 sg13g2_buf_1 _15808_ (.A(net150),
    .X(_07175_));
 sg13g2_nand2_1 _15809_ (.Y(_07176_),
    .A(_07066_),
    .B(net61));
 sg13g2_buf_1 _15810_ (.A(_07113_),
    .X(_07177_));
 sg13g2_a21oi_1 _15811_ (.A1(_07174_),
    .A2(_07176_),
    .Y(_00902_),
    .B1(net60));
 sg13g2_nand2_1 _15812_ (.Y(_07178_),
    .A(_06794_),
    .B(net203));
 sg13g2_nand2_1 _15813_ (.Y(_07179_),
    .A(_07073_),
    .B(net61));
 sg13g2_a21oi_1 _15814_ (.A1(_07178_),
    .A2(_07179_),
    .Y(_00903_),
    .B1(net60));
 sg13g2_nand2_1 _15815_ (.Y(_07180_),
    .A(_06807_),
    .B(net203));
 sg13g2_nand2_1 _15816_ (.Y(_07181_),
    .A(\am_sdr0.cic3.comb2_in_del[17] ),
    .B(net61));
 sg13g2_a21oi_1 _15817_ (.A1(_07180_),
    .A2(_07181_),
    .Y(_00904_),
    .B1(net60));
 sg13g2_nand2_1 _15818_ (.Y(_07182_),
    .A(_06825_),
    .B(net203));
 sg13g2_nand2_1 _15819_ (.Y(_07183_),
    .A(_07097_),
    .B(net61));
 sg13g2_a21oi_1 _15820_ (.A1(_07182_),
    .A2(_07183_),
    .Y(_00905_),
    .B1(net60));
 sg13g2_buf_1 _15821_ (.A(_06675_),
    .X(_07184_));
 sg13g2_nand2_1 _15822_ (.Y(_07185_),
    .A(\am_sdr0.cic3.comb1[19] ),
    .B(_07184_));
 sg13g2_nand2_1 _15823_ (.Y(_07186_),
    .A(\am_sdr0.cic3.comb2_in_del[19] ),
    .B(net61));
 sg13g2_a21oi_1 _15824_ (.A1(_07185_),
    .A2(_07186_),
    .Y(_00906_),
    .B1(net60));
 sg13g2_nand2_1 _15825_ (.Y(_07187_),
    .A(_06833_),
    .B(net202));
 sg13g2_nand2_1 _15826_ (.Y(_07188_),
    .A(_06960_),
    .B(net61));
 sg13g2_a21oi_1 _15827_ (.A1(_07187_),
    .A2(_07188_),
    .Y(_00907_),
    .B1(net60));
 sg13g2_nand2_1 _15828_ (.Y(_07189_),
    .A(_06838_),
    .B(net202));
 sg13g2_nand2_1 _15829_ (.Y(_07190_),
    .A(_06957_),
    .B(net61));
 sg13g2_a21oi_1 _15830_ (.A1(_07189_),
    .A2(_07190_),
    .Y(_00908_),
    .B1(net60));
 sg13g2_nand2_1 _15831_ (.Y(_07191_),
    .A(_06845_),
    .B(net202));
 sg13g2_nand2_1 _15832_ (.Y(_07192_),
    .A(\am_sdr0.cic3.comb2_in_del[3] ),
    .B(net61));
 sg13g2_a21oi_1 _15833_ (.A1(_07191_),
    .A2(_07192_),
    .Y(_00909_),
    .B1(net60));
 sg13g2_nand2_1 _15834_ (.Y(_07193_),
    .A(_06851_),
    .B(net202));
 sg13g2_nand2_1 _15835_ (.Y(_07194_),
    .A(_06952_),
    .B(_07175_));
 sg13g2_a21oi_1 _15836_ (.A1(_07193_),
    .A2(_07194_),
    .Y(_00910_),
    .B1(_07177_));
 sg13g2_nand2_1 _15837_ (.Y(_07195_),
    .A(_06856_),
    .B(net202));
 sg13g2_nand2_1 _15838_ (.Y(_07196_),
    .A(_06950_),
    .B(_07175_));
 sg13g2_a21oi_1 _15839_ (.A1(_07195_),
    .A2(_07196_),
    .Y(_00911_),
    .B1(_07177_));
 sg13g2_nand2_1 _15840_ (.Y(_07197_),
    .A(_06863_),
    .B(net202));
 sg13g2_buf_1 _15841_ (.A(_06671_),
    .X(_07198_));
 sg13g2_nand2_1 _15842_ (.Y(_07199_),
    .A(\am_sdr0.cic3.comb2_in_del[6] ),
    .B(net148));
 sg13g2_buf_1 _15843_ (.A(_07113_),
    .X(_07200_));
 sg13g2_a21oi_1 _15844_ (.A1(_07197_),
    .A2(_07199_),
    .Y(_00912_),
    .B1(net59));
 sg13g2_nand2_1 _15845_ (.Y(_07201_),
    .A(_06873_),
    .B(_07184_));
 sg13g2_nand2_1 _15846_ (.Y(_07202_),
    .A(_06977_),
    .B(net148));
 sg13g2_a21oi_1 _15847_ (.A1(_07201_),
    .A2(_07202_),
    .Y(_00913_),
    .B1(net59));
 sg13g2_nand2_1 _15848_ (.Y(_07203_),
    .A(_06882_),
    .B(net202));
 sg13g2_nand2_1 _15849_ (.Y(_07204_),
    .A(_06946_),
    .B(net148));
 sg13g2_a21oi_1 _15850_ (.A1(_07203_),
    .A2(_07204_),
    .Y(_00914_),
    .B1(net59));
 sg13g2_nand2_1 _15851_ (.Y(_07205_),
    .A(_06890_),
    .B(net202));
 sg13g2_nand2_1 _15852_ (.Y(_07206_),
    .A(_06947_),
    .B(net148));
 sg13g2_a21oi_1 _15853_ (.A1(_07205_),
    .A2(_07206_),
    .Y(_00915_),
    .B1(net59));
 sg13g2_buf_1 _15854_ (.A(\am_sdr0.cic3.comb3_in_del[8] ),
    .X(_07207_));
 sg13g2_inv_1 _15855_ (.Y(_07208_),
    .A(_07149_));
 sg13g2_inv_1 _15856_ (.Y(_07209_),
    .A(\am_sdr0.cic3.comb3_in_del[7] ));
 sg13g2_inv_1 _15857_ (.Y(_07210_),
    .A(\am_sdr0.cic3.comb2[5] ));
 sg13g2_inv_1 _15858_ (.Y(_07211_),
    .A(\am_sdr0.cic3.comb2[3] ));
 sg13g2_nand2b_1 _15859_ (.Y(_07212_),
    .B(_07115_),
    .A_N(\am_sdr0.cic3.comb3_in_del[2] ));
 sg13g2_nand2b_1 _15860_ (.Y(_07213_),
    .B(\am_sdr0.cic3.comb3_in_del[2] ),
    .A_N(_07115_));
 sg13g2_inv_1 _15861_ (.Y(_07214_),
    .A(\am_sdr0.cic3.comb2[1] ));
 sg13g2_nor2b_1 _15862_ (.A(\am_sdr0.cic3.comb2[0] ),
    .B_N(\am_sdr0.cic3.comb3_in_del[0] ),
    .Y(_07215_));
 sg13g2_nand2_1 _15863_ (.Y(_07216_),
    .A(_07214_),
    .B(_07215_));
 sg13g2_o21ai_1 _15864_ (.B1(\am_sdr0.cic3.comb3_in_del[1] ),
    .Y(_07217_),
    .A1(_07214_),
    .A2(_07215_));
 sg13g2_nand3_1 _15865_ (.B(_07216_),
    .C(_07217_),
    .A(_07213_),
    .Y(_07218_));
 sg13g2_a22oi_1 _15866_ (.Y(_07219_),
    .B1(_07212_),
    .B2(_07218_),
    .A2(_07211_),
    .A1(\am_sdr0.cic3.comb3_in_del[3] ));
 sg13g2_nand2b_1 _15867_ (.Y(_07220_),
    .B(_07126_),
    .A_N(\am_sdr0.cic3.comb3_in_del[4] ));
 sg13g2_o21ai_1 _15868_ (.B1(_07220_),
    .Y(_07221_),
    .A1(\am_sdr0.cic3.comb3_in_del[3] ),
    .A2(_07211_));
 sg13g2_nand2b_1 _15869_ (.Y(_07222_),
    .B(\am_sdr0.cic3.comb3_in_del[4] ),
    .A_N(_07126_));
 sg13g2_o21ai_1 _15870_ (.B1(_07222_),
    .Y(_07223_),
    .A1(_07219_),
    .A2(_07221_));
 sg13g2_o21ai_1 _15871_ (.B1(_07223_),
    .Y(_07224_),
    .A1(\am_sdr0.cic3.comb3_in_del[5] ),
    .A2(_07210_));
 sg13g2_inv_1 _15872_ (.Y(_07225_),
    .A(\am_sdr0.cic3.comb2[6] ));
 sg13g2_a22oi_1 _15873_ (.Y(_07226_),
    .B1(\am_sdr0.cic3.comb3_in_del[5] ),
    .B2(_07210_),
    .A2(_07225_),
    .A1(\am_sdr0.cic3.comb3_in_del[6] ));
 sg13g2_nor2_1 _15874_ (.A(\am_sdr0.cic3.comb3_in_del[6] ),
    .B(_07225_),
    .Y(_07227_));
 sg13g2_a21o_1 _15875_ (.A2(_07226_),
    .A1(_07224_),
    .B1(_07227_),
    .X(_07228_));
 sg13g2_o21ai_1 _15876_ (.B1(_07228_),
    .Y(_07229_),
    .A1(_07209_),
    .A2(_07143_));
 sg13g2_inv_1 _15877_ (.Y(_07230_),
    .A(_07207_));
 sg13g2_a22oi_1 _15878_ (.Y(_07231_),
    .B1(_07209_),
    .B2(_07143_),
    .A2(_07149_),
    .A1(_07230_));
 sg13g2_nor2b_1 _15879_ (.A(_06996_),
    .B_N(\am_sdr0.cic3.comb3_in_del[11] ),
    .Y(_07232_));
 sg13g2_nand2b_1 _15880_ (.Y(_07233_),
    .B(_06996_),
    .A_N(\am_sdr0.cic3.comb3_in_del[11] ));
 sg13g2_nand2b_1 _15881_ (.Y(_07234_),
    .B(_07233_),
    .A_N(_07232_));
 sg13g2_xor2_1 _15882_ (.B(_06944_),
    .A(\am_sdr0.cic3.comb3_in_del[10] ),
    .X(_07235_));
 sg13g2_nor2b_1 _15883_ (.A(\am_sdr0.cic3.comb3_in_del[9] ),
    .B_N(_07158_),
    .Y(_07236_));
 sg13g2_nor2b_1 _15884_ (.A(_07158_),
    .B_N(\am_sdr0.cic3.comb3_in_del[9] ),
    .Y(_07237_));
 sg13g2_or3_1 _15885_ (.A(_07235_),
    .B(_07236_),
    .C(_07237_),
    .X(_07238_));
 sg13g2_or2_1 _15886_ (.X(_07239_),
    .B(_07238_),
    .A(_07234_));
 sg13g2_a221oi_1 _15887_ (.B2(_07231_),
    .C1(_07239_),
    .B1(_07229_),
    .A1(_07207_),
    .Y(_07240_),
    .A2(_07208_));
 sg13g2_nand2_1 _15888_ (.Y(_07241_),
    .A(_06944_),
    .B(_07236_));
 sg13g2_nand2_1 _15889_ (.Y(_07242_),
    .A(\am_sdr0.cic3.comb3_in_del[10] ),
    .B(_07241_));
 sg13g2_o21ai_1 _15890_ (.B1(_07242_),
    .Y(_07243_),
    .A1(_06944_),
    .A2(_07236_));
 sg13g2_a21oi_1 _15891_ (.A1(_07233_),
    .A2(_07243_),
    .Y(_07244_),
    .B1(_07232_));
 sg13g2_nor2_1 _15892_ (.A(_07240_),
    .B(_07244_),
    .Y(_07245_));
 sg13g2_buf_1 _15893_ (.A(\am_sdr0.cic3.comb3_in_del[12] ),
    .X(_07246_));
 sg13g2_xor2_1 _15894_ (.B(_07246_),
    .A(_07008_),
    .X(_07247_));
 sg13g2_xnor2_1 _15895_ (.Y(_07248_),
    .A(_07245_),
    .B(_07247_));
 sg13g2_nand2_1 _15896_ (.Y(_07249_),
    .A(net269),
    .B(_07248_));
 sg13g2_o21ai_1 _15897_ (.B1(_07249_),
    .Y(_07250_),
    .A1(net268),
    .A2(\am_sdr0.cic3.comb3[12] ));
 sg13g2_nor2_1 _15898_ (.A(net67),
    .B(_07250_),
    .Y(_00916_));
 sg13g2_or3_1 _15899_ (.A(_07234_),
    .B(_07238_),
    .C(_07247_),
    .X(_07251_));
 sg13g2_a221oi_1 _15900_ (.B2(_07231_),
    .C1(_07251_),
    .B1(_07229_),
    .A1(_07207_),
    .Y(_07252_),
    .A2(_07208_));
 sg13g2_buf_1 _15901_ (.A(_07252_),
    .X(_07253_));
 sg13g2_nor2b_1 _15902_ (.A(_07246_),
    .B_N(_07008_),
    .Y(_07254_));
 sg13g2_nand2b_1 _15903_ (.Y(_07255_),
    .B(_07246_),
    .A_N(_07008_));
 sg13g2_o21ai_1 _15904_ (.B1(_07255_),
    .Y(_07256_),
    .A1(_07244_),
    .A2(_07254_));
 sg13g2_nor2b_1 _15905_ (.A(_07253_),
    .B_N(_07256_),
    .Y(_07257_));
 sg13g2_buf_1 _15906_ (.A(\am_sdr0.cic3.comb3_in_del[13] ),
    .X(_07258_));
 sg13g2_xor2_1 _15907_ (.B(_07258_),
    .A(_07020_),
    .X(_07259_));
 sg13g2_xnor2_1 _15908_ (.Y(_07260_),
    .A(_07257_),
    .B(_07259_));
 sg13g2_nand2_1 _15909_ (.Y(_07261_),
    .A(_06663_),
    .B(_07260_));
 sg13g2_o21ai_1 _15910_ (.B1(_07261_),
    .Y(_07262_),
    .A1(net268),
    .A2(\am_sdr0.cic3.comb3[13] ));
 sg13g2_nor2_1 _15911_ (.A(net67),
    .B(_07262_),
    .Y(_00917_));
 sg13g2_nand2_1 _15912_ (.Y(_07263_),
    .A(_07258_),
    .B(_07256_));
 sg13g2_o21ai_1 _15913_ (.B1(_07020_),
    .Y(_07264_),
    .A1(_07253_),
    .A2(_07263_));
 sg13g2_o21ai_1 _15914_ (.B1(_07264_),
    .Y(_07265_),
    .A1(_07258_),
    .A2(_07257_));
 sg13g2_buf_1 _15915_ (.A(\am_sdr0.cic3.comb3_in_del[14] ),
    .X(_07266_));
 sg13g2_xor2_1 _15916_ (.B(_07266_),
    .A(_07033_),
    .X(_07267_));
 sg13g2_xnor2_1 _15917_ (.Y(_07268_),
    .A(_07265_),
    .B(_07267_));
 sg13g2_nor2b_1 _15918_ (.A(net271),
    .B_N(\am_sdr0.cic3.comb3[14] ),
    .Y(_07269_));
 sg13g2_a21oi_1 _15919_ (.A1(_06786_),
    .A2(_07268_),
    .Y(_07270_),
    .B1(_07269_));
 sg13g2_nor2_1 _15920_ (.A(net67),
    .B(_07270_),
    .Y(_00918_));
 sg13g2_buf_1 _15921_ (.A(_06365_),
    .X(_07271_));
 sg13g2_inv_1 _15922_ (.Y(_07272_),
    .A(_07020_));
 sg13g2_nand2_1 _15923_ (.Y(_07273_),
    .A(_07272_),
    .B(_07256_));
 sg13g2_a21o_1 _15924_ (.A2(_07273_),
    .A1(_07263_),
    .B1(_07253_),
    .X(_07274_));
 sg13g2_inv_1 _15925_ (.Y(_07275_),
    .A(_07033_));
 sg13g2_a22oi_1 _15926_ (.Y(_07276_),
    .B1(_07275_),
    .B2(_07266_),
    .A2(_07258_),
    .A1(_07272_));
 sg13g2_nor2_1 _15927_ (.A(_07275_),
    .B(_07266_),
    .Y(_07277_));
 sg13g2_a21oi_2 _15928_ (.B1(_07277_),
    .Y(_07278_),
    .A2(_07276_),
    .A1(_07274_));
 sg13g2_buf_1 _15929_ (.A(\am_sdr0.cic3.comb3_in_del[15] ),
    .X(_07279_));
 sg13g2_xnor2_1 _15930_ (.Y(_07280_),
    .A(_07049_),
    .B(_07279_));
 sg13g2_xnor2_1 _15931_ (.Y(_07281_),
    .A(_07278_),
    .B(_07280_));
 sg13g2_nor2b_1 _15932_ (.A(net271),
    .B_N(\am_sdr0.cic3.comb3[15] ),
    .Y(_07282_));
 sg13g2_a21oi_1 _15933_ (.A1(net206),
    .A2(_07281_),
    .Y(_07283_),
    .B1(_07282_));
 sg13g2_nor2_1 _15934_ (.A(_07271_),
    .B(_07283_),
    .Y(_00919_));
 sg13g2_nor2_1 _15935_ (.A(_07279_),
    .B(_07278_),
    .Y(_07284_));
 sg13g2_nand2_1 _15936_ (.Y(_07285_),
    .A(_07279_),
    .B(_07278_));
 sg13g2_o21ai_1 _15937_ (.B1(_07285_),
    .Y(_07286_),
    .A1(_07049_),
    .A2(_07284_));
 sg13g2_nor2b_1 _15938_ (.A(\am_sdr0.cic3.comb3_in_del[16] ),
    .B_N(_07076_),
    .Y(_07287_));
 sg13g2_nand2b_1 _15939_ (.Y(_07288_),
    .B(\am_sdr0.cic3.comb3_in_del[16] ),
    .A_N(_07076_));
 sg13g2_nor2b_1 _15940_ (.A(_07287_),
    .B_N(_07288_),
    .Y(_07289_));
 sg13g2_xnor2_1 _15941_ (.Y(_07290_),
    .A(_07286_),
    .B(_07289_));
 sg13g2_nor2b_1 _15942_ (.A(net271),
    .B_N(\am_sdr0.cic3.comb3[16] ),
    .Y(_07291_));
 sg13g2_a21oi_1 _15943_ (.A1(net206),
    .A2(_07290_),
    .Y(_07292_),
    .B1(_07291_));
 sg13g2_nor2_1 _15944_ (.A(_07271_),
    .B(_07292_),
    .Y(_00920_));
 sg13g2_nor2_1 _15945_ (.A(_07277_),
    .B(_07287_),
    .Y(_07293_));
 sg13g2_nand2_1 _15946_ (.Y(_07294_),
    .A(_07279_),
    .B(_07293_));
 sg13g2_nand2b_1 _15947_ (.Y(_07295_),
    .B(_07293_),
    .A_N(_07049_));
 sg13g2_a22oi_1 _15948_ (.Y(_07296_),
    .B1(_07294_),
    .B2(_07295_),
    .A2(_07276_),
    .A1(_07274_));
 sg13g2_nand2b_1 _15949_ (.Y(_07297_),
    .B(_07279_),
    .A_N(_07049_));
 sg13g2_o21ai_1 _15950_ (.B1(_07288_),
    .Y(_07298_),
    .A1(_07297_),
    .A2(_07287_));
 sg13g2_nor2_1 _15951_ (.A(_07296_),
    .B(_07298_),
    .Y(_07299_));
 sg13g2_buf_1 _15952_ (.A(\am_sdr0.cic3.comb3_in_del[17] ),
    .X(_07300_));
 sg13g2_xnor2_1 _15953_ (.Y(_07301_),
    .A(_07078_),
    .B(_07300_));
 sg13g2_xnor2_1 _15954_ (.Y(_07302_),
    .A(_07299_),
    .B(_07301_));
 sg13g2_o21ai_1 _15955_ (.B1(_05549_),
    .Y(_07303_),
    .A1(net268),
    .A2(\am_sdr0.cic3.comb3[17] ));
 sg13g2_a21oi_1 _15956_ (.A1(net209),
    .A2(_07302_),
    .Y(_00921_),
    .B1(_07303_));
 sg13g2_nor3_1 _15957_ (.A(_07300_),
    .B(_07296_),
    .C(_07298_),
    .Y(_07304_));
 sg13g2_o21ai_1 _15958_ (.B1(_07300_),
    .Y(_07305_),
    .A1(_07296_),
    .A2(_07298_));
 sg13g2_o21ai_1 _15959_ (.B1(_07305_),
    .Y(_07306_),
    .A1(_07078_),
    .A2(_07304_));
 sg13g2_nor2b_1 _15960_ (.A(_07095_),
    .B_N(\am_sdr0.cic3.comb3_in_del[18] ),
    .Y(_07307_));
 sg13g2_nand2b_1 _15961_ (.Y(_07308_),
    .B(_07095_),
    .A_N(\am_sdr0.cic3.comb3_in_del[18] ));
 sg13g2_nand2b_1 _15962_ (.Y(_07309_),
    .B(_07308_),
    .A_N(_07307_));
 sg13g2_xnor2_1 _15963_ (.Y(_07310_),
    .A(_07306_),
    .B(_07309_));
 sg13g2_nor2_1 _15964_ (.A(net271),
    .B(\am_sdr0.cic3.comb3[18] ),
    .Y(_07311_));
 sg13g2_a21oi_1 _15965_ (.A1(net268),
    .A2(_07310_),
    .Y(_07312_),
    .B1(_07311_));
 sg13g2_and2_1 _15966_ (.A(net210),
    .B(_07312_),
    .X(_00922_));
 sg13g2_a21oi_1 _15967_ (.A1(_07306_),
    .A2(_07308_),
    .Y(_07313_),
    .B1(_07307_));
 sg13g2_xnor2_1 _15968_ (.Y(_07314_),
    .A(\am_sdr0.cic3.comb2[19] ),
    .B(\am_sdr0.cic3.comb3_in_del[19] ));
 sg13g2_xnor2_1 _15969_ (.Y(_07315_),
    .A(_07313_),
    .B(_07314_));
 sg13g2_o21ai_1 _15970_ (.B1(net254),
    .Y(_07316_),
    .A1(net268),
    .A2(\am_sdr0.cic3.comb3[19] ));
 sg13g2_a21oi_1 _15971_ (.A1(net209),
    .A2(_07315_),
    .Y(_00923_),
    .B1(_07316_));
 sg13g2_buf_1 _15972_ (.A(_06675_),
    .X(_07317_));
 sg13g2_nand2_1 _15973_ (.Y(_07318_),
    .A(\am_sdr0.cic3.comb2[0] ),
    .B(net201));
 sg13g2_nand2_1 _15974_ (.Y(_07319_),
    .A(\am_sdr0.cic3.comb3_in_del[0] ),
    .B(_07198_));
 sg13g2_a21oi_1 _15975_ (.A1(_07318_),
    .A2(_07319_),
    .Y(_00924_),
    .B1(_07200_));
 sg13g2_nand2_1 _15976_ (.Y(_07320_),
    .A(_06944_),
    .B(net201));
 sg13g2_nand2_1 _15977_ (.Y(_07321_),
    .A(\am_sdr0.cic3.comb3_in_del[10] ),
    .B(net148));
 sg13g2_a21oi_1 _15978_ (.A1(_07320_),
    .A2(_07321_),
    .Y(_00925_),
    .B1(net59));
 sg13g2_nand2_1 _15979_ (.Y(_07322_),
    .A(_06996_),
    .B(net201));
 sg13g2_nand2_1 _15980_ (.Y(_07323_),
    .A(\am_sdr0.cic3.comb3_in_del[11] ),
    .B(net148));
 sg13g2_a21oi_1 _15981_ (.A1(_07322_),
    .A2(_07323_),
    .Y(_00926_),
    .B1(net59));
 sg13g2_nand2_1 _15982_ (.Y(_07324_),
    .A(_07008_),
    .B(_07317_));
 sg13g2_nand2_1 _15983_ (.Y(_07325_),
    .A(_07246_),
    .B(net148));
 sg13g2_a21oi_1 _15984_ (.A1(_07324_),
    .A2(_07325_),
    .Y(_00927_),
    .B1(net59));
 sg13g2_nand2_1 _15985_ (.Y(_07326_),
    .A(_07020_),
    .B(net201));
 sg13g2_nand2_1 _15986_ (.Y(_07327_),
    .A(_07258_),
    .B(net148));
 sg13g2_a21oi_1 _15987_ (.A1(_07326_),
    .A2(_07327_),
    .Y(_00928_),
    .B1(net59));
 sg13g2_nand2_1 _15988_ (.Y(_07328_),
    .A(_07033_),
    .B(_07317_));
 sg13g2_nand2_1 _15989_ (.Y(_07329_),
    .A(_07266_),
    .B(_07198_));
 sg13g2_a21oi_1 _15990_ (.A1(_07328_),
    .A2(_07329_),
    .Y(_00929_),
    .B1(_07200_));
 sg13g2_nand2_1 _15991_ (.Y(_07330_),
    .A(_07049_),
    .B(net201));
 sg13g2_buf_1 _15992_ (.A(_06671_),
    .X(_07331_));
 sg13g2_nand2_1 _15993_ (.Y(_07332_),
    .A(_07279_),
    .B(net147));
 sg13g2_buf_1 _15994_ (.A(_07113_),
    .X(_07333_));
 sg13g2_a21oi_1 _15995_ (.A1(_07330_),
    .A2(_07332_),
    .Y(_00930_),
    .B1(net57));
 sg13g2_nand2_1 _15996_ (.Y(_07334_),
    .A(_07076_),
    .B(net201));
 sg13g2_nand2_1 _15997_ (.Y(_07335_),
    .A(\am_sdr0.cic3.comb3_in_del[16] ),
    .B(net147));
 sg13g2_a21oi_1 _15998_ (.A1(_07334_),
    .A2(_07335_),
    .Y(_00931_),
    .B1(net57));
 sg13g2_nand2_1 _15999_ (.Y(_07336_),
    .A(_07078_),
    .B(net201));
 sg13g2_nand2_1 _16000_ (.Y(_07337_),
    .A(_07300_),
    .B(net147));
 sg13g2_a21oi_1 _16001_ (.A1(_07336_),
    .A2(_07337_),
    .Y(_00932_),
    .B1(net57));
 sg13g2_nand2_1 _16002_ (.Y(_07338_),
    .A(_07095_),
    .B(net201));
 sg13g2_nand2_1 _16003_ (.Y(_07339_),
    .A(\am_sdr0.cic3.comb3_in_del[18] ),
    .B(net147));
 sg13g2_a21oi_1 _16004_ (.A1(_07338_),
    .A2(_07339_),
    .Y(_00933_),
    .B1(net57));
 sg13g2_buf_1 _16005_ (.A(_06675_),
    .X(_07340_));
 sg13g2_nand2_1 _16006_ (.Y(_07341_),
    .A(\am_sdr0.cic3.comb2[19] ),
    .B(_07340_));
 sg13g2_nand2_1 _16007_ (.Y(_07342_),
    .A(\am_sdr0.cic3.comb3_in_del[19] ),
    .B(net147));
 sg13g2_a21oi_1 _16008_ (.A1(_07341_),
    .A2(_07342_),
    .Y(_00934_),
    .B1(net57));
 sg13g2_nand2_1 _16009_ (.Y(_07343_),
    .A(\am_sdr0.cic3.comb2[1] ),
    .B(net200));
 sg13g2_nand2_1 _16010_ (.Y(_07344_),
    .A(\am_sdr0.cic3.comb3_in_del[1] ),
    .B(net147));
 sg13g2_a21oi_1 _16011_ (.A1(_07343_),
    .A2(_07344_),
    .Y(_00935_),
    .B1(net57));
 sg13g2_nand2_1 _16012_ (.Y(_07345_),
    .A(_07115_),
    .B(net200));
 sg13g2_nand2_1 _16013_ (.Y(_07346_),
    .A(\am_sdr0.cic3.comb3_in_del[2] ),
    .B(net147));
 sg13g2_a21oi_1 _16014_ (.A1(_07345_),
    .A2(_07346_),
    .Y(_00936_),
    .B1(net57));
 sg13g2_nand2_1 _16015_ (.Y(_07347_),
    .A(\am_sdr0.cic3.comb2[3] ),
    .B(net200));
 sg13g2_nand2_1 _16016_ (.Y(_07348_),
    .A(\am_sdr0.cic3.comb3_in_del[3] ),
    .B(net147));
 sg13g2_a21oi_1 _16017_ (.A1(_07347_),
    .A2(_07348_),
    .Y(_00937_),
    .B1(net57));
 sg13g2_nand2_1 _16018_ (.Y(_07349_),
    .A(_07126_),
    .B(net200));
 sg13g2_nand2_1 _16019_ (.Y(_07350_),
    .A(\am_sdr0.cic3.comb3_in_del[4] ),
    .B(_07331_));
 sg13g2_a21oi_1 _16020_ (.A1(_07349_),
    .A2(_07350_),
    .Y(_00938_),
    .B1(_07333_));
 sg13g2_nand2_1 _16021_ (.Y(_07351_),
    .A(\am_sdr0.cic3.comb2[5] ),
    .B(_07340_));
 sg13g2_nand2_1 _16022_ (.Y(_07352_),
    .A(\am_sdr0.cic3.comb3_in_del[5] ),
    .B(_07331_));
 sg13g2_a21oi_1 _16023_ (.A1(_07351_),
    .A2(_07352_),
    .Y(_00939_),
    .B1(_07333_));
 sg13g2_nand2_1 _16024_ (.Y(_07353_),
    .A(\am_sdr0.cic3.comb2[6] ),
    .B(net200));
 sg13g2_buf_1 _16025_ (.A(_06671_),
    .X(_07354_));
 sg13g2_nand2_1 _16026_ (.Y(_07355_),
    .A(\am_sdr0.cic3.comb3_in_del[6] ),
    .B(net146));
 sg13g2_buf_1 _16027_ (.A(_07113_),
    .X(_07356_));
 sg13g2_a21oi_1 _16028_ (.A1(_07353_),
    .A2(_07355_),
    .Y(_00940_),
    .B1(net56));
 sg13g2_nand2_1 _16029_ (.Y(_07357_),
    .A(_07143_),
    .B(net200));
 sg13g2_nand2_1 _16030_ (.Y(_07358_),
    .A(\am_sdr0.cic3.comb3_in_del[7] ),
    .B(net146));
 sg13g2_a21oi_1 _16031_ (.A1(_07357_),
    .A2(_07358_),
    .Y(_00941_),
    .B1(net56));
 sg13g2_nand2_1 _16032_ (.Y(_07359_),
    .A(_07149_),
    .B(net200));
 sg13g2_nand2_1 _16033_ (.Y(_07360_),
    .A(_07207_),
    .B(_07354_));
 sg13g2_a21oi_1 _16034_ (.A1(_07359_),
    .A2(_07360_),
    .Y(_00942_),
    .B1(_07356_));
 sg13g2_nand2_1 _16035_ (.Y(_07361_),
    .A(_07158_),
    .B(net200));
 sg13g2_nand2_1 _16036_ (.Y(_07362_),
    .A(\am_sdr0.cic3.comb3_in_del[9] ),
    .B(_07354_));
 sg13g2_a21oi_1 _16037_ (.A1(_07361_),
    .A2(_07362_),
    .Y(_00943_),
    .B1(_07356_));
 sg13g2_buf_1 _16038_ (.A(_02425_),
    .X(_07363_));
 sg13g2_buf_1 _16039_ (.A(net267),
    .X(_07364_));
 sg13g2_xnor2_1 _16040_ (.Y(_07365_),
    .A(\am_sdr0.cic3.count[0] ),
    .B(_07364_));
 sg13g2_nor2_1 _16041_ (.A(net58),
    .B(_07365_),
    .Y(_00944_));
 sg13g2_buf_1 _16042_ (.A(net267),
    .X(_07366_));
 sg13g2_nand2_1 _16043_ (.Y(_07367_),
    .A(\am_sdr0.cic3.count[0] ),
    .B(net198));
 sg13g2_xor2_1 _16044_ (.B(_07367_),
    .A(\am_sdr0.cic3.count[1] ),
    .X(_07368_));
 sg13g2_nor2_1 _16045_ (.A(net58),
    .B(_07368_),
    .Y(_00945_));
 sg13g2_xnor2_1 _16046_ (.Y(_07369_),
    .A(_02424_),
    .B(_02426_));
 sg13g2_nor2_1 _16047_ (.A(net58),
    .B(_07369_),
    .Y(_00946_));
 sg13g2_xnor2_1 _16048_ (.Y(_07370_),
    .A(_02423_),
    .B(_02427_));
 sg13g2_nor2_1 _16049_ (.A(net58),
    .B(_07370_),
    .Y(_00947_));
 sg13g2_nand2_1 _16050_ (.Y(_07371_),
    .A(_02423_),
    .B(_02427_));
 sg13g2_xor2_1 _16051_ (.B(_07371_),
    .A(\am_sdr0.cic3.count[4] ),
    .X(_07372_));
 sg13g2_nor2_1 _16052_ (.A(net58),
    .B(_07372_),
    .Y(_00948_));
 sg13g2_nand3_1 _16053_ (.B(\am_sdr0.cic3.count[4] ),
    .C(_02427_),
    .A(_02423_),
    .Y(_07373_));
 sg13g2_xor2_1 _16054_ (.B(_07373_),
    .A(\am_sdr0.cic3.count[5] ),
    .X(_07374_));
 sg13g2_nor2_1 _16055_ (.A(net58),
    .B(_07374_),
    .Y(_00949_));
 sg13g2_inv_1 _16056_ (.Y(_07375_),
    .A(\am_sdr0.cic3.count[7] ));
 sg13g2_nor3_1 _16057_ (.A(_07375_),
    .B(_02422_),
    .C(_02429_),
    .Y(_07376_));
 sg13g2_a21oi_1 _16058_ (.A1(_02422_),
    .A2(_02429_),
    .Y(_07377_),
    .B1(_07376_));
 sg13g2_nor2_1 _16059_ (.A(net58),
    .B(_07377_),
    .Y(_00950_));
 sg13g2_inv_1 _16060_ (.Y(_07378_),
    .A(_02422_));
 sg13g2_nor2_1 _16061_ (.A(_07378_),
    .B(_02429_),
    .Y(_07379_));
 sg13g2_xnor2_1 _16062_ (.Y(_07380_),
    .A(\am_sdr0.cic3.count[7] ),
    .B(_07379_));
 sg13g2_nor2_1 _16063_ (.A(net58),
    .B(_07380_),
    .Y(_00951_));
 sg13g2_buf_1 _16064_ (.A(_06365_),
    .X(_07381_));
 sg13g2_buf_1 _16065_ (.A(net267),
    .X(_07382_));
 sg13g2_nand2_1 _16066_ (.Y(_07383_),
    .A(net197),
    .B(_05267_));
 sg13g2_xor2_1 _16067_ (.B(_07383_),
    .A(\am_sdr0.cic3.integ1[0] ),
    .X(_07384_));
 sg13g2_nor2_1 _16068_ (.A(net55),
    .B(_07384_),
    .Y(_00952_));
 sg13g2_buf_1 _16069_ (.A(\am_sdr0.cic3.integ1[10] ),
    .X(_07385_));
 sg13g2_inv_1 _16070_ (.Y(_07386_),
    .A(_05262_));
 sg13g2_buf_1 _16071_ (.A(_07386_),
    .X(_07387_));
 sg13g2_buf_2 _16072_ (.A(\am_sdr0.cic3.integ1[6] ),
    .X(_07388_));
 sg13g2_inv_1 _16073_ (.Y(_07389_),
    .A(\am_sdr0.cic3.integ1[5] ));
 sg13g2_buf_2 _16074_ (.A(\am_sdr0.cic3.integ1[4] ),
    .X(_07390_));
 sg13g2_inv_1 _16075_ (.Y(_07391_),
    .A(\am_sdr0.cic1.x_out[11] ));
 sg13g2_nor2_1 _16076_ (.A(_05270_),
    .B(\am_sdr0.cic3.integ1[1] ),
    .Y(_07392_));
 sg13g2_a22oi_1 _16077_ (.Y(_07393_),
    .B1(_05270_),
    .B2(\am_sdr0.cic3.integ1[1] ),
    .A2(\am_sdr0.cic3.integ1[0] ),
    .A1(_05267_));
 sg13g2_nand2_1 _16078_ (.Y(_07394_),
    .A(_05250_),
    .B(\am_sdr0.cic3.integ1[2] ));
 sg13g2_o21ai_1 _16079_ (.B1(_07394_),
    .Y(_07395_),
    .A1(_07392_),
    .A2(_07393_));
 sg13g2_or2_1 _16080_ (.X(_07396_),
    .B(\am_sdr0.cic3.integ1[2] ),
    .A(_05250_));
 sg13g2_buf_1 _16081_ (.A(_07396_),
    .X(_07397_));
 sg13g2_buf_2 _16082_ (.A(\am_sdr0.cic3.integ1[3] ),
    .X(_07398_));
 sg13g2_a21oi_1 _16083_ (.A1(_07395_),
    .A2(_07397_),
    .Y(_07399_),
    .B1(_07398_));
 sg13g2_nand3_1 _16084_ (.B(_07395_),
    .C(_07397_),
    .A(_07398_),
    .Y(_07400_));
 sg13g2_o21ai_1 _16085_ (.B1(_07400_),
    .Y(_07401_),
    .A1(_07391_),
    .A2(_07399_));
 sg13g2_buf_1 _16086_ (.A(_07401_),
    .X(_07402_));
 sg13g2_nand2_1 _16087_ (.Y(_07403_),
    .A(_07390_),
    .B(_07402_));
 sg13g2_o21ai_1 _16088_ (.B1(\am_sdr0.cic1.x_out[12] ),
    .Y(_07404_),
    .A1(_07390_),
    .A2(_07402_));
 sg13g2_nand3_1 _16089_ (.B(_07403_),
    .C(_07404_),
    .A(_07389_),
    .Y(_07405_));
 sg13g2_a21oi_1 _16090_ (.A1(_07403_),
    .A2(_07404_),
    .Y(_07406_),
    .B1(_07389_));
 sg13g2_a21o_1 _16091_ (.A2(_07405_),
    .A1(\am_sdr0.cic1.x_out[13] ),
    .B1(_07406_),
    .X(_07407_));
 sg13g2_buf_1 _16092_ (.A(_07407_),
    .X(_07408_));
 sg13g2_nor2_1 _16093_ (.A(_07388_),
    .B(_07408_),
    .Y(_07409_));
 sg13g2_a21oi_1 _16094_ (.A1(_07388_),
    .A2(_07408_),
    .Y(_07410_),
    .B1(\am_sdr0.cic1.x_out[14] ));
 sg13g2_nor2_1 _16095_ (.A(_07409_),
    .B(_07410_),
    .Y(_07411_));
 sg13g2_buf_2 _16096_ (.A(_07411_),
    .X(_07412_));
 sg13g2_buf_2 _16097_ (.A(\am_sdr0.cic3.integ1[8] ),
    .X(_07413_));
 sg13g2_inv_1 _16098_ (.Y(_07414_),
    .A(_07413_));
 sg13g2_buf_2 _16099_ (.A(\am_sdr0.cic3.integ1[9] ),
    .X(_07415_));
 sg13g2_inv_1 _16100_ (.Y(_07416_),
    .A(_07415_));
 sg13g2_nand2_1 _16101_ (.Y(_07417_),
    .A(_07414_),
    .B(_07416_));
 sg13g2_o21ai_1 _16102_ (.B1(net286),
    .Y(_07418_),
    .A1(_07412_),
    .A2(_07417_));
 sg13g2_nor4_1 _16103_ (.A(_07414_),
    .B(_07416_),
    .C(_07409_),
    .D(_07410_),
    .Y(_07419_));
 sg13g2_buf_1 _16104_ (.A(\am_sdr0.cic3.integ1[7] ),
    .X(_07420_));
 sg13g2_buf_1 _16105_ (.A(_07420_),
    .X(_07421_));
 sg13g2_o21ai_1 _16106_ (.B1(net266),
    .Y(_07422_),
    .A1(_05262_),
    .A2(_07419_));
 sg13g2_nand2_2 _16107_ (.Y(_07423_),
    .A(_07418_),
    .B(_07422_));
 sg13g2_xnor2_1 _16108_ (.Y(_07424_),
    .A(net196),
    .B(_07423_));
 sg13g2_nand2_1 _16109_ (.Y(_07425_),
    .A(net197),
    .B(_07424_));
 sg13g2_xor2_1 _16110_ (.B(_07425_),
    .A(net325),
    .X(_07426_));
 sg13g2_nor2_1 _16111_ (.A(net55),
    .B(_07426_),
    .Y(_00953_));
 sg13g2_nand2b_1 _16112_ (.Y(_07427_),
    .B(net226),
    .A_N(net325));
 sg13g2_nand4_1 _16113_ (.B(net266),
    .C(net325),
    .A(_07386_),
    .Y(_07428_),
    .D(_07419_));
 sg13g2_buf_2 _16114_ (.A(_07428_),
    .X(_07429_));
 sg13g2_o21ai_1 _16115_ (.B1(_07429_),
    .Y(_07430_),
    .A1(_07423_),
    .A2(_07427_));
 sg13g2_buf_1 _16116_ (.A(\am_sdr0.cic3.integ1[11] ),
    .X(_07431_));
 sg13g2_inv_1 _16117_ (.Y(_07432_),
    .A(net324));
 sg13g2_a21o_1 _16118_ (.A2(_07430_),
    .A1(net199),
    .B1(_07432_),
    .X(_07433_));
 sg13g2_nand3_1 _16119_ (.B(_07432_),
    .C(_07430_),
    .A(net199),
    .Y(_07434_));
 sg13g2_a21oi_1 _16120_ (.A1(_07433_),
    .A2(_07434_),
    .Y(_00954_),
    .B1(net56));
 sg13g2_buf_2 _16121_ (.A(\am_sdr0.cic3.integ1[12] ),
    .X(_07435_));
 sg13g2_inv_2 _16122_ (.Y(_07436_),
    .A(_07435_));
 sg13g2_or2_1 _16123_ (.X(_07437_),
    .B(net324),
    .A(net325));
 sg13g2_nor4_1 _16124_ (.A(net266),
    .B(_07415_),
    .C(_07412_),
    .D(_07437_),
    .Y(_07438_));
 sg13g2_nand4_1 _16125_ (.B(_07415_),
    .C(net325),
    .A(_07420_),
    .Y(_07439_),
    .D(net324));
 sg13g2_nor3_1 _16126_ (.A(_07409_),
    .B(_07410_),
    .C(_07439_),
    .Y(_07440_));
 sg13g2_o21ai_1 _16127_ (.B1(_07413_),
    .Y(_07441_),
    .A1(net286),
    .A2(_07440_));
 sg13g2_o21ai_1 _16128_ (.B1(_07441_),
    .Y(_07442_),
    .A1(_07386_),
    .A2(_07438_));
 sg13g2_buf_1 _16129_ (.A(_07442_),
    .X(_07443_));
 sg13g2_xnor2_1 _16130_ (.Y(_07444_),
    .A(net196),
    .B(_07443_));
 sg13g2_nand2_1 _16131_ (.Y(_07445_),
    .A(net199),
    .B(_07444_));
 sg13g2_xnor2_1 _16132_ (.Y(_07446_),
    .A(_07436_),
    .B(_07445_));
 sg13g2_nor2_1 _16133_ (.A(net55),
    .B(_07446_),
    .Y(_00955_));
 sg13g2_buf_1 _16134_ (.A(\am_sdr0.cic3.integ1[13] ),
    .X(_07447_));
 sg13g2_inv_1 _16135_ (.Y(_07448_),
    .A(_02425_));
 sg13g2_buf_2 _16136_ (.A(_07448_),
    .X(_07449_));
 sg13g2_buf_1 _16137_ (.A(_07449_),
    .X(_07450_));
 sg13g2_nand2b_1 _16138_ (.Y(_07451_),
    .B(_07436_),
    .A_N(_07437_));
 sg13g2_nor4_2 _16139_ (.A(net266),
    .B(_07412_),
    .C(_07417_),
    .Y(_07452_),
    .D(_07451_));
 sg13g2_nor3_2 _16140_ (.A(_07432_),
    .B(_07436_),
    .C(_07429_),
    .Y(_07453_));
 sg13g2_a21oi_1 _16141_ (.A1(net226),
    .A2(_07452_),
    .Y(_07454_),
    .B1(_07453_));
 sg13g2_nor2_1 _16142_ (.A(net145),
    .B(_07454_),
    .Y(_07455_));
 sg13g2_xnor2_1 _16143_ (.Y(_07456_),
    .A(net323),
    .B(_07455_));
 sg13g2_nor2_1 _16144_ (.A(net55),
    .B(_07456_),
    .Y(_00956_));
 sg13g2_buf_1 _16145_ (.A(\am_sdr0.cic3.integ1[14] ),
    .X(_07457_));
 sg13g2_nor4_1 _16146_ (.A(net196),
    .B(net323),
    .C(_07423_),
    .D(_07451_),
    .Y(_07458_));
 sg13g2_a21oi_1 _16147_ (.A1(net323),
    .A2(_07453_),
    .Y(_07459_),
    .B1(_07458_));
 sg13g2_nor2_1 _16148_ (.A(net145),
    .B(_07459_),
    .Y(_07460_));
 sg13g2_xnor2_1 _16149_ (.Y(_07461_),
    .A(net322),
    .B(_07460_));
 sg13g2_nor2_1 _16150_ (.A(net55),
    .B(_07461_),
    .Y(_00957_));
 sg13g2_buf_1 _16151_ (.A(\am_sdr0.cic3.integ1[15] ),
    .X(_07462_));
 sg13g2_nor2_1 _16152_ (.A(net323),
    .B(net322),
    .Y(_07463_));
 sg13g2_nor2_1 _16153_ (.A(net286),
    .B(net324),
    .Y(_07464_));
 sg13g2_a21oi_1 _16154_ (.A1(_07452_),
    .A2(_07463_),
    .Y(_07465_),
    .B1(_07464_));
 sg13g2_inv_1 _16155_ (.Y(_07466_),
    .A(net322));
 sg13g2_nand2_1 _16156_ (.Y(_07467_),
    .A(_07435_),
    .B(net323));
 sg13g2_or4_1 _16157_ (.A(_07466_),
    .B(_07429_),
    .C(_07467_),
    .D(_07464_),
    .X(_07468_));
 sg13g2_o21ai_1 _16158_ (.B1(_07468_),
    .Y(_07469_),
    .A1(net196),
    .A2(_07465_));
 sg13g2_nand2_1 _16159_ (.Y(_07470_),
    .A(net197),
    .B(_07469_));
 sg13g2_xor2_1 _16160_ (.B(_07470_),
    .A(net321),
    .X(_07471_));
 sg13g2_nor2_1 _16161_ (.A(net55),
    .B(_07471_),
    .Y(_00958_));
 sg13g2_buf_1 _16162_ (.A(\am_sdr0.cic3.integ1[16] ),
    .X(_07472_));
 sg13g2_inv_1 _16163_ (.Y(_07473_),
    .A(net320));
 sg13g2_nand2b_1 _16164_ (.Y(_07474_),
    .B(net286),
    .A_N(net321));
 sg13g2_nor4_1 _16165_ (.A(_07435_),
    .B(net323),
    .C(net322),
    .D(_07474_),
    .Y(_07475_));
 sg13g2_nand2_1 _16166_ (.Y(_07476_),
    .A(net322),
    .B(net321));
 sg13g2_nor3_1 _16167_ (.A(net226),
    .B(_07467_),
    .C(_07476_),
    .Y(_07477_));
 sg13g2_mux2_1 _16168_ (.A0(_07475_),
    .A1(_07477_),
    .S(_07443_),
    .X(_07478_));
 sg13g2_nand2_1 _16169_ (.Y(_07479_),
    .A(net199),
    .B(_07478_));
 sg13g2_xnor2_1 _16170_ (.Y(_07480_),
    .A(_07473_),
    .B(_07479_));
 sg13g2_nor2_1 _16171_ (.A(net55),
    .B(_07480_),
    .Y(_00959_));
 sg13g2_buf_1 _16172_ (.A(\am_sdr0.cic3.integ1[17] ),
    .X(_07481_));
 sg13g2_nor4_2 _16173_ (.A(net323),
    .B(net322),
    .C(net321),
    .Y(_07482_),
    .D(net320));
 sg13g2_nand2_1 _16174_ (.Y(_07483_),
    .A(_05264_),
    .B(_07482_));
 sg13g2_nor2_1 _16175_ (.A(net196),
    .B(_07452_),
    .Y(_07484_));
 sg13g2_inv_1 _16176_ (.Y(_07485_),
    .A(_07447_));
 sg13g2_nor3_1 _16177_ (.A(_05262_),
    .B(_07485_),
    .C(_07476_),
    .Y(_07486_));
 sg13g2_a22oi_1 _16178_ (.Y(_07487_),
    .B1(_07486_),
    .B2(net320),
    .A2(_07482_),
    .A1(net286));
 sg13g2_inv_1 _16179_ (.Y(_07488_),
    .A(_07487_));
 sg13g2_o21ai_1 _16180_ (.B1(_07488_),
    .Y(_07489_),
    .A1(_07453_),
    .A2(_07484_));
 sg13g2_buf_1 _16181_ (.A(_07489_),
    .X(_07490_));
 sg13g2_mux2_1 _16182_ (.A0(net226),
    .A1(_07483_),
    .S(_07490_),
    .X(_07491_));
 sg13g2_nor2_1 _16183_ (.A(_07450_),
    .B(_07491_),
    .Y(_07492_));
 sg13g2_xnor2_1 _16184_ (.Y(_07493_),
    .A(net319),
    .B(_07492_));
 sg13g2_nor2_1 _16185_ (.A(_07381_),
    .B(_07493_),
    .Y(_00960_));
 sg13g2_inv_1 _16186_ (.Y(_07494_),
    .A(_07482_));
 sg13g2_or4_1 _16187_ (.A(net319),
    .B(_07423_),
    .C(_07451_),
    .D(_07494_),
    .X(_07495_));
 sg13g2_nand2_1 _16188_ (.Y(_07496_),
    .A(net320),
    .B(net319));
 sg13g2_nor3_1 _16189_ (.A(_07467_),
    .B(_07476_),
    .C(_07496_),
    .Y(_07497_));
 sg13g2_and3_1 _16190_ (.X(_07498_),
    .A(net325),
    .B(net324),
    .C(_07423_));
 sg13g2_a22oi_1 _16191_ (.Y(_07499_),
    .B1(_07497_),
    .B2(_07498_),
    .A2(_07495_),
    .A1(net286));
 sg13g2_xnor2_1 _16192_ (.Y(_07500_),
    .A(net226),
    .B(_07499_));
 sg13g2_buf_1 _16193_ (.A(\am_sdr0.cic3.integ1[18] ),
    .X(_07501_));
 sg13g2_buf_1 _16194_ (.A(_07501_),
    .X(_07502_));
 sg13g2_nand2_1 _16195_ (.Y(_07503_),
    .A(_01559_),
    .B(_07502_));
 sg13g2_a21oi_1 _16196_ (.A1(net199),
    .A2(_07500_),
    .Y(_07504_),
    .B1(_07503_));
 sg13g2_inv_1 _16197_ (.Y(_07505_),
    .A(_07502_));
 sg13g2_nand4_1 _16198_ (.B(net199),
    .C(_07505_),
    .A(_01743_),
    .Y(_07506_),
    .D(_07500_));
 sg13g2_nand2b_1 _16199_ (.Y(_00961_),
    .B(_07506_),
    .A_N(_07504_));
 sg13g2_buf_1 _16200_ (.A(\am_sdr0.cic3.integ1[19] ),
    .X(_07507_));
 sg13g2_nor4_1 _16201_ (.A(net320),
    .B(net319),
    .C(net265),
    .D(_07474_),
    .Y(_07508_));
 sg13g2_nand4_1 _16202_ (.B(net320),
    .C(net319),
    .A(net321),
    .Y(_07509_),
    .D(net265));
 sg13g2_nor4_1 _16203_ (.A(_07466_),
    .B(_07429_),
    .C(_07467_),
    .D(_07509_),
    .Y(_07510_));
 sg13g2_o21ai_1 _16204_ (.B1(_07465_),
    .Y(_07511_),
    .A1(_07508_),
    .A2(_07510_));
 sg13g2_mux2_1 _16205_ (.A0(_07387_),
    .A1(_07508_),
    .S(_07511_),
    .X(_07512_));
 sg13g2_nand2_1 _16206_ (.Y(_07513_),
    .A(net267),
    .B(_07512_));
 sg13g2_xnor2_1 _16207_ (.Y(_07514_),
    .A(net318),
    .B(_07513_));
 sg13g2_and2_1 _16208_ (.A(_06552_),
    .B(_07514_),
    .X(_00962_));
 sg13g2_nand2_1 _16209_ (.Y(_07515_),
    .A(_05267_),
    .B(\am_sdr0.cic3.integ1[0] ));
 sg13g2_xnor2_1 _16210_ (.Y(_07516_),
    .A(_05270_),
    .B(_07515_));
 sg13g2_nand2_1 _16211_ (.Y(_07517_),
    .A(net197),
    .B(_07516_));
 sg13g2_xor2_1 _16212_ (.B(_07517_),
    .A(\am_sdr0.cic3.integ1[1] ),
    .X(_07518_));
 sg13g2_nor2_1 _16213_ (.A(net55),
    .B(_07518_),
    .Y(_00963_));
 sg13g2_buf_1 _16214_ (.A(\am_sdr0.cic3.integ1[20] ),
    .X(_07519_));
 sg13g2_buf_1 _16215_ (.A(_07519_),
    .X(_07520_));
 sg13g2_nor3_1 _16216_ (.A(net319),
    .B(net265),
    .C(net318),
    .Y(_07521_));
 sg13g2_nand3_1 _16217_ (.B(_07482_),
    .C(_07521_),
    .A(_07436_),
    .Y(_07522_));
 sg13g2_or2_1 _16218_ (.X(_07523_),
    .B(_07522_),
    .A(_07443_));
 sg13g2_nand3_1 _16219_ (.B(net318),
    .C(_07497_),
    .A(net265),
    .Y(_07524_));
 sg13g2_nor2_1 _16220_ (.A(_07441_),
    .B(_07524_),
    .Y(_07525_));
 sg13g2_nor2_1 _16221_ (.A(net286),
    .B(_07525_),
    .Y(_07526_));
 sg13g2_a21oi_1 _16222_ (.A1(net226),
    .A2(_07523_),
    .Y(_07527_),
    .B1(_07526_));
 sg13g2_and2_1 _16223_ (.A(net267),
    .B(_07527_),
    .X(_07528_));
 sg13g2_xnor2_1 _16224_ (.Y(_07529_),
    .A(net264),
    .B(_07528_));
 sg13g2_nor2_1 _16225_ (.A(_07381_),
    .B(_07529_),
    .Y(_00964_));
 sg13g2_buf_2 _16226_ (.A(_02778_),
    .X(_07530_));
 sg13g2_buf_1 _16227_ (.A(_07530_),
    .X(_07531_));
 sg13g2_buf_1 _16228_ (.A(\am_sdr0.cic3.integ1[21] ),
    .X(_07532_));
 sg13g2_buf_1 _16229_ (.A(net317),
    .X(_07533_));
 sg13g2_nor2_1 _16230_ (.A(net196),
    .B(net264),
    .Y(_07534_));
 sg13g2_nand2_1 _16231_ (.Y(_07535_),
    .A(_02425_),
    .B(_07534_));
 sg13g2_nor4_2 _16232_ (.A(net319),
    .B(net265),
    .C(net318),
    .Y(_07536_),
    .D(_07535_));
 sg13g2_and2_1 _16233_ (.A(_07482_),
    .B(_07490_),
    .X(_07537_));
 sg13g2_nand2_1 _16234_ (.Y(_07538_),
    .A(_02425_),
    .B(_07387_));
 sg13g2_inv_1 _16235_ (.Y(_07539_),
    .A(net264));
 sg13g2_nand2_1 _16236_ (.Y(_07540_),
    .A(net265),
    .B(net318));
 sg13g2_nor3_1 _16237_ (.A(_05263_),
    .B(_07539_),
    .C(_07540_),
    .Y(_07541_));
 sg13g2_a22oi_1 _16238_ (.Y(_07542_),
    .B1(_07541_),
    .B2(net319),
    .A2(_07534_),
    .A1(_07521_));
 sg13g2_nor3_1 _16239_ (.A(_07487_),
    .B(_07538_),
    .C(_07542_),
    .Y(_07543_));
 sg13g2_a22oi_1 _16240_ (.Y(_07544_),
    .B1(_07543_),
    .B2(_07453_),
    .A2(_07537_),
    .A1(_07536_));
 sg13g2_xor2_1 _16241_ (.B(_07544_),
    .A(net263),
    .X(_07545_));
 sg13g2_nor2_1 _16242_ (.A(net54),
    .B(_07545_),
    .Y(_00965_));
 sg13g2_buf_1 _16243_ (.A(\am_sdr0.cic3.integ1[22] ),
    .X(_07546_));
 sg13g2_nand2_1 _16244_ (.Y(_07547_),
    .A(net264),
    .B(net263));
 sg13g2_nor3_1 _16245_ (.A(_07540_),
    .B(_07538_),
    .C(_07547_),
    .Y(_07548_));
 sg13g2_nor4_1 _16246_ (.A(net265),
    .B(net318),
    .C(net263),
    .D(_07535_),
    .Y(_07549_));
 sg13g2_mux2_1 _16247_ (.A0(_07548_),
    .A1(_07549_),
    .S(_07499_),
    .X(_07550_));
 sg13g2_xnor2_1 _16248_ (.Y(_07551_),
    .A(net316),
    .B(_07550_));
 sg13g2_nor2_1 _16249_ (.A(net54),
    .B(_07551_),
    .Y(_00966_));
 sg13g2_buf_2 _16250_ (.A(\am_sdr0.cic3.integ1[23] ),
    .X(_07552_));
 sg13g2_nor2_1 _16251_ (.A(_07538_),
    .B(_07547_),
    .Y(_07553_));
 sg13g2_nand3_1 _16252_ (.B(net316),
    .C(_07553_),
    .A(net318),
    .Y(_07554_));
 sg13g2_nor4_1 _16253_ (.A(net321),
    .B(net320),
    .C(net263),
    .D(net316),
    .Y(_07555_));
 sg13g2_nand2_1 _16254_ (.Y(_07556_),
    .A(_07536_),
    .B(_07555_));
 sg13g2_mux2_1 _16255_ (.A0(_07554_),
    .A1(_07556_),
    .S(_07511_),
    .X(_07557_));
 sg13g2_xor2_1 _16256_ (.B(_07557_),
    .A(_07552_),
    .X(_07558_));
 sg13g2_nor2_1 _16257_ (.A(_07531_),
    .B(_07558_),
    .Y(_00967_));
 sg13g2_buf_2 _16258_ (.A(\am_sdr0.cic3.integ1[24] ),
    .X(_07559_));
 sg13g2_nand3_1 _16259_ (.B(_07552_),
    .C(_07553_),
    .A(net316),
    .Y(_07560_));
 sg13g2_nor4_1 _16260_ (.A(net263),
    .B(net316),
    .C(_07552_),
    .D(_07535_),
    .Y(_07561_));
 sg13g2_nand2b_1 _16261_ (.Y(_07562_),
    .B(_07561_),
    .A_N(_07523_));
 sg13g2_o21ai_1 _16262_ (.B1(_07562_),
    .Y(_07563_),
    .A1(_07526_),
    .A2(_07560_));
 sg13g2_xnor2_1 _16263_ (.Y(_07564_),
    .A(_07559_),
    .B(_07563_));
 sg13g2_nor2_1 _16264_ (.A(_07531_),
    .B(_07564_),
    .Y(_00968_));
 sg13g2_buf_1 _16265_ (.A(\am_sdr0.cic3.integ1[25] ),
    .X(_07565_));
 sg13g2_and2_1 _16266_ (.A(net297),
    .B(_07565_),
    .X(_07566_));
 sg13g2_nor2_1 _16267_ (.A(net251),
    .B(_07565_),
    .Y(_07567_));
 sg13g2_nand4_1 _16268_ (.B(net316),
    .C(_07552_),
    .A(net263),
    .Y(_07568_),
    .D(_07559_));
 sg13g2_or4_1 _16269_ (.A(_07449_),
    .B(_05264_),
    .C(_07542_),
    .D(_07568_),
    .X(_07569_));
 sg13g2_nor4_1 _16270_ (.A(net263),
    .B(net316),
    .C(_07552_),
    .D(_07559_),
    .Y(_07570_));
 sg13g2_nand3_1 _16271_ (.B(_07537_),
    .C(_07570_),
    .A(_07536_),
    .Y(_07571_));
 sg13g2_o21ai_1 _16272_ (.B1(_07571_),
    .Y(_07572_),
    .A1(_07490_),
    .A2(_07569_));
 sg13g2_mux2_1 _16273_ (.A0(_07566_),
    .A1(_07567_),
    .S(_07572_),
    .X(_00969_));
 sg13g2_nor2_1 _16274_ (.A(_07392_),
    .B(_07393_),
    .Y(_07573_));
 sg13g2_xor2_1 _16275_ (.B(_07573_),
    .A(_05250_),
    .X(_07574_));
 sg13g2_nand2_1 _16276_ (.Y(_07575_),
    .A(net197),
    .B(_07574_));
 sg13g2_xor2_1 _16277_ (.B(_07575_),
    .A(\am_sdr0.cic3.integ1[2] ),
    .X(_07576_));
 sg13g2_nor2_1 _16278_ (.A(net54),
    .B(_07576_),
    .Y(_00970_));
 sg13g2_nand2_1 _16279_ (.Y(_07577_),
    .A(_07395_),
    .B(_07397_));
 sg13g2_xnor2_1 _16280_ (.Y(_07578_),
    .A(_07391_),
    .B(_07577_));
 sg13g2_nor2_1 _16281_ (.A(net145),
    .B(_07578_),
    .Y(_07579_));
 sg13g2_xnor2_1 _16282_ (.Y(_07580_),
    .A(_07398_),
    .B(_07579_));
 sg13g2_nor2_1 _16283_ (.A(net54),
    .B(_07580_),
    .Y(_00971_));
 sg13g2_xnor2_1 _16284_ (.Y(_07581_),
    .A(\am_sdr0.cic1.x_out[12] ),
    .B(_07402_));
 sg13g2_nor2_1 _16285_ (.A(net145),
    .B(_07581_),
    .Y(_07582_));
 sg13g2_xnor2_1 _16286_ (.Y(_07583_),
    .A(_07390_),
    .B(_07582_));
 sg13g2_nor2_1 _16287_ (.A(net54),
    .B(_07583_),
    .Y(_00972_));
 sg13g2_nand2_1 _16288_ (.Y(_07584_),
    .A(_07403_),
    .B(_07404_));
 sg13g2_xor2_1 _16289_ (.B(_07584_),
    .A(\am_sdr0.cic1.x_out[13] ),
    .X(_07585_));
 sg13g2_nand2_1 _16290_ (.Y(_07586_),
    .A(net199),
    .B(_07585_));
 sg13g2_xnor2_1 _16291_ (.Y(_07587_),
    .A(_07389_),
    .B(_07586_));
 sg13g2_nor2_1 _16292_ (.A(net54),
    .B(_07587_),
    .Y(_00973_));
 sg13g2_xnor2_1 _16293_ (.Y(_07588_),
    .A(\am_sdr0.cic1.x_out[14] ),
    .B(_07408_));
 sg13g2_nor2_1 _16294_ (.A(net145),
    .B(_07588_),
    .Y(_07589_));
 sg13g2_xnor2_1 _16295_ (.Y(_07590_),
    .A(_07388_),
    .B(_07589_));
 sg13g2_nor2_1 _16296_ (.A(net54),
    .B(_07590_),
    .Y(_00974_));
 sg13g2_xnor2_1 _16297_ (.Y(_07591_),
    .A(net226),
    .B(_07412_));
 sg13g2_nor2_1 _16298_ (.A(net145),
    .B(_07591_),
    .Y(_07592_));
 sg13g2_xnor2_1 _16299_ (.Y(_07593_),
    .A(net266),
    .B(_07592_));
 sg13g2_nor2_1 _16300_ (.A(net54),
    .B(_07593_),
    .Y(_00975_));
 sg13g2_buf_1 _16301_ (.A(_07530_),
    .X(_07594_));
 sg13g2_nor2b_1 _16302_ (.A(net286),
    .B_N(net266),
    .Y(_07595_));
 sg13g2_and2_1 _16303_ (.A(_07412_),
    .B(_07595_),
    .X(_07596_));
 sg13g2_nor3_1 _16304_ (.A(net196),
    .B(net266),
    .C(_07412_),
    .Y(_07597_));
 sg13g2_o21ai_1 _16305_ (.B1(net198),
    .Y(_07598_),
    .A1(_07596_),
    .A2(_07597_));
 sg13g2_xnor2_1 _16306_ (.Y(_07599_),
    .A(_07414_),
    .B(_07598_));
 sg13g2_nor2_1 _16307_ (.A(net53),
    .B(_07599_),
    .Y(_00976_));
 sg13g2_nand3_1 _16308_ (.B(_07412_),
    .C(_07595_),
    .A(_07413_),
    .Y(_07600_));
 sg13g2_or4_1 _16309_ (.A(net196),
    .B(net266),
    .C(_07413_),
    .D(_07412_),
    .X(_07601_));
 sg13g2_a21oi_1 _16310_ (.A1(_07600_),
    .A2(_07601_),
    .Y(_07602_),
    .B1(_07449_));
 sg13g2_xnor2_1 _16311_ (.Y(_07603_),
    .A(_07415_),
    .B(_07602_));
 sg13g2_nor2_1 _16312_ (.A(net53),
    .B(_07603_),
    .Y(_00977_));
 sg13g2_buf_1 _16313_ (.A(net267),
    .X(_07604_));
 sg13g2_nand2_1 _16314_ (.Y(_07605_),
    .A(net195),
    .B(_07398_));
 sg13g2_xor2_1 _16315_ (.B(_07605_),
    .A(\am_sdr0.cic3.integ2[0] ),
    .X(_07606_));
 sg13g2_nor2_1 _16316_ (.A(net53),
    .B(_07606_),
    .Y(_00978_));
 sg13g2_buf_1 _16317_ (.A(\am_sdr0.cic3.integ2[10] ),
    .X(_07607_));
 sg13g2_buf_2 _16318_ (.A(\am_sdr0.cic3.integ2[9] ),
    .X(_07608_));
 sg13g2_inv_1 _16319_ (.Y(_07609_),
    .A(_07608_));
 sg13g2_buf_2 _16320_ (.A(\am_sdr0.cic3.integ2[7] ),
    .X(_07610_));
 sg13g2_nor2_1 _16321_ (.A(net325),
    .B(_07610_),
    .Y(_07611_));
 sg13g2_buf_2 _16322_ (.A(\am_sdr0.cic3.integ2[5] ),
    .X(_07612_));
 sg13g2_nor2_1 _16323_ (.A(_07413_),
    .B(_07612_),
    .Y(_07613_));
 sg13g2_buf_2 _16324_ (.A(\am_sdr0.cic3.integ2[4] ),
    .X(_07614_));
 sg13g2_nor2_1 _16325_ (.A(_07420_),
    .B(_07614_),
    .Y(_07615_));
 sg13g2_or2_1 _16326_ (.X(_07616_),
    .B(_07615_),
    .A(_07613_));
 sg13g2_buf_1 _16327_ (.A(\am_sdr0.cic3.integ2[3] ),
    .X(_07617_));
 sg13g2_inv_1 _16328_ (.Y(_07618_),
    .A(_07617_));
 sg13g2_nand2_1 _16329_ (.Y(_07619_),
    .A(\am_sdr0.cic3.integ1[5] ),
    .B(\am_sdr0.cic3.integ2[2] ));
 sg13g2_nor2_1 _16330_ (.A(\am_sdr0.cic3.integ1[5] ),
    .B(\am_sdr0.cic3.integ2[2] ),
    .Y(_07620_));
 sg13g2_nor2_1 _16331_ (.A(_07390_),
    .B(\am_sdr0.cic3.integ2[1] ),
    .Y(_07621_));
 sg13g2_a22oi_1 _16332_ (.Y(_07622_),
    .B1(\am_sdr0.cic3.integ2[1] ),
    .B2(_07390_),
    .A2(\am_sdr0.cic3.integ2[0] ),
    .A1(_07398_));
 sg13g2_or3_1 _16333_ (.A(_07620_),
    .B(_07621_),
    .C(_07622_),
    .X(_07623_));
 sg13g2_buf_1 _16334_ (.A(_07623_),
    .X(_07624_));
 sg13g2_nand3_1 _16335_ (.B(_07619_),
    .C(_07624_),
    .A(_07618_),
    .Y(_07625_));
 sg13g2_a21oi_1 _16336_ (.A1(_07619_),
    .A2(_07624_),
    .Y(_07626_),
    .B1(_07618_));
 sg13g2_a221oi_1 _16337_ (.B2(_07388_),
    .C1(_07626_),
    .B1(_07625_),
    .A1(_07420_),
    .Y(_07627_),
    .A2(_07614_));
 sg13g2_nand2_1 _16338_ (.Y(_07628_),
    .A(_07413_),
    .B(_07612_));
 sg13g2_o21ai_1 _16339_ (.B1(_07628_),
    .Y(_07629_),
    .A1(_07616_),
    .A2(_07627_));
 sg13g2_buf_2 _16340_ (.A(\am_sdr0.cic3.integ2[6] ),
    .X(_07630_));
 sg13g2_or2_1 _16341_ (.X(_07631_),
    .B(_07630_),
    .A(_07415_));
 sg13g2_and2_1 _16342_ (.A(_07415_),
    .B(_07630_),
    .X(_07632_));
 sg13g2_a221oi_1 _16343_ (.B2(_07631_),
    .C1(_07632_),
    .B1(_07629_),
    .A1(net325),
    .Y(_07633_),
    .A2(_07610_));
 sg13g2_buf_1 _16344_ (.A(_07633_),
    .X(_07634_));
 sg13g2_buf_2 _16345_ (.A(\am_sdr0.cic3.integ2[8] ),
    .X(_07635_));
 sg13g2_inv_1 _16346_ (.Y(_07636_),
    .A(_07635_));
 sg13g2_o21ai_1 _16347_ (.B1(_07636_),
    .Y(_07637_),
    .A1(_07611_),
    .A2(_07634_));
 sg13g2_nor3_1 _16348_ (.A(_07636_),
    .B(_07611_),
    .C(_07634_),
    .Y(_07638_));
 sg13g2_a21oi_2 _16349_ (.B1(_07638_),
    .Y(_07639_),
    .A2(_07637_),
    .A1(net324));
 sg13g2_o21ai_1 _16350_ (.B1(_07436_),
    .Y(_07640_),
    .A1(_07609_),
    .A2(_07639_));
 sg13g2_nand2_1 _16351_ (.Y(_07641_),
    .A(_07609_),
    .B(_07639_));
 sg13g2_nand2_1 _16352_ (.Y(_07642_),
    .A(_07640_),
    .B(_07641_));
 sg13g2_xnor2_1 _16353_ (.Y(_07643_),
    .A(net323),
    .B(_07642_));
 sg13g2_nand2_1 _16354_ (.Y(_07644_),
    .A(net195),
    .B(_07643_));
 sg13g2_xor2_1 _16355_ (.B(_07644_),
    .A(net315),
    .X(_07645_));
 sg13g2_nor2_1 _16356_ (.A(net53),
    .B(_07645_),
    .Y(_00979_));
 sg13g2_buf_1 _16357_ (.A(\am_sdr0.cic3.integ2[11] ),
    .X(_07646_));
 sg13g2_a21oi_1 _16358_ (.A1(_07640_),
    .A2(_07641_),
    .Y(_07647_),
    .B1(net315));
 sg13g2_nand3_1 _16359_ (.B(_07640_),
    .C(_07641_),
    .A(net315),
    .Y(_07648_));
 sg13g2_o21ai_1 _16360_ (.B1(_07648_),
    .Y(_07649_),
    .A1(_07485_),
    .A2(_07647_));
 sg13g2_xnor2_1 _16361_ (.Y(_07650_),
    .A(net322),
    .B(_07649_));
 sg13g2_nor2_1 _16362_ (.A(net145),
    .B(_07650_),
    .Y(_07651_));
 sg13g2_xnor2_1 _16363_ (.Y(_07652_),
    .A(net314),
    .B(_07651_));
 sg13g2_nor2_1 _16364_ (.A(net53),
    .B(_07652_),
    .Y(_00980_));
 sg13g2_buf_2 _16365_ (.A(\am_sdr0.cic3.integ2[12] ),
    .X(_07653_));
 sg13g2_or2_1 _16366_ (.X(_07654_),
    .B(net314),
    .A(net322));
 sg13g2_and2_1 _16367_ (.A(_07457_),
    .B(net314),
    .X(_07655_));
 sg13g2_a21oi_1 _16368_ (.A1(_07649_),
    .A2(_07654_),
    .Y(_07656_),
    .B1(_07655_));
 sg13g2_xnor2_1 _16369_ (.Y(_07657_),
    .A(net321),
    .B(_07656_));
 sg13g2_nand2_1 _16370_ (.Y(_07658_),
    .A(net195),
    .B(_07657_));
 sg13g2_xor2_1 _16371_ (.B(_07658_),
    .A(_07653_),
    .X(_07659_));
 sg13g2_nor2_1 _16372_ (.A(net53),
    .B(_07659_),
    .Y(_00981_));
 sg13g2_buf_2 _16373_ (.A(\am_sdr0.cic3.integ2[13] ),
    .X(_07660_));
 sg13g2_buf_1 _16374_ (.A(_07449_),
    .X(_07661_));
 sg13g2_nor2_1 _16375_ (.A(\am_sdr0.cic3.integ1[13] ),
    .B(net315),
    .Y(_07662_));
 sg13g2_or2_1 _16376_ (.X(_07663_),
    .B(_07608_),
    .A(_07435_));
 sg13g2_or2_1 _16377_ (.X(_07664_),
    .B(_07635_),
    .A(net324));
 sg13g2_and2_1 _16378_ (.A(_07435_),
    .B(_07608_),
    .X(_07665_));
 sg13g2_a21oi_1 _16379_ (.A1(_07663_),
    .A2(_07664_),
    .Y(_07666_),
    .B1(_07665_));
 sg13g2_nand2_1 _16380_ (.Y(_07667_),
    .A(_07447_),
    .B(net315));
 sg13g2_o21ai_1 _16381_ (.B1(_07667_),
    .Y(_07668_),
    .A1(_07662_),
    .A2(_07666_));
 sg13g2_nand2_1 _16382_ (.Y(_07669_),
    .A(net314),
    .B(_07668_));
 sg13g2_o21ai_1 _16383_ (.B1(_07457_),
    .Y(_07670_),
    .A1(net314),
    .A2(_07668_));
 sg13g2_nor2_1 _16384_ (.A(net321),
    .B(_07653_),
    .Y(_07671_));
 sg13g2_a21oi_1 _16385_ (.A1(_07669_),
    .A2(_07670_),
    .Y(_07672_),
    .B1(_07671_));
 sg13g2_a21oi_2 _16386_ (.B1(_07672_),
    .Y(_07673_),
    .A2(_07653_),
    .A1(_07462_));
 sg13g2_nand2_1 _16387_ (.Y(_07674_),
    .A(_07435_),
    .B(_07608_));
 sg13g2_a21oi_1 _16388_ (.A1(_07674_),
    .A2(_07667_),
    .Y(_07675_),
    .B1(_07662_));
 sg13g2_a221oi_1 _16389_ (.B2(_07462_),
    .C1(_07655_),
    .B1(_07653_),
    .A1(net324),
    .Y(_07676_),
    .A2(_07635_));
 sg13g2_nor2b_1 _16390_ (.A(_07675_),
    .B_N(_07676_),
    .Y(_07677_));
 sg13g2_o21ai_1 _16391_ (.B1(_07677_),
    .Y(_07678_),
    .A1(_07611_),
    .A2(_07634_));
 sg13g2_nand2b_1 _16392_ (.Y(_07679_),
    .B(_07678_),
    .A_N(_07673_));
 sg13g2_xnor2_1 _16393_ (.Y(_07680_),
    .A(_07473_),
    .B(_07679_));
 sg13g2_nor2_1 _16394_ (.A(net144),
    .B(_07680_),
    .Y(_07681_));
 sg13g2_xnor2_1 _16395_ (.Y(_07682_),
    .A(_07660_),
    .B(_07681_));
 sg13g2_nor2_1 _16396_ (.A(net53),
    .B(_07682_),
    .Y(_00982_));
 sg13g2_buf_2 _16397_ (.A(\am_sdr0.cic3.integ2[14] ),
    .X(_07683_));
 sg13g2_nor2_1 _16398_ (.A(net320),
    .B(_07660_),
    .Y(_07684_));
 sg13g2_nand2_1 _16399_ (.Y(_07685_),
    .A(_07472_),
    .B(_07660_));
 sg13g2_o21ai_1 _16400_ (.B1(_07685_),
    .Y(_07686_),
    .A1(_07679_),
    .A2(_07684_));
 sg13g2_xnor2_1 _16401_ (.Y(_07687_),
    .A(_07481_),
    .B(_07686_));
 sg13g2_nor2_1 _16402_ (.A(_07661_),
    .B(_07687_),
    .Y(_07688_));
 sg13g2_xnor2_1 _16403_ (.Y(_07689_),
    .A(_07683_),
    .B(_07688_));
 sg13g2_nor2_1 _16404_ (.A(net53),
    .B(_07689_),
    .Y(_00983_));
 sg13g2_buf_1 _16405_ (.A(\am_sdr0.cic3.integ2[15] ),
    .X(_07690_));
 sg13g2_inv_1 _16406_ (.Y(_07691_),
    .A(_07660_));
 sg13g2_nor2_1 _16407_ (.A(\am_sdr0.cic3.integ1[17] ),
    .B(_07683_),
    .Y(_07692_));
 sg13g2_buf_1 _16408_ (.A(_07692_),
    .X(_07693_));
 sg13g2_nor3_1 _16409_ (.A(_07691_),
    .B(_07673_),
    .C(_07693_),
    .Y(_07694_));
 sg13g2_nor3_1 _16410_ (.A(_07473_),
    .B(_07673_),
    .C(_07693_),
    .Y(_07695_));
 sg13g2_o21ai_1 _16411_ (.B1(_07678_),
    .Y(_07696_),
    .A1(_07694_),
    .A2(_07695_));
 sg13g2_and2_1 _16412_ (.A(_07481_),
    .B(_07683_),
    .X(_07697_));
 sg13g2_nor2_1 _16413_ (.A(_07685_),
    .B(_07693_),
    .Y(_07698_));
 sg13g2_nor2_1 _16414_ (.A(_07697_),
    .B(_07698_),
    .Y(_07699_));
 sg13g2_nand2_1 _16415_ (.Y(_07700_),
    .A(_07696_),
    .B(_07699_));
 sg13g2_xnor2_1 _16416_ (.Y(_07701_),
    .A(_07505_),
    .B(_07700_));
 sg13g2_nand2_1 _16417_ (.Y(_07702_),
    .A(_07604_),
    .B(_07701_));
 sg13g2_xor2_1 _16418_ (.B(_07702_),
    .A(net313),
    .X(_07703_));
 sg13g2_nor2_1 _16419_ (.A(_07594_),
    .B(_07703_),
    .Y(_00984_));
 sg13g2_buf_1 _16420_ (.A(\am_sdr0.cic3.integ2[16] ),
    .X(_07704_));
 sg13g2_or2_1 _16421_ (.X(_07705_),
    .B(net313),
    .A(_07501_));
 sg13g2_buf_1 _16422_ (.A(_07705_),
    .X(_07706_));
 sg13g2_and2_1 _16423_ (.A(_07501_),
    .B(net313),
    .X(_07707_));
 sg13g2_a21oi_1 _16424_ (.A1(_07700_),
    .A2(_07706_),
    .Y(_07708_),
    .B1(_07707_));
 sg13g2_xnor2_1 _16425_ (.Y(_07709_),
    .A(net318),
    .B(_07708_));
 sg13g2_nand2_1 _16426_ (.Y(_07710_),
    .A(net195),
    .B(_07709_));
 sg13g2_xor2_1 _16427_ (.B(_07710_),
    .A(net312),
    .X(_07711_));
 sg13g2_nor2_1 _16428_ (.A(_07594_),
    .B(_07711_),
    .Y(_00985_));
 sg13g2_buf_1 _16429_ (.A(_07530_),
    .X(_07712_));
 sg13g2_buf_1 _16430_ (.A(\am_sdr0.cic3.integ2[17] ),
    .X(_07713_));
 sg13g2_buf_1 _16431_ (.A(_07713_),
    .X(_07714_));
 sg13g2_inv_2 _16432_ (.Y(_07715_),
    .A(_07714_));
 sg13g2_nand2_1 _16433_ (.Y(_07716_),
    .A(net312),
    .B(_07706_));
 sg13g2_nor4_1 _16434_ (.A(_07691_),
    .B(_07673_),
    .C(_07693_),
    .D(_07716_),
    .Y(_07717_));
 sg13g2_nor4_1 _16435_ (.A(_07473_),
    .B(_07673_),
    .C(_07693_),
    .D(_07716_),
    .Y(_07718_));
 sg13g2_o21ai_1 _16436_ (.B1(_07678_),
    .Y(_07719_),
    .A1(_07717_),
    .A2(_07718_));
 sg13g2_or3_1 _16437_ (.A(_07685_),
    .B(_07693_),
    .C(_07716_),
    .X(_07720_));
 sg13g2_a21o_1 _16438_ (.A2(_07706_),
    .A1(_07697_),
    .B1(_07707_),
    .X(_07721_));
 sg13g2_a21oi_1 _16439_ (.A1(net312),
    .A2(_07721_),
    .Y(_07722_),
    .B1(_07507_));
 sg13g2_nand3_1 _16440_ (.B(_07720_),
    .C(_07722_),
    .A(_07719_),
    .Y(_07723_));
 sg13g2_nor2_1 _16441_ (.A(net313),
    .B(net312),
    .Y(_07724_));
 sg13g2_nand3_1 _16442_ (.B(_07699_),
    .C(_07724_),
    .A(_07696_),
    .Y(_07725_));
 sg13g2_nor2_1 _16443_ (.A(net265),
    .B(net312),
    .Y(_07726_));
 sg13g2_nand3_1 _16444_ (.B(_07699_),
    .C(_07726_),
    .A(_07696_),
    .Y(_07727_));
 sg13g2_or2_1 _16445_ (.X(_07728_),
    .B(_07706_),
    .A(net312));
 sg13g2_nand4_1 _16446_ (.B(_07725_),
    .C(_07727_),
    .A(_07723_),
    .Y(_07729_),
    .D(_07728_));
 sg13g2_buf_2 _16447_ (.A(_07729_),
    .X(_07730_));
 sg13g2_xnor2_1 _16448_ (.Y(_07731_),
    .A(net264),
    .B(_07730_));
 sg13g2_nand2_1 _16449_ (.Y(_07732_),
    .A(net197),
    .B(_07731_));
 sg13g2_xnor2_1 _16450_ (.Y(_07733_),
    .A(_07715_),
    .B(_07732_));
 sg13g2_nor2_1 _16451_ (.A(_07712_),
    .B(_07733_),
    .Y(_00986_));
 sg13g2_buf_1 _16452_ (.A(\am_sdr0.cic3.integ2[18] ),
    .X(_07734_));
 sg13g2_buf_1 _16453_ (.A(_07734_),
    .X(_07735_));
 sg13g2_nand2_1 _16454_ (.Y(_07736_),
    .A(_07715_),
    .B(_07730_));
 sg13g2_nor2_1 _16455_ (.A(_07715_),
    .B(_07730_),
    .Y(_07737_));
 sg13g2_a21oi_1 _16456_ (.A1(net264),
    .A2(_07736_),
    .Y(_07738_),
    .B1(_07737_));
 sg13g2_xnor2_1 _16457_ (.Y(_07739_),
    .A(_07533_),
    .B(_07738_));
 sg13g2_nand2_1 _16458_ (.Y(_07740_),
    .A(_07604_),
    .B(_07739_));
 sg13g2_xor2_1 _16459_ (.B(_07740_),
    .A(net261),
    .X(_07741_));
 sg13g2_nor2_1 _16460_ (.A(net52),
    .B(_07741_),
    .Y(_00987_));
 sg13g2_nand2_1 _16461_ (.Y(_07742_),
    .A(net263),
    .B(net261));
 sg13g2_nor2_1 _16462_ (.A(_07533_),
    .B(_07735_),
    .Y(_07743_));
 sg13g2_a21oi_1 _16463_ (.A1(_07738_),
    .A2(_07742_),
    .Y(_07744_),
    .B1(_07743_));
 sg13g2_xor2_1 _16464_ (.B(_07744_),
    .A(net316),
    .X(_07745_));
 sg13g2_buf_1 _16465_ (.A(\am_sdr0.cic3.integ2[19] ),
    .X(_07746_));
 sg13g2_buf_1 _16466_ (.A(_07746_),
    .X(_07747_));
 sg13g2_nand2_1 _16467_ (.Y(_07748_),
    .A(_01559_),
    .B(net260));
 sg13g2_a21oi_1 _16468_ (.A1(_07364_),
    .A2(_07745_),
    .Y(_07749_),
    .B1(_07748_));
 sg13g2_inv_1 _16469_ (.Y(_07750_),
    .A(net260));
 sg13g2_nand4_1 _16470_ (.B(net199),
    .C(_07750_),
    .A(_01743_),
    .Y(_07751_),
    .D(_07745_));
 sg13g2_nand2b_1 _16471_ (.Y(_00988_),
    .B(_07751_),
    .A_N(_07749_));
 sg13g2_nand2_1 _16472_ (.Y(_07752_),
    .A(_07398_),
    .B(\am_sdr0.cic3.integ2[0] ));
 sg13g2_xnor2_1 _16473_ (.Y(_07753_),
    .A(_07390_),
    .B(_07752_));
 sg13g2_nand2_1 _16474_ (.Y(_07754_),
    .A(net195),
    .B(_07753_));
 sg13g2_xor2_1 _16475_ (.B(_07754_),
    .A(\am_sdr0.cic3.integ2[1] ),
    .X(_07755_));
 sg13g2_nor2_1 _16476_ (.A(net52),
    .B(_07755_),
    .Y(_00989_));
 sg13g2_buf_2 _16477_ (.A(\am_sdr0.cic3.integ2[20] ),
    .X(_07756_));
 sg13g2_and2_1 _16478_ (.A(_02808_),
    .B(_07756_),
    .X(_07757_));
 sg13g2_nor2_1 _16479_ (.A(_01968_),
    .B(_07756_),
    .Y(_07758_));
 sg13g2_nand3_1 _16480_ (.B(net261),
    .C(net260),
    .A(net262),
    .Y(_07759_));
 sg13g2_nand3_1 _16481_ (.B(net261),
    .C(_07746_),
    .A(net264),
    .Y(_07760_));
 sg13g2_a21oi_1 _16482_ (.A1(_07759_),
    .A2(_07760_),
    .Y(_07761_),
    .B1(_07730_));
 sg13g2_nand3_1 _16483_ (.B(net262),
    .C(net260),
    .A(net317),
    .Y(_07762_));
 sg13g2_nand3_1 _16484_ (.B(net317),
    .C(net311),
    .A(net264),
    .Y(_07763_));
 sg13g2_a21oi_1 _16485_ (.A1(_07762_),
    .A2(_07763_),
    .Y(_07764_),
    .B1(_07730_));
 sg13g2_nand4_1 _16486_ (.B(net262),
    .C(net261),
    .A(_07520_),
    .Y(_07765_),
    .D(net260));
 sg13g2_nand3_1 _16487_ (.B(net261),
    .C(net260),
    .A(net317),
    .Y(_07766_));
 sg13g2_nand4_1 _16488_ (.B(_07532_),
    .C(net262),
    .A(_07520_),
    .Y(_07767_),
    .D(net260));
 sg13g2_nand3_1 _16489_ (.B(_07766_),
    .C(_07767_),
    .A(_07765_),
    .Y(_07768_));
 sg13g2_nor3_1 _16490_ (.A(_07761_),
    .B(_07764_),
    .C(_07768_),
    .Y(_07769_));
 sg13g2_nor3_1 _16491_ (.A(net262),
    .B(_07734_),
    .C(net311),
    .Y(_07770_));
 sg13g2_nor3_1 _16492_ (.A(_07519_),
    .B(net261),
    .C(net311),
    .Y(_07771_));
 sg13g2_o21ai_1 _16493_ (.B1(_07730_),
    .Y(_07772_),
    .A1(_07770_),
    .A2(_07771_));
 sg13g2_nor3_1 _16494_ (.A(net317),
    .B(net262),
    .C(net311),
    .Y(_07773_));
 sg13g2_nor3_1 _16495_ (.A(_07519_),
    .B(net317),
    .C(net311),
    .Y(_07774_));
 sg13g2_o21ai_1 _16496_ (.B1(_07730_),
    .Y(_07775_),
    .A1(_07773_),
    .A2(_07774_));
 sg13g2_nor4_1 _16497_ (.A(_07519_),
    .B(net262),
    .C(_07734_),
    .D(net311),
    .Y(_07776_));
 sg13g2_nor3_1 _16498_ (.A(net317),
    .B(net261),
    .C(net311),
    .Y(_07777_));
 sg13g2_nor4_1 _16499_ (.A(_07519_),
    .B(net317),
    .C(net262),
    .D(net311),
    .Y(_07778_));
 sg13g2_nor3_1 _16500_ (.A(_07776_),
    .B(_07777_),
    .C(_07778_),
    .Y(_07779_));
 sg13g2_nand4_1 _16501_ (.B(_07772_),
    .C(_07775_),
    .A(_07546_),
    .Y(_07780_),
    .D(_07779_));
 sg13g2_nand2_1 _16502_ (.Y(_07781_),
    .A(_07769_),
    .B(_07780_));
 sg13g2_xnor2_1 _16503_ (.Y(_07782_),
    .A(_07552_),
    .B(_07781_));
 sg13g2_nor2_1 _16504_ (.A(_07450_),
    .B(_07782_),
    .Y(_07783_));
 sg13g2_mux2_1 _16505_ (.A0(_07757_),
    .A1(_07758_),
    .S(_07783_),
    .X(_00990_));
 sg13g2_buf_2 _16506_ (.A(\am_sdr0.cic3.integ2[21] ),
    .X(_07784_));
 sg13g2_nand2_1 _16507_ (.Y(_07785_),
    .A(_07552_),
    .B(_07756_));
 sg13g2_nand3_1 _16508_ (.B(_07559_),
    .C(_07785_),
    .A(_02425_),
    .Y(_07786_));
 sg13g2_nor2_1 _16509_ (.A(_07552_),
    .B(_07756_),
    .Y(_07787_));
 sg13g2_nor2_1 _16510_ (.A(_07449_),
    .B(_07559_),
    .Y(_07788_));
 sg13g2_nand2b_1 _16511_ (.Y(_07789_),
    .B(_07788_),
    .A_N(_07787_));
 sg13g2_mux2_1 _16512_ (.A0(_07786_),
    .A1(_07789_),
    .S(_07781_),
    .X(_07790_));
 sg13g2_nand3_1 _16513_ (.B(_07559_),
    .C(_07787_),
    .A(net267),
    .Y(_07791_));
 sg13g2_nand2b_1 _16514_ (.Y(_07792_),
    .B(_07788_),
    .A_N(_07785_));
 sg13g2_and2_1 _16515_ (.A(_07791_),
    .B(_07792_),
    .X(_07793_));
 sg13g2_nand3_1 _16516_ (.B(_07790_),
    .C(_07793_),
    .A(_07784_),
    .Y(_07794_));
 sg13g2_a21o_1 _16517_ (.A2(_07793_),
    .A1(_07790_),
    .B1(_07784_),
    .X(_07795_));
 sg13g2_a21oi_1 _16518_ (.A1(_07794_),
    .A2(_07795_),
    .Y(_00991_),
    .B1(net56));
 sg13g2_nand2_1 _16519_ (.Y(_07796_),
    .A(net267),
    .B(_07565_));
 sg13g2_nand2b_1 _16520_ (.Y(_07797_),
    .B(_07363_),
    .A_N(_07565_));
 sg13g2_nand2_1 _16521_ (.Y(_07798_),
    .A(_07559_),
    .B(_07784_));
 sg13g2_nand2_1 _16522_ (.Y(_07799_),
    .A(_07785_),
    .B(_07798_));
 sg13g2_nor4_1 _16523_ (.A(_07761_),
    .B(_07764_),
    .C(_07768_),
    .D(_07799_),
    .Y(_07800_));
 sg13g2_nor2_1 _16524_ (.A(_07559_),
    .B(_07784_),
    .Y(_07801_));
 sg13g2_a221oi_1 _16525_ (.B2(_07780_),
    .C1(_07801_),
    .B1(_07800_),
    .A1(_07787_),
    .Y(_07802_),
    .A2(_07798_));
 sg13g2_mux2_1 _16526_ (.A0(_07796_),
    .A1(_07797_),
    .S(_07802_),
    .X(_07803_));
 sg13g2_xor2_1 _16527_ (.B(_07803_),
    .A(\am_sdr0.cic3.integ2[22] ),
    .X(_07804_));
 sg13g2_nor2_1 _16528_ (.A(_07712_),
    .B(_07804_),
    .Y(_00992_));
 sg13g2_nor2_1 _16529_ (.A(_07621_),
    .B(_07622_),
    .Y(_07805_));
 sg13g2_xnor2_1 _16530_ (.Y(_07806_),
    .A(_07389_),
    .B(_07805_));
 sg13g2_nand2_1 _16531_ (.Y(_07807_),
    .A(net195),
    .B(_07806_));
 sg13g2_xor2_1 _16532_ (.B(_07807_),
    .A(\am_sdr0.cic3.integ2[2] ),
    .X(_07808_));
 sg13g2_nor2_1 _16533_ (.A(net52),
    .B(_07808_),
    .Y(_00993_));
 sg13g2_nand2_1 _16534_ (.Y(_07809_),
    .A(_07619_),
    .B(_07624_));
 sg13g2_xnor2_1 _16535_ (.Y(_07810_),
    .A(_07388_),
    .B(_07809_));
 sg13g2_nor2_1 _16536_ (.A(net144),
    .B(_07810_),
    .Y(_07811_));
 sg13g2_xnor2_1 _16537_ (.Y(_07812_),
    .A(_07617_),
    .B(_07811_));
 sg13g2_nor2_1 _16538_ (.A(net52),
    .B(_07812_),
    .Y(_00994_));
 sg13g2_a21oi_1 _16539_ (.A1(_07388_),
    .A2(_07625_),
    .Y(_07813_),
    .B1(_07626_));
 sg13g2_xnor2_1 _16540_ (.Y(_07814_),
    .A(_07421_),
    .B(_07813_));
 sg13g2_nand2_1 _16541_ (.Y(_07815_),
    .A(net195),
    .B(_07814_));
 sg13g2_xor2_1 _16542_ (.B(_07815_),
    .A(_07614_),
    .X(_07816_));
 sg13g2_nor2_1 _16543_ (.A(net52),
    .B(_07816_),
    .Y(_00995_));
 sg13g2_nand2_1 _16544_ (.Y(_07817_),
    .A(_07421_),
    .B(_07614_));
 sg13g2_o21ai_1 _16545_ (.B1(_07817_),
    .Y(_07818_),
    .A1(_07615_),
    .A2(_07813_));
 sg13g2_xnor2_1 _16546_ (.Y(_07819_),
    .A(_07413_),
    .B(_07818_));
 sg13g2_nor2_1 _16547_ (.A(net144),
    .B(_07819_),
    .Y(_07820_));
 sg13g2_xnor2_1 _16548_ (.Y(_07821_),
    .A(_07612_),
    .B(_07820_));
 sg13g2_nor2_1 _16549_ (.A(net52),
    .B(_07821_),
    .Y(_00996_));
 sg13g2_xnor2_1 _16550_ (.Y(_07822_),
    .A(_07415_),
    .B(_07629_));
 sg13g2_nor2_1 _16551_ (.A(net144),
    .B(_07822_),
    .Y(_07823_));
 sg13g2_xnor2_1 _16552_ (.Y(_07824_),
    .A(_07630_),
    .B(_07823_));
 sg13g2_nor2_1 _16553_ (.A(net52),
    .B(_07824_),
    .Y(_00997_));
 sg13g2_a21oi_1 _16554_ (.A1(_07629_),
    .A2(_07631_),
    .Y(_07825_),
    .B1(_07632_));
 sg13g2_xnor2_1 _16555_ (.Y(_07826_),
    .A(_07385_),
    .B(_07825_));
 sg13g2_nand2_1 _16556_ (.Y(_07827_),
    .A(net195),
    .B(_07826_));
 sg13g2_xor2_1 _16557_ (.B(_07827_),
    .A(_07610_),
    .X(_07828_));
 sg13g2_nor2_1 _16558_ (.A(net52),
    .B(_07828_),
    .Y(_00998_));
 sg13g2_buf_1 _16559_ (.A(_07530_),
    .X(_07829_));
 sg13g2_nor2_1 _16560_ (.A(_07611_),
    .B(_07634_),
    .Y(_07830_));
 sg13g2_xnor2_1 _16561_ (.Y(_07831_),
    .A(_07431_),
    .B(_07830_));
 sg13g2_nor2_1 _16562_ (.A(net144),
    .B(_07831_),
    .Y(_07832_));
 sg13g2_xnor2_1 _16563_ (.Y(_07833_),
    .A(_07635_),
    .B(_07832_));
 sg13g2_nor2_1 _16564_ (.A(net51),
    .B(_07833_),
    .Y(_00999_));
 sg13g2_xnor2_1 _16565_ (.Y(_07834_),
    .A(_07435_),
    .B(_07639_));
 sg13g2_nand2_1 _16566_ (.Y(_07835_),
    .A(net197),
    .B(_07834_));
 sg13g2_xnor2_1 _16567_ (.Y(_07836_),
    .A(_07609_),
    .B(_07835_));
 sg13g2_nor2_1 _16568_ (.A(net51),
    .B(_07836_),
    .Y(_01000_));
 sg13g2_nand2_1 _16569_ (.Y(_07837_),
    .A(net198),
    .B(_07617_));
 sg13g2_xor2_1 _16570_ (.B(_07837_),
    .A(_02420_),
    .X(_07838_));
 sg13g2_nor2_1 _16571_ (.A(net51),
    .B(_07838_),
    .Y(_01001_));
 sg13g2_nand2_1 _16572_ (.Y(_07839_),
    .A(_07612_),
    .B(_02465_));
 sg13g2_nor2_1 _16573_ (.A(_07612_),
    .B(_02465_),
    .Y(_07840_));
 sg13g2_nor2_1 _16574_ (.A(_07614_),
    .B(_02462_),
    .Y(_07841_));
 sg13g2_a22oi_1 _16575_ (.Y(_07842_),
    .B1(_02462_),
    .B2(_07614_),
    .A2(_02420_),
    .A1(_07617_));
 sg13g2_or3_1 _16576_ (.A(_07840_),
    .B(_07841_),
    .C(_07842_),
    .X(_07843_));
 sg13g2_buf_1 _16577_ (.A(_07843_),
    .X(_07844_));
 sg13g2_nand3_1 _16578_ (.B(_07839_),
    .C(_07844_),
    .A(_02467_),
    .Y(_07845_));
 sg13g2_a21oi_1 _16579_ (.A1(_07839_),
    .A2(_07844_),
    .Y(_07846_),
    .B1(_02467_));
 sg13g2_a221oi_1 _16580_ (.B2(_07630_),
    .C1(_07846_),
    .B1(_07845_),
    .A1(_07610_),
    .Y(_07847_),
    .A2(_02470_));
 sg13g2_buf_1 _16581_ (.A(_07847_),
    .X(_07848_));
 sg13g2_nor2_1 _16582_ (.A(_07610_),
    .B(_02470_),
    .Y(_07849_));
 sg13g2_o21ai_1 _16583_ (.B1(_02472_),
    .Y(_07850_),
    .A1(_07848_),
    .A2(_07849_));
 sg13g2_nor3_1 _16584_ (.A(_02472_),
    .B(_07848_),
    .C(_07849_),
    .Y(_07851_));
 sg13g2_a21oi_2 _16585_ (.B1(_07851_),
    .Y(_07852_),
    .A2(_07850_),
    .A1(_07635_));
 sg13g2_nor2_1 _16586_ (.A(_07608_),
    .B(_02475_),
    .Y(_07853_));
 sg13g2_nand2_1 _16587_ (.Y(_07854_),
    .A(_07608_),
    .B(_02475_));
 sg13g2_o21ai_1 _16588_ (.B1(_07854_),
    .Y(_07855_),
    .A1(_07852_),
    .A2(_07853_));
 sg13g2_buf_1 _16589_ (.A(_07855_),
    .X(_07856_));
 sg13g2_nor2_1 _16590_ (.A(_02477_),
    .B(_07856_),
    .Y(_07857_));
 sg13g2_a21oi_1 _16591_ (.A1(_02477_),
    .A2(_07856_),
    .Y(_07858_),
    .B1(net315));
 sg13g2_nor2_1 _16592_ (.A(_07857_),
    .B(_07858_),
    .Y(_07859_));
 sg13g2_a21o_1 _16593_ (.A2(_07859_),
    .A1(_02481_),
    .B1(net314),
    .X(_07860_));
 sg13g2_o21ai_1 _16594_ (.B1(_07860_),
    .Y(_07861_),
    .A1(_02481_),
    .A2(_07859_));
 sg13g2_nor2_1 _16595_ (.A(_07653_),
    .B(_02485_),
    .Y(_07862_));
 sg13g2_nand2_1 _16596_ (.Y(_07863_),
    .A(_07653_),
    .B(_02485_));
 sg13g2_o21ai_1 _16597_ (.B1(_07863_),
    .Y(_07864_),
    .A1(_07861_),
    .A2(_07862_));
 sg13g2_xnor2_1 _16598_ (.Y(_07865_),
    .A(_07660_),
    .B(_07864_));
 sg13g2_nor2_1 _16599_ (.A(_07661_),
    .B(_07865_),
    .Y(_07866_));
 sg13g2_xnor2_1 _16600_ (.Y(_07867_),
    .A(_02436_),
    .B(_07866_));
 sg13g2_nor2_1 _16601_ (.A(net51),
    .B(_07867_),
    .Y(_01002_));
 sg13g2_xnor2_1 _16602_ (.Y(_07868_),
    .A(_07660_),
    .B(_02436_));
 sg13g2_xnor2_1 _16603_ (.Y(_07869_),
    .A(net315),
    .B(_02477_));
 sg13g2_xnor2_1 _16604_ (.Y(_07870_),
    .A(net314),
    .B(_02481_));
 sg13g2_nand2b_1 _16605_ (.Y(_07871_),
    .B(_07863_),
    .A_N(_07862_));
 sg13g2_nor4_1 _16606_ (.A(_07868_),
    .B(_07869_),
    .C(_07870_),
    .D(_07871_),
    .Y(_07872_));
 sg13g2_nand2b_1 _16607_ (.Y(_07873_),
    .B(_07872_),
    .A_N(_07853_));
 sg13g2_nor2_1 _16608_ (.A(net314),
    .B(_02481_),
    .Y(_07874_));
 sg13g2_a22oi_1 _16609_ (.Y(_07875_),
    .B1(_02481_),
    .B2(_07646_),
    .A2(_02477_),
    .A1(net315));
 sg13g2_nor2_1 _16610_ (.A(_07874_),
    .B(_07875_),
    .Y(_07876_));
 sg13g2_a21oi_1 _16611_ (.A1(_02485_),
    .A2(_07876_),
    .Y(_07877_),
    .B1(_07653_));
 sg13g2_nor2_1 _16612_ (.A(_02485_),
    .B(_07876_),
    .Y(_07878_));
 sg13g2_nand2_1 _16613_ (.Y(_07879_),
    .A(_07660_),
    .B(_02436_));
 sg13g2_o21ai_1 _16614_ (.B1(_07879_),
    .Y(_07880_),
    .A1(_07877_),
    .A2(_07878_));
 sg13g2_o21ai_1 _16615_ (.B1(_07880_),
    .Y(_07881_),
    .A1(_07660_),
    .A2(_02436_));
 sg13g2_nand2b_1 _16616_ (.Y(_07882_),
    .B(_07872_),
    .A_N(_07854_));
 sg13g2_and2_1 _16617_ (.A(_07881_),
    .B(_07882_),
    .X(_07883_));
 sg13g2_o21ai_1 _16618_ (.B1(_07883_),
    .Y(_07884_),
    .A1(_07852_),
    .A2(_07873_));
 sg13g2_buf_2 _16619_ (.A(_07884_),
    .X(_07885_));
 sg13g2_xnor2_1 _16620_ (.Y(_07886_),
    .A(_07683_),
    .B(_07885_));
 sg13g2_nor2_1 _16621_ (.A(net144),
    .B(_07886_),
    .Y(_07887_));
 sg13g2_xnor2_1 _16622_ (.Y(_07888_),
    .A(_02438_),
    .B(_07887_));
 sg13g2_nor2_1 _16623_ (.A(net51),
    .B(_07888_),
    .Y(_01003_));
 sg13g2_nor2_1 _16624_ (.A(_02438_),
    .B(_07885_),
    .Y(_07889_));
 sg13g2_a21oi_1 _16625_ (.A1(_02438_),
    .A2(_07885_),
    .Y(_07890_),
    .B1(_07683_));
 sg13g2_nor2_1 _16626_ (.A(_07889_),
    .B(_07890_),
    .Y(_07891_));
 sg13g2_xnor2_1 _16627_ (.Y(_07892_),
    .A(net313),
    .B(_07891_));
 sg13g2_nor2_1 _16628_ (.A(net144),
    .B(_07892_),
    .Y(_07893_));
 sg13g2_xnor2_1 _16629_ (.Y(_07894_),
    .A(_02440_),
    .B(_07893_));
 sg13g2_nor2_1 _16630_ (.A(net51),
    .B(_07894_),
    .Y(_01004_));
 sg13g2_or2_1 _16631_ (.X(_07895_),
    .B(_02440_),
    .A(net313));
 sg13g2_and2_1 _16632_ (.A(net313),
    .B(_02440_),
    .X(_07896_));
 sg13g2_a21oi_1 _16633_ (.A1(_07891_),
    .A2(_07895_),
    .Y(_07897_),
    .B1(_07896_));
 sg13g2_xnor2_1 _16634_ (.Y(_07898_),
    .A(net312),
    .B(_07897_));
 sg13g2_nand2_1 _16635_ (.Y(_07899_),
    .A(_07366_),
    .B(_07898_));
 sg13g2_xor2_1 _16636_ (.B(_07899_),
    .A(_02444_),
    .X(_07900_));
 sg13g2_nor2_1 _16637_ (.A(net51),
    .B(_07900_),
    .Y(_01005_));
 sg13g2_or2_1 _16638_ (.X(_07901_),
    .B(_02444_),
    .A(net312));
 sg13g2_buf_1 _16639_ (.A(_07901_),
    .X(_07902_));
 sg13g2_and3_1 _16640_ (.X(_07903_),
    .A(_02438_),
    .B(_02440_),
    .C(_07902_));
 sg13g2_and3_1 _16641_ (.X(_07904_),
    .A(_07683_),
    .B(_02440_),
    .C(_07902_));
 sg13g2_o21ai_1 _16642_ (.B1(_07885_),
    .Y(_07905_),
    .A1(_07903_),
    .A2(_07904_));
 sg13g2_and3_1 _16643_ (.X(_07906_),
    .A(net313),
    .B(_02438_),
    .C(_07902_));
 sg13g2_and3_1 _16644_ (.X(_07907_),
    .A(_07683_),
    .B(_07690_),
    .C(_07902_));
 sg13g2_o21ai_1 _16645_ (.B1(_07885_),
    .Y(_07908_),
    .A1(_07906_),
    .A2(_07907_));
 sg13g2_and4_1 _16646_ (.A(_07683_),
    .B(_02438_),
    .C(_02440_),
    .D(_07902_),
    .X(_07909_));
 sg13g2_a221oi_1 _16647_ (.B2(_02438_),
    .C1(_07909_),
    .B1(_07907_),
    .A1(_07896_),
    .Y(_07910_),
    .A2(_07902_));
 sg13g2_buf_1 _16648_ (.A(_07910_),
    .X(_07911_));
 sg13g2_nand2_1 _16649_ (.Y(_07912_),
    .A(_07704_),
    .B(_02444_));
 sg13g2_nand4_1 _16650_ (.B(_07908_),
    .C(_07911_),
    .A(_07905_),
    .Y(_07913_),
    .D(_07912_));
 sg13g2_xnor2_1 _16651_ (.Y(_07914_),
    .A(_07715_),
    .B(_07913_));
 sg13g2_nand2_1 _16652_ (.Y(_07915_),
    .A(net197),
    .B(_07914_));
 sg13g2_xnor2_1 _16653_ (.Y(_07916_),
    .A(_02447_),
    .B(_07915_));
 sg13g2_nor2_1 _16654_ (.A(_07829_),
    .B(_07916_),
    .Y(_01006_));
 sg13g2_o21ai_1 _16655_ (.B1(_07913_),
    .Y(_07917_),
    .A1(_07714_),
    .A2(_02446_));
 sg13g2_o21ai_1 _16656_ (.B1(_07917_),
    .Y(_07918_),
    .A1(_07715_),
    .A2(_02447_));
 sg13g2_xor2_1 _16657_ (.B(_07918_),
    .A(_07735_),
    .X(_07919_));
 sg13g2_nand2_1 _16658_ (.Y(_07920_),
    .A(_07363_),
    .B(_07919_));
 sg13g2_xnor2_1 _16659_ (.Y(_07921_),
    .A(_02451_),
    .B(_07920_));
 sg13g2_and2_1 _16660_ (.A(_06552_),
    .B(_07921_),
    .X(_01007_));
 sg13g2_nand2_1 _16661_ (.Y(_07922_),
    .A(_07734_),
    .B(_02451_));
 sg13g2_nand2_1 _16662_ (.Y(_07923_),
    .A(_07912_),
    .B(_07922_));
 sg13g2_nor2_1 _16663_ (.A(_02446_),
    .B(_07923_),
    .Y(_07924_));
 sg13g2_nand4_1 _16664_ (.B(_07908_),
    .C(_07911_),
    .A(_07905_),
    .Y(_07925_),
    .D(_07924_));
 sg13g2_nor2_1 _16665_ (.A(_07713_),
    .B(_07923_),
    .Y(_07926_));
 sg13g2_nand4_1 _16666_ (.B(_07908_),
    .C(_07911_),
    .A(_07905_),
    .Y(_07927_),
    .D(_07926_));
 sg13g2_nor2_1 _16667_ (.A(_07713_),
    .B(_02446_),
    .Y(_07928_));
 sg13g2_nor2_1 _16668_ (.A(_07734_),
    .B(_02451_),
    .Y(_07929_));
 sg13g2_a21oi_1 _16669_ (.A1(_07928_),
    .A2(_07922_),
    .Y(_07930_),
    .B1(_07929_));
 sg13g2_nand3_1 _16670_ (.B(_07927_),
    .C(_07930_),
    .A(_07925_),
    .Y(_07931_));
 sg13g2_buf_1 _16671_ (.A(_07931_),
    .X(_07932_));
 sg13g2_xnor2_1 _16672_ (.Y(_07933_),
    .A(net260),
    .B(_07932_));
 sg13g2_nand2_1 _16673_ (.Y(_07934_),
    .A(_07382_),
    .B(_07933_));
 sg13g2_xnor2_1 _16674_ (.Y(_07935_),
    .A(_02453_),
    .B(_07934_));
 sg13g2_nor2_1 _16675_ (.A(_07829_),
    .B(_07935_),
    .Y(_01008_));
 sg13g2_o21ai_1 _16676_ (.B1(_07750_),
    .Y(_07936_),
    .A1(_02453_),
    .A2(_07932_));
 sg13g2_nand2_1 _16677_ (.Y(_07937_),
    .A(_02453_),
    .B(_07932_));
 sg13g2_nand2_1 _16678_ (.Y(_07938_),
    .A(_07936_),
    .B(_07937_));
 sg13g2_xnor2_1 _16679_ (.Y(_07939_),
    .A(_07756_),
    .B(_07938_));
 sg13g2_nand2_1 _16680_ (.Y(_07940_),
    .A(_07382_),
    .B(_07939_));
 sg13g2_xnor2_1 _16681_ (.Y(_07941_),
    .A(_02457_),
    .B(_07940_));
 sg13g2_nor2_1 _16682_ (.A(net51),
    .B(_07941_),
    .Y(_01009_));
 sg13g2_buf_1 _16683_ (.A(_07530_),
    .X(_07942_));
 sg13g2_a21oi_1 _16684_ (.A1(_02453_),
    .A2(_07932_),
    .Y(_07943_),
    .B1(_02457_));
 sg13g2_nor2_1 _16685_ (.A(\am_sdr0.cic3.integ3[16] ),
    .B(_02456_),
    .Y(_07944_));
 sg13g2_nor2_1 _16686_ (.A(_07747_),
    .B(_02456_),
    .Y(_07945_));
 sg13g2_o21ai_1 _16687_ (.B1(_07932_),
    .Y(_07946_),
    .A1(_07944_),
    .A2(_07945_));
 sg13g2_nor3_1 _16688_ (.A(_07747_),
    .B(\am_sdr0.cic3.integ3[16] ),
    .C(_02456_),
    .Y(_07947_));
 sg13g2_nor2b_1 _16689_ (.A(_07947_),
    .B_N(_07756_),
    .Y(_07948_));
 sg13g2_a22oi_1 _16690_ (.Y(_07949_),
    .B1(_07946_),
    .B2(_07948_),
    .A2(_07943_),
    .A1(_07936_));
 sg13g2_xnor2_1 _16691_ (.Y(_07950_),
    .A(_07784_),
    .B(_07949_));
 sg13g2_nand2_1 _16692_ (.Y(_07951_),
    .A(_07366_),
    .B(_07950_));
 sg13g2_xor2_1 _16693_ (.B(_07951_),
    .A(_02460_),
    .X(_07952_));
 sg13g2_nor2_1 _16694_ (.A(_07942_),
    .B(_07952_),
    .Y(_01010_));
 sg13g2_and2_1 _16695_ (.A(_02808_),
    .B(\am_sdr0.cic3.integ3[19] ),
    .X(_07953_));
 sg13g2_nor2_1 _16696_ (.A(_01968_),
    .B(\am_sdr0.cic3.integ3[19] ),
    .Y(_07954_));
 sg13g2_or2_1 _16697_ (.X(_07955_),
    .B(_02460_),
    .A(_07784_));
 sg13g2_o21ai_1 _16698_ (.B1(_07955_),
    .Y(_07956_),
    .A1(_07756_),
    .A2(_02456_));
 sg13g2_a22oi_1 _16699_ (.Y(_07957_),
    .B1(_07936_),
    .B2(_07937_),
    .A2(_02456_),
    .A1(_07756_));
 sg13g2_nand2_1 _16700_ (.Y(_07958_),
    .A(_07784_),
    .B(_02460_));
 sg13g2_o21ai_1 _16701_ (.B1(_07958_),
    .Y(_07959_),
    .A1(_07956_),
    .A2(_07957_));
 sg13g2_xnor2_1 _16702_ (.Y(_07960_),
    .A(\am_sdr0.cic3.integ2[22] ),
    .B(_07959_));
 sg13g2_nor2_1 _16703_ (.A(net145),
    .B(_07960_),
    .Y(_07961_));
 sg13g2_mux2_1 _16704_ (.A0(_07953_),
    .A1(_07954_),
    .S(_07961_),
    .X(_01011_));
 sg13g2_nand2_1 _16705_ (.Y(_07962_),
    .A(_07617_),
    .B(_02420_));
 sg13g2_xnor2_1 _16706_ (.Y(_07963_),
    .A(_07614_),
    .B(_07962_));
 sg13g2_nand2_1 _16707_ (.Y(_07964_),
    .A(net198),
    .B(_07963_));
 sg13g2_xor2_1 _16708_ (.B(_07964_),
    .A(_02462_),
    .X(_07965_));
 sg13g2_nor2_1 _16709_ (.A(net50),
    .B(_07965_),
    .Y(_01012_));
 sg13g2_nor2_1 _16710_ (.A(_07841_),
    .B(_07842_),
    .Y(_07966_));
 sg13g2_xor2_1 _16711_ (.B(_07966_),
    .A(_07612_),
    .X(_07967_));
 sg13g2_nand2_1 _16712_ (.Y(_07968_),
    .A(net198),
    .B(_07967_));
 sg13g2_xor2_1 _16713_ (.B(_07968_),
    .A(_02465_),
    .X(_07969_));
 sg13g2_nor2_1 _16714_ (.A(net50),
    .B(_07969_),
    .Y(_01013_));
 sg13g2_nand2_1 _16715_ (.Y(_07970_),
    .A(_07839_),
    .B(_07844_));
 sg13g2_xnor2_1 _16716_ (.Y(_07971_),
    .A(_07630_),
    .B(_07970_));
 sg13g2_nor2_1 _16717_ (.A(net144),
    .B(_07971_),
    .Y(_07972_));
 sg13g2_xnor2_1 _16718_ (.Y(_07973_),
    .A(\am_sdr0.cic3.integ3[3] ),
    .B(_07972_));
 sg13g2_nor2_1 _16719_ (.A(net50),
    .B(_07973_),
    .Y(_01014_));
 sg13g2_a21oi_1 _16720_ (.A1(_07630_),
    .A2(_07845_),
    .Y(_07974_),
    .B1(_07846_));
 sg13g2_xnor2_1 _16721_ (.Y(_07975_),
    .A(_07610_),
    .B(_07974_));
 sg13g2_nand2_1 _16722_ (.Y(_07976_),
    .A(net198),
    .B(_07975_));
 sg13g2_xor2_1 _16723_ (.B(_07976_),
    .A(_02470_),
    .X(_07977_));
 sg13g2_nor2_1 _16724_ (.A(net50),
    .B(_07977_),
    .Y(_01015_));
 sg13g2_nor2_1 _16725_ (.A(_07848_),
    .B(_07849_),
    .Y(_07978_));
 sg13g2_xnor2_1 _16726_ (.Y(_07979_),
    .A(_07635_),
    .B(_07978_));
 sg13g2_nor2_1 _16727_ (.A(_07449_),
    .B(_07979_),
    .Y(_07980_));
 sg13g2_xnor2_1 _16728_ (.Y(_07981_),
    .A(\am_sdr0.cic3.integ3[5] ),
    .B(_07980_));
 sg13g2_nor2_1 _16729_ (.A(net50),
    .B(_07981_),
    .Y(_01016_));
 sg13g2_xnor2_1 _16730_ (.Y(_07982_),
    .A(_07608_),
    .B(_07852_));
 sg13g2_nand2_1 _16731_ (.Y(_07983_),
    .A(net198),
    .B(_07982_));
 sg13g2_xor2_1 _16732_ (.B(_07983_),
    .A(_02475_),
    .X(_07984_));
 sg13g2_nor2_1 _16733_ (.A(net50),
    .B(_07984_),
    .Y(_01017_));
 sg13g2_xnor2_1 _16734_ (.Y(_07985_),
    .A(_07607_),
    .B(_07856_));
 sg13g2_nor2_1 _16735_ (.A(_07449_),
    .B(_07985_),
    .Y(_07986_));
 sg13g2_xnor2_1 _16736_ (.Y(_07987_),
    .A(_02477_),
    .B(_07986_));
 sg13g2_nor2_1 _16737_ (.A(net50),
    .B(_07987_),
    .Y(_01018_));
 sg13g2_xnor2_1 _16738_ (.Y(_07988_),
    .A(_07646_),
    .B(_07859_));
 sg13g2_nor2_1 _16739_ (.A(_07449_),
    .B(_07988_),
    .Y(_07989_));
 sg13g2_xnor2_1 _16740_ (.Y(_07990_),
    .A(_02481_),
    .B(_07989_));
 sg13g2_nor2_1 _16741_ (.A(net50),
    .B(_07990_),
    .Y(_01019_));
 sg13g2_xnor2_1 _16742_ (.Y(_07991_),
    .A(_07653_),
    .B(_07861_));
 sg13g2_nand2_1 _16743_ (.Y(_07992_),
    .A(net198),
    .B(_07991_));
 sg13g2_xor2_1 _16744_ (.B(_07992_),
    .A(_02485_),
    .X(_07993_));
 sg13g2_nor2_1 _16745_ (.A(_07942_),
    .B(_07993_),
    .Y(_01020_));
 sg13g2_nand2_1 _16746_ (.Y(_07994_),
    .A(net209),
    .B(\am_sdr0.cic3.comb3[14] ));
 sg13g2_nand2_1 _16747_ (.Y(_07995_),
    .A(\am_sdr0.am0.Q_in[2] ),
    .B(net146));
 sg13g2_a21oi_1 _16748_ (.A1(_07994_),
    .A2(_07995_),
    .Y(_01042_),
    .B1(net56));
 sg13g2_nand2_1 _16749_ (.Y(_07996_),
    .A(_06664_),
    .B(\am_sdr0.cic3.comb3[15] ));
 sg13g2_nand2_1 _16750_ (.Y(_07997_),
    .A(\am_sdr0.am0.Q_in[3] ),
    .B(net146));
 sg13g2_a21oi_1 _16751_ (.A1(_07996_),
    .A2(_07997_),
    .Y(_01043_),
    .B1(net56));
 sg13g2_nand2_1 _16752_ (.Y(_07998_),
    .A(_06664_),
    .B(\am_sdr0.cic3.comb3[16] ));
 sg13g2_nand2_1 _16753_ (.Y(_07999_),
    .A(\am_sdr0.am0.Q_in[4] ),
    .B(net146));
 sg13g2_a21oi_1 _16754_ (.A1(_07998_),
    .A2(_07999_),
    .Y(_01044_),
    .B1(net56));
 sg13g2_nand2_1 _16755_ (.Y(_08000_),
    .A(net206),
    .B(\am_sdr0.cic3.comb3[17] ));
 sg13g2_nand2_1 _16756_ (.Y(_08001_),
    .A(\am_sdr0.am0.Q_in[5] ),
    .B(net146));
 sg13g2_a21oi_1 _16757_ (.A1(_08000_),
    .A2(_08001_),
    .Y(_01045_),
    .B1(net56));
 sg13g2_nand2_1 _16758_ (.Y(_08002_),
    .A(net206),
    .B(\am_sdr0.cic3.comb3[18] ));
 sg13g2_nand2_1 _16759_ (.Y(_08003_),
    .A(\am_sdr0.am0.Q_in[6] ),
    .B(net146));
 sg13g2_buf_1 _16760_ (.A(_07113_),
    .X(_08004_));
 sg13g2_a21oi_1 _16761_ (.A1(_08002_),
    .A2(_08003_),
    .Y(_01046_),
    .B1(net49));
 sg13g2_nand2_1 _16762_ (.Y(_08005_),
    .A(net206),
    .B(\am_sdr0.cic3.comb3[19] ));
 sg13g2_nand2_1 _16763_ (.Y(_08006_),
    .A(\am_sdr0.am0.Q_in[7] ),
    .B(net146));
 sg13g2_a21oi_1 _16764_ (.A1(_08005_),
    .A2(_08006_),
    .Y(_01047_),
    .B1(net49));
 sg13g2_nand2_1 _16765_ (.Y(_08007_),
    .A(net206),
    .B(\am_sdr0.cic3.comb3[12] ));
 sg13g2_nand2_1 _16766_ (.Y(_08008_),
    .A(\am_sdr0.am0.Q_in[0] ),
    .B(net149));
 sg13g2_a21oi_1 _16767_ (.A1(_08007_),
    .A2(_08008_),
    .Y(_01048_),
    .B1(_08004_));
 sg13g2_nand2_1 _16768_ (.Y(_08009_),
    .A(net206),
    .B(\am_sdr0.cic3.comb3[13] ));
 sg13g2_nand2_1 _16769_ (.Y(_08010_),
    .A(\am_sdr0.am0.Q_in[1] ),
    .B(net149));
 sg13g2_a21oi_1 _16770_ (.A1(_08009_),
    .A2(_08010_),
    .Y(_01049_),
    .B1(_08004_));
 sg13g2_and2_1 _16771_ (.A(net210),
    .B(_00068_),
    .X(_01050_));
 sg13g2_buf_1 _16772_ (.A(_07530_),
    .X(_08011_));
 sg13g2_xnor2_1 _16773_ (.Y(_08012_),
    .A(_02626_),
    .B(_02666_));
 sg13g2_nor2_1 _16774_ (.A(net48),
    .B(_08012_),
    .Y(_01051_));
 sg13g2_nand2_1 _16775_ (.Y(_08013_),
    .A(_02626_),
    .B(_02666_));
 sg13g2_xnor2_1 _16776_ (.Y(_08014_),
    .A(_02665_),
    .B(_08013_));
 sg13g2_nor2_1 _16777_ (.A(net48),
    .B(_08014_),
    .Y(_01052_));
 sg13g2_nand3_1 _16778_ (.B(_02626_),
    .C(_02666_),
    .A(_02601_),
    .Y(_08015_));
 sg13g2_xnor2_1 _16779_ (.Y(_08016_),
    .A(_02605_),
    .B(_08015_));
 sg13g2_nor2_1 _16780_ (.A(net48),
    .B(_08016_),
    .Y(_01053_));
 sg13g2_nor2_1 _16781_ (.A(_02605_),
    .B(_08015_),
    .Y(_08017_));
 sg13g2_xnor2_1 _16782_ (.Y(_08018_),
    .A(net298),
    .B(_08017_));
 sg13g2_nor2_1 _16783_ (.A(net48),
    .B(_08018_),
    .Y(_01054_));
 sg13g2_nand2_1 _16784_ (.Y(_08019_),
    .A(net298),
    .B(_08017_));
 sg13g2_xnor2_1 _16785_ (.Y(_08020_),
    .A(_02625_),
    .B(_08019_));
 sg13g2_nor2_1 _16786_ (.A(_08011_),
    .B(_08020_),
    .Y(_01055_));
 sg13g2_nand3_1 _16787_ (.B(net298),
    .C(_08017_),
    .A(_02611_),
    .Y(_08021_));
 sg13g2_xnor2_1 _16788_ (.Y(_08022_),
    .A(_02593_),
    .B(_08021_));
 sg13g2_nor2_1 _16789_ (.A(_08011_),
    .B(_08022_),
    .Y(_01056_));
 sg13g2_or2_1 _16790_ (.X(_08023_),
    .B(_08021_),
    .A(_02593_));
 sg13g2_xnor2_1 _16791_ (.Y(_08024_),
    .A(_02617_),
    .B(_08023_));
 sg13g2_nor2_1 _16792_ (.A(net48),
    .B(_08024_),
    .Y(_01057_));
 sg13g2_and2_1 _16793_ (.A(net210),
    .B(net1),
    .X(_01058_));
 sg13g2_and2_1 _16794_ (.A(net210),
    .B(\am_sdr0.mix0.RF_in_q ),
    .X(_01059_));
 sg13g2_and2_1 _16795_ (.A(net210),
    .B(_01469_),
    .X(_01060_));
 sg13g2_and2_1 _16796_ (.A(net210),
    .B(\am_sdr0.cos[0] ),
    .X(_01061_));
 sg13g2_buf_1 _16797_ (.A(net297),
    .X(_08025_));
 sg13g2_and2_1 _16798_ (.A(net194),
    .B(\am_sdr0.cos[1] ),
    .X(_01062_));
 sg13g2_and2_1 _16799_ (.A(net194),
    .B(\am_sdr0.cos[2] ),
    .X(_01063_));
 sg13g2_and2_1 _16800_ (.A(net194),
    .B(\am_sdr0.cos[3] ),
    .X(_01064_));
 sg13g2_and2_1 _16801_ (.A(net194),
    .B(\am_sdr0.cos[4] ),
    .X(_01065_));
 sg13g2_and2_1 _16802_ (.A(net194),
    .B(\am_sdr0.cos[5] ),
    .X(_01066_));
 sg13g2_and2_1 _16803_ (.A(net194),
    .B(\am_sdr0.cos[6] ),
    .X(_01067_));
 sg13g2_and2_1 _16804_ (.A(net194),
    .B(\am_sdr0.cos[7] ),
    .X(_01068_));
 sg13g2_and2_1 _16805_ (.A(net194),
    .B(\am_sdr0.mix0.sin_in[0] ),
    .X(_01069_));
 sg13g2_and2_1 _16806_ (.A(_08025_),
    .B(\am_sdr0.mix0.sin_in[1] ),
    .X(_01070_));
 sg13g2_and2_1 _16807_ (.A(_08025_),
    .B(\am_sdr0.mix0.sin_in[2] ),
    .X(_01071_));
 sg13g2_buf_1 _16808_ (.A(net297),
    .X(_08026_));
 sg13g2_and2_1 _16809_ (.A(net193),
    .B(\am_sdr0.mix0.sin_in[3] ),
    .X(_01072_));
 sg13g2_and2_1 _16810_ (.A(net193),
    .B(\am_sdr0.mix0.sin_in[4] ),
    .X(_01073_));
 sg13g2_and2_1 _16811_ (.A(net193),
    .B(\am_sdr0.mix0.sin_in[5] ),
    .X(_01074_));
 sg13g2_and2_1 _16812_ (.A(net193),
    .B(\am_sdr0.mix0.sin_in[6] ),
    .X(_01075_));
 sg13g2_and2_1 _16813_ (.A(net193),
    .B(\am_sdr0.mix0.sin_in[7] ),
    .X(_01076_));
 sg13g2_xnor2_1 _16814_ (.Y(_08027_),
    .A(\am_sdr0.nco0.phase[0] ),
    .B(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_nor2_1 _16815_ (.A(net48),
    .B(_08027_),
    .Y(_01077_));
 sg13g2_buf_2 _16816_ (.A(\am_sdr0.nco0.phase[9] ),
    .X(_08028_));
 sg13g2_buf_1 _16817_ (.A(\am_sdr0.nco0.phase_inc[9] ),
    .X(_08029_));
 sg13g2_buf_1 _16818_ (.A(\am_sdr0.nco0.phase[7] ),
    .X(_08030_));
 sg13g2_inv_1 _16819_ (.Y(_08031_),
    .A(_08030_));
 sg13g2_buf_1 _16820_ (.A(\am_sdr0.nco0.phase_inc[7] ),
    .X(_08032_));
 sg13g2_inv_1 _16821_ (.Y(_08033_),
    .A(_08032_));
 sg13g2_buf_1 _16822_ (.A(\am_sdr0.nco0.phase_inc[5] ),
    .X(_08034_));
 sg13g2_buf_1 _16823_ (.A(\am_sdr0.nco0.phase[3] ),
    .X(_08035_));
 sg13g2_buf_1 _16824_ (.A(\am_sdr0.nco0.phase_inc[3] ),
    .X(_08036_));
 sg13g2_buf_1 _16825_ (.A(\am_sdr0.nco0.phase_inc[2] ),
    .X(_08037_));
 sg13g2_or2_1 _16826_ (.X(_08038_),
    .B(_08037_),
    .A(\am_sdr0.nco0.phase[2] ));
 sg13g2_buf_1 _16827_ (.A(\am_sdr0.nco0.phase_inc[1] ),
    .X(_08039_));
 sg13g2_nor2_1 _16828_ (.A(\am_sdr0.nco0.phase[1] ),
    .B(_08039_),
    .Y(_08040_));
 sg13g2_nand2_1 _16829_ (.Y(_08041_),
    .A(\am_sdr0.nco0.phase[0] ),
    .B(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_nand2_1 _16830_ (.Y(_08042_),
    .A(\am_sdr0.nco0.phase[1] ),
    .B(_08039_));
 sg13g2_o21ai_1 _16831_ (.B1(_08042_),
    .Y(_08043_),
    .A1(_08040_),
    .A2(_08041_));
 sg13g2_buf_1 _16832_ (.A(_08043_),
    .X(_08044_));
 sg13g2_and2_1 _16833_ (.A(\am_sdr0.nco0.phase[2] ),
    .B(_08037_),
    .X(_08045_));
 sg13g2_a221oi_1 _16834_ (.B2(_08044_),
    .C1(_08045_),
    .B1(_08038_),
    .A1(_08035_),
    .Y(_08046_),
    .A2(_08036_));
 sg13g2_or2_1 _16835_ (.X(_08047_),
    .B(\am_sdr0.nco0.phase_inc[4] ),
    .A(\am_sdr0.nco0.phase[4] ));
 sg13g2_o21ai_1 _16836_ (.B1(_08047_),
    .Y(_08048_),
    .A1(_08035_),
    .A2(_08036_));
 sg13g2_nand2_1 _16837_ (.Y(_08049_),
    .A(\am_sdr0.nco0.phase[4] ),
    .B(\am_sdr0.nco0.phase_inc[4] ));
 sg13g2_o21ai_1 _16838_ (.B1(_08049_),
    .Y(_08050_),
    .A1(_08046_),
    .A2(_08048_));
 sg13g2_buf_1 _16839_ (.A(_08050_),
    .X(_08051_));
 sg13g2_nor2_1 _16840_ (.A(_08034_),
    .B(_08051_),
    .Y(_08052_));
 sg13g2_a21oi_1 _16841_ (.A1(_08034_),
    .A2(_08051_),
    .Y(_08053_),
    .B1(\am_sdr0.nco0.phase[5] ));
 sg13g2_buf_1 _16842_ (.A(\am_sdr0.nco0.phase[6] ),
    .X(_08054_));
 sg13g2_buf_1 _16843_ (.A(\am_sdr0.nco0.phase_inc[6] ),
    .X(_08055_));
 sg13g2_nor2_1 _16844_ (.A(_08054_),
    .B(_08055_),
    .Y(_08056_));
 sg13g2_or3_1 _16845_ (.A(_08052_),
    .B(_08053_),
    .C(_08056_),
    .X(_08057_));
 sg13g2_buf_1 _16846_ (.A(_08057_),
    .X(_08058_));
 sg13g2_a22oi_1 _16847_ (.Y(_08059_),
    .B1(_08030_),
    .B2(_08032_),
    .A2(_08055_),
    .A1(_08054_));
 sg13g2_buf_1 _16848_ (.A(\am_sdr0.nco0.phase_inc[8] ),
    .X(_08060_));
 sg13g2_inv_1 _16849_ (.Y(_01172_),
    .A(_08060_));
 sg13g2_a221oi_1 _16850_ (.B2(_08059_),
    .C1(_01172_),
    .B1(_08058_),
    .A1(_08031_),
    .Y(_01173_),
    .A2(_08033_));
 sg13g2_a22oi_1 _16851_ (.Y(_01174_),
    .B1(_08058_),
    .B2(_08059_),
    .A2(_08033_),
    .A1(_08031_));
 sg13g2_buf_1 _16852_ (.A(_01174_),
    .X(_01175_));
 sg13g2_buf_1 _16853_ (.A(\am_sdr0.nco0.phase[8] ),
    .X(_01176_));
 sg13g2_o21ai_1 _16854_ (.B1(_01176_),
    .Y(_01177_),
    .A1(_08060_),
    .A2(_01175_));
 sg13g2_nand2b_1 _16855_ (.Y(_01178_),
    .B(_01177_),
    .A_N(_01173_));
 sg13g2_o21ai_1 _16856_ (.B1(_01178_),
    .Y(_01179_),
    .A1(_08028_),
    .A2(_08029_));
 sg13g2_nand2_1 _16857_ (.Y(_01180_),
    .A(_08028_),
    .B(_08029_));
 sg13g2_buf_1 _16858_ (.A(\am_sdr0.nco0.phase[10] ),
    .X(_01181_));
 sg13g2_buf_1 _16859_ (.A(\am_sdr0.nco0.phase_inc[10] ),
    .X(_01182_));
 sg13g2_xor2_1 _16860_ (.B(_01182_),
    .A(_01181_),
    .X(_01183_));
 sg13g2_a21o_1 _16861_ (.A2(_01180_),
    .A1(_01179_),
    .B1(_01183_),
    .X(_01184_));
 sg13g2_nand3_1 _16862_ (.B(_01179_),
    .C(_01180_),
    .A(_01183_),
    .Y(_01185_));
 sg13g2_a21oi_1 _16863_ (.A1(_01184_),
    .A2(_01185_),
    .Y(_01078_),
    .B1(net49));
 sg13g2_o21ai_1 _16864_ (.B1(_08029_),
    .Y(_01186_),
    .A1(_01181_),
    .A2(_01182_));
 sg13g2_inv_1 _16865_ (.Y(_01187_),
    .A(_01186_));
 sg13g2_o21ai_1 _16866_ (.B1(_01176_),
    .Y(_01188_),
    .A1(_08030_),
    .A2(_08032_));
 sg13g2_a21o_1 _16867_ (.A2(_08059_),
    .A1(_08058_),
    .B1(_01188_),
    .X(_01189_));
 sg13g2_a21oi_1 _16868_ (.A1(_01176_),
    .A2(_08060_),
    .Y(_01190_),
    .B1(_08028_));
 sg13g2_nand2_1 _16869_ (.Y(_01191_),
    .A(_01189_),
    .B(_01190_));
 sg13g2_and2_1 _16870_ (.A(_08028_),
    .B(_01182_),
    .X(_01192_));
 sg13g2_inv_1 _16871_ (.Y(_01193_),
    .A(_01176_));
 sg13g2_o21ai_1 _16872_ (.B1(_08028_),
    .Y(_01194_),
    .A1(_01181_),
    .A2(_01182_));
 sg13g2_nor2_1 _16873_ (.A(_01193_),
    .B(_01194_),
    .Y(_01195_));
 sg13g2_a21o_1 _16874_ (.A2(_01192_),
    .A1(_01175_),
    .B1(_01195_),
    .X(_01196_));
 sg13g2_nand2_1 _16875_ (.Y(_01197_),
    .A(_01172_),
    .B(_01189_));
 sg13g2_a21o_1 _16876_ (.A2(_01181_),
    .A1(_08028_),
    .B1(_01187_),
    .X(_01198_));
 sg13g2_and2_1 _16877_ (.A(_01181_),
    .B(_01182_),
    .X(_01199_));
 sg13g2_a21o_1 _16878_ (.A2(_01198_),
    .A1(_01173_),
    .B1(_01199_),
    .X(_01200_));
 sg13g2_a221oi_1 _16879_ (.B2(_01197_),
    .C1(_01200_),
    .B1(_01196_),
    .A1(_01187_),
    .Y(_01201_),
    .A2(_01191_));
 sg13g2_buf_1 _16880_ (.A(_01201_),
    .X(_01202_));
 sg13g2_buf_1 _16881_ (.A(\am_sdr0.nco0.phase[11] ),
    .X(_01203_));
 sg13g2_buf_1 _16882_ (.A(\am_sdr0.nco0.phase_inc[11] ),
    .X(_01204_));
 sg13g2_xnor2_1 _16883_ (.Y(_01205_),
    .A(_01203_),
    .B(_01204_));
 sg13g2_xnor2_1 _16884_ (.Y(_01206_),
    .A(_01202_),
    .B(_01205_));
 sg13g2_nor2_1 _16885_ (.A(net48),
    .B(_01206_),
    .Y(_01079_));
 sg13g2_nand2b_1 _16886_ (.Y(_01207_),
    .B(_01202_),
    .A_N(_01204_));
 sg13g2_nor2b_1 _16887_ (.A(_01202_),
    .B_N(_01204_),
    .Y(_01208_));
 sg13g2_a21o_1 _16888_ (.A2(_01207_),
    .A1(_01203_),
    .B1(_01208_),
    .X(_01209_));
 sg13g2_buf_1 _16889_ (.A(\am_sdr0.nco0.phase[12] ),
    .X(_01210_));
 sg13g2_buf_1 _16890_ (.A(\am_sdr0.nco0.phase_inc[12] ),
    .X(_01211_));
 sg13g2_xor2_1 _16891_ (.B(_01211_),
    .A(_01210_),
    .X(_01212_));
 sg13g2_xnor2_1 _16892_ (.Y(_01213_),
    .A(_01209_),
    .B(_01212_));
 sg13g2_nor2_1 _16893_ (.A(net48),
    .B(_01213_),
    .Y(_01080_));
 sg13g2_buf_1 _16894_ (.A(_07530_),
    .X(_01214_));
 sg13g2_buf_1 _16895_ (.A(\am_sdr0.nco0.phase[13] ),
    .X(_01215_));
 sg13g2_buf_1 _16896_ (.A(\am_sdr0.nco0.phase_inc[13] ),
    .X(_01216_));
 sg13g2_xnor2_1 _16897_ (.Y(_01217_),
    .A(_01215_),
    .B(_01216_));
 sg13g2_or2_1 _16898_ (.X(_01218_),
    .B(_01211_),
    .A(_01210_));
 sg13g2_and2_1 _16899_ (.A(_01210_),
    .B(_01211_),
    .X(_01219_));
 sg13g2_a21oi_1 _16900_ (.A1(_01209_),
    .A2(_01218_),
    .Y(_01220_),
    .B1(_01219_));
 sg13g2_xnor2_1 _16901_ (.Y(_01221_),
    .A(_01217_),
    .B(_01220_));
 sg13g2_nor2_1 _16902_ (.A(net47),
    .B(_01221_),
    .Y(_01081_));
 sg13g2_nor2_1 _16903_ (.A(_01215_),
    .B(_01216_),
    .Y(_01222_));
 sg13g2_nand2_1 _16904_ (.Y(_01223_),
    .A(_01215_),
    .B(_01216_));
 sg13g2_o21ai_1 _16905_ (.B1(_01223_),
    .Y(_01224_),
    .A1(_01222_),
    .A2(_01220_));
 sg13g2_buf_1 _16906_ (.A(\am_sdr0.nco0.phase[14] ),
    .X(_01225_));
 sg13g2_buf_1 _16907_ (.A(\am_sdr0.nco0.phase_inc[14] ),
    .X(_01226_));
 sg13g2_xor2_1 _16908_ (.B(_01226_),
    .A(_01225_),
    .X(_01227_));
 sg13g2_xnor2_1 _16909_ (.Y(_01228_),
    .A(_01224_),
    .B(_01227_));
 sg13g2_nor2_1 _16910_ (.A(net47),
    .B(_01228_),
    .Y(_01082_));
 sg13g2_nand2_1 _16911_ (.Y(_01229_),
    .A(_01210_),
    .B(_01211_));
 sg13g2_nand2_1 _16912_ (.Y(_01230_),
    .A(_01203_),
    .B(_01204_));
 sg13g2_nand3_1 _16913_ (.B(_01229_),
    .C(_01230_),
    .A(_01223_),
    .Y(_01231_));
 sg13g2_nor2_1 _16914_ (.A(_01226_),
    .B(_01231_),
    .Y(_01232_));
 sg13g2_nor2_1 _16915_ (.A(_01225_),
    .B(_01231_),
    .Y(_01233_));
 sg13g2_o21ai_1 _16916_ (.B1(_01202_),
    .Y(_01234_),
    .A1(_01232_),
    .A2(_01233_));
 sg13g2_o21ai_1 _16917_ (.B1(_01218_),
    .Y(_01235_),
    .A1(_01203_),
    .A2(_01204_));
 sg13g2_a21oi_1 _16918_ (.A1(_01229_),
    .A2(_01235_),
    .Y(_01236_),
    .B1(_01222_));
 sg13g2_a221oi_1 _16919_ (.B2(_01226_),
    .C1(_01236_),
    .B1(_01225_),
    .A1(_01215_),
    .Y(_01237_),
    .A2(_01216_));
 sg13g2_nor2_1 _16920_ (.A(_01225_),
    .B(_01226_),
    .Y(_01238_));
 sg13g2_nor2_1 _16921_ (.A(_01237_),
    .B(_01238_),
    .Y(_01239_));
 sg13g2_nand2_2 _16922_ (.Y(_01240_),
    .A(_01234_),
    .B(_01239_));
 sg13g2_buf_1 _16923_ (.A(\am_sdr0.nco0.phase[15] ),
    .X(_01241_));
 sg13g2_buf_1 _16924_ (.A(\am_sdr0.nco0.phase_inc[15] ),
    .X(_01242_));
 sg13g2_xnor2_1 _16925_ (.Y(_01243_),
    .A(_01241_),
    .B(_01242_));
 sg13g2_xnor2_1 _16926_ (.Y(_01244_),
    .A(_01240_),
    .B(_01243_));
 sg13g2_nor2_1 _16927_ (.A(net47),
    .B(_01244_),
    .Y(_01083_));
 sg13g2_buf_1 _16928_ (.A(\am_sdr0.nco0.phase[16] ),
    .X(_01245_));
 sg13g2_buf_1 _16929_ (.A(\am_sdr0.nco0.phase_inc[16] ),
    .X(_01246_));
 sg13g2_xnor2_1 _16930_ (.Y(_01247_),
    .A(_01245_),
    .B(_01246_));
 sg13g2_nand2_1 _16931_ (.Y(_01248_),
    .A(_01241_),
    .B(_01242_));
 sg13g2_nor2_1 _16932_ (.A(_01241_),
    .B(_01242_),
    .Y(_01249_));
 sg13g2_nand3b_1 _16933_ (.B(_01239_),
    .C(_01234_),
    .Y(_01250_),
    .A_N(_01249_));
 sg13g2_nand2_1 _16934_ (.Y(_01251_),
    .A(_01248_),
    .B(_01250_));
 sg13g2_xor2_1 _16935_ (.B(_01251_),
    .A(_01247_),
    .X(_01252_));
 sg13g2_nor2_1 _16936_ (.A(_01214_),
    .B(_01252_),
    .Y(_01084_));
 sg13g2_buf_1 _16937_ (.A(\am_sdr0.nco0.phase[17] ),
    .X(_01253_));
 sg13g2_buf_2 _16938_ (.A(\am_sdr0.nco0.phase_inc[17] ),
    .X(_01254_));
 sg13g2_xor2_1 _16939_ (.B(_01254_),
    .A(_01253_),
    .X(_01255_));
 sg13g2_or2_1 _16940_ (.X(_01256_),
    .B(_01246_),
    .A(_01245_));
 sg13g2_nand2_1 _16941_ (.Y(_01257_),
    .A(_01245_),
    .B(_01246_));
 sg13g2_nand3_1 _16942_ (.B(_01250_),
    .C(_01257_),
    .A(_01248_),
    .Y(_01258_));
 sg13g2_nand2_1 _16943_ (.Y(_01259_),
    .A(_01256_),
    .B(_01258_));
 sg13g2_xor2_1 _16944_ (.B(_01259_),
    .A(_01255_),
    .X(_01260_));
 sg13g2_nor2_1 _16945_ (.A(net47),
    .B(_01260_),
    .Y(_01085_));
 sg13g2_a221oi_1 _16946_ (.B2(_01246_),
    .C1(_01254_),
    .B1(_01245_),
    .A1(_01241_),
    .Y(_01261_),
    .A2(_01242_));
 sg13g2_nor2_1 _16947_ (.A(_01245_),
    .B(_01246_),
    .Y(_01262_));
 sg13g2_a21oi_1 _16948_ (.A1(_01249_),
    .A2(_01257_),
    .Y(_01263_),
    .B1(_01262_));
 sg13g2_o21ai_1 _16949_ (.B1(_01253_),
    .Y(_01264_),
    .A1(_01254_),
    .A2(_01263_));
 sg13g2_a21oi_1 _16950_ (.A1(_01240_),
    .A2(_01261_),
    .Y(_01265_),
    .B1(_01264_));
 sg13g2_nand3_1 _16951_ (.B(_01256_),
    .C(_01258_),
    .A(_01254_),
    .Y(_01266_));
 sg13g2_nor2b_1 _16952_ (.A(_01265_),
    .B_N(_01266_),
    .Y(_01267_));
 sg13g2_buf_1 _16953_ (.A(\am_sdr0.nco0.phase[18] ),
    .X(_01268_));
 sg13g2_buf_2 _16954_ (.A(\am_sdr0.nco0.phase_inc[18] ),
    .X(_01269_));
 sg13g2_xnor2_1 _16955_ (.Y(_01270_),
    .A(_01268_),
    .B(_01269_));
 sg13g2_xnor2_1 _16956_ (.Y(_01271_),
    .A(_01267_),
    .B(_01270_));
 sg13g2_nor2_1 _16957_ (.A(net47),
    .B(_01271_),
    .Y(_01086_));
 sg13g2_buf_1 _16958_ (.A(\am_sdr0.nco0.phase_inc[19] ),
    .X(_01272_));
 sg13g2_xnor2_1 _16959_ (.Y(_01273_),
    .A(\am_sdr0.nco0.phase[19] ),
    .B(_01272_));
 sg13g2_a21oi_1 _16960_ (.A1(_01268_),
    .A2(_01269_),
    .Y(_01274_),
    .B1(_01265_));
 sg13g2_nor2_1 _16961_ (.A(_01268_),
    .B(_01269_),
    .Y(_01275_));
 sg13g2_a21oi_1 _16962_ (.A1(_01266_),
    .A2(_01274_),
    .Y(_01276_),
    .B1(_01275_));
 sg13g2_xor2_1 _16963_ (.B(_01276_),
    .A(_01273_),
    .X(_01277_));
 sg13g2_nor2_1 _16964_ (.A(net47),
    .B(_01277_),
    .Y(_01087_));
 sg13g2_xnor2_1 _16965_ (.Y(_01278_),
    .A(\am_sdr0.nco0.phase[1] ),
    .B(_08039_));
 sg13g2_xnor2_1 _16966_ (.Y(_01279_),
    .A(_08041_),
    .B(_01278_));
 sg13g2_nor2_1 _16967_ (.A(_01214_),
    .B(_01279_),
    .Y(_01088_));
 sg13g2_nor2_1 _16968_ (.A(_01270_),
    .B(_01273_),
    .Y(_01280_));
 sg13g2_nand2_1 _16969_ (.Y(_01281_),
    .A(_01255_),
    .B(_01280_));
 sg13g2_nor2_1 _16970_ (.A(_01247_),
    .B(_01281_),
    .Y(_01282_));
 sg13g2_nor2_1 _16971_ (.A(\am_sdr0.nco0.phase[19] ),
    .B(_01272_),
    .Y(_01283_));
 sg13g2_nand2_1 _16972_ (.Y(_01284_),
    .A(_01253_),
    .B(_01254_));
 sg13g2_nor2_1 _16973_ (.A(_01253_),
    .B(_01254_),
    .Y(_01285_));
 sg13g2_a21oi_1 _16974_ (.A1(_01257_),
    .A2(_01284_),
    .Y(_01286_),
    .B1(_01285_));
 sg13g2_a21o_1 _16975_ (.A2(_01286_),
    .A1(_01269_),
    .B1(_01268_),
    .X(_01287_));
 sg13g2_o21ai_1 _16976_ (.B1(_01287_),
    .Y(_01288_),
    .A1(_01269_),
    .A2(_01286_));
 sg13g2_nand2_1 _16977_ (.Y(_01289_),
    .A(\am_sdr0.nco0.phase[19] ),
    .B(_01272_));
 sg13g2_o21ai_1 _16978_ (.B1(_01289_),
    .Y(_01290_),
    .A1(_01283_),
    .A2(_01288_));
 sg13g2_a21oi_1 _16979_ (.A1(_01251_),
    .A2(_01282_),
    .Y(_01291_),
    .B1(_01290_));
 sg13g2_buf_1 _16980_ (.A(\am_sdr0.nco0.phase[20] ),
    .X(_01292_));
 sg13g2_buf_2 _16981_ (.A(\am_sdr0.nco0.phase_inc[20] ),
    .X(_01293_));
 sg13g2_xnor2_1 _16982_ (.Y(_01294_),
    .A(_01292_),
    .B(_01293_));
 sg13g2_xnor2_1 _16983_ (.Y(_01295_),
    .A(_01291_),
    .B(_01294_));
 sg13g2_nor2_1 _16984_ (.A(net47),
    .B(_01295_),
    .Y(_01089_));
 sg13g2_inv_1 _16985_ (.Y(_01296_),
    .A(_01292_));
 sg13g2_nor2_1 _16986_ (.A(_01275_),
    .B(_01284_),
    .Y(_01297_));
 sg13g2_a21oi_1 _16987_ (.A1(_01268_),
    .A2(_01269_),
    .Y(_01298_),
    .B1(_01297_));
 sg13g2_a21oi_1 _16988_ (.A1(_01289_),
    .A2(_01298_),
    .Y(_01299_),
    .B1(_01283_));
 sg13g2_nor2_1 _16989_ (.A(_01293_),
    .B(_01299_),
    .Y(_01300_));
 sg13g2_nand2_1 _16990_ (.Y(_01301_),
    .A(_01281_),
    .B(_01300_));
 sg13g2_o21ai_1 _16991_ (.B1(_01301_),
    .Y(_01302_),
    .A1(_01292_),
    .A2(_01293_));
 sg13g2_a221oi_1 _16992_ (.B2(_01259_),
    .C1(_01302_),
    .B1(_01300_),
    .A1(_01296_),
    .Y(_01303_),
    .A2(_01291_));
 sg13g2_buf_1 _16993_ (.A(\am_sdr0.nco0.phase[21] ),
    .X(_01304_));
 sg13g2_buf_1 _16994_ (.A(\am_sdr0.nco0.phase_inc[21] ),
    .X(_01305_));
 sg13g2_xor2_1 _16995_ (.B(_01305_),
    .A(_01304_),
    .X(_01306_));
 sg13g2_xnor2_1 _16996_ (.Y(_01307_),
    .A(_01303_),
    .B(_01306_));
 sg13g2_nor2_1 _16997_ (.A(net47),
    .B(_01307_),
    .Y(_01090_));
 sg13g2_buf_1 _16998_ (.A(_02779_),
    .X(_01308_));
 sg13g2_a221oi_1 _16999_ (.B2(_01305_),
    .C1(_01290_),
    .B1(_01304_),
    .A1(_01292_),
    .Y(_01309_),
    .A2(_01293_));
 sg13g2_buf_1 _17000_ (.A(_01309_),
    .X(_01310_));
 sg13g2_and2_1 _17001_ (.A(_01248_),
    .B(_01310_),
    .X(_01311_));
 sg13g2_or2_1 _17002_ (.X(_01312_),
    .B(_01282_),
    .A(_01290_));
 sg13g2_o21ai_1 _17003_ (.B1(_01292_),
    .Y(_01313_),
    .A1(_01293_),
    .A2(_01312_));
 sg13g2_nand2_1 _17004_ (.Y(_01314_),
    .A(_01293_),
    .B(_01312_));
 sg13g2_nor2_1 _17005_ (.A(_01304_),
    .B(_01305_),
    .Y(_01315_));
 sg13g2_a21oi_1 _17006_ (.A1(_01313_),
    .A2(_01314_),
    .Y(_01316_),
    .B1(_01315_));
 sg13g2_a21oi_1 _17007_ (.A1(_01304_),
    .A2(_01305_),
    .Y(_01317_),
    .B1(_01316_));
 sg13g2_a221oi_1 _17008_ (.B2(_01240_),
    .C1(_01317_),
    .B1(_01311_),
    .A1(_01249_),
    .Y(_01318_),
    .A2(_01310_));
 sg13g2_buf_1 _17009_ (.A(_01318_),
    .X(_01319_));
 sg13g2_buf_1 _17010_ (.A(\am_sdr0.nco0.phase_inc[22] ),
    .X(_01320_));
 sg13g2_xor2_1 _17011_ (.B(_01320_),
    .A(net365),
    .X(_01321_));
 sg13g2_xnor2_1 _17012_ (.Y(_01322_),
    .A(_01319_),
    .B(_01321_));
 sg13g2_nor2_1 _17013_ (.A(net46),
    .B(_01322_),
    .Y(_01091_));
 sg13g2_and2_1 _17014_ (.A(_01501_),
    .B(\am_sdr0.nco0.phase_inc[23] ),
    .X(_01323_));
 sg13g2_buf_1 _17015_ (.A(_01323_),
    .X(_01324_));
 sg13g2_nor2_1 _17016_ (.A(_01501_),
    .B(\am_sdr0.nco0.phase_inc[23] ),
    .Y(_01325_));
 sg13g2_nor2_1 _17017_ (.A(_01324_),
    .B(_01325_),
    .Y(_01326_));
 sg13g2_inv_1 _17018_ (.Y(_01327_),
    .A(_01320_));
 sg13g2_o21ai_1 _17019_ (.B1(_01319_),
    .Y(_01328_),
    .A1(_01502_),
    .A2(_01320_));
 sg13g2_o21ai_1 _17020_ (.B1(_01328_),
    .Y(_01329_),
    .A1(_01511_),
    .A2(_01327_));
 sg13g2_xnor2_1 _17021_ (.Y(_01330_),
    .A(_01326_),
    .B(_01329_));
 sg13g2_nor2_1 _17022_ (.A(net46),
    .B(_01330_),
    .Y(_01092_));
 sg13g2_nand3b_1 _17023_ (.B(_01319_),
    .C(_01320_),
    .Y(_01331_),
    .A_N(_01325_));
 sg13g2_nand4_1 _17024_ (.B(_01240_),
    .C(_01248_),
    .A(_01327_),
    .Y(_01332_),
    .D(_01310_));
 sg13g2_a21oi_1 _17025_ (.A1(_01249_),
    .A2(_01310_),
    .Y(_01333_),
    .B1(_01317_));
 sg13g2_nor2_1 _17026_ (.A(_01320_),
    .B(_01333_),
    .Y(_01334_));
 sg13g2_nor3_1 _17027_ (.A(_01511_),
    .B(_01325_),
    .C(_01334_),
    .Y(_01335_));
 sg13g2_a21oi_1 _17028_ (.A1(_01332_),
    .A2(_01335_),
    .Y(_01336_),
    .B1(_01324_));
 sg13g2_nand2_1 _17029_ (.Y(_01337_),
    .A(_01331_),
    .B(_01336_));
 sg13g2_buf_1 _17030_ (.A(\am_sdr0.nco0.phase_inc[24] ),
    .X(_01338_));
 sg13g2_xor2_1 _17031_ (.B(_01338_),
    .A(net306),
    .X(_01339_));
 sg13g2_xnor2_1 _17032_ (.Y(_01340_),
    .A(_01337_),
    .B(_01339_));
 sg13g2_nor2_1 _17033_ (.A(net46),
    .B(_01340_),
    .Y(_01093_));
 sg13g2_xor2_1 _17034_ (.B(\am_sdr0.nco0.phase_inc[25] ),
    .A(_01495_),
    .X(_01341_));
 sg13g2_a221oi_1 _17035_ (.B2(_01335_),
    .C1(_01324_),
    .B1(_01332_),
    .A1(net306),
    .Y(_01342_),
    .A2(_01338_));
 sg13g2_nor2_1 _17036_ (.A(_01499_),
    .B(_01338_),
    .Y(_01343_));
 sg13g2_a21oi_1 _17037_ (.A1(_01331_),
    .A2(_01342_),
    .Y(_01344_),
    .B1(_01343_));
 sg13g2_xnor2_1 _17038_ (.Y(_01345_),
    .A(_01341_),
    .B(_01344_));
 sg13g2_nor2_1 _17039_ (.A(net46),
    .B(_01345_),
    .Y(_01094_));
 sg13g2_xor2_1 _17040_ (.B(_08037_),
    .A(\am_sdr0.nco0.phase[2] ),
    .X(_01346_));
 sg13g2_xnor2_1 _17041_ (.Y(_01347_),
    .A(_08044_),
    .B(_01346_));
 sg13g2_nor2_1 _17042_ (.A(net46),
    .B(_01347_),
    .Y(_01095_));
 sg13g2_a21oi_1 _17043_ (.A1(_08038_),
    .A2(_08044_),
    .Y(_01348_),
    .B1(_08045_));
 sg13g2_xnor2_1 _17044_ (.Y(_01349_),
    .A(_08035_),
    .B(_08036_));
 sg13g2_xnor2_1 _17045_ (.Y(_01350_),
    .A(_01348_),
    .B(_01349_));
 sg13g2_nor2_1 _17046_ (.A(net46),
    .B(_01350_),
    .Y(_01096_));
 sg13g2_nor2_1 _17047_ (.A(_08035_),
    .B(_08036_),
    .Y(_01351_));
 sg13g2_nand2_1 _17048_ (.Y(_01352_),
    .A(_08035_),
    .B(_08036_));
 sg13g2_o21ai_1 _17049_ (.B1(_01352_),
    .Y(_01353_),
    .A1(_01348_),
    .A2(_01351_));
 sg13g2_and2_1 _17050_ (.A(_08047_),
    .B(_08049_),
    .X(_01354_));
 sg13g2_xnor2_1 _17051_ (.Y(_01355_),
    .A(_01353_),
    .B(_01354_));
 sg13g2_nor2_1 _17052_ (.A(net46),
    .B(_01355_),
    .Y(_01097_));
 sg13g2_xor2_1 _17053_ (.B(_08034_),
    .A(\am_sdr0.nco0.phase[5] ),
    .X(_01356_));
 sg13g2_xnor2_1 _17054_ (.Y(_01357_),
    .A(_08051_),
    .B(_01356_));
 sg13g2_nor2_1 _17055_ (.A(net46),
    .B(_01357_),
    .Y(_01098_));
 sg13g2_nor2_1 _17056_ (.A(_08052_),
    .B(_08053_),
    .Y(_01358_));
 sg13g2_xor2_1 _17057_ (.B(_08055_),
    .A(_08054_),
    .X(_01359_));
 sg13g2_xnor2_1 _17058_ (.Y(_01360_),
    .A(_01358_),
    .B(_01359_));
 sg13g2_nor2_1 _17059_ (.A(_01308_),
    .B(_01360_),
    .Y(_01099_));
 sg13g2_nand2_1 _17060_ (.Y(_01361_),
    .A(_08054_),
    .B(_08055_));
 sg13g2_nand2_1 _17061_ (.Y(_01362_),
    .A(_08058_),
    .B(_01361_));
 sg13g2_xor2_1 _17062_ (.B(_08032_),
    .A(_08030_),
    .X(_01363_));
 sg13g2_xnor2_1 _17063_ (.Y(_01364_),
    .A(_01362_),
    .B(_01363_));
 sg13g2_nor2_1 _17064_ (.A(_01308_),
    .B(_01364_),
    .Y(_01100_));
 sg13g2_xor2_1 _17065_ (.B(_08060_),
    .A(_01176_),
    .X(_01365_));
 sg13g2_xnor2_1 _17066_ (.Y(_01366_),
    .A(_01175_),
    .B(_01365_));
 sg13g2_nor2_1 _17067_ (.A(net181),
    .B(_01366_),
    .Y(_01101_));
 sg13g2_xor2_1 _17068_ (.B(_08029_),
    .A(_08028_),
    .X(_01367_));
 sg13g2_xnor2_1 _17069_ (.Y(_01368_),
    .A(_01178_),
    .B(_01367_));
 sg13g2_nor2_1 _17070_ (.A(net181),
    .B(_01368_),
    .Y(_01102_));
 sg13g2_a21oi_1 _17071_ (.A1(_01508_),
    .A2(_01541_),
    .Y(_01103_),
    .B1(_01514_));
 sg13g2_and2_1 _17072_ (.A(net193),
    .B(net4),
    .X(_01104_));
 sg13g2_and2_1 _17073_ (.A(net193),
    .B(\am_sdr0.spi0.CS_q ),
    .X(_01105_));
 sg13g2_nor2_1 _17074_ (.A(net259),
    .B(_02490_),
    .Y(_01106_));
 sg13g2_and2_1 _17075_ (.A(net193),
    .B(net2),
    .X(_01107_));
 sg13g2_and2_1 _17076_ (.A(_08026_),
    .B(\am_sdr0.spi0.MOSI_q ),
    .X(_01108_));
 sg13g2_and2_1 _17077_ (.A(_08026_),
    .B(net3),
    .X(_01109_));
 sg13g2_and2_1 _17078_ (.A(net257),
    .B(\am_sdr0.spi0.SCK_q ),
    .X(_01110_));
 sg13g2_and2_1 _17079_ (.A(net257),
    .B(\am_sdr0.spi0.SCK_qq ),
    .X(_01111_));
 sg13g2_nor2b_1 _17080_ (.A(_02488_),
    .B_N(_02492_),
    .Y(_01369_));
 sg13g2_buf_1 _17081_ (.A(_01369_),
    .X(_01370_));
 sg13g2_buf_1 _17082_ (.A(_01370_),
    .X(_01371_));
 sg13g2_nand2_1 _17083_ (.Y(_01372_),
    .A(\am_sdr0.spi0.shift_reg[26] ),
    .B(net143));
 sg13g2_nand2b_1 _17084_ (.Y(_01373_),
    .B(_02492_),
    .A_N(_02488_));
 sg13g2_buf_1 _17085_ (.A(_01373_),
    .X(_01374_));
 sg13g2_buf_1 _17086_ (.A(_01374_),
    .X(_01375_));
 sg13g2_nand2_1 _17087_ (.Y(_01376_),
    .A(_02588_),
    .B(net142));
 sg13g2_a21oi_1 _17088_ (.A1(_01372_),
    .A2(_01376_),
    .Y(_01112_),
    .B1(net49));
 sg13g2_buf_1 _17089_ (.A(net301),
    .X(_01377_));
 sg13g2_buf_1 _17090_ (.A(_01374_),
    .X(_01378_));
 sg13g2_buf_1 _17091_ (.A(net141),
    .X(_01379_));
 sg13g2_nand2_1 _17092_ (.Y(_01380_),
    .A(_02619_),
    .B(net45));
 sg13g2_buf_1 _17093_ (.A(_01370_),
    .X(_01381_));
 sg13g2_buf_1 _17094_ (.A(net140),
    .X(_01382_));
 sg13g2_nand2_1 _17095_ (.Y(_01383_),
    .A(\am_sdr0.spi0.shift_reg[27] ),
    .B(_01382_));
 sg13g2_nand3_1 _17096_ (.B(_01380_),
    .C(_01383_),
    .A(net192),
    .Y(_01113_));
 sg13g2_nand2_1 _17097_ (.Y(_01384_),
    .A(\am_sdr0.spi0.shift_reg[28] ),
    .B(net143));
 sg13g2_nand2_1 _17098_ (.Y(_01385_),
    .A(_02643_),
    .B(net142));
 sg13g2_a21oi_1 _17099_ (.A1(_01384_),
    .A2(_01385_),
    .Y(_01114_),
    .B1(net49));
 sg13g2_nand2_1 _17100_ (.Y(_01386_),
    .A(\am_sdr0.nco0.phase_inc[0] ),
    .B(net45));
 sg13g2_nand2_1 _17101_ (.Y(_01387_),
    .A(\am_sdr0.spi0.shift_reg[0] ),
    .B(_01382_));
 sg13g2_nand3_1 _17102_ (.B(_01386_),
    .C(_01387_),
    .A(net192),
    .Y(_01115_));
 sg13g2_nand2_1 _17103_ (.Y(_01388_),
    .A(\am_sdr0.spi0.shift_reg[10] ),
    .B(net143));
 sg13g2_nand2_1 _17104_ (.Y(_01389_),
    .A(_01182_),
    .B(net142));
 sg13g2_a21oi_1 _17105_ (.A1(_01388_),
    .A2(_01389_),
    .Y(_01116_),
    .B1(net49));
 sg13g2_nand2_1 _17106_ (.Y(_01390_),
    .A(\am_sdr0.spi0.shift_reg[11] ),
    .B(net143));
 sg13g2_nand2_1 _17107_ (.Y(_01391_),
    .A(_01204_),
    .B(net142));
 sg13g2_a21oi_1 _17108_ (.A1(_01390_),
    .A2(_01391_),
    .Y(_01117_),
    .B1(net49));
 sg13g2_nand2_1 _17109_ (.Y(_01392_),
    .A(_01211_),
    .B(net45));
 sg13g2_nand2_1 _17110_ (.Y(_01393_),
    .A(\am_sdr0.spi0.shift_reg[12] ),
    .B(net44));
 sg13g2_nand3_1 _17111_ (.B(_01392_),
    .C(_01393_),
    .A(net192),
    .Y(_01118_));
 sg13g2_nand2_1 _17112_ (.Y(_01394_),
    .A(\am_sdr0.spi0.shift_reg[13] ),
    .B(net143));
 sg13g2_nand2_1 _17113_ (.Y(_01395_),
    .A(_01216_),
    .B(net142));
 sg13g2_a21oi_1 _17114_ (.A1(_01394_),
    .A2(_01395_),
    .Y(_01119_),
    .B1(net49));
 sg13g2_nand2_1 _17115_ (.Y(_01396_),
    .A(\am_sdr0.spi0.shift_reg[14] ),
    .B(net143));
 sg13g2_nand2_1 _17116_ (.Y(_01397_),
    .A(_01226_),
    .B(net142));
 sg13g2_buf_1 _17117_ (.A(_07113_),
    .X(_01398_));
 sg13g2_a21oi_1 _17118_ (.A1(_01396_),
    .A2(_01397_),
    .Y(_01120_),
    .B1(net43));
 sg13g2_nand2_1 _17119_ (.Y(_01399_),
    .A(\am_sdr0.spi0.shift_reg[15] ),
    .B(net143));
 sg13g2_nand2_1 _17120_ (.Y(_01400_),
    .A(_01242_),
    .B(net142));
 sg13g2_a21oi_1 _17121_ (.A1(_01399_),
    .A2(_01400_),
    .Y(_01121_),
    .B1(_01398_));
 sg13g2_nand2_1 _17122_ (.Y(_01401_),
    .A(_01246_),
    .B(net45));
 sg13g2_nand2_1 _17123_ (.Y(_01402_),
    .A(\am_sdr0.spi0.shift_reg[16] ),
    .B(net44));
 sg13g2_nand3_1 _17124_ (.B(_01401_),
    .C(_01402_),
    .A(net192),
    .Y(_01122_));
 sg13g2_nand2_1 _17125_ (.Y(_01403_),
    .A(_01254_),
    .B(net45));
 sg13g2_nand2_1 _17126_ (.Y(_01404_),
    .A(\am_sdr0.spi0.shift_reg[17] ),
    .B(net44));
 sg13g2_nand3_1 _17127_ (.B(_01403_),
    .C(_01404_),
    .A(net192),
    .Y(_01123_));
 sg13g2_nand2_1 _17128_ (.Y(_01405_),
    .A(\am_sdr0.spi0.shift_reg[18] ),
    .B(net143));
 sg13g2_nand2_1 _17129_ (.Y(_01406_),
    .A(_01269_),
    .B(net142));
 sg13g2_a21oi_1 _17130_ (.A1(_01405_),
    .A2(_01406_),
    .Y(_01124_),
    .B1(_01398_));
 sg13g2_nand2_1 _17131_ (.Y(_01407_),
    .A(\am_sdr0.spi0.shift_reg[19] ),
    .B(net140));
 sg13g2_nand2_1 _17132_ (.Y(_01408_),
    .A(_01272_),
    .B(net141));
 sg13g2_a21oi_1 _17133_ (.A1(_01407_),
    .A2(_01408_),
    .Y(_01125_),
    .B1(net43));
 sg13g2_nand2_1 _17134_ (.Y(_01409_),
    .A(_08039_),
    .B(net45));
 sg13g2_nand2_1 _17135_ (.Y(_01410_),
    .A(\am_sdr0.spi0.shift_reg[1] ),
    .B(net44));
 sg13g2_nand3_1 _17136_ (.B(_01409_),
    .C(_01410_),
    .A(net192),
    .Y(_01126_));
 sg13g2_nand2_1 _17137_ (.Y(_01411_),
    .A(_01293_),
    .B(net45));
 sg13g2_nand2_1 _17138_ (.Y(_01412_),
    .A(\am_sdr0.spi0.shift_reg[20] ),
    .B(net44));
 sg13g2_nand3_1 _17139_ (.B(_01411_),
    .C(_01412_),
    .A(net192),
    .Y(_01127_));
 sg13g2_nand2_1 _17140_ (.Y(_01413_),
    .A(\am_sdr0.spi0.shift_reg[21] ),
    .B(net140));
 sg13g2_nand2_1 _17141_ (.Y(_01414_),
    .A(_01305_),
    .B(net141));
 sg13g2_a21oi_1 _17142_ (.A1(_01413_),
    .A2(_01414_),
    .Y(_01128_),
    .B1(net43));
 sg13g2_nand2_1 _17143_ (.Y(_01415_),
    .A(\am_sdr0.spi0.shift_reg[22] ),
    .B(net140));
 sg13g2_nand2_1 _17144_ (.Y(_01416_),
    .A(_01320_),
    .B(net141));
 sg13g2_a21oi_1 _17145_ (.A1(_01415_),
    .A2(_01416_),
    .Y(_01129_),
    .B1(net43));
 sg13g2_nand2_1 _17146_ (.Y(_01417_),
    .A(\am_sdr0.spi0.shift_reg[23] ),
    .B(net140));
 sg13g2_nand2_1 _17147_ (.Y(_01418_),
    .A(\am_sdr0.nco0.phase_inc[23] ),
    .B(net141));
 sg13g2_a21oi_1 _17148_ (.A1(_01417_),
    .A2(_01418_),
    .Y(_01130_),
    .B1(net43));
 sg13g2_nand2_1 _17149_ (.Y(_01419_),
    .A(\am_sdr0.spi0.shift_reg[24] ),
    .B(net140));
 sg13g2_nand2_1 _17150_ (.Y(_01420_),
    .A(_01338_),
    .B(net141));
 sg13g2_a21oi_1 _17151_ (.A1(_01419_),
    .A2(_01420_),
    .Y(_01131_),
    .B1(net43));
 sg13g2_nand2_1 _17152_ (.Y(_01421_),
    .A(\am_sdr0.spi0.shift_reg[25] ),
    .B(net140));
 sg13g2_nand2_1 _17153_ (.Y(_01422_),
    .A(\am_sdr0.nco0.phase_inc[25] ),
    .B(net141));
 sg13g2_a21oi_1 _17154_ (.A1(_01421_),
    .A2(_01422_),
    .Y(_01132_),
    .B1(net43));
 sg13g2_nand2_1 _17155_ (.Y(_01423_),
    .A(\am_sdr0.spi0.shift_reg[2] ),
    .B(_01381_));
 sg13g2_nand2_1 _17156_ (.Y(_01424_),
    .A(_08037_),
    .B(_01378_));
 sg13g2_a21oi_1 _17157_ (.A1(_01423_),
    .A2(_01424_),
    .Y(_01133_),
    .B1(net43));
 sg13g2_nand2_1 _17158_ (.Y(_01425_),
    .A(_08036_),
    .B(net45));
 sg13g2_nand2_1 _17159_ (.Y(_01426_),
    .A(\am_sdr0.spi0.shift_reg[3] ),
    .B(net44));
 sg13g2_nand3_1 _17160_ (.B(_01425_),
    .C(_01426_),
    .A(net192),
    .Y(_01134_));
 sg13g2_nand2_1 _17161_ (.Y(_01427_),
    .A(\am_sdr0.spi0.shift_reg[4] ),
    .B(_01381_));
 sg13g2_nand2_1 _17162_ (.Y(_01428_),
    .A(\am_sdr0.nco0.phase_inc[4] ),
    .B(net141));
 sg13g2_a21oi_1 _17163_ (.A1(_01427_),
    .A2(_01428_),
    .Y(_01135_),
    .B1(net177));
 sg13g2_nand2_1 _17164_ (.Y(_01429_),
    .A(_08034_),
    .B(_01379_));
 sg13g2_nand2_1 _17165_ (.Y(_01430_),
    .A(\am_sdr0.spi0.shift_reg[5] ),
    .B(net44));
 sg13g2_nand3_1 _17166_ (.B(_01429_),
    .C(_01430_),
    .A(_01377_),
    .Y(_01136_));
 sg13g2_nand2_1 _17167_ (.Y(_01431_),
    .A(_08055_),
    .B(_01379_));
 sg13g2_nand2_1 _17168_ (.Y(_01432_),
    .A(\am_sdr0.spi0.shift_reg[6] ),
    .B(net44));
 sg13g2_nand3_1 _17169_ (.B(_01431_),
    .C(_01432_),
    .A(_01377_),
    .Y(_01137_));
 sg13g2_nand2_1 _17170_ (.Y(_01433_),
    .A(_08032_),
    .B(_01375_));
 sg13g2_nand2_1 _17171_ (.Y(_01434_),
    .A(\am_sdr0.spi0.shift_reg[7] ),
    .B(_01371_));
 sg13g2_nand3_1 _17172_ (.B(_01433_),
    .C(_01434_),
    .A(_02809_),
    .Y(_01138_));
 sg13g2_nand2_1 _17173_ (.Y(_01435_),
    .A(\am_sdr0.spi0.shift_reg[8] ),
    .B(net140));
 sg13g2_nand2_1 _17174_ (.Y(_01436_),
    .A(_08060_),
    .B(_01378_));
 sg13g2_a21oi_1 _17175_ (.A1(_01435_),
    .A2(_01436_),
    .Y(_01139_),
    .B1(net177));
 sg13g2_nand2_1 _17176_ (.Y(_01437_),
    .A(_08029_),
    .B(_01375_));
 sg13g2_nand2_1 _17177_ (.Y(_01438_),
    .A(\am_sdr0.spi0.shift_reg[9] ),
    .B(_01371_));
 sg13g2_nand3_1 _17178_ (.B(_01437_),
    .C(_01438_),
    .A(net246),
    .Y(_01140_));
 sg13g2_o21ai_1 _17179_ (.B1(\am_sdr0.spi0.CS_qqq ),
    .Y(_01439_),
    .A1(_02488_),
    .A2(_02490_));
 sg13g2_nand2_1 _17180_ (.Y(_01440_),
    .A(_02488_),
    .B(_02490_));
 sg13g2_a21oi_1 _17181_ (.A1(_01439_),
    .A2(_01440_),
    .Y(_01170_),
    .B1(_02493_));
 sg13g2_inv_1 _17182_ (.Y(_01441_),
    .A(\am_sdr0.spi0.CS_qqq ));
 sg13g2_and3_1 _17183_ (.X(_01171_),
    .A(_01441_),
    .B(net184),
    .C(_01106_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_tiehi \am_sdr0.PWM_OUT$_SDFF_PN0__390  (.L_HI(net390));
 sg13g2_buf_1 _17186_ (.A(net368),
    .X(uio_oe[0]));
 sg13g2_buf_1 _17187_ (.A(net369),
    .X(uio_oe[1]));
 sg13g2_buf_1 _17188_ (.A(net370),
    .X(uio_oe[2]));
 sg13g2_buf_1 _17189_ (.A(net371),
    .X(uio_oe[3]));
 sg13g2_buf_1 _17190_ (.A(net372),
    .X(uio_oe[4]));
 sg13g2_buf_1 _17191_ (.A(net373),
    .X(uio_oe[5]));
 sg13g2_buf_1 _17192_ (.A(net374),
    .X(uio_oe[6]));
 sg13g2_buf_1 _17193_ (.A(net375),
    .X(uio_oe[7]));
 sg13g2_buf_1 _17194_ (.A(net376),
    .X(uio_out[0]));
 sg13g2_buf_1 _17195_ (.A(net377),
    .X(uio_out[1]));
 sg13g2_buf_1 _17196_ (.A(net378),
    .X(uio_out[2]));
 sg13g2_buf_1 _17197_ (.A(net379),
    .X(uio_out[3]));
 sg13g2_buf_1 _17198_ (.A(net380),
    .X(uio_out[4]));
 sg13g2_buf_1 _17199_ (.A(net381),
    .X(uio_out[5]));
 sg13g2_buf_1 _17200_ (.A(net382),
    .X(uio_out[6]));
 sg13g2_buf_1 _17201_ (.A(net383),
    .X(uio_out[7]));
 sg13g2_buf_1 _17202_ (.A(COMP_OUT),
    .X(net5));
 sg13g2_buf_1 _17203_ (.A(PWM_OUT),
    .X(net6));
 sg13g2_buf_1 _17204_ (.A(net384),
    .X(uo_out[2]));
 sg13g2_buf_1 _17205_ (.A(net385),
    .X(uo_out[3]));
 sg13g2_buf_1 _17206_ (.A(net386),
    .X(uo_out[4]));
 sg13g2_buf_1 _17207_ (.A(net387),
    .X(uo_out[5]));
 sg13g2_buf_1 _17208_ (.A(net388),
    .X(uo_out[6]));
 sg13g2_buf_1 _17209_ (.A(net389),
    .X(uo_out[7]));
 sg13g2_dfrbp_1 \am_sdr0.PWM_OUT$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net390),
    .D(_00074_),
    .Q_N(_09120_),
    .Q(PWM_OUT));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net391),
    .D(_00075_),
    .Q_N(_09119_),
    .Q(\am_sdr0.am0.a[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[10]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net392),
    .D(_00076_),
    .Q_N(_09118_),
    .Q(\am_sdr0.am0.a[10] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[11]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net393),
    .D(_00077_),
    .Q_N(_09117_),
    .Q(\am_sdr0.am0.a[11] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[12]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net394),
    .D(_00078_),
    .Q_N(_09116_),
    .Q(\am_sdr0.am0.a[12] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[13]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net395),
    .D(_00079_),
    .Q_N(_09115_),
    .Q(\am_sdr0.am0.a[13] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[14]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net396),
    .D(_00080_),
    .Q_N(_09114_),
    .Q(\am_sdr0.am0.a[14] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[15]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net397),
    .D(_00081_),
    .Q_N(_09113_),
    .Q(\am_sdr0.am0.a[15] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net398),
    .D(_00082_),
    .Q_N(_09112_),
    .Q(\am_sdr0.am0.a[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net399),
    .D(_00083_),
    .Q_N(_09111_),
    .Q(\am_sdr0.am0.a[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[3]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net400),
    .D(_00084_),
    .Q_N(_09110_),
    .Q(\am_sdr0.am0.a[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[4]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net401),
    .D(_00085_),
    .Q_N(_09109_),
    .Q(\am_sdr0.am0.a[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[5]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net402),
    .D(_00086_),
    .Q_N(_09108_),
    .Q(\am_sdr0.am0.a[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net403),
    .D(_00087_),
    .Q_N(_09107_),
    .Q(\am_sdr0.am0.a[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[7]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net404),
    .D(_00088_),
    .Q_N(_09106_),
    .Q(\am_sdr0.am0.a[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[8]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net405),
    .D(_00089_),
    .Q_N(_09105_),
    .Q(\am_sdr0.am0.a[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.a[9]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net406),
    .D(_00090_),
    .Q_N(_09104_),
    .Q(\am_sdr0.am0.a[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count2[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net407),
    .D(_00091_),
    .Q_N(_00070_),
    .Q(\am_sdr0.am0.count2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count2[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net408),
    .D(_00092_),
    .Q_N(_09103_),
    .Q(\am_sdr0.am0.count2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count2[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net409),
    .D(_00093_),
    .Q_N(_09102_),
    .Q(\am_sdr0.am0.count2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count2[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net410),
    .D(_00094_),
    .Q_N(_09101_),
    .Q(\am_sdr0.am0.count2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net411),
    .D(_00095_),
    .Q_N(_00069_),
    .Q(\am_sdr0.am0.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.count[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net412),
    .D(_00096_),
    .Q_N(_09100_),
    .Q(\am_sdr0.am0.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net413),
    .D(_00097_),
    .Q_N(_09099_),
    .Q(\am_sdr0.am0.demod_out[10] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net414),
    .D(_00098_),
    .Q_N(_09098_),
    .Q(\am_sdr0.am0.demod_out[11] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net415),
    .D(_00099_),
    .Q_N(_09097_),
    .Q(\am_sdr0.am0.demod_out[12] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net416),
    .D(_00100_),
    .Q_N(_09096_),
    .Q(\am_sdr0.am0.demod_out[13] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net417),
    .D(_00101_),
    .Q_N(_09095_),
    .Q(\am_sdr0.am0.demod_out[14] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net418),
    .D(_00102_),
    .Q_N(_09094_),
    .Q(\am_sdr0.am0.demod_out[15] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net419),
    .D(_00103_),
    .Q_N(_09093_),
    .Q(\am_sdr0.am0.demod_out[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.demod_out[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net420),
    .D(_00104_),
    .Q_N(_09092_),
    .Q(\am_sdr0.am0.demod_out[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net421),
    .D(_00105_),
    .Q_N(_09091_),
    .Q(\am_sdr0.am0.left[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net422),
    .D(_00106_),
    .Q_N(_09090_),
    .Q(\am_sdr0.am0.left[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net423),
    .D(_00107_),
    .Q_N(_00042_),
    .Q(\am_sdr0.am0.left[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net424),
    .D(_00108_),
    .Q_N(_09089_),
    .Q(\am_sdr0.am0.left[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net425),
    .D(_00109_),
    .Q_N(_09088_),
    .Q(\am_sdr0.am0.left[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net426),
    .D(_00110_),
    .Q_N(_09087_),
    .Q(\am_sdr0.am0.left[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net427),
    .D(_00111_),
    .Q_N(_09086_),
    .Q(\am_sdr0.am0.left[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net428),
    .D(_00112_),
    .Q_N(_09085_),
    .Q(\am_sdr0.am0.left[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net429),
    .D(_00113_),
    .Q_N(_09084_),
    .Q(\am_sdr0.am0.left[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.left[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net430),
    .D(_00114_),
    .Q_N(_09083_),
    .Q(\am_sdr0.am0.left[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.m_count[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net431),
    .D(_00115_),
    .Q_N(_00071_),
    .Q(\am_sdr0.am0.m_count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.m_count[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net432),
    .D(_00116_),
    .Q_N(_09082_),
    .Q(\am_sdr0.am0.m_count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.m_count[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net433),
    .D(_00117_),
    .Q_N(_09081_),
    .Q(\am_sdr0.am0.m_count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.m_count[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net434),
    .D(_00118_),
    .Q_N(_09080_),
    .Q(\am_sdr0.am0.m_count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net435),
    .D(_00119_),
    .Q_N(_00055_),
    .Q(\am_sdr0.am0.multA[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[10]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net436),
    .D(_00120_),
    .Q_N(_00062_),
    .Q(\am_sdr0.am0.multA[10] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[11]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net437),
    .D(_00121_),
    .Q_N(_00063_),
    .Q(\am_sdr0.am0.multA[11] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[12]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net438),
    .D(_00122_),
    .Q_N(_00064_),
    .Q(\am_sdr0.am0.multA[12] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[13]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net439),
    .D(_00123_),
    .Q_N(_00065_),
    .Q(\am_sdr0.am0.multA[13] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[14]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net440),
    .D(_00124_),
    .Q_N(_00066_),
    .Q(\am_sdr0.am0.multA[14] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[15]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net441),
    .D(_00125_),
    .Q_N(_00067_),
    .Q(\am_sdr0.am0.multA[15] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[16]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net442),
    .D(_00126_),
    .Q_N(_09079_),
    .Q(\am_sdr0.am0.multA[16] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net443),
    .D(_00127_),
    .Q_N(_00052_),
    .Q(\am_sdr0.am0.multA[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net444),
    .D(_00128_),
    .Q_N(_00053_),
    .Q(\am_sdr0.am0.multA[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net445),
    .D(_00129_),
    .Q_N(_00054_),
    .Q(\am_sdr0.am0.multA[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net446),
    .D(_00130_),
    .Q_N(_00056_),
    .Q(\am_sdr0.am0.multA[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net447),
    .D(_00131_),
    .Q_N(_00057_),
    .Q(\am_sdr0.am0.multA[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[6]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net448),
    .D(_00132_),
    .Q_N(_00058_),
    .Q(\am_sdr0.am0.multA[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[7]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net449),
    .D(_00133_),
    .Q_N(_00059_),
    .Q(\am_sdr0.am0.multA[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[8]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net450),
    .D(_00134_),
    .Q_N(_00060_),
    .Q(\am_sdr0.am0.multA[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multA[9]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net451),
    .D(_00135_),
    .Q_N(_00061_),
    .Q(\am_sdr0.am0.multA[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net452),
    .D(_00136_),
    .Q_N(_09078_),
    .Q(\am_sdr0.am0.multB[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net453),
    .D(_00137_),
    .Q_N(_09077_),
    .Q(\am_sdr0.am0.multB[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net454),
    .D(_00138_),
    .Q_N(_09076_),
    .Q(\am_sdr0.am0.multB[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net455),
    .D(_00139_),
    .Q_N(_09075_),
    .Q(\am_sdr0.am0.multB[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[4]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net456),
    .D(_00140_),
    .Q_N(_09074_),
    .Q(\am_sdr0.am0.multB[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[5]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net457),
    .D(_00141_),
    .Q_N(_09073_),
    .Q(\am_sdr0.am0.multB[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[6]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net458),
    .D(_00142_),
    .Q_N(_09072_),
    .Q(\am_sdr0.am0.multB[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.multB[7]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net459),
    .D(_00143_),
    .Q_N(_09071_),
    .Q(\am_sdr0.am0.multB[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net460),
    .D(_00144_),
    .Q_N(_09070_),
    .Q(\am_sdr0.am0.q[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net461),
    .D(_00145_),
    .Q_N(_09069_),
    .Q(\am_sdr0.am0.q[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net462),
    .D(_00146_),
    .Q_N(_09068_),
    .Q(\am_sdr0.am0.q[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net463),
    .D(_00147_),
    .Q_N(_09067_),
    .Q(\am_sdr0.am0.q[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net464),
    .D(_00148_),
    .Q_N(_09066_),
    .Q(\am_sdr0.am0.q[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net465),
    .D(_00149_),
    .Q_N(_09065_),
    .Q(\am_sdr0.am0.q[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net466),
    .D(_00150_),
    .Q_N(_09064_),
    .Q(\am_sdr0.am0.q[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.q[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net467),
    .D(_00151_),
    .Q_N(_09063_),
    .Q(\am_sdr0.am0.q[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net468),
    .D(_00152_),
    .Q_N(_09062_),
    .Q(\am_sdr0.am0.r[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net469),
    .D(_00153_),
    .Q_N(_09061_),
    .Q(\am_sdr0.am0.r[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net470),
    .D(_00154_),
    .Q_N(_09060_),
    .Q(\am_sdr0.am0.r[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net471),
    .D(_00155_),
    .Q_N(_09059_),
    .Q(\am_sdr0.am0.r[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net472),
    .D(_00156_),
    .Q_N(_09058_),
    .Q(\am_sdr0.am0.r[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net473),
    .D(_00157_),
    .Q_N(_09057_),
    .Q(\am_sdr0.am0.r[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net474),
    .D(_00158_),
    .Q_N(_09056_),
    .Q(\am_sdr0.am0.r[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net475),
    .D(_00159_),
    .Q_N(_09055_),
    .Q(\am_sdr0.am0.r[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.r[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net476),
    .D(_00160_),
    .Q_N(_00022_),
    .Q(\am_sdr0.am0.r[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net477),
    .D(_00161_),
    .Q_N(_00045_),
    .Q(\am_sdr0.am0.right[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net478),
    .D(_00162_),
    .Q_N(_00041_),
    .Q(\am_sdr0.am0.right[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net479),
    .D(_00163_),
    .Q_N(_00043_),
    .Q(\am_sdr0.am0.right[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net480),
    .D(_00164_),
    .Q_N(_00044_),
    .Q(\am_sdr0.am0.right[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net481),
    .D(_00165_),
    .Q_N(_00046_),
    .Q(\am_sdr0.am0.right[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net482),
    .D(_00166_),
    .Q_N(_00047_),
    .Q(\am_sdr0.am0.right[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net483),
    .D(_00167_),
    .Q_N(_00048_),
    .Q(\am_sdr0.am0.right[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net484),
    .D(_00168_),
    .Q_N(_00049_),
    .Q(\am_sdr0.am0.right[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net485),
    .D(_00169_),
    .Q_N(_00051_),
    .Q(\am_sdr0.am0.right[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.right[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net486),
    .D(_00170_),
    .Q_N(_00050_),
    .Q(\am_sdr0.am0.right[9] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sqrt_done$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net487),
    .D(_00171_),
    .Q_N(_09054_),
    .Q(\am_sdr0.am0.sqrt_done ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sqrt_state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net488),
    .D(_00172_),
    .Q_N(_09053_),
    .Q(\am_sdr0.am0.sqrt_state[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sqrt_state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net489),
    .D(_00173_),
    .Q_N(_09121_),
    .Q(\am_sdr0.am0.sqrt_state[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[0]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net490),
    .D(_00018_),
    .Q_N(_09122_),
    .Q(\am_sdr0.am0.state[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[1]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net491),
    .D(_00019_),
    .Q_N(_09123_),
    .Q(\am_sdr0.am0.state[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[2]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net492),
    .D(_00020_),
    .Q_N(_09124_),
    .Q(\am_sdr0.am0.state[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[3]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net493),
    .D(_00015_),
    .Q_N(_09125_),
    .Q(\am_sdr0.am0.state[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[4]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net494),
    .D(_00016_),
    .Q_N(_09126_),
    .Q(\am_sdr0.am0.state[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[5]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net495),
    .D(_00017_),
    .Q_N(_09127_),
    .Q(\am_sdr0.am0.state[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.state[6]$_DFF_P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net496),
    .D(_00021_),
    .Q_N(_09052_),
    .Q(\am_sdr0.am0.state[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net497),
    .D(_00174_),
    .Q_N(_09051_),
    .Q(\am_sdr0.am0.sum[0] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[10]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net498),
    .D(_00175_),
    .Q_N(_09050_),
    .Q(\am_sdr0.am0.sum[10] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[11]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net499),
    .D(_00176_),
    .Q_N(_09049_),
    .Q(\am_sdr0.am0.sum[11] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[12]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net500),
    .D(_00177_),
    .Q_N(_09048_),
    .Q(\am_sdr0.am0.sum[12] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[13]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net501),
    .D(_00178_),
    .Q_N(_09047_),
    .Q(\am_sdr0.am0.sum[13] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[14]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net502),
    .D(_00179_),
    .Q_N(_09046_),
    .Q(\am_sdr0.am0.sum[14] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[15]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net503),
    .D(_00180_),
    .Q_N(_09045_),
    .Q(\am_sdr0.am0.sum[15] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[16]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net504),
    .D(_00181_),
    .Q_N(_09044_),
    .Q(\am_sdr0.am0.sum[16] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net505),
    .D(_00182_),
    .Q_N(_09043_),
    .Q(\am_sdr0.am0.sum[1] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net506),
    .D(_00183_),
    .Q_N(_09042_),
    .Q(\am_sdr0.am0.sum[2] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net507),
    .D(_00184_),
    .Q_N(_09041_),
    .Q(\am_sdr0.am0.sum[3] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net508),
    .D(_00185_),
    .Q_N(_09040_),
    .Q(\am_sdr0.am0.sum[4] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net509),
    .D(_00186_),
    .Q_N(_09039_),
    .Q(\am_sdr0.am0.sum[5] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net510),
    .D(_00187_),
    .Q_N(_09038_),
    .Q(\am_sdr0.am0.sum[6] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net511),
    .D(_00188_),
    .Q_N(_09037_),
    .Q(\am_sdr0.am0.sum[7] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net512),
    .D(_00189_),
    .Q_N(_09036_),
    .Q(\am_sdr0.am0.sum[8] ));
 sg13g2_dfrbp_1 \am_sdr0.am0.sum[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net513),
    .D(_00190_),
    .Q_N(_09035_),
    .Q(\am_sdr0.am0.sum[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net514),
    .D(_00191_),
    .Q_N(_09034_),
    .Q(\am_sdr0.cic0.comb1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net515),
    .D(_00192_),
    .Q_N(_09033_),
    .Q(\am_sdr0.cic0.comb1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net516),
    .D(_00193_),
    .Q_N(_09032_),
    .Q(\am_sdr0.cic0.comb1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net517),
    .D(_00194_),
    .Q_N(_09031_),
    .Q(\am_sdr0.cic0.comb1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net518),
    .D(_00195_),
    .Q_N(_09030_),
    .Q(\am_sdr0.cic0.comb1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net519),
    .D(_00196_),
    .Q_N(_09029_),
    .Q(\am_sdr0.cic0.comb1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net520),
    .D(_00197_),
    .Q_N(_09028_),
    .Q(\am_sdr0.cic0.comb1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net521),
    .D(_00198_),
    .Q_N(_09027_),
    .Q(\am_sdr0.cic0.comb1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net522),
    .D(_00199_),
    .Q_N(_09026_),
    .Q(\am_sdr0.cic0.comb1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net523),
    .D(_00200_),
    .Q_N(_09025_),
    .Q(\am_sdr0.cic0.comb1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net524),
    .D(_00201_),
    .Q_N(_09024_),
    .Q(\am_sdr0.cic0.comb1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net525),
    .D(_00202_),
    .Q_N(_09023_),
    .Q(\am_sdr0.cic0.comb1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net526),
    .D(_00203_),
    .Q_N(_09022_),
    .Q(\am_sdr0.cic0.comb1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net527),
    .D(_00204_),
    .Q_N(_09021_),
    .Q(\am_sdr0.cic0.comb1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net528),
    .D(_00205_),
    .Q_N(_09020_),
    .Q(\am_sdr0.cic0.comb1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net529),
    .D(_00206_),
    .Q_N(_09019_),
    .Q(\am_sdr0.cic0.comb1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net530),
    .D(_00207_),
    .Q_N(_09018_),
    .Q(\am_sdr0.cic0.comb1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net531),
    .D(_00208_),
    .Q_N(_09017_),
    .Q(\am_sdr0.cic0.comb1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net532),
    .D(_00209_),
    .Q_N(_09016_),
    .Q(\am_sdr0.cic0.comb1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net533),
    .D(_00210_),
    .Q_N(_09015_),
    .Q(\am_sdr0.cic0.comb1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net534),
    .D(_00211_),
    .Q_N(_09014_),
    .Q(\am_sdr0.cic0.comb1_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net535),
    .D(_00212_),
    .Q_N(_09013_),
    .Q(\am_sdr0.cic0.comb1_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net536),
    .D(_00213_),
    .Q_N(_09012_),
    .Q(\am_sdr0.cic0.comb1_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net537),
    .D(_00214_),
    .Q_N(_09011_),
    .Q(\am_sdr0.cic0.comb1_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net538),
    .D(_00215_),
    .Q_N(_09010_),
    .Q(\am_sdr0.cic0.comb1_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net539),
    .D(_00216_),
    .Q_N(_09009_),
    .Q(\am_sdr0.cic0.comb1_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net540),
    .D(_00217_),
    .Q_N(_09008_),
    .Q(\am_sdr0.cic0.comb1_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net541),
    .D(_00218_),
    .Q_N(_09007_),
    .Q(\am_sdr0.cic0.comb1_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net542),
    .D(_00219_),
    .Q_N(_09006_),
    .Q(\am_sdr0.cic0.comb1_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net543),
    .D(_00220_),
    .Q_N(_09005_),
    .Q(\am_sdr0.cic0.comb1_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net544),
    .D(_00221_),
    .Q_N(_09004_),
    .Q(\am_sdr0.cic0.comb1_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net545),
    .D(_00222_),
    .Q_N(_09003_),
    .Q(\am_sdr0.cic0.comb1_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net546),
    .D(_00223_),
    .Q_N(_09002_),
    .Q(\am_sdr0.cic0.comb1_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net547),
    .D(_00224_),
    .Q_N(_09001_),
    .Q(\am_sdr0.cic0.comb1_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net548),
    .D(_00225_),
    .Q_N(_09000_),
    .Q(\am_sdr0.cic0.comb1_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net549),
    .D(_00226_),
    .Q_N(_08999_),
    .Q(\am_sdr0.cic0.comb1_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net550),
    .D(_00227_),
    .Q_N(_08998_),
    .Q(\am_sdr0.cic0.comb1_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net551),
    .D(_00228_),
    .Q_N(_08997_),
    .Q(\am_sdr0.cic0.comb1_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net552),
    .D(_00229_),
    .Q_N(_08996_),
    .Q(\am_sdr0.cic0.comb1_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb1_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net553),
    .D(_00230_),
    .Q_N(_08995_),
    .Q(\am_sdr0.cic0.comb1_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net554),
    .D(_00231_),
    .Q_N(_08994_),
    .Q(\am_sdr0.cic0.comb2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net555),
    .D(_00232_),
    .Q_N(_08993_),
    .Q(\am_sdr0.cic0.comb2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net556),
    .D(_00233_),
    .Q_N(_08992_),
    .Q(\am_sdr0.cic0.comb2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net557),
    .D(_00234_),
    .Q_N(_08991_),
    .Q(\am_sdr0.cic0.comb2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net558),
    .D(_00235_),
    .Q_N(_08990_),
    .Q(\am_sdr0.cic0.comb2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net559),
    .D(_00236_),
    .Q_N(_08989_),
    .Q(\am_sdr0.cic0.comb2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net560),
    .D(_00237_),
    .Q_N(_08988_),
    .Q(\am_sdr0.cic0.comb2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net561),
    .D(_00238_),
    .Q_N(_08987_),
    .Q(\am_sdr0.cic0.comb2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net562),
    .D(_00239_),
    .Q_N(_08986_),
    .Q(\am_sdr0.cic0.comb2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net563),
    .D(_00240_),
    .Q_N(_08985_),
    .Q(\am_sdr0.cic0.comb2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net564),
    .D(_00241_),
    .Q_N(_08984_),
    .Q(\am_sdr0.cic0.comb2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net565),
    .D(_00242_),
    .Q_N(_08983_),
    .Q(\am_sdr0.cic0.comb2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net566),
    .D(_00243_),
    .Q_N(_08982_),
    .Q(\am_sdr0.cic0.comb2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net567),
    .D(_00244_),
    .Q_N(_08981_),
    .Q(\am_sdr0.cic0.comb2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net568),
    .D(_00245_),
    .Q_N(_08980_),
    .Q(\am_sdr0.cic0.comb2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net569),
    .D(_00246_),
    .Q_N(_08979_),
    .Q(\am_sdr0.cic0.comb2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net570),
    .D(_00247_),
    .Q_N(_08978_),
    .Q(\am_sdr0.cic0.comb2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net571),
    .D(_00248_),
    .Q_N(_08977_),
    .Q(\am_sdr0.cic0.comb2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net572),
    .D(_00249_),
    .Q_N(_08976_),
    .Q(\am_sdr0.cic0.comb2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net573),
    .D(_00250_),
    .Q_N(_08975_),
    .Q(\am_sdr0.cic0.comb2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net574),
    .D(_00251_),
    .Q_N(_08974_),
    .Q(\am_sdr0.cic0.comb2_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net575),
    .D(_00252_),
    .Q_N(_08973_),
    .Q(\am_sdr0.cic0.comb2_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net576),
    .D(_00253_),
    .Q_N(_08972_),
    .Q(\am_sdr0.cic0.comb2_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net577),
    .D(_00254_),
    .Q_N(_08971_),
    .Q(\am_sdr0.cic0.comb2_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net578),
    .D(_00255_),
    .Q_N(_08970_),
    .Q(\am_sdr0.cic0.comb2_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net579),
    .D(_00256_),
    .Q_N(_08969_),
    .Q(\am_sdr0.cic0.comb2_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net580),
    .D(_00257_),
    .Q_N(_08968_),
    .Q(\am_sdr0.cic0.comb2_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net581),
    .D(_00258_),
    .Q_N(_08967_),
    .Q(\am_sdr0.cic0.comb2_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net582),
    .D(_00259_),
    .Q_N(_08966_),
    .Q(\am_sdr0.cic0.comb2_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net583),
    .D(_00260_),
    .Q_N(_08965_),
    .Q(\am_sdr0.cic0.comb2_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net584),
    .D(_00261_),
    .Q_N(_08964_),
    .Q(\am_sdr0.cic0.comb2_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net585),
    .D(_00262_),
    .Q_N(_08963_),
    .Q(\am_sdr0.cic0.comb2_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net586),
    .D(_00263_),
    .Q_N(_08962_),
    .Q(\am_sdr0.cic0.comb2_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net587),
    .D(_00264_),
    .Q_N(_08961_),
    .Q(\am_sdr0.cic0.comb2_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net588),
    .D(_00265_),
    .Q_N(_08960_),
    .Q(\am_sdr0.cic0.comb2_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net589),
    .D(_00266_),
    .Q_N(_08959_),
    .Q(\am_sdr0.cic0.comb2_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net590),
    .D(_00267_),
    .Q_N(_08958_),
    .Q(\am_sdr0.cic0.comb2_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net591),
    .D(_00268_),
    .Q_N(_08957_),
    .Q(\am_sdr0.cic0.comb2_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net592),
    .D(_00269_),
    .Q_N(_08956_),
    .Q(\am_sdr0.cic0.comb2_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb2_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net593),
    .D(_00270_),
    .Q_N(_08955_),
    .Q(\am_sdr0.cic0.comb2_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net594),
    .D(_00271_),
    .Q_N(_08954_),
    .Q(\am_sdr0.cic0.comb3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net595),
    .D(_00272_),
    .Q_N(_08953_),
    .Q(\am_sdr0.cic0.comb3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net596),
    .D(_00273_),
    .Q_N(_08952_),
    .Q(\am_sdr0.cic0.comb3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net597),
    .D(_00274_),
    .Q_N(_08951_),
    .Q(\am_sdr0.cic0.comb3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net598),
    .D(_00275_),
    .Q_N(_08950_),
    .Q(\am_sdr0.cic0.comb3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net599),
    .D(_00276_),
    .Q_N(_08949_),
    .Q(\am_sdr0.cic0.comb3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net600),
    .D(_00277_),
    .Q_N(_08948_),
    .Q(\am_sdr0.cic0.comb3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net601),
    .D(_00278_),
    .Q_N(_08947_),
    .Q(\am_sdr0.cic0.comb3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net602),
    .D(_00279_),
    .Q_N(_08946_),
    .Q(\am_sdr0.cic0.comb3_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net603),
    .D(_00280_),
    .Q_N(_08945_),
    .Q(\am_sdr0.cic0.comb3_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net604),
    .D(_00281_),
    .Q_N(_08944_),
    .Q(\am_sdr0.cic0.comb3_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net605),
    .D(_00282_),
    .Q_N(_08943_),
    .Q(\am_sdr0.cic0.comb3_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net606),
    .D(_00283_),
    .Q_N(_08942_),
    .Q(\am_sdr0.cic0.comb3_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net607),
    .D(_00284_),
    .Q_N(_08941_),
    .Q(\am_sdr0.cic0.comb3_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net608),
    .D(_00285_),
    .Q_N(_08940_),
    .Q(\am_sdr0.cic0.comb3_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net609),
    .D(_00286_),
    .Q_N(_08939_),
    .Q(\am_sdr0.cic0.comb3_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net610),
    .D(_00287_),
    .Q_N(_08938_),
    .Q(\am_sdr0.cic0.comb3_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net611),
    .D(_00288_),
    .Q_N(_08937_),
    .Q(\am_sdr0.cic0.comb3_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net612),
    .D(_00289_),
    .Q_N(_08936_),
    .Q(\am_sdr0.cic0.comb3_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net613),
    .D(_00290_),
    .Q_N(_08935_),
    .Q(\am_sdr0.cic0.comb3_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net614),
    .D(_00291_),
    .Q_N(_08934_),
    .Q(\am_sdr0.cic0.comb3_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net615),
    .D(_00292_),
    .Q_N(_08933_),
    .Q(\am_sdr0.cic0.comb3_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net616),
    .D(_00293_),
    .Q_N(_08932_),
    .Q(\am_sdr0.cic0.comb3_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net617),
    .D(_00294_),
    .Q_N(_08931_),
    .Q(\am_sdr0.cic0.comb3_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net618),
    .D(_00295_),
    .Q_N(_08930_),
    .Q(\am_sdr0.cic0.comb3_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net619),
    .D(_00296_),
    .Q_N(_08929_),
    .Q(\am_sdr0.cic0.comb3_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net620),
    .D(_00297_),
    .Q_N(_08928_),
    .Q(\am_sdr0.cic0.comb3_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.comb3_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net621),
    .D(_00298_),
    .Q_N(_08927_),
    .Q(\am_sdr0.cic0.comb3_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[0]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net622),
    .D(_00299_),
    .Q_N(_00072_),
    .Q(\am_sdr0.cic0.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[1]$_SDFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net623),
    .D(_00300_),
    .Q_N(_08926_),
    .Q(\am_sdr0.cic0.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[2]$_SDFF_PP0_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net624),
    .D(_00301_),
    .Q_N(_08925_),
    .Q(\am_sdr0.cic0.count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[3]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net625),
    .D(_00302_),
    .Q_N(_08924_),
    .Q(\am_sdr0.cic0.count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[4]$_SDFF_PP0_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net626),
    .D(_00303_),
    .Q_N(_08923_),
    .Q(\am_sdr0.cic0.count[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[5]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net627),
    .D(_00304_),
    .Q_N(_08922_),
    .Q(\am_sdr0.cic0.count[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[6]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net628),
    .D(_00305_),
    .Q_N(_08921_),
    .Q(\am_sdr0.cic0.count[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.count[7]$_SDFF_PP0_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net629),
    .D(_00306_),
    .Q_N(_08920_),
    .Q(\am_sdr0.cic0.count[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[0]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net630),
    .D(_00307_),
    .Q_N(_08919_),
    .Q(\am_sdr0.cic0.integ1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[10]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net631),
    .D(_00308_),
    .Q_N(_08918_),
    .Q(\am_sdr0.cic0.integ1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[11]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net632),
    .D(_00309_),
    .Q_N(_08917_),
    .Q(\am_sdr0.cic0.integ1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[12]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net633),
    .D(_00310_),
    .Q_N(_08916_),
    .Q(\am_sdr0.cic0.integ1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[13]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net634),
    .D(_00311_),
    .Q_N(_08915_),
    .Q(\am_sdr0.cic0.integ1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[14]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net635),
    .D(_00312_),
    .Q_N(_08914_),
    .Q(\am_sdr0.cic0.integ1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[15]$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net636),
    .D(_00313_),
    .Q_N(_08913_),
    .Q(\am_sdr0.cic0.integ1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[16]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net637),
    .D(_00314_),
    .Q_N(_08912_),
    .Q(\am_sdr0.cic0.integ1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[17]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net638),
    .D(_00315_),
    .Q_N(_08911_),
    .Q(\am_sdr0.cic0.integ1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[18]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net639),
    .D(_00316_),
    .Q_N(_08910_),
    .Q(\am_sdr0.cic0.integ1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[19]$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net640),
    .D(_00317_),
    .Q_N(_08909_),
    .Q(\am_sdr0.cic0.integ1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[1]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net641),
    .D(_00318_),
    .Q_N(_08908_),
    .Q(\am_sdr0.cic0.integ1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[20]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net642),
    .D(_00319_),
    .Q_N(_08907_),
    .Q(\am_sdr0.cic0.integ1[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[21]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net643),
    .D(_00320_),
    .Q_N(_08906_),
    .Q(\am_sdr0.cic0.integ1[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[22]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net644),
    .D(_00321_),
    .Q_N(_08905_),
    .Q(\am_sdr0.cic0.integ1[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[23]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net645),
    .D(_00322_),
    .Q_N(_08904_),
    .Q(\am_sdr0.cic0.integ1[23] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[24]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net646),
    .D(_00323_),
    .Q_N(_08903_),
    .Q(\am_sdr0.cic0.integ1[24] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[25]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net647),
    .D(_00324_),
    .Q_N(_08902_),
    .Q(\am_sdr0.cic0.integ1[25] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[2]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net648),
    .D(_00325_),
    .Q_N(_08901_),
    .Q(\am_sdr0.cic0.integ1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[3]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net649),
    .D(_00326_),
    .Q_N(_08900_),
    .Q(\am_sdr0.cic0.integ1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[4]$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net650),
    .D(_00327_),
    .Q_N(_08899_),
    .Q(\am_sdr0.cic0.integ1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[5]$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net651),
    .D(_00328_),
    .Q_N(_08898_),
    .Q(\am_sdr0.cic0.integ1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[6]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net652),
    .D(_00329_),
    .Q_N(_08897_),
    .Q(\am_sdr0.cic0.integ1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[7]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net653),
    .D(_00330_),
    .Q_N(_08896_),
    .Q(\am_sdr0.cic0.integ1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[8]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net654),
    .D(_00331_),
    .Q_N(_08895_),
    .Q(\am_sdr0.cic0.integ1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ1[9]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net655),
    .D(_00332_),
    .Q_N(_08894_),
    .Q(\am_sdr0.cic0.integ1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[0]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net656),
    .D(_00333_),
    .Q_N(_08893_),
    .Q(\am_sdr0.cic0.integ2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[10]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net657),
    .D(_00334_),
    .Q_N(_08892_),
    .Q(\am_sdr0.cic0.integ2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[11]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net658),
    .D(_00335_),
    .Q_N(_08891_),
    .Q(\am_sdr0.cic0.integ2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[12]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net659),
    .D(_00336_),
    .Q_N(_08890_),
    .Q(\am_sdr0.cic0.integ2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[13]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net660),
    .D(_00337_),
    .Q_N(_08889_),
    .Q(\am_sdr0.cic0.integ2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[14]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net661),
    .D(_00338_),
    .Q_N(_08888_),
    .Q(\am_sdr0.cic0.integ2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[15]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net662),
    .D(_00339_),
    .Q_N(_08887_),
    .Q(\am_sdr0.cic0.integ2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[16]$_SDFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net663),
    .D(_00340_),
    .Q_N(_08886_),
    .Q(\am_sdr0.cic0.integ2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[17]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net664),
    .D(_00341_),
    .Q_N(_08885_),
    .Q(\am_sdr0.cic0.integ2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[18]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net665),
    .D(_00342_),
    .Q_N(_08884_),
    .Q(\am_sdr0.cic0.integ2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[19]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net666),
    .D(_00343_),
    .Q_N(_08883_),
    .Q(\am_sdr0.cic0.integ2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[1]$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net667),
    .D(_00344_),
    .Q_N(_08882_),
    .Q(\am_sdr0.cic0.integ2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[20]$_SDFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net668),
    .D(_00345_),
    .Q_N(_08881_),
    .Q(\am_sdr0.cic0.integ2[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[21]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net669),
    .D(_00346_),
    .Q_N(_08880_),
    .Q(\am_sdr0.cic0.integ2[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[22]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net670),
    .D(_00347_),
    .Q_N(_08879_),
    .Q(\am_sdr0.cic0.integ2[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[2]$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net671),
    .D(_00348_),
    .Q_N(_08878_),
    .Q(\am_sdr0.cic0.integ2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[3]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net672),
    .D(_00349_),
    .Q_N(_08877_),
    .Q(\am_sdr0.cic0.integ2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[4]$_SDFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net673),
    .D(_00350_),
    .Q_N(_08876_),
    .Q(\am_sdr0.cic0.integ2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[5]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net674),
    .D(_00351_),
    .Q_N(_08875_),
    .Q(\am_sdr0.cic0.integ2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[6]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net675),
    .D(_00352_),
    .Q_N(_08874_),
    .Q(\am_sdr0.cic0.integ2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[7]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net676),
    .D(_00353_),
    .Q_N(_08873_),
    .Q(\am_sdr0.cic0.integ2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[8]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net677),
    .D(_00354_),
    .Q_N(_08872_),
    .Q(\am_sdr0.cic0.integ2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ2[9]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net678),
    .D(_00355_),
    .Q_N(_08871_),
    .Q(\am_sdr0.cic0.integ2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[0]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net679),
    .D(_00356_),
    .Q_N(_08870_),
    .Q(\am_sdr0.cic0.integ3[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[10]$_SDFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net680),
    .D(_00357_),
    .Q_N(_08869_),
    .Q(\am_sdr0.cic0.integ3[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[11]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net681),
    .D(_00358_),
    .Q_N(_08868_),
    .Q(\am_sdr0.cic0.integ3[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[12]$_SDFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net682),
    .D(_00359_),
    .Q_N(_08867_),
    .Q(\am_sdr0.cic0.integ3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[13]$_SDFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net683),
    .D(_00360_),
    .Q_N(_08866_),
    .Q(\am_sdr0.cic0.integ3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[14]$_SDFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net684),
    .D(_00361_),
    .Q_N(_08865_),
    .Q(\am_sdr0.cic0.integ3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[15]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net685),
    .D(_00362_),
    .Q_N(_08864_),
    .Q(\am_sdr0.cic0.integ3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[16]$_SDFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net686),
    .D(_00363_),
    .Q_N(_08863_),
    .Q(\am_sdr0.cic0.integ3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[17]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net687),
    .D(_00364_),
    .Q_N(_08862_),
    .Q(\am_sdr0.cic0.integ3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[18]$_SDFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net688),
    .D(_00365_),
    .Q_N(_08861_),
    .Q(\am_sdr0.cic0.integ3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[19]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net689),
    .D(_00366_),
    .Q_N(_08860_),
    .Q(\am_sdr0.cic0.integ3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[1]$_SDFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net690),
    .D(_00367_),
    .Q_N(_08859_),
    .Q(\am_sdr0.cic0.integ3[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[2]$_SDFF_PN0_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net691),
    .D(_00368_),
    .Q_N(_08858_),
    .Q(\am_sdr0.cic0.integ3[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[3]$_SDFF_PN0_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net692),
    .D(_00369_),
    .Q_N(_08857_),
    .Q(\am_sdr0.cic0.integ3[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[4]$_SDFF_PN0_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net693),
    .D(_00370_),
    .Q_N(_08856_),
    .Q(\am_sdr0.cic0.integ3[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[5]$_SDFF_PN0_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net694),
    .D(_00371_),
    .Q_N(_08855_),
    .Q(\am_sdr0.cic0.integ3[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[6]$_SDFF_PN0_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net695),
    .D(_00372_),
    .Q_N(_08854_),
    .Q(\am_sdr0.cic0.integ3[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[7]$_SDFF_PN0_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net696),
    .D(_00373_),
    .Q_N(_08853_),
    .Q(\am_sdr0.cic0.integ3[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[8]$_SDFF_PN0_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net697),
    .D(_00374_),
    .Q_N(_08852_),
    .Q(\am_sdr0.cic0.integ3[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ3[9]$_SDFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net698),
    .D(_00375_),
    .Q_N(_08851_),
    .Q(\am_sdr0.cic0.integ3[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[0]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net699),
    .D(_00376_),
    .Q_N(_08850_),
    .Q(\am_sdr0.cic0.integ_sample[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net700),
    .D(_00377_),
    .Q_N(_08849_),
    .Q(\am_sdr0.cic0.integ_sample[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net701),
    .D(_00378_),
    .Q_N(_08848_),
    .Q(\am_sdr0.cic0.integ_sample[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[12]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net702),
    .D(_00379_),
    .Q_N(_08847_),
    .Q(\am_sdr0.cic0.integ_sample[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[13]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net703),
    .D(_00380_),
    .Q_N(_08846_),
    .Q(\am_sdr0.cic0.integ_sample[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[14]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net704),
    .D(_00381_),
    .Q_N(_08845_),
    .Q(\am_sdr0.cic0.integ_sample[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[15]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net705),
    .D(_00382_),
    .Q_N(_08844_),
    .Q(\am_sdr0.cic0.integ_sample[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net706),
    .D(_00383_),
    .Q_N(_08843_),
    .Q(\am_sdr0.cic0.integ_sample[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[17]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net707),
    .D(_00384_),
    .Q_N(_08842_),
    .Q(\am_sdr0.cic0.integ_sample[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[18]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net708),
    .D(_00385_),
    .Q_N(_08841_),
    .Q(\am_sdr0.cic0.integ_sample[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[19]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net709),
    .D(_00386_),
    .Q_N(_08840_),
    .Q(\am_sdr0.cic0.integ_sample[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[1]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net710),
    .D(_00387_),
    .Q_N(_08839_),
    .Q(\am_sdr0.cic0.integ_sample[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[2]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net711),
    .D(_00388_),
    .Q_N(_08838_),
    .Q(\am_sdr0.cic0.integ_sample[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[3]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net712),
    .D(_00389_),
    .Q_N(_08837_),
    .Q(\am_sdr0.cic0.integ_sample[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net713),
    .D(_00390_),
    .Q_N(_08836_),
    .Q(\am_sdr0.cic0.integ_sample[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[5]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net714),
    .D(_00391_),
    .Q_N(_08835_),
    .Q(\am_sdr0.cic0.integ_sample[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[6]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net715),
    .D(_00392_),
    .Q_N(_08834_),
    .Q(\am_sdr0.cic0.integ_sample[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[7]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net716),
    .D(_00393_),
    .Q_N(_08833_),
    .Q(\am_sdr0.cic0.integ_sample[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[8]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net717),
    .D(_00394_),
    .Q_N(_08832_),
    .Q(\am_sdr0.cic0.integ_sample[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.integ_sample[9]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net718),
    .D(_00395_),
    .Q_N(_08831_),
    .Q(\am_sdr0.cic0.integ_sample[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.out_tick$_SDFF_PN0_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net719),
    .D(_00396_),
    .Q_N(_08830_),
    .Q(\am_sdr0.cic0.out_tick ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.sample$_SDFF_PN0_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net720),
    .D(net21),
    .Q_N(_08829_),
    .Q(\am_sdr0.cic0.sample ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net721),
    .D(_00398_),
    .Q_N(_08828_),
    .Q(\am_sdr0.cic0.x_out[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net722),
    .D(_00399_),
    .Q_N(_08827_),
    .Q(\am_sdr0.cic0.x_out[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net723),
    .D(_00400_),
    .Q_N(_08826_),
    .Q(\am_sdr0.cic0.x_out[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net724),
    .D(_00401_),
    .Q_N(_08825_),
    .Q(\am_sdr0.cic0.x_out[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net725),
    .D(_00402_),
    .Q_N(_08824_),
    .Q(\am_sdr0.cic0.x_out[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net726),
    .D(_00403_),
    .Q_N(_08823_),
    .Q(\am_sdr0.cic0.x_out[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net727),
    .D(_00404_),
    .Q_N(_08822_),
    .Q(\am_sdr0.cic0.x_out[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic0.x_out[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net728),
    .D(_00405_),
    .Q_N(_08821_),
    .Q(\am_sdr0.cic0.x_out[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net729),
    .D(_00406_),
    .Q_N(_08820_),
    .Q(\am_sdr0.cic1.comb1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net730),
    .D(_00407_),
    .Q_N(_08819_),
    .Q(\am_sdr0.cic1.comb1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net731),
    .D(_00408_),
    .Q_N(_08818_),
    .Q(\am_sdr0.cic1.comb1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net732),
    .D(_00409_),
    .Q_N(_08817_),
    .Q(\am_sdr0.cic1.comb1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net733),
    .D(_00410_),
    .Q_N(_08816_),
    .Q(\am_sdr0.cic1.comb1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net734),
    .D(_00411_),
    .Q_N(_08815_),
    .Q(\am_sdr0.cic1.comb1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net735),
    .D(_00412_),
    .Q_N(_08814_),
    .Q(\am_sdr0.cic1.comb1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net736),
    .D(_00413_),
    .Q_N(_08813_),
    .Q(\am_sdr0.cic1.comb1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net737),
    .D(_00414_),
    .Q_N(_08812_),
    .Q(\am_sdr0.cic1.comb1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net738),
    .D(_00415_),
    .Q_N(_08811_),
    .Q(\am_sdr0.cic1.comb1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net739),
    .D(_00416_),
    .Q_N(_08810_),
    .Q(\am_sdr0.cic1.comb1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net740),
    .D(_00417_),
    .Q_N(_08809_),
    .Q(\am_sdr0.cic1.comb1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net741),
    .D(_00418_),
    .Q_N(_08808_),
    .Q(\am_sdr0.cic1.comb1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net742),
    .D(_00419_),
    .Q_N(_08807_),
    .Q(\am_sdr0.cic1.comb1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net743),
    .D(_00420_),
    .Q_N(_08806_),
    .Q(\am_sdr0.cic1.comb1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net744),
    .D(_00421_),
    .Q_N(_08805_),
    .Q(\am_sdr0.cic1.comb1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net745),
    .D(_00422_),
    .Q_N(_08804_),
    .Q(\am_sdr0.cic1.comb1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net746),
    .D(_00423_),
    .Q_N(_08803_),
    .Q(\am_sdr0.cic1.comb1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net747),
    .D(_00424_),
    .Q_N(_08802_),
    .Q(\am_sdr0.cic1.comb1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net748),
    .D(_00425_),
    .Q_N(_08801_),
    .Q(\am_sdr0.cic1.comb1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net749),
    .D(_00426_),
    .Q_N(_08800_),
    .Q(\am_sdr0.cic1.comb1_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net750),
    .D(_00427_),
    .Q_N(_08799_),
    .Q(\am_sdr0.cic1.comb1_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net751),
    .D(_00428_),
    .Q_N(_08798_),
    .Q(\am_sdr0.cic1.comb1_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net752),
    .D(_00429_),
    .Q_N(_08797_),
    .Q(\am_sdr0.cic1.comb1_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net753),
    .D(_00430_),
    .Q_N(_08796_),
    .Q(\am_sdr0.cic1.comb1_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net754),
    .D(_00431_),
    .Q_N(_08795_),
    .Q(\am_sdr0.cic1.comb1_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net755),
    .D(_00432_),
    .Q_N(_08794_),
    .Q(\am_sdr0.cic1.comb1_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net756),
    .D(_00433_),
    .Q_N(_08793_),
    .Q(\am_sdr0.cic1.comb1_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net757),
    .D(_00434_),
    .Q_N(_08792_),
    .Q(\am_sdr0.cic1.comb1_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net758),
    .D(_00435_),
    .Q_N(_08791_),
    .Q(\am_sdr0.cic1.comb1_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net759),
    .D(_00436_),
    .Q_N(_08790_),
    .Q(\am_sdr0.cic1.comb1_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net760),
    .D(_00437_),
    .Q_N(_08789_),
    .Q(\am_sdr0.cic1.comb1_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net761),
    .D(_00438_),
    .Q_N(_08788_),
    .Q(\am_sdr0.cic1.comb1_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net762),
    .D(_00439_),
    .Q_N(_08787_),
    .Q(\am_sdr0.cic1.comb1_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net763),
    .D(_00440_),
    .Q_N(_08786_),
    .Q(\am_sdr0.cic1.comb1_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net764),
    .D(_00441_),
    .Q_N(_08785_),
    .Q(\am_sdr0.cic1.comb1_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net765),
    .D(_00442_),
    .Q_N(_08784_),
    .Q(\am_sdr0.cic1.comb1_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net766),
    .D(_00443_),
    .Q_N(_08783_),
    .Q(\am_sdr0.cic1.comb1_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net767),
    .D(_00444_),
    .Q_N(_08782_),
    .Q(\am_sdr0.cic1.comb1_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb1_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net768),
    .D(_00445_),
    .Q_N(_08781_),
    .Q(\am_sdr0.cic1.comb1_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net769),
    .D(_00446_),
    .Q_N(_08780_),
    .Q(\am_sdr0.cic1.comb2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net770),
    .D(_00447_),
    .Q_N(_08779_),
    .Q(\am_sdr0.cic1.comb2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net771),
    .D(_00448_),
    .Q_N(_08778_),
    .Q(\am_sdr0.cic1.comb2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net772),
    .D(_00449_),
    .Q_N(_08777_),
    .Q(\am_sdr0.cic1.comb2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net773),
    .D(_00450_),
    .Q_N(_08776_),
    .Q(\am_sdr0.cic1.comb2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net774),
    .D(_00451_),
    .Q_N(_08775_),
    .Q(\am_sdr0.cic1.comb2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net775),
    .D(_00452_),
    .Q_N(_08774_),
    .Q(\am_sdr0.cic1.comb2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net776),
    .D(_00453_),
    .Q_N(_08773_),
    .Q(\am_sdr0.cic1.comb2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net777),
    .D(_00454_),
    .Q_N(_08772_),
    .Q(\am_sdr0.cic1.comb2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net778),
    .D(_00455_),
    .Q_N(_08771_),
    .Q(\am_sdr0.cic1.comb2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net779),
    .D(_00456_),
    .Q_N(_08770_),
    .Q(\am_sdr0.cic1.comb2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net780),
    .D(_00457_),
    .Q_N(_08769_),
    .Q(\am_sdr0.cic1.comb2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net781),
    .D(_00458_),
    .Q_N(_08768_),
    .Q(\am_sdr0.cic1.comb2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net782),
    .D(_00459_),
    .Q_N(_08767_),
    .Q(\am_sdr0.cic1.comb2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net783),
    .D(_00460_),
    .Q_N(_08766_),
    .Q(\am_sdr0.cic1.comb2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net784),
    .D(_00461_),
    .Q_N(_08765_),
    .Q(\am_sdr0.cic1.comb2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net785),
    .D(_00462_),
    .Q_N(_08764_),
    .Q(\am_sdr0.cic1.comb2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net786),
    .D(_00463_),
    .Q_N(_08763_),
    .Q(\am_sdr0.cic1.comb2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net787),
    .D(_00464_),
    .Q_N(_08762_),
    .Q(\am_sdr0.cic1.comb2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net788),
    .D(_00465_),
    .Q_N(_08761_),
    .Q(\am_sdr0.cic1.comb2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net789),
    .D(_00466_),
    .Q_N(_08760_),
    .Q(\am_sdr0.cic1.comb2_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net790),
    .D(_00467_),
    .Q_N(_08759_),
    .Q(\am_sdr0.cic1.comb2_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net791),
    .D(_00468_),
    .Q_N(_08758_),
    .Q(\am_sdr0.cic1.comb2_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net792),
    .D(_00469_),
    .Q_N(_08757_),
    .Q(\am_sdr0.cic1.comb2_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net793),
    .D(_00470_),
    .Q_N(_08756_),
    .Q(\am_sdr0.cic1.comb2_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net794),
    .D(_00471_),
    .Q_N(_08755_),
    .Q(\am_sdr0.cic1.comb2_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net795),
    .D(_00472_),
    .Q_N(_08754_),
    .Q(\am_sdr0.cic1.comb2_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net796),
    .D(_00473_),
    .Q_N(_08753_),
    .Q(\am_sdr0.cic1.comb2_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net797),
    .D(_00474_),
    .Q_N(_08752_),
    .Q(\am_sdr0.cic1.comb2_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net798),
    .D(_00475_),
    .Q_N(_08751_),
    .Q(\am_sdr0.cic1.comb2_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net799),
    .D(_00476_),
    .Q_N(_08750_),
    .Q(\am_sdr0.cic1.comb2_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net800),
    .D(_00477_),
    .Q_N(_08749_),
    .Q(\am_sdr0.cic1.comb2_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net801),
    .D(_00478_),
    .Q_N(_08748_),
    .Q(\am_sdr0.cic1.comb2_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net802),
    .D(_00479_),
    .Q_N(_08747_),
    .Q(\am_sdr0.cic1.comb2_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net803),
    .D(_00480_),
    .Q_N(_08746_),
    .Q(\am_sdr0.cic1.comb2_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net804),
    .D(_00481_),
    .Q_N(_08745_),
    .Q(\am_sdr0.cic1.comb2_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net805),
    .D(_00482_),
    .Q_N(_08744_),
    .Q(\am_sdr0.cic1.comb2_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net806),
    .D(_00483_),
    .Q_N(_08743_),
    .Q(\am_sdr0.cic1.comb2_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net807),
    .D(_00484_),
    .Q_N(_08742_),
    .Q(\am_sdr0.cic1.comb2_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb2_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net808),
    .D(_00485_),
    .Q_N(_08741_),
    .Q(\am_sdr0.cic1.comb2_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net809),
    .D(_00486_),
    .Q_N(_08740_),
    .Q(\am_sdr0.cic1.comb3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net810),
    .D(_00487_),
    .Q_N(_08739_),
    .Q(\am_sdr0.cic1.comb3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net811),
    .D(_00488_),
    .Q_N(_08738_),
    .Q(\am_sdr0.cic1.comb3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net812),
    .D(_00489_),
    .Q_N(_08737_),
    .Q(\am_sdr0.cic1.comb3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net813),
    .D(_00490_),
    .Q_N(_08736_),
    .Q(\am_sdr0.cic1.comb3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net814),
    .D(_00491_),
    .Q_N(_08735_),
    .Q(\am_sdr0.cic1.comb3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net815),
    .D(_00492_),
    .Q_N(_08734_),
    .Q(\am_sdr0.cic1.comb3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net816),
    .D(_00493_),
    .Q_N(_08733_),
    .Q(\am_sdr0.cic1.comb3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net817),
    .D(_00494_),
    .Q_N(_08732_),
    .Q(\am_sdr0.cic1.comb3_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net818),
    .D(_00495_),
    .Q_N(_08731_),
    .Q(\am_sdr0.cic1.comb3_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net819),
    .D(_00496_),
    .Q_N(_08730_),
    .Q(\am_sdr0.cic1.comb3_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net820),
    .D(_00497_),
    .Q_N(_08729_),
    .Q(\am_sdr0.cic1.comb3_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net821),
    .D(_00498_),
    .Q_N(_08728_),
    .Q(\am_sdr0.cic1.comb3_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net822),
    .D(_00499_),
    .Q_N(_08727_),
    .Q(\am_sdr0.cic1.comb3_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net823),
    .D(_00500_),
    .Q_N(_08726_),
    .Q(\am_sdr0.cic1.comb3_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net824),
    .D(_00501_),
    .Q_N(_08725_),
    .Q(\am_sdr0.cic1.comb3_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net825),
    .D(_00502_),
    .Q_N(_08724_),
    .Q(\am_sdr0.cic1.comb3_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net826),
    .D(_00503_),
    .Q_N(_08723_),
    .Q(\am_sdr0.cic1.comb3_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net827),
    .D(_00504_),
    .Q_N(_08722_),
    .Q(\am_sdr0.cic1.comb3_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net828),
    .D(_00505_),
    .Q_N(_08721_),
    .Q(\am_sdr0.cic1.comb3_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net829),
    .D(_00506_),
    .Q_N(_08720_),
    .Q(\am_sdr0.cic1.comb3_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net830),
    .D(_00507_),
    .Q_N(_08719_),
    .Q(\am_sdr0.cic1.comb3_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net831),
    .D(_00508_),
    .Q_N(_08718_),
    .Q(\am_sdr0.cic1.comb3_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net832),
    .D(_00509_),
    .Q_N(_08717_),
    .Q(\am_sdr0.cic1.comb3_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net833),
    .D(_00510_),
    .Q_N(_08716_),
    .Q(\am_sdr0.cic1.comb3_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net834),
    .D(_00511_),
    .Q_N(_08715_),
    .Q(\am_sdr0.cic1.comb3_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net835),
    .D(_00512_),
    .Q_N(_08714_),
    .Q(\am_sdr0.cic1.comb3_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.comb3_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net836),
    .D(_00513_),
    .Q_N(_08713_),
    .Q(\am_sdr0.cic1.comb3_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[0]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net837),
    .D(_00514_),
    .Q_N(_00073_),
    .Q(\am_sdr0.cic1.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[1]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net838),
    .D(_00515_),
    .Q_N(_08712_),
    .Q(\am_sdr0.cic1.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[2]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net839),
    .D(_00516_),
    .Q_N(_08711_),
    .Q(\am_sdr0.cic1.count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[3]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net840),
    .D(_00517_),
    .Q_N(_08710_),
    .Q(\am_sdr0.cic1.count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[4]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net841),
    .D(_00518_),
    .Q_N(_08709_),
    .Q(\am_sdr0.cic1.count[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[5]$_SDFF_PP0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net842),
    .D(_00519_),
    .Q_N(_08708_),
    .Q(\am_sdr0.cic1.count[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[6]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net843),
    .D(_00520_),
    .Q_N(_08707_),
    .Q(\am_sdr0.cic1.count[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.count[7]$_SDFF_PP0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net844),
    .D(_00521_),
    .Q_N(_08706_),
    .Q(\am_sdr0.cic1.count[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[0]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net845),
    .D(_00522_),
    .Q_N(_08705_),
    .Q(\am_sdr0.cic1.integ1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[10]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net846),
    .D(_00523_),
    .Q_N(_08704_),
    .Q(\am_sdr0.cic1.integ1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[11]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net847),
    .D(_00524_),
    .Q_N(_08703_),
    .Q(\am_sdr0.cic1.integ1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[12]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net848),
    .D(_00525_),
    .Q_N(_08702_),
    .Q(\am_sdr0.cic1.integ1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[13]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net849),
    .D(_00526_),
    .Q_N(_08701_),
    .Q(\am_sdr0.cic1.integ1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[14]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net850),
    .D(_00527_),
    .Q_N(_08700_),
    .Q(\am_sdr0.cic1.integ1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[15]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net851),
    .D(_00528_),
    .Q_N(_08699_),
    .Q(\am_sdr0.cic1.integ1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[16]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net852),
    .D(_00529_),
    .Q_N(_08698_),
    .Q(\am_sdr0.cic1.integ1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[17]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net853),
    .D(_00530_),
    .Q_N(_08697_),
    .Q(\am_sdr0.cic1.integ1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[18]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net854),
    .D(_00531_),
    .Q_N(_08696_),
    .Q(\am_sdr0.cic1.integ1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[19]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net855),
    .D(_00532_),
    .Q_N(_08695_),
    .Q(\am_sdr0.cic1.integ1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[1]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net856),
    .D(_00533_),
    .Q_N(_08694_),
    .Q(\am_sdr0.cic1.integ1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[20]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net857),
    .D(_00534_),
    .Q_N(_08693_),
    .Q(\am_sdr0.cic1.integ1[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[21]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net858),
    .D(_00535_),
    .Q_N(_08692_),
    .Q(\am_sdr0.cic1.integ1[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[22]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net859),
    .D(_00536_),
    .Q_N(_08691_),
    .Q(\am_sdr0.cic1.integ1[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[23]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net860),
    .D(_00537_),
    .Q_N(_08690_),
    .Q(\am_sdr0.cic1.integ1[23] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[24]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net861),
    .D(_00538_),
    .Q_N(_08689_),
    .Q(\am_sdr0.cic1.integ1[24] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[25]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net862),
    .D(_00539_),
    .Q_N(_08688_),
    .Q(\am_sdr0.cic1.integ1[25] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[2]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net863),
    .D(_00540_),
    .Q_N(_08687_),
    .Q(\am_sdr0.cic1.integ1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[3]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net864),
    .D(_00541_),
    .Q_N(_08686_),
    .Q(\am_sdr0.cic1.integ1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[4]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net865),
    .D(_00542_),
    .Q_N(_08685_),
    .Q(\am_sdr0.cic1.integ1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[5]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net866),
    .D(_00543_),
    .Q_N(_08684_),
    .Q(\am_sdr0.cic1.integ1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[6]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net867),
    .D(_00544_),
    .Q_N(_08683_),
    .Q(\am_sdr0.cic1.integ1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[7]$_SDFF_PN0_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net868),
    .D(_00545_),
    .Q_N(_08682_),
    .Q(\am_sdr0.cic1.integ1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[8]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net869),
    .D(_00546_),
    .Q_N(_08681_),
    .Q(\am_sdr0.cic1.integ1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ1[9]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net870),
    .D(_00547_),
    .Q_N(_08680_),
    .Q(\am_sdr0.cic1.integ1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[0]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net871),
    .D(_00548_),
    .Q_N(_08679_),
    .Q(\am_sdr0.cic1.integ2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[10]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net872),
    .D(_00549_),
    .Q_N(_08678_),
    .Q(\am_sdr0.cic1.integ2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[11]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net873),
    .D(_00550_),
    .Q_N(_08677_),
    .Q(\am_sdr0.cic1.integ2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[12]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net874),
    .D(_00551_),
    .Q_N(_08676_),
    .Q(\am_sdr0.cic1.integ2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[13]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net875),
    .D(_00552_),
    .Q_N(_08675_),
    .Q(\am_sdr0.cic1.integ2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[14]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net876),
    .D(_00553_),
    .Q_N(_08674_),
    .Q(\am_sdr0.cic1.integ2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[15]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net877),
    .D(_00554_),
    .Q_N(_08673_),
    .Q(\am_sdr0.cic1.integ2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[16]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net878),
    .D(_00555_),
    .Q_N(_08672_),
    .Q(\am_sdr0.cic1.integ2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[17]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net879),
    .D(_00556_),
    .Q_N(_08671_),
    .Q(\am_sdr0.cic1.integ2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[18]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net880),
    .D(_00557_),
    .Q_N(_08670_),
    .Q(\am_sdr0.cic1.integ2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[19]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net881),
    .D(_00558_),
    .Q_N(_08669_),
    .Q(\am_sdr0.cic1.integ2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[1]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net882),
    .D(_00559_),
    .Q_N(_08668_),
    .Q(\am_sdr0.cic1.integ2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[20]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net883),
    .D(_00560_),
    .Q_N(_08667_),
    .Q(\am_sdr0.cic1.integ2[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[21]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net884),
    .D(_00561_),
    .Q_N(_08666_),
    .Q(\am_sdr0.cic1.integ2[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[22]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net885),
    .D(_00562_),
    .Q_N(_08665_),
    .Q(\am_sdr0.cic1.integ2[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[2]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net886),
    .D(_00563_),
    .Q_N(_08664_),
    .Q(\am_sdr0.cic1.integ2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[3]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net887),
    .D(_00564_),
    .Q_N(_08663_),
    .Q(\am_sdr0.cic1.integ2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[4]$_SDFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net888),
    .D(_00565_),
    .Q_N(_08662_),
    .Q(\am_sdr0.cic1.integ2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[5]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net889),
    .D(_00566_),
    .Q_N(_08661_),
    .Q(\am_sdr0.cic1.integ2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[6]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net890),
    .D(_00567_),
    .Q_N(_08660_),
    .Q(\am_sdr0.cic1.integ2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[7]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net891),
    .D(_00568_),
    .Q_N(_08659_),
    .Q(\am_sdr0.cic1.integ2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[8]$_SDFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net892),
    .D(_00569_),
    .Q_N(_08658_),
    .Q(\am_sdr0.cic1.integ2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ2[9]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net893),
    .D(_00570_),
    .Q_N(_08657_),
    .Q(\am_sdr0.cic1.integ2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[0]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net894),
    .D(_00571_),
    .Q_N(_08656_),
    .Q(\am_sdr0.cic1.integ3[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[10]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net895),
    .D(_00572_),
    .Q_N(_08655_),
    .Q(\am_sdr0.cic1.integ3[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[11]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net896),
    .D(_00573_),
    .Q_N(_08654_),
    .Q(\am_sdr0.cic1.integ3[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[12]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net897),
    .D(_00574_),
    .Q_N(_08653_),
    .Q(\am_sdr0.cic1.integ3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[13]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net898),
    .D(_00575_),
    .Q_N(_08652_),
    .Q(\am_sdr0.cic1.integ3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[14]$_SDFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net899),
    .D(_00576_),
    .Q_N(_08651_),
    .Q(\am_sdr0.cic1.integ3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[15]$_SDFF_PN0_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net900),
    .D(_00577_),
    .Q_N(_08650_),
    .Q(\am_sdr0.cic1.integ3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[16]$_SDFF_PN0_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net901),
    .D(_00578_),
    .Q_N(_08649_),
    .Q(\am_sdr0.cic1.integ3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[17]$_SDFF_PN0_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net902),
    .D(_00579_),
    .Q_N(_08648_),
    .Q(\am_sdr0.cic1.integ3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[18]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net903),
    .D(_00580_),
    .Q_N(_08647_),
    .Q(\am_sdr0.cic1.integ3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[19]$_SDFF_PN0_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net904),
    .D(_00581_),
    .Q_N(_08646_),
    .Q(\am_sdr0.cic1.integ3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[1]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net905),
    .D(_00582_),
    .Q_N(_08645_),
    .Q(\am_sdr0.cic1.integ3[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[2]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net906),
    .D(_00583_),
    .Q_N(_08644_),
    .Q(\am_sdr0.cic1.integ3[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[3]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net907),
    .D(_00584_),
    .Q_N(_08643_),
    .Q(\am_sdr0.cic1.integ3[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[4]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net908),
    .D(_00585_),
    .Q_N(_08642_),
    .Q(\am_sdr0.cic1.integ3[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[5]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net909),
    .D(_00586_),
    .Q_N(_08641_),
    .Q(\am_sdr0.cic1.integ3[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[6]$_SDFF_PN0_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net910),
    .D(_00587_),
    .Q_N(_08640_),
    .Q(\am_sdr0.cic1.integ3[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[7]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net911),
    .D(_00588_),
    .Q_N(_08639_),
    .Q(\am_sdr0.cic1.integ3[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[8]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net912),
    .D(_00589_),
    .Q_N(_08638_),
    .Q(\am_sdr0.cic1.integ3[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ3[9]$_SDFF_PN0_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net913),
    .D(_00590_),
    .Q_N(_08637_),
    .Q(\am_sdr0.cic1.integ3[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net914),
    .D(_00591_),
    .Q_N(_08636_),
    .Q(\am_sdr0.cic1.integ_sample[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[10]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net915),
    .D(_00592_),
    .Q_N(_08635_),
    .Q(\am_sdr0.cic1.integ_sample[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[11]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net916),
    .D(_00593_),
    .Q_N(_08634_),
    .Q(\am_sdr0.cic1.integ_sample[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[12]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net917),
    .D(_00594_),
    .Q_N(_08633_),
    .Q(\am_sdr0.cic1.integ_sample[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[13]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net918),
    .D(_00595_),
    .Q_N(_08632_),
    .Q(\am_sdr0.cic1.integ_sample[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[14]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net919),
    .D(_00596_),
    .Q_N(_08631_),
    .Q(\am_sdr0.cic1.integ_sample[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[15]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net920),
    .D(_00597_),
    .Q_N(_08630_),
    .Q(\am_sdr0.cic1.integ_sample[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[16]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net921),
    .D(_00598_),
    .Q_N(_08629_),
    .Q(\am_sdr0.cic1.integ_sample[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[17]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net922),
    .D(_00599_),
    .Q_N(_08628_),
    .Q(\am_sdr0.cic1.integ_sample[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[18]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net923),
    .D(_00600_),
    .Q_N(_08627_),
    .Q(\am_sdr0.cic1.integ_sample[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[19]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net924),
    .D(_00601_),
    .Q_N(_08626_),
    .Q(\am_sdr0.cic1.integ_sample[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net925),
    .D(_00602_),
    .Q_N(_08625_),
    .Q(\am_sdr0.cic1.integ_sample[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net926),
    .D(_00603_),
    .Q_N(_08624_),
    .Q(\am_sdr0.cic1.integ_sample[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net927),
    .D(_00604_),
    .Q_N(_08623_),
    .Q(\am_sdr0.cic1.integ_sample[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[4]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net928),
    .D(_00605_),
    .Q_N(_08622_),
    .Q(\am_sdr0.cic1.integ_sample[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net929),
    .D(_00606_),
    .Q_N(_08621_),
    .Q(\am_sdr0.cic1.integ_sample[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net930),
    .D(_00607_),
    .Q_N(_08620_),
    .Q(\am_sdr0.cic1.integ_sample[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net931),
    .D(_00608_),
    .Q_N(_08619_),
    .Q(\am_sdr0.cic1.integ_sample[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[8]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net932),
    .D(_00609_),
    .Q_N(_08618_),
    .Q(\am_sdr0.cic1.integ_sample[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.integ_sample[9]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net933),
    .D(_00610_),
    .Q_N(_08617_),
    .Q(\am_sdr0.cic1.integ_sample[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.out_tick$_SDFF_PN0_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net934),
    .D(_00611_),
    .Q_N(_08616_),
    .Q(\am_sdr0.cic1.out_tick ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.sample$_SDFF_PN0_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net935),
    .D(net27),
    .Q_N(_08615_),
    .Q(\am_sdr0.cic1.sample ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net936),
    .D(_00613_),
    .Q_N(_08614_),
    .Q(\am_sdr0.cic1.x_out[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net937),
    .D(_00614_),
    .Q_N(_08613_),
    .Q(\am_sdr0.cic1.x_out[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net938),
    .D(_00615_),
    .Q_N(_08612_),
    .Q(\am_sdr0.cic1.x_out[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net939),
    .D(_00616_),
    .Q_N(_08611_),
    .Q(\am_sdr0.cic1.x_out[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net940),
    .D(_00617_),
    .Q_N(_08610_),
    .Q(\am_sdr0.cic1.x_out[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net941),
    .D(_00618_),
    .Q_N(_08609_),
    .Q(\am_sdr0.cic1.x_out[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net942),
    .D(_00619_),
    .Q_N(_08608_),
    .Q(\am_sdr0.cic1.x_out[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic1.x_out[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net943),
    .D(_00620_),
    .Q_N(_08607_),
    .Q(\am_sdr0.cic1.x_out[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net944),
    .D(_00621_),
    .Q_N(_08606_),
    .Q(\am_sdr0.cic2.comb1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net945),
    .D(_00622_),
    .Q_N(_08605_),
    .Q(\am_sdr0.cic2.comb1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net946),
    .D(_00623_),
    .Q_N(_08604_),
    .Q(\am_sdr0.cic2.comb1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net947),
    .D(_00624_),
    .Q_N(_08603_),
    .Q(\am_sdr0.cic2.comb1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net948),
    .D(_00625_),
    .Q_N(_08602_),
    .Q(\am_sdr0.cic2.comb1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net949),
    .D(_00626_),
    .Q_N(_08601_),
    .Q(\am_sdr0.cic2.comb1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net950),
    .D(_00627_),
    .Q_N(_08600_),
    .Q(\am_sdr0.cic2.comb1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net951),
    .D(_00628_),
    .Q_N(_08599_),
    .Q(\am_sdr0.cic2.comb1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net952),
    .D(_00629_),
    .Q_N(_08598_),
    .Q(\am_sdr0.cic2.comb1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net953),
    .D(_00630_),
    .Q_N(_08597_),
    .Q(\am_sdr0.cic2.comb1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net954),
    .D(_00631_),
    .Q_N(_08596_),
    .Q(\am_sdr0.cic2.comb1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net955),
    .D(_00632_),
    .Q_N(_08595_),
    .Q(\am_sdr0.cic2.comb1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net956),
    .D(_00633_),
    .Q_N(_08594_),
    .Q(\am_sdr0.cic2.comb1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net957),
    .D(_00634_),
    .Q_N(_08593_),
    .Q(\am_sdr0.cic2.comb1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net958),
    .D(_00635_),
    .Q_N(_08592_),
    .Q(\am_sdr0.cic2.comb1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net959),
    .D(_00636_),
    .Q_N(_08591_),
    .Q(\am_sdr0.cic2.comb1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net960),
    .D(_00637_),
    .Q_N(_08590_),
    .Q(\am_sdr0.cic2.comb1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net961),
    .D(_00638_),
    .Q_N(_08589_),
    .Q(\am_sdr0.cic2.comb1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net962),
    .D(_00639_),
    .Q_N(_08588_),
    .Q(\am_sdr0.cic2.comb1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net963),
    .D(_00640_),
    .Q_N(_08587_),
    .Q(\am_sdr0.cic2.comb1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net964),
    .D(_00641_),
    .Q_N(_08586_),
    .Q(\am_sdr0.cic2.comb1_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net965),
    .D(_00642_),
    .Q_N(_08585_),
    .Q(\am_sdr0.cic2.comb1_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net966),
    .D(_00643_),
    .Q_N(_08584_),
    .Q(\am_sdr0.cic2.comb1_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net967),
    .D(_00644_),
    .Q_N(_08583_),
    .Q(\am_sdr0.cic2.comb1_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net968),
    .D(_00645_),
    .Q_N(_08582_),
    .Q(\am_sdr0.cic2.comb1_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net969),
    .D(_00646_),
    .Q_N(_08581_),
    .Q(\am_sdr0.cic2.comb1_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net970),
    .D(_00647_),
    .Q_N(_08580_),
    .Q(\am_sdr0.cic2.comb1_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net971),
    .D(_00648_),
    .Q_N(_08579_),
    .Q(\am_sdr0.cic2.comb1_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net972),
    .D(_00649_),
    .Q_N(_08578_),
    .Q(\am_sdr0.cic2.comb1_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net973),
    .D(_00650_),
    .Q_N(_08577_),
    .Q(\am_sdr0.cic2.comb1_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net974),
    .D(_00651_),
    .Q_N(_08576_),
    .Q(\am_sdr0.cic2.comb1_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net975),
    .D(_00652_),
    .Q_N(_08575_),
    .Q(\am_sdr0.cic2.comb1_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net976),
    .D(_00653_),
    .Q_N(_08574_),
    .Q(\am_sdr0.cic2.comb1_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net977),
    .D(_00654_),
    .Q_N(_08573_),
    .Q(\am_sdr0.cic2.comb1_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net978),
    .D(_00655_),
    .Q_N(_08572_),
    .Q(\am_sdr0.cic2.comb1_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net979),
    .D(_00656_),
    .Q_N(_08571_),
    .Q(\am_sdr0.cic2.comb1_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net980),
    .D(_00657_),
    .Q_N(_08570_),
    .Q(\am_sdr0.cic2.comb1_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net981),
    .D(_00658_),
    .Q_N(_08569_),
    .Q(\am_sdr0.cic2.comb1_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net982),
    .D(_00659_),
    .Q_N(_08568_),
    .Q(\am_sdr0.cic2.comb1_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb1_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net983),
    .D(_00660_),
    .Q_N(_08567_),
    .Q(\am_sdr0.cic2.comb1_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net984),
    .D(_00661_),
    .Q_N(_08566_),
    .Q(\am_sdr0.cic2.comb2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net985),
    .D(_00662_),
    .Q_N(_08565_),
    .Q(\am_sdr0.cic2.comb2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net986),
    .D(_00663_),
    .Q_N(_08564_),
    .Q(\am_sdr0.cic2.comb2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net987),
    .D(_00664_),
    .Q_N(_08563_),
    .Q(\am_sdr0.cic2.comb2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net988),
    .D(_00665_),
    .Q_N(_08562_),
    .Q(\am_sdr0.cic2.comb2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net989),
    .D(_00666_),
    .Q_N(_08561_),
    .Q(\am_sdr0.cic2.comb2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net990),
    .D(_00667_),
    .Q_N(_08560_),
    .Q(\am_sdr0.cic2.comb2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net991),
    .D(_00668_),
    .Q_N(_08559_),
    .Q(\am_sdr0.cic2.comb2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net992),
    .D(_00669_),
    .Q_N(_08558_),
    .Q(\am_sdr0.cic2.comb2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net993),
    .D(_00670_),
    .Q_N(_08557_),
    .Q(\am_sdr0.cic2.comb2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net994),
    .D(_00671_),
    .Q_N(_08556_),
    .Q(\am_sdr0.cic2.comb2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net995),
    .D(_00672_),
    .Q_N(_08555_),
    .Q(\am_sdr0.cic2.comb2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net996),
    .D(_00673_),
    .Q_N(_08554_),
    .Q(\am_sdr0.cic2.comb2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net997),
    .D(_00674_),
    .Q_N(_08553_),
    .Q(\am_sdr0.cic2.comb2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net998),
    .D(_00675_),
    .Q_N(_08552_),
    .Q(\am_sdr0.cic2.comb2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net999),
    .D(_00676_),
    .Q_N(_08551_),
    .Q(\am_sdr0.cic2.comb2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1000),
    .D(_00677_),
    .Q_N(_08550_),
    .Q(\am_sdr0.cic2.comb2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1001),
    .D(_00678_),
    .Q_N(_08549_),
    .Q(\am_sdr0.cic2.comb2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1002),
    .D(_00679_),
    .Q_N(_08548_),
    .Q(\am_sdr0.cic2.comb2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1003),
    .D(_00680_),
    .Q_N(_08547_),
    .Q(\am_sdr0.cic2.comb2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1004),
    .D(_00681_),
    .Q_N(_08546_),
    .Q(\am_sdr0.cic2.comb2_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1005),
    .D(_00682_),
    .Q_N(_08545_),
    .Q(\am_sdr0.cic2.comb2_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1006),
    .D(_00683_),
    .Q_N(_08544_),
    .Q(\am_sdr0.cic2.comb2_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1007),
    .D(_00684_),
    .Q_N(_08543_),
    .Q(\am_sdr0.cic2.comb2_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1008),
    .D(_00685_),
    .Q_N(_08542_),
    .Q(\am_sdr0.cic2.comb2_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1009),
    .D(_00686_),
    .Q_N(_08541_),
    .Q(\am_sdr0.cic2.comb2_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1010),
    .D(_00687_),
    .Q_N(_08540_),
    .Q(\am_sdr0.cic2.comb2_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1011),
    .D(_00688_),
    .Q_N(_08539_),
    .Q(\am_sdr0.cic2.comb2_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1012),
    .D(_00689_),
    .Q_N(_08538_),
    .Q(\am_sdr0.cic2.comb2_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1013),
    .D(_00690_),
    .Q_N(_08537_),
    .Q(\am_sdr0.cic2.comb2_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1014),
    .D(_00691_),
    .Q_N(_08536_),
    .Q(\am_sdr0.cic2.comb2_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1015),
    .D(_00692_),
    .Q_N(_08535_),
    .Q(\am_sdr0.cic2.comb2_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1016),
    .D(_00693_),
    .Q_N(_08534_),
    .Q(\am_sdr0.cic2.comb2_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1017),
    .D(_00694_),
    .Q_N(_08533_),
    .Q(\am_sdr0.cic2.comb2_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1018),
    .D(_00695_),
    .Q_N(_08532_),
    .Q(\am_sdr0.cic2.comb2_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1019),
    .D(_00696_),
    .Q_N(_08531_),
    .Q(\am_sdr0.cic2.comb2_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1020),
    .D(_00697_),
    .Q_N(_08530_),
    .Q(\am_sdr0.cic2.comb2_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1021),
    .D(_00698_),
    .Q_N(_08529_),
    .Q(\am_sdr0.cic2.comb2_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1022),
    .D(_00699_),
    .Q_N(_08528_),
    .Q(\am_sdr0.cic2.comb2_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb2_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1023),
    .D(_00700_),
    .Q_N(_08527_),
    .Q(\am_sdr0.cic2.comb2_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1024),
    .D(_00701_),
    .Q_N(_08526_),
    .Q(\am_sdr0.cic2.comb3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1025),
    .D(_00702_),
    .Q_N(_08525_),
    .Q(\am_sdr0.cic2.comb3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1026),
    .D(_00703_),
    .Q_N(_08524_),
    .Q(\am_sdr0.cic2.comb3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1027),
    .D(_00704_),
    .Q_N(_08523_),
    .Q(\am_sdr0.cic2.comb3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1028),
    .D(_00705_),
    .Q_N(_08522_),
    .Q(\am_sdr0.cic2.comb3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1029),
    .D(_00706_),
    .Q_N(_08521_),
    .Q(\am_sdr0.cic2.comb3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1030),
    .D(_00707_),
    .Q_N(_08520_),
    .Q(\am_sdr0.cic2.comb3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1031),
    .D(_00708_),
    .Q_N(_08519_),
    .Q(\am_sdr0.cic2.comb3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1032),
    .D(_00709_),
    .Q_N(_08518_),
    .Q(\am_sdr0.cic2.comb3_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1033),
    .D(_00710_),
    .Q_N(_08517_),
    .Q(\am_sdr0.cic2.comb3_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1034),
    .D(_00711_),
    .Q_N(_08516_),
    .Q(\am_sdr0.cic2.comb3_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1035),
    .D(_00712_),
    .Q_N(_08515_),
    .Q(\am_sdr0.cic2.comb3_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1036),
    .D(_00713_),
    .Q_N(_08514_),
    .Q(\am_sdr0.cic2.comb3_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1037),
    .D(_00714_),
    .Q_N(_08513_),
    .Q(\am_sdr0.cic2.comb3_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1038),
    .D(_00715_),
    .Q_N(_08512_),
    .Q(\am_sdr0.cic2.comb3_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1039),
    .D(_00716_),
    .Q_N(_08511_),
    .Q(\am_sdr0.cic2.comb3_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1040),
    .D(_00717_),
    .Q_N(_08510_),
    .Q(\am_sdr0.cic2.comb3_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1041),
    .D(_00718_),
    .Q_N(_08509_),
    .Q(\am_sdr0.cic2.comb3_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1042),
    .D(_00719_),
    .Q_N(_08508_),
    .Q(\am_sdr0.cic2.comb3_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1043),
    .D(_00720_),
    .Q_N(_08507_),
    .Q(\am_sdr0.cic2.comb3_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1044),
    .D(_00721_),
    .Q_N(_08506_),
    .Q(\am_sdr0.cic2.comb3_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1045),
    .D(_00722_),
    .Q_N(_08505_),
    .Q(\am_sdr0.cic2.comb3_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1046),
    .D(_00723_),
    .Q_N(_08504_),
    .Q(\am_sdr0.cic2.comb3_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1047),
    .D(_00724_),
    .Q_N(_08503_),
    .Q(\am_sdr0.cic2.comb3_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1048),
    .D(_00725_),
    .Q_N(_08502_),
    .Q(\am_sdr0.cic2.comb3_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1049),
    .D(_00726_),
    .Q_N(_08501_),
    .Q(\am_sdr0.cic2.comb3_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1050),
    .D(_00727_),
    .Q_N(_08500_),
    .Q(\am_sdr0.cic2.comb3_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.comb3_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1051),
    .D(_00728_),
    .Q_N(_08499_),
    .Q(\am_sdr0.cic2.comb3_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1052),
    .D(_00729_),
    .Q_N(_08498_),
    .Q(\am_sdr0.cic2.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1053),
    .D(_00730_),
    .Q_N(_08497_),
    .Q(\am_sdr0.cic2.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1054),
    .D(_00731_),
    .Q_N(_08496_),
    .Q(\am_sdr0.cic2.count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1055),
    .D(_00732_),
    .Q_N(_08495_),
    .Q(\am_sdr0.cic2.count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1056),
    .D(_00733_),
    .Q_N(_08494_),
    .Q(\am_sdr0.cic2.count[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1057),
    .D(_00734_),
    .Q_N(_08493_),
    .Q(\am_sdr0.cic2.count[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1058),
    .D(_00735_),
    .Q_N(_08492_),
    .Q(\am_sdr0.cic2.count[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1059),
    .D(_00736_),
    .Q_N(_08491_),
    .Q(\am_sdr0.cic2.count[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1060),
    .D(_00737_),
    .Q_N(_08490_),
    .Q(\am_sdr0.cic2.integ1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1061),
    .D(_00738_),
    .Q_N(_08489_),
    .Q(\am_sdr0.cic2.integ1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1062),
    .D(_00739_),
    .Q_N(_08488_),
    .Q(\am_sdr0.cic2.integ1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1063),
    .D(_00740_),
    .Q_N(_08487_),
    .Q(\am_sdr0.cic2.integ1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1064),
    .D(_00741_),
    .Q_N(_08486_),
    .Q(\am_sdr0.cic2.integ1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1065),
    .D(_00742_),
    .Q_N(_08485_),
    .Q(\am_sdr0.cic2.integ1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1066),
    .D(_00743_),
    .Q_N(_08484_),
    .Q(\am_sdr0.cic2.integ1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1067),
    .D(_00744_),
    .Q_N(_08483_),
    .Q(\am_sdr0.cic2.integ1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1068),
    .D(_00745_),
    .Q_N(_08482_),
    .Q(\am_sdr0.cic2.integ1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1069),
    .D(_00746_),
    .Q_N(_08481_),
    .Q(\am_sdr0.cic2.integ1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1070),
    .D(_00747_),
    .Q_N(_08480_),
    .Q(\am_sdr0.cic2.integ1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1071),
    .D(_00748_),
    .Q_N(_08479_),
    .Q(\am_sdr0.cic2.integ1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1072),
    .D(_00749_),
    .Q_N(_08478_),
    .Q(\am_sdr0.cic2.integ1[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1073),
    .D(_00750_),
    .Q_N(_08477_),
    .Q(\am_sdr0.cic2.integ1[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1074),
    .D(_00751_),
    .Q_N(_08476_),
    .Q(\am_sdr0.cic2.integ1[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1075),
    .D(_00752_),
    .Q_N(_08475_),
    .Q(\am_sdr0.cic2.integ1[23] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1076),
    .D(_00753_),
    .Q_N(_08474_),
    .Q(\am_sdr0.cic2.integ1[24] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1077),
    .D(_00754_),
    .Q_N(_08473_),
    .Q(\am_sdr0.cic2.integ1[25] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1078),
    .D(_00755_),
    .Q_N(_08472_),
    .Q(\am_sdr0.cic2.integ1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1079),
    .D(_00756_),
    .Q_N(_08471_),
    .Q(\am_sdr0.cic2.integ1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1080),
    .D(_00757_),
    .Q_N(_08470_),
    .Q(\am_sdr0.cic2.integ1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1081),
    .D(_00758_),
    .Q_N(_08469_),
    .Q(\am_sdr0.cic2.integ1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1082),
    .D(_00759_),
    .Q_N(_08468_),
    .Q(\am_sdr0.cic2.integ1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1083),
    .D(_00760_),
    .Q_N(_08467_),
    .Q(\am_sdr0.cic2.integ1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1084),
    .D(_00761_),
    .Q_N(_08466_),
    .Q(\am_sdr0.cic2.integ1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1085),
    .D(_00762_),
    .Q_N(_08465_),
    .Q(\am_sdr0.cic2.integ1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1086),
    .D(_00763_),
    .Q_N(_08464_),
    .Q(\am_sdr0.cic2.integ2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1087),
    .D(_00764_),
    .Q_N(_08463_),
    .Q(\am_sdr0.cic2.integ2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1088),
    .D(_00765_),
    .Q_N(_08462_),
    .Q(\am_sdr0.cic2.integ2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1089),
    .D(_00766_),
    .Q_N(_08461_),
    .Q(\am_sdr0.cic2.integ2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1090),
    .D(_00767_),
    .Q_N(_08460_),
    .Q(\am_sdr0.cic2.integ2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1091),
    .D(_00768_),
    .Q_N(_08459_),
    .Q(\am_sdr0.cic2.integ2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1092),
    .D(_00769_),
    .Q_N(_08458_),
    .Q(\am_sdr0.cic2.integ2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1093),
    .D(_00770_),
    .Q_N(_08457_),
    .Q(\am_sdr0.cic2.integ2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1094),
    .D(_00771_),
    .Q_N(_08456_),
    .Q(\am_sdr0.cic2.integ2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1095),
    .D(_00772_),
    .Q_N(_08455_),
    .Q(\am_sdr0.cic2.integ2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1096),
    .D(_00773_),
    .Q_N(_08454_),
    .Q(\am_sdr0.cic2.integ2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1097),
    .D(_00774_),
    .Q_N(_08453_),
    .Q(\am_sdr0.cic2.integ2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1098),
    .D(_00775_),
    .Q_N(_08452_),
    .Q(\am_sdr0.cic2.integ2[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1099),
    .D(_00776_),
    .Q_N(_08451_),
    .Q(\am_sdr0.cic2.integ2[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1100),
    .D(_00777_),
    .Q_N(_08450_),
    .Q(\am_sdr0.cic2.integ2[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1101),
    .D(_00778_),
    .Q_N(_08449_),
    .Q(\am_sdr0.cic2.integ2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1102),
    .D(_00779_),
    .Q_N(_08448_),
    .Q(\am_sdr0.cic2.integ2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1103),
    .D(_00780_),
    .Q_N(_08447_),
    .Q(\am_sdr0.cic2.integ2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1104),
    .D(_00781_),
    .Q_N(_08446_),
    .Q(\am_sdr0.cic2.integ2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1105),
    .D(_00782_),
    .Q_N(_08445_),
    .Q(\am_sdr0.cic2.integ2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1106),
    .D(_00783_),
    .Q_N(_08444_),
    .Q(\am_sdr0.cic2.integ2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1107),
    .D(_00784_),
    .Q_N(_08443_),
    .Q(\am_sdr0.cic2.integ2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1108),
    .D(_00785_),
    .Q_N(_08442_),
    .Q(\am_sdr0.cic2.integ2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1109),
    .D(_00786_),
    .Q_N(_08441_),
    .Q(\am_sdr0.cic2.integ3[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1110),
    .D(_00787_),
    .Q_N(_08440_),
    .Q(\am_sdr0.cic2.integ3[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1111),
    .D(_00788_),
    .Q_N(_08439_),
    .Q(\am_sdr0.cic2.integ3[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1112),
    .D(_00789_),
    .Q_N(_08438_),
    .Q(\am_sdr0.cic2.integ3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1113),
    .D(_00790_),
    .Q_N(_08437_),
    .Q(\am_sdr0.cic2.integ3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1114),
    .D(_00791_),
    .Q_N(_08436_),
    .Q(\am_sdr0.cic2.integ3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1115),
    .D(_00792_),
    .Q_N(_08435_),
    .Q(\am_sdr0.cic2.integ3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1116),
    .D(_00793_),
    .Q_N(_08434_),
    .Q(\am_sdr0.cic2.integ3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1117),
    .D(_00794_),
    .Q_N(_08433_),
    .Q(\am_sdr0.cic2.integ3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1118),
    .D(_00795_),
    .Q_N(_08432_),
    .Q(\am_sdr0.cic2.integ3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1119),
    .D(_00796_),
    .Q_N(_08431_),
    .Q(\am_sdr0.cic2.integ3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1120),
    .D(_00797_),
    .Q_N(_08430_),
    .Q(\am_sdr0.cic2.integ3[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1121),
    .D(_00798_),
    .Q_N(_08429_),
    .Q(\am_sdr0.cic2.integ3[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1122),
    .D(_00799_),
    .Q_N(_08428_),
    .Q(\am_sdr0.cic2.integ3[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1123),
    .D(_00800_),
    .Q_N(_08427_),
    .Q(\am_sdr0.cic2.integ3[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1124),
    .D(_00801_),
    .Q_N(_08426_),
    .Q(\am_sdr0.cic2.integ3[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1125),
    .D(_00802_),
    .Q_N(_08425_),
    .Q(\am_sdr0.cic2.integ3[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1126),
    .D(_00803_),
    .Q_N(_08424_),
    .Q(\am_sdr0.cic2.integ3[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1127),
    .D(_00804_),
    .Q_N(_08423_),
    .Q(\am_sdr0.cic2.integ3[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ3[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1128),
    .D(_00805_),
    .Q_N(_08422_),
    .Q(\am_sdr0.cic2.integ3[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[0]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1129),
    .D(_00806_),
    .Q_N(_08421_),
    .Q(\am_sdr0.cic2.integ_sample[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[10]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1130),
    .D(_00807_),
    .Q_N(_08420_),
    .Q(\am_sdr0.cic2.integ_sample[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[11]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1131),
    .D(_00808_),
    .Q_N(_08419_),
    .Q(\am_sdr0.cic2.integ_sample[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[12]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1132),
    .D(_00809_),
    .Q_N(_08418_),
    .Q(\am_sdr0.cic2.integ_sample[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[13]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1133),
    .D(_00810_),
    .Q_N(_08417_),
    .Q(\am_sdr0.cic2.integ_sample[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[14]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1134),
    .D(_00811_),
    .Q_N(_08416_),
    .Q(\am_sdr0.cic2.integ_sample[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[15]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1135),
    .D(_00812_),
    .Q_N(_08415_),
    .Q(\am_sdr0.cic2.integ_sample[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[16]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1136),
    .D(_00813_),
    .Q_N(_08414_),
    .Q(\am_sdr0.cic2.integ_sample[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[17]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1137),
    .D(_00814_),
    .Q_N(_08413_),
    .Q(\am_sdr0.cic2.integ_sample[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[18]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1138),
    .D(_00815_),
    .Q_N(_08412_),
    .Q(\am_sdr0.cic2.integ_sample[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[19]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1139),
    .D(_00816_),
    .Q_N(_08411_),
    .Q(\am_sdr0.cic2.integ_sample[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[1]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1140),
    .D(_00817_),
    .Q_N(_08410_),
    .Q(\am_sdr0.cic2.integ_sample[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[2]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1141),
    .D(_00818_),
    .Q_N(_08409_),
    .Q(\am_sdr0.cic2.integ_sample[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1142),
    .D(_00819_),
    .Q_N(_08408_),
    .Q(\am_sdr0.cic2.integ_sample[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[4]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1143),
    .D(_00820_),
    .Q_N(_08407_),
    .Q(\am_sdr0.cic2.integ_sample[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[5]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1144),
    .D(_00821_),
    .Q_N(_08406_),
    .Q(\am_sdr0.cic2.integ_sample[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[6]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1145),
    .D(_00822_),
    .Q_N(_08405_),
    .Q(\am_sdr0.cic2.integ_sample[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1146),
    .D(_00823_),
    .Q_N(_08404_),
    .Q(\am_sdr0.cic2.integ_sample[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[8]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1147),
    .D(_00824_),
    .Q_N(_08403_),
    .Q(\am_sdr0.cic2.integ_sample[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.integ_sample[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1148),
    .D(_00825_),
    .Q_N(_08402_),
    .Q(\am_sdr0.cic2.integ_sample[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.out_tick$_SDFF_PN0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1149),
    .D(_00826_),
    .Q_N(_08401_),
    .Q(\am_sdr0.am0.load_tick ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.sample$_SDFF_PN0_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1150),
    .D(_00827_),
    .Q_N(_08400_),
    .Q(\am_sdr0.cic2.sample ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1151),
    .D(_00828_),
    .Q_N(_08399_),
    .Q(\am_sdr0.am0.I_in[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1152),
    .D(_00829_),
    .Q_N(_08398_),
    .Q(\am_sdr0.am0.I_in[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1153),
    .D(_00830_),
    .Q_N(_08397_),
    .Q(\am_sdr0.am0.I_in[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1154),
    .D(_00831_),
    .Q_N(_08396_),
    .Q(\am_sdr0.am0.I_in[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1155),
    .D(_00832_),
    .Q_N(_08395_),
    .Q(\am_sdr0.am0.I_in[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1156),
    .D(_00833_),
    .Q_N(_08394_),
    .Q(\am_sdr0.am0.I_in[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1157),
    .D(_00834_),
    .Q_N(_08393_),
    .Q(\am_sdr0.am0.I_in[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic2.x_out[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1158),
    .D(_00835_),
    .Q_N(_08392_),
    .Q(\am_sdr0.am0.I_in[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1159),
    .D(_00836_),
    .Q_N(_08391_),
    .Q(\am_sdr0.cic3.comb1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1160),
    .D(_00837_),
    .Q_N(_08390_),
    .Q(\am_sdr0.cic3.comb1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1161),
    .D(_00838_),
    .Q_N(_08389_),
    .Q(\am_sdr0.cic3.comb1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1162),
    .D(_00839_),
    .Q_N(_08388_),
    .Q(\am_sdr0.cic3.comb1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1163),
    .D(_00840_),
    .Q_N(_08387_),
    .Q(\am_sdr0.cic3.comb1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1164),
    .D(_00841_),
    .Q_N(_08386_),
    .Q(\am_sdr0.cic3.comb1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1165),
    .D(_00842_),
    .Q_N(_08385_),
    .Q(\am_sdr0.cic3.comb1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1166),
    .D(_00843_),
    .Q_N(_08384_),
    .Q(\am_sdr0.cic3.comb1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1167),
    .D(_00844_),
    .Q_N(_08383_),
    .Q(\am_sdr0.cic3.comb1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1168),
    .D(_00845_),
    .Q_N(_08382_),
    .Q(\am_sdr0.cic3.comb1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1169),
    .D(_00846_),
    .Q_N(_08381_),
    .Q(\am_sdr0.cic3.comb1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1170),
    .D(_00847_),
    .Q_N(_08380_),
    .Q(\am_sdr0.cic3.comb1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1171),
    .D(_00848_),
    .Q_N(_08379_),
    .Q(\am_sdr0.cic3.comb1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1172),
    .D(_00849_),
    .Q_N(_08378_),
    .Q(\am_sdr0.cic3.comb1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1173),
    .D(_00850_),
    .Q_N(_08377_),
    .Q(\am_sdr0.cic3.comb1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1174),
    .D(_00851_),
    .Q_N(_08376_),
    .Q(\am_sdr0.cic3.comb1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1175),
    .D(_00852_),
    .Q_N(_08375_),
    .Q(\am_sdr0.cic3.comb1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1176),
    .D(_00853_),
    .Q_N(_08374_),
    .Q(\am_sdr0.cic3.comb1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1177),
    .D(_00854_),
    .Q_N(_08373_),
    .Q(\am_sdr0.cic3.comb1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1178),
    .D(_00855_),
    .Q_N(_08372_),
    .Q(\am_sdr0.cic3.comb1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1179),
    .D(_00856_),
    .Q_N(_08371_),
    .Q(\am_sdr0.cic3.comb1_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1180),
    .D(_00857_),
    .Q_N(_08370_),
    .Q(\am_sdr0.cic3.comb1_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1181),
    .D(_00858_),
    .Q_N(_08369_),
    .Q(\am_sdr0.cic3.comb1_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1182),
    .D(_00859_),
    .Q_N(_08368_),
    .Q(\am_sdr0.cic3.comb1_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1183),
    .D(_00860_),
    .Q_N(_08367_),
    .Q(\am_sdr0.cic3.comb1_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1184),
    .D(_00861_),
    .Q_N(_08366_),
    .Q(\am_sdr0.cic3.comb1_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1185),
    .D(_00862_),
    .Q_N(_08365_),
    .Q(\am_sdr0.cic3.comb1_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1186),
    .D(_00863_),
    .Q_N(_08364_),
    .Q(\am_sdr0.cic3.comb1_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1187),
    .D(_00864_),
    .Q_N(_08363_),
    .Q(\am_sdr0.cic3.comb1_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1188),
    .D(_00865_),
    .Q_N(_08362_),
    .Q(\am_sdr0.cic3.comb1_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1189),
    .D(_00866_),
    .Q_N(_08361_),
    .Q(\am_sdr0.cic3.comb1_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1190),
    .D(_00867_),
    .Q_N(_08360_),
    .Q(\am_sdr0.cic3.comb1_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1191),
    .D(_00868_),
    .Q_N(_08359_),
    .Q(\am_sdr0.cic3.comb1_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1192),
    .D(_00869_),
    .Q_N(_08358_),
    .Q(\am_sdr0.cic3.comb1_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1193),
    .D(_00870_),
    .Q_N(_08357_),
    .Q(\am_sdr0.cic3.comb1_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1194),
    .D(_00871_),
    .Q_N(_08356_),
    .Q(\am_sdr0.cic3.comb1_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net1195),
    .D(_00872_),
    .Q_N(_08355_),
    .Q(\am_sdr0.cic3.comb1_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1196),
    .D(_00873_),
    .Q_N(_08354_),
    .Q(\am_sdr0.cic3.comb1_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1197),
    .D(_00874_),
    .Q_N(_08353_),
    .Q(\am_sdr0.cic3.comb1_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb1_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1198),
    .D(_00875_),
    .Q_N(_08352_),
    .Q(\am_sdr0.cic3.comb1_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1199),
    .D(_00876_),
    .Q_N(_08351_),
    .Q(\am_sdr0.cic3.comb2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1200),
    .D(_00877_),
    .Q_N(_08350_),
    .Q(\am_sdr0.cic3.comb2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1201),
    .D(_00878_),
    .Q_N(_08349_),
    .Q(\am_sdr0.cic3.comb2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1202),
    .D(_00879_),
    .Q_N(_08348_),
    .Q(\am_sdr0.cic3.comb2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1203),
    .D(_00880_),
    .Q_N(_08347_),
    .Q(\am_sdr0.cic3.comb2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1204),
    .D(_00881_),
    .Q_N(_08346_),
    .Q(\am_sdr0.cic3.comb2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1205),
    .D(_00882_),
    .Q_N(_08345_),
    .Q(\am_sdr0.cic3.comb2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1206),
    .D(_00883_),
    .Q_N(_08344_),
    .Q(\am_sdr0.cic3.comb2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1207),
    .D(_00884_),
    .Q_N(_08343_),
    .Q(\am_sdr0.cic3.comb2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1208),
    .D(_00885_),
    .Q_N(_08342_),
    .Q(\am_sdr0.cic3.comb2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1209),
    .D(_00886_),
    .Q_N(_08341_),
    .Q(\am_sdr0.cic3.comb2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1210),
    .D(_00887_),
    .Q_N(_08340_),
    .Q(\am_sdr0.cic3.comb2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1211),
    .D(_00888_),
    .Q_N(_08339_),
    .Q(\am_sdr0.cic3.comb2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1212),
    .D(_00889_),
    .Q_N(_08338_),
    .Q(\am_sdr0.cic3.comb2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1213),
    .D(_00890_),
    .Q_N(_08337_),
    .Q(\am_sdr0.cic3.comb2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1214),
    .D(_00891_),
    .Q_N(_08336_),
    .Q(\am_sdr0.cic3.comb2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1215),
    .D(_00892_),
    .Q_N(_08335_),
    .Q(\am_sdr0.cic3.comb2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1216),
    .D(_00893_),
    .Q_N(_08334_),
    .Q(\am_sdr0.cic3.comb2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1217),
    .D(_00894_),
    .Q_N(_08333_),
    .Q(\am_sdr0.cic3.comb2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1218),
    .D(_00895_),
    .Q_N(_08332_),
    .Q(\am_sdr0.cic3.comb2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1219),
    .D(_00896_),
    .Q_N(_08331_),
    .Q(\am_sdr0.cic3.comb2_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1220),
    .D(_00897_),
    .Q_N(_08330_),
    .Q(\am_sdr0.cic3.comb2_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1221),
    .D(_00898_),
    .Q_N(_08329_),
    .Q(\am_sdr0.cic3.comb2_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1222),
    .D(_00899_),
    .Q_N(_08328_),
    .Q(\am_sdr0.cic3.comb2_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1223),
    .D(_00900_),
    .Q_N(_08327_),
    .Q(\am_sdr0.cic3.comb2_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1224),
    .D(_00901_),
    .Q_N(_08326_),
    .Q(\am_sdr0.cic3.comb2_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1225),
    .D(_00902_),
    .Q_N(_08325_),
    .Q(\am_sdr0.cic3.comb2_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1226),
    .D(_00903_),
    .Q_N(_08324_),
    .Q(\am_sdr0.cic3.comb2_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1227),
    .D(_00904_),
    .Q_N(_08323_),
    .Q(\am_sdr0.cic3.comb2_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1228),
    .D(_00905_),
    .Q_N(_08322_),
    .Q(\am_sdr0.cic3.comb2_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1229),
    .D(_00906_),
    .Q_N(_08321_),
    .Q(\am_sdr0.cic3.comb2_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1230),
    .D(_00907_),
    .Q_N(_08320_),
    .Q(\am_sdr0.cic3.comb2_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1231),
    .D(_00908_),
    .Q_N(_08319_),
    .Q(\am_sdr0.cic3.comb2_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1232),
    .D(_00909_),
    .Q_N(_08318_),
    .Q(\am_sdr0.cic3.comb2_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1233),
    .D(_00910_),
    .Q_N(_08317_),
    .Q(\am_sdr0.cic3.comb2_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1234),
    .D(_00911_),
    .Q_N(_08316_),
    .Q(\am_sdr0.cic3.comb2_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1235),
    .D(_00912_),
    .Q_N(_08315_),
    .Q(\am_sdr0.cic3.comb2_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1236),
    .D(_00913_),
    .Q_N(_08314_),
    .Q(\am_sdr0.cic3.comb2_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1237),
    .D(_00914_),
    .Q_N(_08313_),
    .Q(\am_sdr0.cic3.comb2_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb2_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1238),
    .D(_00915_),
    .Q_N(_08312_),
    .Q(\am_sdr0.cic3.comb2_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1239),
    .D(_00916_),
    .Q_N(_08311_),
    .Q(\am_sdr0.cic3.comb3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1240),
    .D(_00917_),
    .Q_N(_08310_),
    .Q(\am_sdr0.cic3.comb3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1241),
    .D(_00918_),
    .Q_N(_08309_),
    .Q(\am_sdr0.cic3.comb3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1242),
    .D(_00919_),
    .Q_N(_08308_),
    .Q(\am_sdr0.cic3.comb3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1243),
    .D(_00920_),
    .Q_N(_08307_),
    .Q(\am_sdr0.cic3.comb3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1244),
    .D(_00921_),
    .Q_N(_08306_),
    .Q(\am_sdr0.cic3.comb3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1245),
    .D(_00922_),
    .Q_N(_08305_),
    .Q(\am_sdr0.cic3.comb3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1246),
    .D(_00923_),
    .Q_N(_08304_),
    .Q(\am_sdr0.cic3.comb3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1247),
    .D(_00924_),
    .Q_N(_08303_),
    .Q(\am_sdr0.cic3.comb3_in_del[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1248),
    .D(_00925_),
    .Q_N(_08302_),
    .Q(\am_sdr0.cic3.comb3_in_del[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1249),
    .D(_00926_),
    .Q_N(_08301_),
    .Q(\am_sdr0.cic3.comb3_in_del[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1250),
    .D(_00927_),
    .Q_N(_08300_),
    .Q(\am_sdr0.cic3.comb3_in_del[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1251),
    .D(_00928_),
    .Q_N(_08299_),
    .Q(\am_sdr0.cic3.comb3_in_del[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1252),
    .D(_00929_),
    .Q_N(_08298_),
    .Q(\am_sdr0.cic3.comb3_in_del[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1253),
    .D(_00930_),
    .Q_N(_08297_),
    .Q(\am_sdr0.cic3.comb3_in_del[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1254),
    .D(_00931_),
    .Q_N(_08296_),
    .Q(\am_sdr0.cic3.comb3_in_del[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1255),
    .D(_00932_),
    .Q_N(_08295_),
    .Q(\am_sdr0.cic3.comb3_in_del[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1256),
    .D(_00933_),
    .Q_N(_08294_),
    .Q(\am_sdr0.cic3.comb3_in_del[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1257),
    .D(_00934_),
    .Q_N(_08293_),
    .Q(\am_sdr0.cic3.comb3_in_del[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1258),
    .D(_00935_),
    .Q_N(_08292_),
    .Q(\am_sdr0.cic3.comb3_in_del[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1259),
    .D(_00936_),
    .Q_N(_08291_),
    .Q(\am_sdr0.cic3.comb3_in_del[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1260),
    .D(_00937_),
    .Q_N(_08290_),
    .Q(\am_sdr0.cic3.comb3_in_del[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1261),
    .D(_00938_),
    .Q_N(_08289_),
    .Q(\am_sdr0.cic3.comb3_in_del[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1262),
    .D(_00939_),
    .Q_N(_08288_),
    .Q(\am_sdr0.cic3.comb3_in_del[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1263),
    .D(_00940_),
    .Q_N(_08287_),
    .Q(\am_sdr0.cic3.comb3_in_del[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1264),
    .D(_00941_),
    .Q_N(_08286_),
    .Q(\am_sdr0.cic3.comb3_in_del[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1265),
    .D(_00942_),
    .Q_N(_08285_),
    .Q(\am_sdr0.cic3.comb3_in_del[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.comb3_in_del[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1266),
    .D(_00943_),
    .Q_N(_08284_),
    .Q(\am_sdr0.cic3.comb3_in_del[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1267),
    .D(_00944_),
    .Q_N(_08283_),
    .Q(\am_sdr0.cic3.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1268),
    .D(_00945_),
    .Q_N(_08282_),
    .Q(\am_sdr0.cic3.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1269),
    .D(_00946_),
    .Q_N(_08281_),
    .Q(\am_sdr0.cic3.count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1270),
    .D(_00947_),
    .Q_N(_08280_),
    .Q(\am_sdr0.cic3.count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1271),
    .D(_00948_),
    .Q_N(_08279_),
    .Q(\am_sdr0.cic3.count[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1272),
    .D(_00949_),
    .Q_N(_08278_),
    .Q(\am_sdr0.cic3.count[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1273),
    .D(_00950_),
    .Q_N(_08277_),
    .Q(\am_sdr0.cic3.count[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.count[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1274),
    .D(_00951_),
    .Q_N(_08276_),
    .Q(\am_sdr0.cic3.count[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1275),
    .D(_00952_),
    .Q_N(_08275_),
    .Q(\am_sdr0.cic3.integ1[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1276),
    .D(_00953_),
    .Q_N(_08274_),
    .Q(\am_sdr0.cic3.integ1[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1277),
    .D(_00954_),
    .Q_N(_08273_),
    .Q(\am_sdr0.cic3.integ1[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1278),
    .D(_00955_),
    .Q_N(_08272_),
    .Q(\am_sdr0.cic3.integ1[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1279),
    .D(_00956_),
    .Q_N(_08271_),
    .Q(\am_sdr0.cic3.integ1[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1280),
    .D(_00957_),
    .Q_N(_08270_),
    .Q(\am_sdr0.cic3.integ1[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1281),
    .D(_00958_),
    .Q_N(_08269_),
    .Q(\am_sdr0.cic3.integ1[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1282),
    .D(_00959_),
    .Q_N(_08268_),
    .Q(\am_sdr0.cic3.integ1[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1283),
    .D(_00960_),
    .Q_N(_08267_),
    .Q(\am_sdr0.cic3.integ1[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1284),
    .D(_00961_),
    .Q_N(_08266_),
    .Q(\am_sdr0.cic3.integ1[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1285),
    .D(_00962_),
    .Q_N(_08265_),
    .Q(\am_sdr0.cic3.integ1[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1286),
    .D(_00963_),
    .Q_N(_08264_),
    .Q(\am_sdr0.cic3.integ1[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1287),
    .D(_00964_),
    .Q_N(_08263_),
    .Q(\am_sdr0.cic3.integ1[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1288),
    .D(_00965_),
    .Q_N(_08262_),
    .Q(\am_sdr0.cic3.integ1[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1289),
    .D(_00966_),
    .Q_N(_08261_),
    .Q(\am_sdr0.cic3.integ1[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1290),
    .D(_00967_),
    .Q_N(_08260_),
    .Q(\am_sdr0.cic3.integ1[23] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1291),
    .D(_00968_),
    .Q_N(_08259_),
    .Q(\am_sdr0.cic3.integ1[24] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1292),
    .D(_00969_),
    .Q_N(_08258_),
    .Q(\am_sdr0.cic3.integ1[25] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1293),
    .D(_00970_),
    .Q_N(_08257_),
    .Q(\am_sdr0.cic3.integ1[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1294),
    .D(_00971_),
    .Q_N(_08256_),
    .Q(\am_sdr0.cic3.integ1[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1295),
    .D(_00972_),
    .Q_N(_08255_),
    .Q(\am_sdr0.cic3.integ1[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1296),
    .D(_00973_),
    .Q_N(_08254_),
    .Q(\am_sdr0.cic3.integ1[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1297),
    .D(_00974_),
    .Q_N(_08253_),
    .Q(\am_sdr0.cic3.integ1[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1298),
    .D(_00975_),
    .Q_N(_08252_),
    .Q(\am_sdr0.cic3.integ1[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1299),
    .D(_00976_),
    .Q_N(_08251_),
    .Q(\am_sdr0.cic3.integ1[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1300),
    .D(_00977_),
    .Q_N(_08250_),
    .Q(\am_sdr0.cic3.integ1[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1301),
    .D(_00978_),
    .Q_N(_08249_),
    .Q(\am_sdr0.cic3.integ2[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1302),
    .D(_00979_),
    .Q_N(_08248_),
    .Q(\am_sdr0.cic3.integ2[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1303),
    .D(_00980_),
    .Q_N(_08247_),
    .Q(\am_sdr0.cic3.integ2[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1304),
    .D(_00981_),
    .Q_N(_08246_),
    .Q(\am_sdr0.cic3.integ2[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1305),
    .D(_00982_),
    .Q_N(_08245_),
    .Q(\am_sdr0.cic3.integ2[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1306),
    .D(_00983_),
    .Q_N(_08244_),
    .Q(\am_sdr0.cic3.integ2[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1307),
    .D(_00984_),
    .Q_N(_08243_),
    .Q(\am_sdr0.cic3.integ2[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1308),
    .D(_00985_),
    .Q_N(_08242_),
    .Q(\am_sdr0.cic3.integ2[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1309),
    .D(_00986_),
    .Q_N(_08241_),
    .Q(\am_sdr0.cic3.integ2[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1310),
    .D(_00987_),
    .Q_N(_08240_),
    .Q(\am_sdr0.cic3.integ2[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1311),
    .D(_00988_),
    .Q_N(_08239_),
    .Q(\am_sdr0.cic3.integ2[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1312),
    .D(_00989_),
    .Q_N(_08238_),
    .Q(\am_sdr0.cic3.integ2[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1313),
    .D(_00990_),
    .Q_N(_08237_),
    .Q(\am_sdr0.cic3.integ2[20] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1314),
    .D(_00991_),
    .Q_N(_08236_),
    .Q(\am_sdr0.cic3.integ2[21] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1315),
    .D(_00992_),
    .Q_N(_08235_),
    .Q(\am_sdr0.cic3.integ2[22] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1316),
    .D(_00993_),
    .Q_N(_08234_),
    .Q(\am_sdr0.cic3.integ2[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1317),
    .D(_00994_),
    .Q_N(_08233_),
    .Q(\am_sdr0.cic3.integ2[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1318),
    .D(_00995_),
    .Q_N(_08232_),
    .Q(\am_sdr0.cic3.integ2[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1319),
    .D(_00996_),
    .Q_N(_08231_),
    .Q(\am_sdr0.cic3.integ2[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1320),
    .D(_00997_),
    .Q_N(_08230_),
    .Q(\am_sdr0.cic3.integ2[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1321),
    .D(_00998_),
    .Q_N(_08229_),
    .Q(\am_sdr0.cic3.integ2[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1322),
    .D(_00999_),
    .Q_N(_08228_),
    .Q(\am_sdr0.cic3.integ2[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1323),
    .D(_01000_),
    .Q_N(_08227_),
    .Q(\am_sdr0.cic3.integ2[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1324),
    .D(_01001_),
    .Q_N(_08226_),
    .Q(\am_sdr0.cic3.integ3[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1325),
    .D(_01002_),
    .Q_N(_08225_),
    .Q(\am_sdr0.cic3.integ3[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1326),
    .D(_01003_),
    .Q_N(_08224_),
    .Q(\am_sdr0.cic3.integ3[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1327),
    .D(_01004_),
    .Q_N(_08223_),
    .Q(\am_sdr0.cic3.integ3[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1328),
    .D(_01005_),
    .Q_N(_08222_),
    .Q(\am_sdr0.cic3.integ3[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1329),
    .D(_01006_),
    .Q_N(_08221_),
    .Q(\am_sdr0.cic3.integ3[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1330),
    .D(_01007_),
    .Q_N(_08220_),
    .Q(\am_sdr0.cic3.integ3[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1331),
    .D(_01008_),
    .Q_N(_08219_),
    .Q(\am_sdr0.cic3.integ3[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1332),
    .D(_01009_),
    .Q_N(_08218_),
    .Q(\am_sdr0.cic3.integ3[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1333),
    .D(_01010_),
    .Q_N(_08217_),
    .Q(\am_sdr0.cic3.integ3[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1334),
    .D(_01011_),
    .Q_N(_08216_),
    .Q(\am_sdr0.cic3.integ3[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1335),
    .D(_01012_),
    .Q_N(_08215_),
    .Q(\am_sdr0.cic3.integ3[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1336),
    .D(_01013_),
    .Q_N(_08214_),
    .Q(\am_sdr0.cic3.integ3[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1337),
    .D(_01014_),
    .Q_N(_08213_),
    .Q(\am_sdr0.cic3.integ3[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1338),
    .D(_01015_),
    .Q_N(_08212_),
    .Q(\am_sdr0.cic3.integ3[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1339),
    .D(_01016_),
    .Q_N(_08211_),
    .Q(\am_sdr0.cic3.integ3[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1340),
    .D(_01017_),
    .Q_N(_08210_),
    .Q(\am_sdr0.cic3.integ3[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1341),
    .D(_01018_),
    .Q_N(_08209_),
    .Q(\am_sdr0.cic3.integ3[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1342),
    .D(_01019_),
    .Q_N(_08208_),
    .Q(\am_sdr0.cic3.integ3[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ3[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1343),
    .D(_01020_),
    .Q_N(_08207_),
    .Q(\am_sdr0.cic3.integ3[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[0]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1344),
    .D(_01021_),
    .Q_N(_08206_),
    .Q(\am_sdr0.cic3.integ_sample[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[10]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1345),
    .D(_01022_),
    .Q_N(_08205_),
    .Q(\am_sdr0.cic3.integ_sample[10] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1346),
    .D(_01023_),
    .Q_N(_08204_),
    .Q(\am_sdr0.cic3.integ_sample[11] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[12]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1347),
    .D(_01024_),
    .Q_N(_08203_),
    .Q(\am_sdr0.cic3.integ_sample[12] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[13]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1348),
    .D(_01025_),
    .Q_N(_08202_),
    .Q(\am_sdr0.cic3.integ_sample[13] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[14]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1349),
    .D(_01026_),
    .Q_N(_08201_),
    .Q(\am_sdr0.cic3.integ_sample[14] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[15]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1350),
    .D(_01027_),
    .Q_N(_08200_),
    .Q(\am_sdr0.cic3.integ_sample[15] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[16]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1351),
    .D(_01028_),
    .Q_N(_08199_),
    .Q(\am_sdr0.cic3.integ_sample[16] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[17]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1352),
    .D(_01029_),
    .Q_N(_08198_),
    .Q(\am_sdr0.cic3.integ_sample[17] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[18]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1353),
    .D(_01030_),
    .Q_N(_08197_),
    .Q(\am_sdr0.cic3.integ_sample[18] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[19]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1354),
    .D(_01031_),
    .Q_N(_08196_),
    .Q(\am_sdr0.cic3.integ_sample[19] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[1]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1355),
    .D(_01032_),
    .Q_N(_08195_),
    .Q(\am_sdr0.cic3.integ_sample[1] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[2]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1356),
    .D(_01033_),
    .Q_N(_08194_),
    .Q(\am_sdr0.cic3.integ_sample[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1357),
    .D(_01034_),
    .Q_N(_08193_),
    .Q(\am_sdr0.cic3.integ_sample[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[4]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1358),
    .D(_01035_),
    .Q_N(_08192_),
    .Q(\am_sdr0.cic3.integ_sample[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[5]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1359),
    .D(_01036_),
    .Q_N(_08191_),
    .Q(\am_sdr0.cic3.integ_sample[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[6]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1360),
    .D(_01037_),
    .Q_N(_08190_),
    .Q(\am_sdr0.cic3.integ_sample[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[7]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1361),
    .D(_01038_),
    .Q_N(_08189_),
    .Q(\am_sdr0.cic3.integ_sample[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[8]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1362),
    .D(_01039_),
    .Q_N(_08188_),
    .Q(\am_sdr0.cic3.integ_sample[8] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.integ_sample[9]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1363),
    .D(_01040_),
    .Q_N(_08187_),
    .Q(\am_sdr0.cic3.integ_sample[9] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.sample$_SDFF_PN0_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1364),
    .D(net11),
    .Q_N(_08186_),
    .Q(\am_sdr0.cic3.sample ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1365),
    .D(_01042_),
    .Q_N(_08185_),
    .Q(\am_sdr0.am0.Q_in[2] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1366),
    .D(_01043_),
    .Q_N(_08184_),
    .Q(\am_sdr0.am0.Q_in[3] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1367),
    .D(_01044_),
    .Q_N(_08183_),
    .Q(\am_sdr0.am0.Q_in[4] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1368),
    .D(_01045_),
    .Q_N(_08182_),
    .Q(\am_sdr0.am0.Q_in[5] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1369),
    .D(_01046_),
    .Q_N(_08181_),
    .Q(\am_sdr0.am0.Q_in[6] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1370),
    .D(_01047_),
    .Q_N(_08180_),
    .Q(\am_sdr0.am0.Q_in[7] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1371),
    .D(_01048_),
    .Q_N(_08179_),
    .Q(\am_sdr0.am0.Q_in[0] ));
 sg13g2_dfrbp_1 \am_sdr0.cic3.x_out[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1372),
    .D(_01049_),
    .Q_N(_08178_),
    .Q(\am_sdr0.am0.Q_in[1] ));
 sg13g2_dfrbp_1 \am_sdr0.count[0]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1373),
    .D(_01050_),
    .Q_N(_00068_),
    .Q(\am_sdr0.count[0] ));
 sg13g2_dfrbp_1 \am_sdr0.count[1]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1374),
    .D(_01051_),
    .Q_N(_08177_),
    .Q(\am_sdr0.count[1] ));
 sg13g2_dfrbp_1 \am_sdr0.count[2]$_SDFF_PN0_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1375),
    .D(_01052_),
    .Q_N(_08176_),
    .Q(\am_sdr0.count[2] ));
 sg13g2_dfrbp_1 \am_sdr0.count[3]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1376),
    .D(_01053_),
    .Q_N(_08175_),
    .Q(\am_sdr0.count[3] ));
 sg13g2_dfrbp_1 \am_sdr0.count[4]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1377),
    .D(_01054_),
    .Q_N(_08174_),
    .Q(\am_sdr0.count[4] ));
 sg13g2_dfrbp_1 \am_sdr0.count[5]$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1378),
    .D(_01055_),
    .Q_N(_08173_),
    .Q(\am_sdr0.count[5] ));
 sg13g2_dfrbp_1 \am_sdr0.count[6]$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1379),
    .D(_01056_),
    .Q_N(_08172_),
    .Q(\am_sdr0.count[6] ));
 sg13g2_dfrbp_1 \am_sdr0.count[7]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1380),
    .D(_01057_),
    .Q_N(_09128_),
    .Q(\am_sdr0.count[7] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[0]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1381),
    .D(\am_sdr0.mix0.cos_q[0] ),
    .Q_N(_09129_),
    .Q(\am_sdr0.I_out[0] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[1]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1382),
    .D(_00023_),
    .Q_N(_09130_),
    .Q(\am_sdr0.I_out[1] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[2]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1383),
    .D(_00024_),
    .Q_N(_09131_),
    .Q(\am_sdr0.I_out[2] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1384),
    .D(_00025_),
    .Q_N(_09132_),
    .Q(\am_sdr0.I_out[3] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[4]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1385),
    .D(_00026_),
    .Q_N(_09133_),
    .Q(\am_sdr0.I_out[4] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[5]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1386),
    .D(_00027_),
    .Q_N(_09134_),
    .Q(\am_sdr0.I_out[5] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[6]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1387),
    .D(_00028_),
    .Q_N(_09135_),
    .Q(\am_sdr0.I_out[6] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.I_out[7]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1388),
    .D(_00029_),
    .Q_N(_09136_),
    .Q(\am_sdr0.I_out[7] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[0]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1389),
    .D(\am_sdr0.mix0.sin_q[0] ),
    .Q_N(_09137_),
    .Q(\am_sdr0.Q_out[0] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[1]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1390),
    .D(_00030_),
    .Q_N(_09138_),
    .Q(\am_sdr0.Q_out[1] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1391),
    .D(_00031_),
    .Q_N(_09139_),
    .Q(\am_sdr0.Q_out[2] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[3]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1392),
    .D(_00032_),
    .Q_N(_09140_),
    .Q(\am_sdr0.Q_out[3] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[4]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1393),
    .D(_00033_),
    .Q_N(_09141_),
    .Q(\am_sdr0.Q_out[4] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[5]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1394),
    .D(_00034_),
    .Q_N(_09142_),
    .Q(\am_sdr0.Q_out[5] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[6]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1395),
    .D(_00035_),
    .Q_N(_09143_),
    .Q(\am_sdr0.Q_out[6] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.Q_out[7]$_DFF_P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1396),
    .D(_00036_),
    .Q_N(_08171_),
    .Q(\am_sdr0.Q_out[7] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.RF_in_q$_SDFF_PN0_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1397),
    .D(_01058_),
    .Q_N(_08170_),
    .Q(\am_sdr0.mix0.RF_in_q ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.RF_in_qq$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1398),
    .D(_01059_),
    .Q_N(_08169_),
    .Q(\am_sdr0.mix0.RF_in_qq ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.RF_out$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1399),
    .D(_01060_),
    .Q_N(_08168_),
    .Q(COMP_OUT));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[0]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1400),
    .D(_01061_),
    .Q_N(_08167_),
    .Q(\am_sdr0.mix0.cos_q[0] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[1]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1401),
    .D(_01062_),
    .Q_N(_08166_),
    .Q(\am_sdr0.mix0.cos_q[1] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[2]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1402),
    .D(_01063_),
    .Q_N(_08165_),
    .Q(\am_sdr0.mix0.cos_q[2] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[3]$_SDFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1403),
    .D(_01064_),
    .Q_N(_08164_),
    .Q(\am_sdr0.mix0.cos_q[3] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[4]$_SDFF_PN0_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1404),
    .D(_01065_),
    .Q_N(_08163_),
    .Q(\am_sdr0.mix0.cos_q[4] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[5]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1405),
    .D(_01066_),
    .Q_N(_08162_),
    .Q(\am_sdr0.mix0.cos_q[5] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[6]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1406),
    .D(_01067_),
    .Q_N(_08161_),
    .Q(\am_sdr0.mix0.cos_q[6] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.cos_q[7]$_SDFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1407),
    .D(_01068_),
    .Q_N(_08160_),
    .Q(\am_sdr0.mix0.cos_q[7] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[0]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1408),
    .D(_01069_),
    .Q_N(_08159_),
    .Q(\am_sdr0.mix0.sin_q[0] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[1]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1409),
    .D(_01070_),
    .Q_N(_08158_),
    .Q(\am_sdr0.mix0.sin_q[1] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[2]$_SDFF_PN0_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1410),
    .D(_01071_),
    .Q_N(_08157_),
    .Q(\am_sdr0.mix0.sin_q[2] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[3]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1411),
    .D(_01072_),
    .Q_N(_08156_),
    .Q(\am_sdr0.mix0.sin_q[3] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[4]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1412),
    .D(_01073_),
    .Q_N(_08155_),
    .Q(\am_sdr0.mix0.sin_q[4] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[5]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1413),
    .D(_01074_),
    .Q_N(_08154_),
    .Q(\am_sdr0.mix0.sin_q[5] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[6]$_SDFF_PN0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1414),
    .D(_01075_),
    .Q_N(_08153_),
    .Q(\am_sdr0.mix0.sin_q[6] ));
 sg13g2_dfrbp_1 \am_sdr0.mix0.sin_q[7]$_SDFF_PN0_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1415),
    .D(_01076_),
    .Q_N(_09144_),
    .Q(\am_sdr0.mix0.sin_q[7] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[0]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1416),
    .D(_00000_),
    .Q_N(_09145_),
    .Q(\am_sdr0.cos[0] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[1]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1417),
    .D(_00001_),
    .Q_N(_09146_),
    .Q(\am_sdr0.cos[1] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[2]$_DFF_P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1418),
    .D(_00002_),
    .Q_N(_09147_),
    .Q(\am_sdr0.cos[2] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1419),
    .D(_00003_),
    .Q_N(_09148_),
    .Q(\am_sdr0.cos[3] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[4]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1420),
    .D(_00004_),
    .Q_N(_09149_),
    .Q(\am_sdr0.cos[4] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[5]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1421),
    .D(_00005_),
    .Q_N(_09150_),
    .Q(\am_sdr0.cos[5] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[6]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1422),
    .D(_00006_),
    .Q_N(_09151_),
    .Q(\am_sdr0.cos[6] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.cos0.data[7]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1423),
    .D(_00007_),
    .Q_N(_08152_),
    .Q(\am_sdr0.cos[7] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[0]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1424),
    .D(_01077_),
    .Q_N(_08151_),
    .Q(\am_sdr0.nco0.phase[0] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[10]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1425),
    .D(_01078_),
    .Q_N(_08150_),
    .Q(\am_sdr0.nco0.phase[10] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[11]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1426),
    .D(_01079_),
    .Q_N(_08149_),
    .Q(\am_sdr0.nco0.phase[11] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[12]$_SDFF_PN0_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1427),
    .D(_01080_),
    .Q_N(_08148_),
    .Q(\am_sdr0.nco0.phase[12] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[13]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1428),
    .D(_01081_),
    .Q_N(_08147_),
    .Q(\am_sdr0.nco0.phase[13] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[14]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1429),
    .D(_01082_),
    .Q_N(_08146_),
    .Q(\am_sdr0.nco0.phase[14] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[15]$_SDFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1430),
    .D(_01083_),
    .Q_N(_08145_),
    .Q(\am_sdr0.nco0.phase[15] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[16]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1431),
    .D(_01084_),
    .Q_N(_08144_),
    .Q(\am_sdr0.nco0.phase[16] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[17]$_SDFF_PN0_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1432),
    .D(_01085_),
    .Q_N(_08143_),
    .Q(\am_sdr0.nco0.phase[17] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[18]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1433),
    .D(_01086_),
    .Q_N(_08142_),
    .Q(\am_sdr0.nco0.phase[18] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[19]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1434),
    .D(_01087_),
    .Q_N(_08141_),
    .Q(\am_sdr0.nco0.phase[19] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[1]$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1435),
    .D(_01088_),
    .Q_N(_08140_),
    .Q(\am_sdr0.nco0.phase[1] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[20]$_SDFF_PN0_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1436),
    .D(_01089_),
    .Q_N(_08139_),
    .Q(\am_sdr0.nco0.phase[20] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[21]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1437),
    .D(_01090_),
    .Q_N(_08138_),
    .Q(\am_sdr0.nco0.phase[21] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[22]$_SDFF_PN0_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1438),
    .D(_01091_),
    .Q_N(_08137_),
    .Q(\am_sdr0.nco0.phase[22] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[23]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1439),
    .D(_01092_),
    .Q_N(_00038_),
    .Q(\am_sdr0.nco0.phase[23] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[24]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1440),
    .D(_01093_),
    .Q_N(_00039_),
    .Q(\am_sdr0.nco0.phase[24] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[25]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1441),
    .D(_01094_),
    .Q_N(_00037_),
    .Q(\am_sdr0.nco0.phase[25] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[2]$_SDFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1442),
    .D(_01095_),
    .Q_N(_08136_),
    .Q(\am_sdr0.nco0.phase[2] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[3]$_SDFF_PN0_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1443),
    .D(_01096_),
    .Q_N(_08135_),
    .Q(\am_sdr0.nco0.phase[3] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[4]$_SDFF_PN0_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1444),
    .D(_01097_),
    .Q_N(_08134_),
    .Q(\am_sdr0.nco0.phase[4] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[5]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1445),
    .D(_01098_),
    .Q_N(_08133_),
    .Q(\am_sdr0.nco0.phase[5] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[6]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1446),
    .D(_01099_),
    .Q_N(_08132_),
    .Q(\am_sdr0.nco0.phase[6] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[7]$_SDFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1447),
    .D(_01100_),
    .Q_N(_08131_),
    .Q(\am_sdr0.nco0.phase[7] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[8]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1448),
    .D(_01101_),
    .Q_N(_08130_),
    .Q(\am_sdr0.nco0.phase[8] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.phase[9]$_SDFF_PN0_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1449),
    .D(_01102_),
    .Q_N(_09152_),
    .Q(\am_sdr0.nco0.phase[9] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[0]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1450),
    .D(_00008_),
    .Q_N(_09153_),
    .Q(\am_sdr0.mix0.sin_in[0] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[1]$_DFF_P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1451),
    .D(_00009_),
    .Q_N(_09154_),
    .Q(\am_sdr0.mix0.sin_in[1] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[2]$_DFF_P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1452),
    .D(_00010_),
    .Q_N(_09155_),
    .Q(\am_sdr0.mix0.sin_in[2] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[3]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1453),
    .D(_00011_),
    .Q_N(_09156_),
    .Q(\am_sdr0.mix0.sin_in[3] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[4]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1454),
    .D(_00012_),
    .Q_N(_09157_),
    .Q(\am_sdr0.mix0.sin_in[4] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[5]$_DFF_P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1455),
    .D(_00013_),
    .Q_N(_09158_),
    .Q(\am_sdr0.mix0.sin_in[5] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[6]$_DFF_P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1456),
    .D(_00014_),
    .Q_N(_08129_),
    .Q(\am_sdr0.mix0.sin_in[6] ));
 sg13g2_dfrbp_1 \am_sdr0.nco0.sin0.data[7]$_SDFF_PN0_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1457),
    .D(_01103_),
    .Q_N(_08128_),
    .Q(\am_sdr0.mix0.sin_in[7] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.CS_q$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1458),
    .D(_01104_),
    .Q_N(_08127_),
    .Q(\am_sdr0.spi0.CS_q ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.CS_qq$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1459),
    .D(_01105_),
    .Q_N(_08126_),
    .Q(\am_sdr0.spi0.CS_qq ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.CS_qqq$_SDFF_PN0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1460),
    .D(_01106_),
    .Q_N(_08125_),
    .Q(\am_sdr0.spi0.CS_qqq ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.MOSI_q$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1461),
    .D(_01107_),
    .Q_N(_08124_),
    .Q(\am_sdr0.spi0.MOSI_q ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.MOSI_qq$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1462),
    .D(_01108_),
    .Q_N(_08123_),
    .Q(\am_sdr0.spi0.MOSI_qq ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.SCK_q$_SDFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1463),
    .D(_01109_),
    .Q_N(_08122_),
    .Q(\am_sdr0.spi0.SCK_q ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.SCK_qq$_SDFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1464),
    .D(_01110_),
    .Q_N(_08121_),
    .Q(\am_sdr0.spi0.SCK_qq ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.SCK_qqq$_SDFF_PN0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1465),
    .D(_01111_),
    .Q_N(_08120_),
    .Q(\am_sdr0.spi0.SCK_qqq ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.gain[0]$_SDFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1466),
    .D(_01112_),
    .Q_N(_08119_),
    .Q(\am_sdr0.gain_spi[0] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.gain[1]$_SDFFE_PN1N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1467),
    .D(_01113_),
    .Q_N(_08118_),
    .Q(\am_sdr0.gain_spi[1] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.gain[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1468),
    .D(_01114_),
    .Q_N(_00040_),
    .Q(\am_sdr0.gain_spi[2] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[0]$_SDFFE_PN1N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1469),
    .D(_01115_),
    .Q_N(_08117_),
    .Q(\am_sdr0.nco0.phase_inc[0] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[10]$_SDFFE_PN0N_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1470),
    .D(_01116_),
    .Q_N(_08116_),
    .Q(\am_sdr0.nco0.phase_inc[10] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[11]$_SDFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1471),
    .D(_01117_),
    .Q_N(_08115_),
    .Q(\am_sdr0.nco0.phase_inc[11] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[12]$_SDFFE_PN1N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1472),
    .D(_01118_),
    .Q_N(_08114_),
    .Q(\am_sdr0.nco0.phase_inc[12] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[13]$_SDFFE_PN0N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1473),
    .D(_01119_),
    .Q_N(_08113_),
    .Q(\am_sdr0.nco0.phase_inc[13] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[14]$_SDFFE_PN0N_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1474),
    .D(_01120_),
    .Q_N(_08112_),
    .Q(\am_sdr0.nco0.phase_inc[14] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[15]$_SDFFE_PN0N_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1475),
    .D(_01121_),
    .Q_N(_08111_),
    .Q(\am_sdr0.nco0.phase_inc[15] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[16]$_SDFFE_PN1N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1476),
    .D(_01122_),
    .Q_N(_08110_),
    .Q(\am_sdr0.nco0.phase_inc[16] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[17]$_SDFFE_PN1N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1477),
    .D(_01123_),
    .Q_N(_08109_),
    .Q(\am_sdr0.nco0.phase_inc[17] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[18]$_SDFFE_PN0N_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1478),
    .D(_01124_),
    .Q_N(_08108_),
    .Q(\am_sdr0.nco0.phase_inc[18] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[19]$_SDFFE_PN0N_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1479),
    .D(_01125_),
    .Q_N(_08107_),
    .Q(\am_sdr0.nco0.phase_inc[19] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[1]$_SDFFE_PN1N_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1480),
    .D(_01126_),
    .Q_N(_08106_),
    .Q(\am_sdr0.nco0.phase_inc[1] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[20]$_SDFFE_PN1N_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1481),
    .D(_01127_),
    .Q_N(_08105_),
    .Q(\am_sdr0.nco0.phase_inc[20] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[21]$_SDFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1482),
    .D(_01128_),
    .Q_N(_08104_),
    .Q(\am_sdr0.nco0.phase_inc[21] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[22]$_SDFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1483),
    .D(_01129_),
    .Q_N(_08103_),
    .Q(\am_sdr0.nco0.phase_inc[22] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[23]$_SDFFE_PN0N_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1484),
    .D(_01130_),
    .Q_N(_08102_),
    .Q(\am_sdr0.nco0.phase_inc[23] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[24]$_SDFFE_PN0N_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1485),
    .D(_01131_),
    .Q_N(_08101_),
    .Q(\am_sdr0.nco0.phase_inc[24] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[25]$_SDFFE_PN0N_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1486),
    .D(_01132_),
    .Q_N(_08100_),
    .Q(\am_sdr0.nco0.phase_inc[25] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1487),
    .D(_01133_),
    .Q_N(_08099_),
    .Q(\am_sdr0.nco0.phase_inc[2] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[3]$_SDFFE_PN1N_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1488),
    .D(_01134_),
    .Q_N(_08098_),
    .Q(\am_sdr0.nco0.phase_inc[3] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[4]$_SDFFE_PN0N_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1489),
    .D(_01135_),
    .Q_N(_08097_),
    .Q(\am_sdr0.nco0.phase_inc[4] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[5]$_SDFFE_PN1N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1490),
    .D(_01136_),
    .Q_N(_08096_),
    .Q(\am_sdr0.nco0.phase_inc[5] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[6]$_SDFFE_PN1N_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1491),
    .D(_01137_),
    .Q_N(_08095_),
    .Q(\am_sdr0.nco0.phase_inc[6] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[7]$_SDFFE_PN1N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1492),
    .D(_01138_),
    .Q_N(_08094_),
    .Q(\am_sdr0.nco0.phase_inc[7] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[8]$_SDFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1493),
    .D(_01139_),
    .Q_N(_08093_),
    .Q(\am_sdr0.nco0.phase_inc[8] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.phase_inc[9]$_SDFFE_PN1N_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1494),
    .D(_01140_),
    .Q_N(_08092_),
    .Q(\am_sdr0.nco0.phase_inc[9] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1495),
    .D(_01141_),
    .Q_N(_08091_),
    .Q(\am_sdr0.spi0.shift_reg[0] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1496),
    .D(_01142_),
    .Q_N(_08090_),
    .Q(\am_sdr0.spi0.shift_reg[10] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1497),
    .D(_01143_),
    .Q_N(_08089_),
    .Q(\am_sdr0.spi0.shift_reg[11] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[12]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1498),
    .D(_01144_),
    .Q_N(_08088_),
    .Q(\am_sdr0.spi0.shift_reg[12] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[13]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1499),
    .D(_01145_),
    .Q_N(_08087_),
    .Q(\am_sdr0.spi0.shift_reg[13] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[14]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1500),
    .D(_01146_),
    .Q_N(_08086_),
    .Q(\am_sdr0.spi0.shift_reg[14] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[15]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1501),
    .D(_01147_),
    .Q_N(_08085_),
    .Q(\am_sdr0.spi0.shift_reg[15] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[16]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1502),
    .D(_01148_),
    .Q_N(_08084_),
    .Q(\am_sdr0.spi0.shift_reg[16] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[17]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1503),
    .D(_01149_),
    .Q_N(_08083_),
    .Q(\am_sdr0.spi0.shift_reg[17] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[18]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1504),
    .D(_01150_),
    .Q_N(_08082_),
    .Q(\am_sdr0.spi0.shift_reg[18] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[19]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1505),
    .D(_01151_),
    .Q_N(_08081_),
    .Q(\am_sdr0.spi0.shift_reg[19] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1506),
    .D(_01152_),
    .Q_N(_08080_),
    .Q(\am_sdr0.spi0.shift_reg[1] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[20]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1507),
    .D(_01153_),
    .Q_N(_08079_),
    .Q(\am_sdr0.spi0.shift_reg[20] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[21]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1508),
    .D(_01154_),
    .Q_N(_08078_),
    .Q(\am_sdr0.spi0.shift_reg[21] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[22]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1509),
    .D(_01155_),
    .Q_N(_08077_),
    .Q(\am_sdr0.spi0.shift_reg[22] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[23]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1510),
    .D(_01156_),
    .Q_N(_08076_),
    .Q(\am_sdr0.spi0.shift_reg[23] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[24]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1511),
    .D(_01157_),
    .Q_N(_08075_),
    .Q(\am_sdr0.spi0.shift_reg[24] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[25]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1512),
    .D(_01158_),
    .Q_N(_08074_),
    .Q(\am_sdr0.spi0.shift_reg[25] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[26]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1513),
    .D(_01159_),
    .Q_N(_08073_),
    .Q(\am_sdr0.spi0.shift_reg[26] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[27]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1514),
    .D(_01160_),
    .Q_N(_08072_),
    .Q(\am_sdr0.spi0.shift_reg[27] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[28]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1515),
    .D(_01161_),
    .Q_N(_08071_),
    .Q(\am_sdr0.spi0.shift_reg[28] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1516),
    .D(_01162_),
    .Q_N(_08070_),
    .Q(\am_sdr0.spi0.shift_reg[2] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1517),
    .D(_01163_),
    .Q_N(_08069_),
    .Q(\am_sdr0.spi0.shift_reg[3] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1518),
    .D(_01164_),
    .Q_N(_08068_),
    .Q(\am_sdr0.spi0.shift_reg[4] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1519),
    .D(_01165_),
    .Q_N(_08067_),
    .Q(\am_sdr0.spi0.shift_reg[5] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1520),
    .D(_01166_),
    .Q_N(_08066_),
    .Q(\am_sdr0.spi0.shift_reg[6] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1521),
    .D(_01167_),
    .Q_N(_08065_),
    .Q(\am_sdr0.spi0.shift_reg[7] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1522),
    .D(_01168_),
    .Q_N(_08064_),
    .Q(\am_sdr0.spi0.shift_reg[8] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.shift_reg[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1523),
    .D(_01169_),
    .Q_N(_08063_),
    .Q(\am_sdr0.spi0.shift_reg[9] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.state[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1524),
    .D(_01170_),
    .Q_N(_08062_),
    .Q(\am_sdr0.spi0.state[0] ));
 sg13g2_dfrbp_1 \am_sdr0.spi0.state[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1525),
    .D(_01171_),
    .Q_N(_08061_),
    .Q(\am_sdr0.spi0.state[1] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[0]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[1]));
 sg13g2_buf_2 fanout7 (.A(_01701_),
    .X(net7));
 sg13g2_buf_2 fanout8 (.A(_01637_),
    .X(net8));
 sg13g2_buf_2 fanout9 (.A(_01588_),
    .X(net9));
 sg13g2_buf_2 fanout10 (.A(_06074_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_01041_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_01667_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_01662_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_01641_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_01595_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_01587_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_02449_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_02432_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_02374_),
    .X(net19));
 sg13g2_buf_4 fanout20 (.X(net20),
    .A(_02269_));
 sg13g2_buf_2 fanout21 (.A(_00397_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_01842_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_01742_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_01684_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_01583_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_02373_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_00612_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_02311_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_02307_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_01984_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_01981_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_01978_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_01566_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02524_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02497_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_01973_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_01733_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_01729_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_01721_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_01714_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_00173_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_01565_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_01398_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_01382_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_01379_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_01308_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_01214_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_08011_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_08004_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_07942_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_07829_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_07712_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_07594_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_07531_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_07381_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_07356_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_07333_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_07271_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_07200_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_07177_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_07175_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_07114_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_06934_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_06928_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_06911_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_06905_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06872_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06839_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_06673_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_06657_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_06635_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_06571_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_06472_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_06366_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_06239_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_06168_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_06068_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_06006_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_06000_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_05977_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_05882_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_05814_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_05806_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_05790_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_05544_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_05542_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_05521_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_05519_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_05491_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_05467_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_05447_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_05370_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_05357_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_05254_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_05246_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_05204_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_05091_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_05036_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04928_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_04842_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04719_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04697_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04617_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_04544_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_04521_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_04363_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_04277_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_04270_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_04254_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_04247_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04220_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_04186_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_04012_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_03989_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_03963_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_03872_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_03792_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_03706_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03614_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_03541_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_03429_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_03405_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_03373_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_03264_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_03241_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_03196_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_03096_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_02992_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_02969_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_02839_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_02780_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_02527_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_02504_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_02498_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_02496_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_01687_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_01598_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_01564_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_01447_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_01381_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_01378_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_01375_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_01371_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_07661_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_07450_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_07354_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_07331_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_07198_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_06737_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_06672_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_06002_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_05979_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_05830_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_05358_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_05356_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04721_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04699_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_04542_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_04519_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_04198_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_04075_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_04011_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03418_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03414_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03395_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03391_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_03254_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_03250_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_03231_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03227_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03004_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_02982_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_02978_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_02959_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_02955_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_02786_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_02781_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_02729_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_02726_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_02718_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_02699_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_02544_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_02521_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_02501_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_01719_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_01716_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_01599_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_01592_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_01589_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_01456_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_01446_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_01377_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_08026_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_08025_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_07604_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_07387_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_07382_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_07366_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_07364_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_07340_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_07317_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_07184_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_07161_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_06919_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_06896_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_06786_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_06728_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_06676_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_06664_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_06552_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_06251_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_06099_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_06071_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_05983_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_05960_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_05810_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_05787_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_05549_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_05525_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_05502_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_05392_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_05372_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_05280_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_05278_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_05274_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_05264_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_04774_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_04691_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_04536_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_04513_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_04271_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_04248_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_04244_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_04143_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_04113_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_04067_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_04066_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_04014_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_04006_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_04002_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_03993_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_03443_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_03098_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_03002_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_02870_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_02809_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_02783_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_02725_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_02721_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_02717_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_01968_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_01847_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_01760_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_01743_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_01723_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_01710_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_01560_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_01500_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_01445_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_07747_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_07735_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_07714_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_07533_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_07520_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_07502_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_07421_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_07363_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_06805_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_06729_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_06667_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_06663_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_06481_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_06400_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_06326_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_06179_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_06170_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_06122_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_06113_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_06097_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_06070_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_06050_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_06008_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_05327_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_05277_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_05273_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_05263_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_04870_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_04858_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_04830_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_04773_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_04001_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_03992_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_03502_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_03498_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_03442_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_03440_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_02808_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_02597_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_01966_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_01846_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_01718_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_01574_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_01559_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_01524_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_01513_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_01499_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_01496_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_01469_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_01463_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_01444_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_07746_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_07704_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_07690_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_07646_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_07607_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_07546_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_07532_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_07507_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_07481_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_07472_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_07462_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_07457_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_07447_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_07431_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_07385_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_06731_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_06390_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_06375_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_06255_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_06151_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_06141_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_06131_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_06125_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_06106_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_06084_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_06069_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_06045_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_06026_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_06007_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_04992_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_04839_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_04818_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_04802_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_04788_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_04775_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_04766_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_03991_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_03768_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_03759_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_03712_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_03703_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_03683_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_03655_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_03634_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_03560_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_03551_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_03542_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_03529_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_03519_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_03490_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_03450_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_03444_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_01736_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_01558_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_01502_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_01495_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_01462_),
    .X(net367));
 sg13g2_tielo _17186__368 (.L_LO(net368));
 sg13g2_tielo _17187__369 (.L_LO(net369));
 sg13g2_tielo _17188__370 (.L_LO(net370));
 sg13g2_tielo _17189__371 (.L_LO(net371));
 sg13g2_tielo _17190__372 (.L_LO(net372));
 sg13g2_tielo _17191__373 (.L_LO(net373));
 sg13g2_tielo _17192__374 (.L_LO(net374));
 sg13g2_tielo _17193__375 (.L_LO(net375));
 sg13g2_tielo _17194__376 (.L_LO(net376));
 sg13g2_tielo _17195__377 (.L_LO(net377));
 sg13g2_tielo _17196__378 (.L_LO(net378));
 sg13g2_tielo _17197__379 (.L_LO(net379));
 sg13g2_tielo _17198__380 (.L_LO(net380));
 sg13g2_tielo _17199__381 (.L_LO(net381));
 sg13g2_tielo _17200__382 (.L_LO(net382));
 sg13g2_tielo _17201__383 (.L_LO(net383));
 sg13g2_tielo _17204__384 (.L_LO(net384));
 sg13g2_tielo _17205__385 (.L_LO(net385));
 sg13g2_tielo _17206__386 (.L_LO(net386));
 sg13g2_tielo _17207__387 (.L_LO(net387));
 sg13g2_tielo _17208__388 (.L_LO(net388));
 sg13g2_tielo _17209__389 (.L_LO(net389));
 sg13g2_tiehi \am_sdr0.am0.a[0]$_SDFFCE_PP0P__391  (.L_HI(net391));
 sg13g2_tiehi \am_sdr0.am0.a[10]$_DFFE_PP__392  (.L_HI(net392));
 sg13g2_tiehi \am_sdr0.am0.a[11]$_DFFE_PP__393  (.L_HI(net393));
 sg13g2_tiehi \am_sdr0.am0.a[12]$_DFFE_PP__394  (.L_HI(net394));
 sg13g2_tiehi \am_sdr0.am0.a[13]$_DFFE_PP__395  (.L_HI(net395));
 sg13g2_tiehi \am_sdr0.am0.a[14]$_DFFE_PP__396  (.L_HI(net396));
 sg13g2_tiehi \am_sdr0.am0.a[15]$_DFFE_PP__397  (.L_HI(net397));
 sg13g2_tiehi \am_sdr0.am0.a[1]$_SDFFCE_PP0P__398  (.L_HI(net398));
 sg13g2_tiehi \am_sdr0.am0.a[2]$_DFFE_PP__399  (.L_HI(net399));
 sg13g2_tiehi \am_sdr0.am0.a[3]$_DFFE_PP__400  (.L_HI(net400));
 sg13g2_tiehi \am_sdr0.am0.a[4]$_DFFE_PP__401  (.L_HI(net401));
 sg13g2_tiehi \am_sdr0.am0.a[5]$_DFFE_PP__402  (.L_HI(net402));
 sg13g2_tiehi \am_sdr0.am0.a[6]$_DFFE_PP__403  (.L_HI(net403));
 sg13g2_tiehi \am_sdr0.am0.a[7]$_DFFE_PP__404  (.L_HI(net404));
 sg13g2_tiehi \am_sdr0.am0.a[8]$_DFFE_PP__405  (.L_HI(net405));
 sg13g2_tiehi \am_sdr0.am0.a[9]$_DFFE_PP__406  (.L_HI(net406));
 sg13g2_tiehi \am_sdr0.am0.count2[0]$_SDFFCE_PN0P__407  (.L_HI(net407));
 sg13g2_tiehi \am_sdr0.am0.count2[1]$_SDFFCE_PN0P__408  (.L_HI(net408));
 sg13g2_tiehi \am_sdr0.am0.count2[2]$_SDFFCE_PN0P__409  (.L_HI(net409));
 sg13g2_tiehi \am_sdr0.am0.count2[3]$_SDFFCE_PN0P__410  (.L_HI(net410));
 sg13g2_tiehi \am_sdr0.am0.count[0]$_SDFFCE_PN0P__411  (.L_HI(net411));
 sg13g2_tiehi \am_sdr0.am0.count[1]$_SDFFCE_PN0P__412  (.L_HI(net412));
 sg13g2_tiehi \am_sdr0.am0.demod_out[10]$_SDFFE_PN0P__413  (.L_HI(net413));
 sg13g2_tiehi \am_sdr0.am0.demod_out[11]$_SDFFE_PN0P__414  (.L_HI(net414));
 sg13g2_tiehi \am_sdr0.am0.demod_out[12]$_SDFFE_PN0P__415  (.L_HI(net415));
 sg13g2_tiehi \am_sdr0.am0.demod_out[13]$_SDFFE_PN0P__416  (.L_HI(net416));
 sg13g2_tiehi \am_sdr0.am0.demod_out[14]$_SDFFE_PN0P__417  (.L_HI(net417));
 sg13g2_tiehi \am_sdr0.am0.demod_out[15]$_SDFFE_PN0P__418  (.L_HI(net418));
 sg13g2_tiehi \am_sdr0.am0.demod_out[8]$_SDFFE_PN0P__419  (.L_HI(net419));
 sg13g2_tiehi \am_sdr0.am0.demod_out[9]$_SDFFE_PN0P__420  (.L_HI(net420));
 sg13g2_tiehi \am_sdr0.am0.left[0]$_SDFFCE_PN0P__421  (.L_HI(net421));
 sg13g2_tiehi \am_sdr0.am0.left[1]$_SDFFCE_PN0P__422  (.L_HI(net422));
 sg13g2_tiehi \am_sdr0.am0.left[2]$_SDFFCE_PN0P__423  (.L_HI(net423));
 sg13g2_tiehi \am_sdr0.am0.left[3]$_SDFFCE_PN0P__424  (.L_HI(net424));
 sg13g2_tiehi \am_sdr0.am0.left[4]$_SDFFCE_PN0P__425  (.L_HI(net425));
 sg13g2_tiehi \am_sdr0.am0.left[5]$_SDFFCE_PN0P__426  (.L_HI(net426));
 sg13g2_tiehi \am_sdr0.am0.left[6]$_SDFFCE_PN0P__427  (.L_HI(net427));
 sg13g2_tiehi \am_sdr0.am0.left[7]$_SDFFCE_PN0P__428  (.L_HI(net428));
 sg13g2_tiehi \am_sdr0.am0.left[8]$_SDFFCE_PN0P__429  (.L_HI(net429));
 sg13g2_tiehi \am_sdr0.am0.left[9]$_SDFFCE_PN0P__430  (.L_HI(net430));
 sg13g2_tiehi \am_sdr0.am0.m_count[0]$_SDFFCE_PP0P__431  (.L_HI(net431));
 sg13g2_tiehi \am_sdr0.am0.m_count[1]$_SDFFCE_PP0P__432  (.L_HI(net432));
 sg13g2_tiehi \am_sdr0.am0.m_count[2]$_SDFFCE_PP0P__433  (.L_HI(net433));
 sg13g2_tiehi \am_sdr0.am0.m_count[3]$_SDFFCE_PP0P__434  (.L_HI(net434));
 sg13g2_tiehi \am_sdr0.am0.multA[0]$_DFFE_PP__435  (.L_HI(net435));
 sg13g2_tiehi \am_sdr0.am0.multA[10]$_DFFE_PP__436  (.L_HI(net436));
 sg13g2_tiehi \am_sdr0.am0.multA[11]$_DFFE_PP__437  (.L_HI(net437));
 sg13g2_tiehi \am_sdr0.am0.multA[12]$_DFFE_PP__438  (.L_HI(net438));
 sg13g2_tiehi \am_sdr0.am0.multA[13]$_DFFE_PP__439  (.L_HI(net439));
 sg13g2_tiehi \am_sdr0.am0.multA[14]$_DFFE_PP__440  (.L_HI(net440));
 sg13g2_tiehi \am_sdr0.am0.multA[15]$_DFFE_PP__441  (.L_HI(net441));
 sg13g2_tiehi \am_sdr0.am0.multA[16]$_DFFE_PP__442  (.L_HI(net442));
 sg13g2_tiehi \am_sdr0.am0.multA[1]$_DFFE_PP__443  (.L_HI(net443));
 sg13g2_tiehi \am_sdr0.am0.multA[2]$_DFFE_PP__444  (.L_HI(net444));
 sg13g2_tiehi \am_sdr0.am0.multA[3]$_DFFE_PP__445  (.L_HI(net445));
 sg13g2_tiehi \am_sdr0.am0.multA[4]$_DFFE_PP__446  (.L_HI(net446));
 sg13g2_tiehi \am_sdr0.am0.multA[5]$_DFFE_PP__447  (.L_HI(net447));
 sg13g2_tiehi \am_sdr0.am0.multA[6]$_DFFE_PP__448  (.L_HI(net448));
 sg13g2_tiehi \am_sdr0.am0.multA[7]$_DFFE_PP__449  (.L_HI(net449));
 sg13g2_tiehi \am_sdr0.am0.multA[8]$_DFFE_PP__450  (.L_HI(net450));
 sg13g2_tiehi \am_sdr0.am0.multA[9]$_DFFE_PP__451  (.L_HI(net451));
 sg13g2_tiehi \am_sdr0.am0.multB[0]$_DFFE_PP__452  (.L_HI(net452));
 sg13g2_tiehi \am_sdr0.am0.multB[1]$_DFFE_PP__453  (.L_HI(net453));
 sg13g2_tiehi \am_sdr0.am0.multB[2]$_DFFE_PP__454  (.L_HI(net454));
 sg13g2_tiehi \am_sdr0.am0.multB[3]$_DFFE_PP__455  (.L_HI(net455));
 sg13g2_tiehi \am_sdr0.am0.multB[4]$_DFFE_PP__456  (.L_HI(net456));
 sg13g2_tiehi \am_sdr0.am0.multB[5]$_DFFE_PP__457  (.L_HI(net457));
 sg13g2_tiehi \am_sdr0.am0.multB[6]$_DFFE_PP__458  (.L_HI(net458));
 sg13g2_tiehi \am_sdr0.am0.multB[7]$_DFFE_PP__459  (.L_HI(net459));
 sg13g2_tiehi \am_sdr0.am0.q[0]$_SDFFCE_PN0P__460  (.L_HI(net460));
 sg13g2_tiehi \am_sdr0.am0.q[1]$_SDFFCE_PN0P__461  (.L_HI(net461));
 sg13g2_tiehi \am_sdr0.am0.q[2]$_SDFFCE_PN0P__462  (.L_HI(net462));
 sg13g2_tiehi \am_sdr0.am0.q[3]$_SDFFCE_PN0P__463  (.L_HI(net463));
 sg13g2_tiehi \am_sdr0.am0.q[4]$_SDFFCE_PN0P__464  (.L_HI(net464));
 sg13g2_tiehi \am_sdr0.am0.q[5]$_SDFFCE_PN0P__465  (.L_HI(net465));
 sg13g2_tiehi \am_sdr0.am0.q[6]$_SDFFCE_PN0P__466  (.L_HI(net466));
 sg13g2_tiehi \am_sdr0.am0.q[7]$_SDFFCE_PN0P__467  (.L_HI(net467));
 sg13g2_tiehi \am_sdr0.am0.r[0]$_SDFFCE_PN0P__468  (.L_HI(net468));
 sg13g2_tiehi \am_sdr0.am0.r[1]$_SDFFCE_PN0P__469  (.L_HI(net469));
 sg13g2_tiehi \am_sdr0.am0.r[2]$_SDFFCE_PN0P__470  (.L_HI(net470));
 sg13g2_tiehi \am_sdr0.am0.r[3]$_SDFFCE_PN0P__471  (.L_HI(net471));
 sg13g2_tiehi \am_sdr0.am0.r[4]$_SDFFCE_PN0P__472  (.L_HI(net472));
 sg13g2_tiehi \am_sdr0.am0.r[5]$_SDFFCE_PN0P__473  (.L_HI(net473));
 sg13g2_tiehi \am_sdr0.am0.r[6]$_SDFFCE_PN0P__474  (.L_HI(net474));
 sg13g2_tiehi \am_sdr0.am0.r[7]$_SDFFCE_PN0P__475  (.L_HI(net475));
 sg13g2_tiehi \am_sdr0.am0.r[9]$_SDFFCE_PN0P__476  (.L_HI(net476));
 sg13g2_tiehi \am_sdr0.am0.right[0]$_SDFFCE_PN0P__477  (.L_HI(net477));
 sg13g2_tiehi \am_sdr0.am0.right[1]$_SDFFCE_PN0P__478  (.L_HI(net478));
 sg13g2_tiehi \am_sdr0.am0.right[2]$_SDFFCE_PN0P__479  (.L_HI(net479));
 sg13g2_tiehi \am_sdr0.am0.right[3]$_SDFFCE_PN0P__480  (.L_HI(net480));
 sg13g2_tiehi \am_sdr0.am0.right[4]$_SDFFCE_PN0P__481  (.L_HI(net481));
 sg13g2_tiehi \am_sdr0.am0.right[5]$_SDFFCE_PN0P__482  (.L_HI(net482));
 sg13g2_tiehi \am_sdr0.am0.right[6]$_SDFFCE_PN0P__483  (.L_HI(net483));
 sg13g2_tiehi \am_sdr0.am0.right[7]$_SDFFCE_PN0P__484  (.L_HI(net484));
 sg13g2_tiehi \am_sdr0.am0.right[8]$_SDFFCE_PN0P__485  (.L_HI(net485));
 sg13g2_tiehi \am_sdr0.am0.right[9]$_SDFFCE_PN0P__486  (.L_HI(net486));
 sg13g2_tiehi \am_sdr0.am0.sqrt_done$_DFFE_PP__487  (.L_HI(net487));
 sg13g2_tiehi \am_sdr0.am0.sqrt_state[0]$_SDFFE_PN0P__488  (.L_HI(net488));
 sg13g2_tiehi \am_sdr0.am0.sqrt_state[1]$_SDFFE_PN0P__489  (.L_HI(net489));
 sg13g2_tiehi \am_sdr0.am0.state[0]$_DFF_P__490  (.L_HI(net490));
 sg13g2_tiehi \am_sdr0.am0.state[1]$_DFF_P__491  (.L_HI(net491));
 sg13g2_tiehi \am_sdr0.am0.state[2]$_DFF_P__492  (.L_HI(net492));
 sg13g2_tiehi \am_sdr0.am0.state[3]$_DFF_P__493  (.L_HI(net493));
 sg13g2_tiehi \am_sdr0.am0.state[4]$_DFF_P__494  (.L_HI(net494));
 sg13g2_tiehi \am_sdr0.am0.state[5]$_DFF_P__495  (.L_HI(net495));
 sg13g2_tiehi \am_sdr0.am0.state[6]$_DFF_P__496  (.L_HI(net496));
 sg13g2_tiehi \am_sdr0.am0.sum[0]$_SDFFCE_PP0P__497  (.L_HI(net497));
 sg13g2_tiehi \am_sdr0.am0.sum[10]$_SDFFCE_PP0P__498  (.L_HI(net498));
 sg13g2_tiehi \am_sdr0.am0.sum[11]$_SDFFCE_PP0P__499  (.L_HI(net499));
 sg13g2_tiehi \am_sdr0.am0.sum[12]$_SDFFCE_PP0P__500  (.L_HI(net500));
 sg13g2_tiehi \am_sdr0.am0.sum[13]$_SDFFCE_PP0P__501  (.L_HI(net501));
 sg13g2_tiehi \am_sdr0.am0.sum[14]$_SDFFCE_PP0P__502  (.L_HI(net502));
 sg13g2_tiehi \am_sdr0.am0.sum[15]$_SDFFCE_PP0P__503  (.L_HI(net503));
 sg13g2_tiehi \am_sdr0.am0.sum[16]$_SDFFCE_PP0P__504  (.L_HI(net504));
 sg13g2_tiehi \am_sdr0.am0.sum[1]$_SDFFCE_PP0P__505  (.L_HI(net505));
 sg13g2_tiehi \am_sdr0.am0.sum[2]$_SDFFCE_PP0P__506  (.L_HI(net506));
 sg13g2_tiehi \am_sdr0.am0.sum[3]$_SDFFCE_PP0P__507  (.L_HI(net507));
 sg13g2_tiehi \am_sdr0.am0.sum[4]$_SDFFCE_PP0P__508  (.L_HI(net508));
 sg13g2_tiehi \am_sdr0.am0.sum[5]$_SDFFCE_PP0P__509  (.L_HI(net509));
 sg13g2_tiehi \am_sdr0.am0.sum[6]$_SDFFCE_PP0P__510  (.L_HI(net510));
 sg13g2_tiehi \am_sdr0.am0.sum[7]$_SDFFCE_PP0P__511  (.L_HI(net511));
 sg13g2_tiehi \am_sdr0.am0.sum[8]$_SDFFCE_PP0P__512  (.L_HI(net512));
 sg13g2_tiehi \am_sdr0.am0.sum[9]$_SDFFCE_PP0P__513  (.L_HI(net513));
 sg13g2_tiehi \am_sdr0.cic0.comb1[0]$_SDFFE_PN0P__514  (.L_HI(net514));
 sg13g2_tiehi \am_sdr0.cic0.comb1[10]$_SDFFE_PN0P__515  (.L_HI(net515));
 sg13g2_tiehi \am_sdr0.cic0.comb1[11]$_SDFFE_PN0P__516  (.L_HI(net516));
 sg13g2_tiehi \am_sdr0.cic0.comb1[12]$_SDFFE_PN0P__517  (.L_HI(net517));
 sg13g2_tiehi \am_sdr0.cic0.comb1[13]$_SDFFE_PN0P__518  (.L_HI(net518));
 sg13g2_tiehi \am_sdr0.cic0.comb1[14]$_SDFFE_PN0P__519  (.L_HI(net519));
 sg13g2_tiehi \am_sdr0.cic0.comb1[15]$_SDFFE_PN0P__520  (.L_HI(net520));
 sg13g2_tiehi \am_sdr0.cic0.comb1[16]$_SDFFE_PN0P__521  (.L_HI(net521));
 sg13g2_tiehi \am_sdr0.cic0.comb1[17]$_SDFFE_PN0P__522  (.L_HI(net522));
 sg13g2_tiehi \am_sdr0.cic0.comb1[18]$_SDFFE_PN0P__523  (.L_HI(net523));
 sg13g2_tiehi \am_sdr0.cic0.comb1[19]$_SDFFE_PN0P__524  (.L_HI(net524));
 sg13g2_tiehi \am_sdr0.cic0.comb1[1]$_SDFFE_PN0P__525  (.L_HI(net525));
 sg13g2_tiehi \am_sdr0.cic0.comb1[2]$_SDFFE_PN0P__526  (.L_HI(net526));
 sg13g2_tiehi \am_sdr0.cic0.comb1[3]$_SDFFE_PN0P__527  (.L_HI(net527));
 sg13g2_tiehi \am_sdr0.cic0.comb1[4]$_SDFFE_PN0P__528  (.L_HI(net528));
 sg13g2_tiehi \am_sdr0.cic0.comb1[5]$_SDFFE_PN0P__529  (.L_HI(net529));
 sg13g2_tiehi \am_sdr0.cic0.comb1[6]$_SDFFE_PN0P__530  (.L_HI(net530));
 sg13g2_tiehi \am_sdr0.cic0.comb1[7]$_SDFFE_PN0P__531  (.L_HI(net531));
 sg13g2_tiehi \am_sdr0.cic0.comb1[8]$_SDFFE_PN0P__532  (.L_HI(net532));
 sg13g2_tiehi \am_sdr0.cic0.comb1[9]$_SDFFE_PN0P__533  (.L_HI(net533));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[0]$_SDFFE_PN0P__534  (.L_HI(net534));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[10]$_SDFFE_PN0P__535  (.L_HI(net535));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[11]$_SDFFE_PN0P__536  (.L_HI(net536));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[12]$_SDFFE_PN0P__537  (.L_HI(net537));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[13]$_SDFFE_PN0P__538  (.L_HI(net538));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[14]$_SDFFE_PN0P__539  (.L_HI(net539));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[15]$_SDFFE_PN0P__540  (.L_HI(net540));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[16]$_SDFFE_PN0P__541  (.L_HI(net541));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[17]$_SDFFE_PN0P__542  (.L_HI(net542));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[18]$_SDFFE_PN0P__543  (.L_HI(net543));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[19]$_SDFFE_PN0P__544  (.L_HI(net544));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[1]$_SDFFE_PN0P__545  (.L_HI(net545));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[2]$_SDFFE_PN0P__546  (.L_HI(net546));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[3]$_SDFFE_PN0P__547  (.L_HI(net547));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[4]$_SDFFE_PN0P__548  (.L_HI(net548));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[5]$_SDFFE_PN0P__549  (.L_HI(net549));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[6]$_SDFFE_PN0P__550  (.L_HI(net550));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[7]$_SDFFE_PN0P__551  (.L_HI(net551));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[8]$_SDFFE_PN0P__552  (.L_HI(net552));
 sg13g2_tiehi \am_sdr0.cic0.comb1_in_del[9]$_SDFFE_PN0P__553  (.L_HI(net553));
 sg13g2_tiehi \am_sdr0.cic0.comb2[0]$_SDFFE_PN0P__554  (.L_HI(net554));
 sg13g2_tiehi \am_sdr0.cic0.comb2[10]$_SDFFE_PN0P__555  (.L_HI(net555));
 sg13g2_tiehi \am_sdr0.cic0.comb2[11]$_SDFFE_PN0P__556  (.L_HI(net556));
 sg13g2_tiehi \am_sdr0.cic0.comb2[12]$_SDFFE_PN0P__557  (.L_HI(net557));
 sg13g2_tiehi \am_sdr0.cic0.comb2[13]$_SDFFE_PN0P__558  (.L_HI(net558));
 sg13g2_tiehi \am_sdr0.cic0.comb2[14]$_SDFFE_PN0P__559  (.L_HI(net559));
 sg13g2_tiehi \am_sdr0.cic0.comb2[15]$_SDFFE_PN0P__560  (.L_HI(net560));
 sg13g2_tiehi \am_sdr0.cic0.comb2[16]$_SDFFE_PN0P__561  (.L_HI(net561));
 sg13g2_tiehi \am_sdr0.cic0.comb2[17]$_SDFFE_PN0P__562  (.L_HI(net562));
 sg13g2_tiehi \am_sdr0.cic0.comb2[18]$_SDFFE_PN0P__563  (.L_HI(net563));
 sg13g2_tiehi \am_sdr0.cic0.comb2[19]$_SDFFE_PN0P__564  (.L_HI(net564));
 sg13g2_tiehi \am_sdr0.cic0.comb2[1]$_SDFFE_PN0P__565  (.L_HI(net565));
 sg13g2_tiehi \am_sdr0.cic0.comb2[2]$_SDFFE_PN0P__566  (.L_HI(net566));
 sg13g2_tiehi \am_sdr0.cic0.comb2[3]$_SDFFE_PN0P__567  (.L_HI(net567));
 sg13g2_tiehi \am_sdr0.cic0.comb2[4]$_SDFFE_PN0P__568  (.L_HI(net568));
 sg13g2_tiehi \am_sdr0.cic0.comb2[5]$_SDFFE_PN0P__569  (.L_HI(net569));
 sg13g2_tiehi \am_sdr0.cic0.comb2[6]$_SDFFE_PN0P__570  (.L_HI(net570));
 sg13g2_tiehi \am_sdr0.cic0.comb2[7]$_SDFFE_PN0P__571  (.L_HI(net571));
 sg13g2_tiehi \am_sdr0.cic0.comb2[8]$_SDFFE_PN0P__572  (.L_HI(net572));
 sg13g2_tiehi \am_sdr0.cic0.comb2[9]$_SDFFE_PN0P__573  (.L_HI(net573));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[0]$_SDFFE_PN0P__574  (.L_HI(net574));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[10]$_SDFFE_PN0P__575  (.L_HI(net575));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[11]$_SDFFE_PN0P__576  (.L_HI(net576));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[12]$_SDFFE_PN0P__577  (.L_HI(net577));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[13]$_SDFFE_PN0P__578  (.L_HI(net578));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[14]$_SDFFE_PN0P__579  (.L_HI(net579));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[15]$_SDFFE_PN0P__580  (.L_HI(net580));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[16]$_SDFFE_PN0P__581  (.L_HI(net581));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[17]$_SDFFE_PN0P__582  (.L_HI(net582));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[18]$_SDFFE_PN0P__583  (.L_HI(net583));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[19]$_SDFFE_PN0P__584  (.L_HI(net584));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[1]$_SDFFE_PN0P__585  (.L_HI(net585));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[2]$_SDFFE_PN0P__586  (.L_HI(net586));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[3]$_SDFFE_PN0P__587  (.L_HI(net587));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[4]$_SDFFE_PN0P__588  (.L_HI(net588));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[5]$_SDFFE_PN0P__589  (.L_HI(net589));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[6]$_SDFFE_PN0P__590  (.L_HI(net590));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[7]$_SDFFE_PN0P__591  (.L_HI(net591));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[8]$_SDFFE_PN0P__592  (.L_HI(net592));
 sg13g2_tiehi \am_sdr0.cic0.comb2_in_del[9]$_SDFFE_PN0P__593  (.L_HI(net593));
 sg13g2_tiehi \am_sdr0.cic0.comb3[12]$_SDFFE_PN0P__594  (.L_HI(net594));
 sg13g2_tiehi \am_sdr0.cic0.comb3[13]$_SDFFE_PN0P__595  (.L_HI(net595));
 sg13g2_tiehi \am_sdr0.cic0.comb3[14]$_SDFFE_PN0P__596  (.L_HI(net596));
 sg13g2_tiehi \am_sdr0.cic0.comb3[15]$_SDFFE_PN0P__597  (.L_HI(net597));
 sg13g2_tiehi \am_sdr0.cic0.comb3[16]$_SDFFE_PN0P__598  (.L_HI(net598));
 sg13g2_tiehi \am_sdr0.cic0.comb3[17]$_SDFFE_PN0P__599  (.L_HI(net599));
 sg13g2_tiehi \am_sdr0.cic0.comb3[18]$_SDFFE_PN0P__600  (.L_HI(net600));
 sg13g2_tiehi \am_sdr0.cic0.comb3[19]$_SDFFE_PN0P__601  (.L_HI(net601));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[0]$_SDFFE_PN0P__602  (.L_HI(net602));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[10]$_SDFFE_PN0P__603  (.L_HI(net603));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[11]$_SDFFE_PN0P__604  (.L_HI(net604));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[12]$_SDFFE_PN0P__605  (.L_HI(net605));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[13]$_SDFFE_PN0P__606  (.L_HI(net606));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[14]$_SDFFE_PN0P__607  (.L_HI(net607));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[15]$_SDFFE_PN0P__608  (.L_HI(net608));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[16]$_SDFFE_PN0P__609  (.L_HI(net609));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[17]$_SDFFE_PN0P__610  (.L_HI(net610));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[18]$_SDFFE_PN0P__611  (.L_HI(net611));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[19]$_SDFFE_PN0P__612  (.L_HI(net612));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[1]$_SDFFE_PN0P__613  (.L_HI(net613));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[2]$_SDFFE_PN0P__614  (.L_HI(net614));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[3]$_SDFFE_PN0P__615  (.L_HI(net615));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[4]$_SDFFE_PN0P__616  (.L_HI(net616));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[5]$_SDFFE_PN0P__617  (.L_HI(net617));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[6]$_SDFFE_PN0P__618  (.L_HI(net618));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[7]$_SDFFE_PN0P__619  (.L_HI(net619));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[8]$_SDFFE_PN0P__620  (.L_HI(net620));
 sg13g2_tiehi \am_sdr0.cic0.comb3_in_del[9]$_SDFFE_PN0P__621  (.L_HI(net621));
 sg13g2_tiehi \am_sdr0.cic0.count[0]$_SDFF_PP0__622  (.L_HI(net622));
 sg13g2_tiehi \am_sdr0.cic0.count[1]$_SDFF_PP0__623  (.L_HI(net623));
 sg13g2_tiehi \am_sdr0.cic0.count[2]$_SDFF_PP0__624  (.L_HI(net624));
 sg13g2_tiehi \am_sdr0.cic0.count[3]$_SDFF_PP0__625  (.L_HI(net625));
 sg13g2_tiehi \am_sdr0.cic0.count[4]$_SDFF_PP0__626  (.L_HI(net626));
 sg13g2_tiehi \am_sdr0.cic0.count[5]$_SDFF_PP0__627  (.L_HI(net627));
 sg13g2_tiehi \am_sdr0.cic0.count[6]$_SDFF_PP0__628  (.L_HI(net628));
 sg13g2_tiehi \am_sdr0.cic0.count[7]$_SDFF_PP0__629  (.L_HI(net629));
 sg13g2_tiehi \am_sdr0.cic0.integ1[0]$_SDFF_PN0__630  (.L_HI(net630));
 sg13g2_tiehi \am_sdr0.cic0.integ1[10]$_SDFF_PN0__631  (.L_HI(net631));
 sg13g2_tiehi \am_sdr0.cic0.integ1[11]$_SDFF_PN0__632  (.L_HI(net632));
 sg13g2_tiehi \am_sdr0.cic0.integ1[12]$_SDFF_PN0__633  (.L_HI(net633));
 sg13g2_tiehi \am_sdr0.cic0.integ1[13]$_SDFF_PN0__634  (.L_HI(net634));
 sg13g2_tiehi \am_sdr0.cic0.integ1[14]$_SDFF_PN0__635  (.L_HI(net635));
 sg13g2_tiehi \am_sdr0.cic0.integ1[15]$_SDFF_PN0__636  (.L_HI(net636));
 sg13g2_tiehi \am_sdr0.cic0.integ1[16]$_SDFF_PN0__637  (.L_HI(net637));
 sg13g2_tiehi \am_sdr0.cic0.integ1[17]$_SDFF_PN0__638  (.L_HI(net638));
 sg13g2_tiehi \am_sdr0.cic0.integ1[18]$_SDFF_PN0__639  (.L_HI(net639));
 sg13g2_tiehi \am_sdr0.cic0.integ1[19]$_SDFF_PN0__640  (.L_HI(net640));
 sg13g2_tiehi \am_sdr0.cic0.integ1[1]$_SDFF_PN0__641  (.L_HI(net641));
 sg13g2_tiehi \am_sdr0.cic0.integ1[20]$_SDFF_PN0__642  (.L_HI(net642));
 sg13g2_tiehi \am_sdr0.cic0.integ1[21]$_SDFF_PN0__643  (.L_HI(net643));
 sg13g2_tiehi \am_sdr0.cic0.integ1[22]$_SDFF_PN0__644  (.L_HI(net644));
 sg13g2_tiehi \am_sdr0.cic0.integ1[23]$_SDFF_PN0__645  (.L_HI(net645));
 sg13g2_tiehi \am_sdr0.cic0.integ1[24]$_SDFF_PN0__646  (.L_HI(net646));
 sg13g2_tiehi \am_sdr0.cic0.integ1[25]$_SDFF_PN0__647  (.L_HI(net647));
 sg13g2_tiehi \am_sdr0.cic0.integ1[2]$_SDFF_PN0__648  (.L_HI(net648));
 sg13g2_tiehi \am_sdr0.cic0.integ1[3]$_SDFF_PN0__649  (.L_HI(net649));
 sg13g2_tiehi \am_sdr0.cic0.integ1[4]$_SDFF_PN0__650  (.L_HI(net650));
 sg13g2_tiehi \am_sdr0.cic0.integ1[5]$_SDFF_PN0__651  (.L_HI(net651));
 sg13g2_tiehi \am_sdr0.cic0.integ1[6]$_SDFF_PN0__652  (.L_HI(net652));
 sg13g2_tiehi \am_sdr0.cic0.integ1[7]$_SDFF_PN0__653  (.L_HI(net653));
 sg13g2_tiehi \am_sdr0.cic0.integ1[8]$_SDFF_PN0__654  (.L_HI(net654));
 sg13g2_tiehi \am_sdr0.cic0.integ1[9]$_SDFF_PN0__655  (.L_HI(net655));
 sg13g2_tiehi \am_sdr0.cic0.integ2[0]$_SDFF_PN0__656  (.L_HI(net656));
 sg13g2_tiehi \am_sdr0.cic0.integ2[10]$_SDFF_PN0__657  (.L_HI(net657));
 sg13g2_tiehi \am_sdr0.cic0.integ2[11]$_SDFF_PN0__658  (.L_HI(net658));
 sg13g2_tiehi \am_sdr0.cic0.integ2[12]$_SDFF_PN0__659  (.L_HI(net659));
 sg13g2_tiehi \am_sdr0.cic0.integ2[13]$_SDFF_PN0__660  (.L_HI(net660));
 sg13g2_tiehi \am_sdr0.cic0.integ2[14]$_SDFF_PN0__661  (.L_HI(net661));
 sg13g2_tiehi \am_sdr0.cic0.integ2[15]$_SDFF_PN0__662  (.L_HI(net662));
 sg13g2_tiehi \am_sdr0.cic0.integ2[16]$_SDFF_PN0__663  (.L_HI(net663));
 sg13g2_tiehi \am_sdr0.cic0.integ2[17]$_SDFF_PN0__664  (.L_HI(net664));
 sg13g2_tiehi \am_sdr0.cic0.integ2[18]$_SDFF_PN0__665  (.L_HI(net665));
 sg13g2_tiehi \am_sdr0.cic0.integ2[19]$_SDFF_PN0__666  (.L_HI(net666));
 sg13g2_tiehi \am_sdr0.cic0.integ2[1]$_SDFF_PN0__667  (.L_HI(net667));
 sg13g2_tiehi \am_sdr0.cic0.integ2[20]$_SDFF_PN0__668  (.L_HI(net668));
 sg13g2_tiehi \am_sdr0.cic0.integ2[21]$_SDFF_PN0__669  (.L_HI(net669));
 sg13g2_tiehi \am_sdr0.cic0.integ2[22]$_SDFF_PN0__670  (.L_HI(net670));
 sg13g2_tiehi \am_sdr0.cic0.integ2[2]$_SDFF_PN0__671  (.L_HI(net671));
 sg13g2_tiehi \am_sdr0.cic0.integ2[3]$_SDFF_PN0__672  (.L_HI(net672));
 sg13g2_tiehi \am_sdr0.cic0.integ2[4]$_SDFF_PN0__673  (.L_HI(net673));
 sg13g2_tiehi \am_sdr0.cic0.integ2[5]$_SDFF_PN0__674  (.L_HI(net674));
 sg13g2_tiehi \am_sdr0.cic0.integ2[6]$_SDFF_PN0__675  (.L_HI(net675));
 sg13g2_tiehi \am_sdr0.cic0.integ2[7]$_SDFF_PN0__676  (.L_HI(net676));
 sg13g2_tiehi \am_sdr0.cic0.integ2[8]$_SDFF_PN0__677  (.L_HI(net677));
 sg13g2_tiehi \am_sdr0.cic0.integ2[9]$_SDFF_PN0__678  (.L_HI(net678));
 sg13g2_tiehi \am_sdr0.cic0.integ3[0]$_SDFF_PN0__679  (.L_HI(net679));
 sg13g2_tiehi \am_sdr0.cic0.integ3[10]$_SDFF_PN0__680  (.L_HI(net680));
 sg13g2_tiehi \am_sdr0.cic0.integ3[11]$_SDFF_PN0__681  (.L_HI(net681));
 sg13g2_tiehi \am_sdr0.cic0.integ3[12]$_SDFF_PN0__682  (.L_HI(net682));
 sg13g2_tiehi \am_sdr0.cic0.integ3[13]$_SDFF_PN0__683  (.L_HI(net683));
 sg13g2_tiehi \am_sdr0.cic0.integ3[14]$_SDFF_PN0__684  (.L_HI(net684));
 sg13g2_tiehi \am_sdr0.cic0.integ3[15]$_SDFF_PN0__685  (.L_HI(net685));
 sg13g2_tiehi \am_sdr0.cic0.integ3[16]$_SDFF_PN0__686  (.L_HI(net686));
 sg13g2_tiehi \am_sdr0.cic0.integ3[17]$_SDFF_PN0__687  (.L_HI(net687));
 sg13g2_tiehi \am_sdr0.cic0.integ3[18]$_SDFF_PN0__688  (.L_HI(net688));
 sg13g2_tiehi \am_sdr0.cic0.integ3[19]$_SDFF_PN0__689  (.L_HI(net689));
 sg13g2_tiehi \am_sdr0.cic0.integ3[1]$_SDFF_PN0__690  (.L_HI(net690));
 sg13g2_tiehi \am_sdr0.cic0.integ3[2]$_SDFF_PN0__691  (.L_HI(net691));
 sg13g2_tiehi \am_sdr0.cic0.integ3[3]$_SDFF_PN0__692  (.L_HI(net692));
 sg13g2_tiehi \am_sdr0.cic0.integ3[4]$_SDFF_PN0__693  (.L_HI(net693));
 sg13g2_tiehi \am_sdr0.cic0.integ3[5]$_SDFF_PN0__694  (.L_HI(net694));
 sg13g2_tiehi \am_sdr0.cic0.integ3[6]$_SDFF_PN0__695  (.L_HI(net695));
 sg13g2_tiehi \am_sdr0.cic0.integ3[7]$_SDFF_PN0__696  (.L_HI(net696));
 sg13g2_tiehi \am_sdr0.cic0.integ3[8]$_SDFF_PN0__697  (.L_HI(net697));
 sg13g2_tiehi \am_sdr0.cic0.integ3[9]$_SDFF_PN0__698  (.L_HI(net698));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[0]$_DFFE_PP__699  (.L_HI(net699));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[10]$_DFFE_PP__700  (.L_HI(net700));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[11]$_DFFE_PP__701  (.L_HI(net701));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[12]$_DFFE_PP__702  (.L_HI(net702));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[13]$_DFFE_PP__703  (.L_HI(net703));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[14]$_DFFE_PP__704  (.L_HI(net704));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[15]$_DFFE_PP__705  (.L_HI(net705));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[16]$_DFFE_PP__706  (.L_HI(net706));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[17]$_DFFE_PP__707  (.L_HI(net707));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[18]$_DFFE_PP__708  (.L_HI(net708));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[19]$_DFFE_PP__709  (.L_HI(net709));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[1]$_DFFE_PP__710  (.L_HI(net710));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[2]$_DFFE_PP__711  (.L_HI(net711));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[3]$_DFFE_PP__712  (.L_HI(net712));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[4]$_DFFE_PP__713  (.L_HI(net713));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[5]$_DFFE_PP__714  (.L_HI(net714));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[6]$_DFFE_PP__715  (.L_HI(net715));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[7]$_DFFE_PP__716  (.L_HI(net716));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[8]$_DFFE_PP__717  (.L_HI(net717));
 sg13g2_tiehi \am_sdr0.cic0.integ_sample[9]$_DFFE_PP__718  (.L_HI(net718));
 sg13g2_tiehi \am_sdr0.cic0.out_tick$_SDFF_PN0__719  (.L_HI(net719));
 sg13g2_tiehi \am_sdr0.cic0.sample$_SDFF_PN0__720  (.L_HI(net720));
 sg13g2_tiehi \am_sdr0.cic0.x_out[10]$_SDFFE_PN0P__721  (.L_HI(net721));
 sg13g2_tiehi \am_sdr0.cic0.x_out[11]$_SDFFE_PN0P__722  (.L_HI(net722));
 sg13g2_tiehi \am_sdr0.cic0.x_out[12]$_SDFFE_PN0P__723  (.L_HI(net723));
 sg13g2_tiehi \am_sdr0.cic0.x_out[13]$_SDFFE_PN0P__724  (.L_HI(net724));
 sg13g2_tiehi \am_sdr0.cic0.x_out[14]$_SDFFE_PN0P__725  (.L_HI(net725));
 sg13g2_tiehi \am_sdr0.cic0.x_out[15]$_SDFFE_PN0P__726  (.L_HI(net726));
 sg13g2_tiehi \am_sdr0.cic0.x_out[8]$_SDFFE_PN0P__727  (.L_HI(net727));
 sg13g2_tiehi \am_sdr0.cic0.x_out[9]$_SDFFE_PN0P__728  (.L_HI(net728));
 sg13g2_tiehi \am_sdr0.cic1.comb1[0]$_SDFFE_PN0P__729  (.L_HI(net729));
 sg13g2_tiehi \am_sdr0.cic1.comb1[10]$_SDFFE_PN0P__730  (.L_HI(net730));
 sg13g2_tiehi \am_sdr0.cic1.comb1[11]$_SDFFE_PN0P__731  (.L_HI(net731));
 sg13g2_tiehi \am_sdr0.cic1.comb1[12]$_SDFFE_PN0P__732  (.L_HI(net732));
 sg13g2_tiehi \am_sdr0.cic1.comb1[13]$_SDFFE_PN0P__733  (.L_HI(net733));
 sg13g2_tiehi \am_sdr0.cic1.comb1[14]$_SDFFE_PN0P__734  (.L_HI(net734));
 sg13g2_tiehi \am_sdr0.cic1.comb1[15]$_SDFFE_PN0P__735  (.L_HI(net735));
 sg13g2_tiehi \am_sdr0.cic1.comb1[16]$_SDFFE_PN0P__736  (.L_HI(net736));
 sg13g2_tiehi \am_sdr0.cic1.comb1[17]$_SDFFE_PN0P__737  (.L_HI(net737));
 sg13g2_tiehi \am_sdr0.cic1.comb1[18]$_SDFFE_PN0P__738  (.L_HI(net738));
 sg13g2_tiehi \am_sdr0.cic1.comb1[19]$_SDFFE_PN0P__739  (.L_HI(net739));
 sg13g2_tiehi \am_sdr0.cic1.comb1[1]$_SDFFE_PN0P__740  (.L_HI(net740));
 sg13g2_tiehi \am_sdr0.cic1.comb1[2]$_SDFFE_PN0P__741  (.L_HI(net741));
 sg13g2_tiehi \am_sdr0.cic1.comb1[3]$_SDFFE_PN0P__742  (.L_HI(net742));
 sg13g2_tiehi \am_sdr0.cic1.comb1[4]$_SDFFE_PN0P__743  (.L_HI(net743));
 sg13g2_tiehi \am_sdr0.cic1.comb1[5]$_SDFFE_PN0P__744  (.L_HI(net744));
 sg13g2_tiehi \am_sdr0.cic1.comb1[6]$_SDFFE_PN0P__745  (.L_HI(net745));
 sg13g2_tiehi \am_sdr0.cic1.comb1[7]$_SDFFE_PN0P__746  (.L_HI(net746));
 sg13g2_tiehi \am_sdr0.cic1.comb1[8]$_SDFFE_PN0P__747  (.L_HI(net747));
 sg13g2_tiehi \am_sdr0.cic1.comb1[9]$_SDFFE_PN0P__748  (.L_HI(net748));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[0]$_SDFFE_PN0P__749  (.L_HI(net749));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[10]$_SDFFE_PN0P__750  (.L_HI(net750));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[11]$_SDFFE_PN0P__751  (.L_HI(net751));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[12]$_SDFFE_PN0P__752  (.L_HI(net752));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[13]$_SDFFE_PN0P__753  (.L_HI(net753));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[14]$_SDFFE_PN0P__754  (.L_HI(net754));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[15]$_SDFFE_PN0P__755  (.L_HI(net755));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[16]$_SDFFE_PN0P__756  (.L_HI(net756));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[17]$_SDFFE_PN0P__757  (.L_HI(net757));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[18]$_SDFFE_PN0P__758  (.L_HI(net758));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[19]$_SDFFE_PN0P__759  (.L_HI(net759));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[1]$_SDFFE_PN0P__760  (.L_HI(net760));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[2]$_SDFFE_PN0P__761  (.L_HI(net761));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[3]$_SDFFE_PN0P__762  (.L_HI(net762));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[4]$_SDFFE_PN0P__763  (.L_HI(net763));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[5]$_SDFFE_PN0P__764  (.L_HI(net764));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[6]$_SDFFE_PN0P__765  (.L_HI(net765));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[7]$_SDFFE_PN0P__766  (.L_HI(net766));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[8]$_SDFFE_PN0P__767  (.L_HI(net767));
 sg13g2_tiehi \am_sdr0.cic1.comb1_in_del[9]$_SDFFE_PN0P__768  (.L_HI(net768));
 sg13g2_tiehi \am_sdr0.cic1.comb2[0]$_SDFFE_PN0P__769  (.L_HI(net769));
 sg13g2_tiehi \am_sdr0.cic1.comb2[10]$_SDFFE_PN0P__770  (.L_HI(net770));
 sg13g2_tiehi \am_sdr0.cic1.comb2[11]$_SDFFE_PN0P__771  (.L_HI(net771));
 sg13g2_tiehi \am_sdr0.cic1.comb2[12]$_SDFFE_PN0P__772  (.L_HI(net772));
 sg13g2_tiehi \am_sdr0.cic1.comb2[13]$_SDFFE_PN0P__773  (.L_HI(net773));
 sg13g2_tiehi \am_sdr0.cic1.comb2[14]$_SDFFE_PN0P__774  (.L_HI(net774));
 sg13g2_tiehi \am_sdr0.cic1.comb2[15]$_SDFFE_PN0P__775  (.L_HI(net775));
 sg13g2_tiehi \am_sdr0.cic1.comb2[16]$_SDFFE_PN0P__776  (.L_HI(net776));
 sg13g2_tiehi \am_sdr0.cic1.comb2[17]$_SDFFE_PN0P__777  (.L_HI(net777));
 sg13g2_tiehi \am_sdr0.cic1.comb2[18]$_SDFFE_PN0P__778  (.L_HI(net778));
 sg13g2_tiehi \am_sdr0.cic1.comb2[19]$_SDFFE_PN0P__779  (.L_HI(net779));
 sg13g2_tiehi \am_sdr0.cic1.comb2[1]$_SDFFE_PN0P__780  (.L_HI(net780));
 sg13g2_tiehi \am_sdr0.cic1.comb2[2]$_SDFFE_PN0P__781  (.L_HI(net781));
 sg13g2_tiehi \am_sdr0.cic1.comb2[3]$_SDFFE_PN0P__782  (.L_HI(net782));
 sg13g2_tiehi \am_sdr0.cic1.comb2[4]$_SDFFE_PN0P__783  (.L_HI(net783));
 sg13g2_tiehi \am_sdr0.cic1.comb2[5]$_SDFFE_PN0P__784  (.L_HI(net784));
 sg13g2_tiehi \am_sdr0.cic1.comb2[6]$_SDFFE_PN0P__785  (.L_HI(net785));
 sg13g2_tiehi \am_sdr0.cic1.comb2[7]$_SDFFE_PN0P__786  (.L_HI(net786));
 sg13g2_tiehi \am_sdr0.cic1.comb2[8]$_SDFFE_PN0P__787  (.L_HI(net787));
 sg13g2_tiehi \am_sdr0.cic1.comb2[9]$_SDFFE_PN0P__788  (.L_HI(net788));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[0]$_SDFFE_PN0P__789  (.L_HI(net789));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[10]$_SDFFE_PN0P__790  (.L_HI(net790));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[11]$_SDFFE_PN0P__791  (.L_HI(net791));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[12]$_SDFFE_PN0P__792  (.L_HI(net792));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[13]$_SDFFE_PN0P__793  (.L_HI(net793));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[14]$_SDFFE_PN0P__794  (.L_HI(net794));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[15]$_SDFFE_PN0P__795  (.L_HI(net795));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[16]$_SDFFE_PN0P__796  (.L_HI(net796));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[17]$_SDFFE_PN0P__797  (.L_HI(net797));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[18]$_SDFFE_PN0P__798  (.L_HI(net798));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[19]$_SDFFE_PN0P__799  (.L_HI(net799));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[1]$_SDFFE_PN0P__800  (.L_HI(net800));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[2]$_SDFFE_PN0P__801  (.L_HI(net801));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[3]$_SDFFE_PN0P__802  (.L_HI(net802));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[4]$_SDFFE_PN0P__803  (.L_HI(net803));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[5]$_SDFFE_PN0P__804  (.L_HI(net804));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[6]$_SDFFE_PN0P__805  (.L_HI(net805));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[7]$_SDFFE_PN0P__806  (.L_HI(net806));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[8]$_SDFFE_PN0P__807  (.L_HI(net807));
 sg13g2_tiehi \am_sdr0.cic1.comb2_in_del[9]$_SDFFE_PN0P__808  (.L_HI(net808));
 sg13g2_tiehi \am_sdr0.cic1.comb3[12]$_SDFFE_PN0P__809  (.L_HI(net809));
 sg13g2_tiehi \am_sdr0.cic1.comb3[13]$_SDFFE_PN0P__810  (.L_HI(net810));
 sg13g2_tiehi \am_sdr0.cic1.comb3[14]$_SDFFE_PN0P__811  (.L_HI(net811));
 sg13g2_tiehi \am_sdr0.cic1.comb3[15]$_SDFFE_PN0P__812  (.L_HI(net812));
 sg13g2_tiehi \am_sdr0.cic1.comb3[16]$_SDFFE_PN0P__813  (.L_HI(net813));
 sg13g2_tiehi \am_sdr0.cic1.comb3[17]$_SDFFE_PN0P__814  (.L_HI(net814));
 sg13g2_tiehi \am_sdr0.cic1.comb3[18]$_SDFFE_PN0P__815  (.L_HI(net815));
 sg13g2_tiehi \am_sdr0.cic1.comb3[19]$_SDFFE_PN0P__816  (.L_HI(net816));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[0]$_SDFFE_PN0P__817  (.L_HI(net817));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[10]$_SDFFE_PN0P__818  (.L_HI(net818));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[11]$_SDFFE_PN0P__819  (.L_HI(net819));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[12]$_SDFFE_PN0P__820  (.L_HI(net820));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[13]$_SDFFE_PN0P__821  (.L_HI(net821));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[14]$_SDFFE_PN0P__822  (.L_HI(net822));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[15]$_SDFFE_PN0P__823  (.L_HI(net823));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[16]$_SDFFE_PN0P__824  (.L_HI(net824));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[17]$_SDFFE_PN0P__825  (.L_HI(net825));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[18]$_SDFFE_PN0P__826  (.L_HI(net826));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[19]$_SDFFE_PN0P__827  (.L_HI(net827));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[1]$_SDFFE_PN0P__828  (.L_HI(net828));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[2]$_SDFFE_PN0P__829  (.L_HI(net829));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[3]$_SDFFE_PN0P__830  (.L_HI(net830));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[4]$_SDFFE_PN0P__831  (.L_HI(net831));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[5]$_SDFFE_PN0P__832  (.L_HI(net832));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[6]$_SDFFE_PN0P__833  (.L_HI(net833));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[7]$_SDFFE_PN0P__834  (.L_HI(net834));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[8]$_SDFFE_PN0P__835  (.L_HI(net835));
 sg13g2_tiehi \am_sdr0.cic1.comb3_in_del[9]$_SDFFE_PN0P__836  (.L_HI(net836));
 sg13g2_tiehi \am_sdr0.cic1.count[0]$_SDFF_PP0__837  (.L_HI(net837));
 sg13g2_tiehi \am_sdr0.cic1.count[1]$_SDFF_PP0__838  (.L_HI(net838));
 sg13g2_tiehi \am_sdr0.cic1.count[2]$_SDFF_PP0__839  (.L_HI(net839));
 sg13g2_tiehi \am_sdr0.cic1.count[3]$_SDFF_PP0__840  (.L_HI(net840));
 sg13g2_tiehi \am_sdr0.cic1.count[4]$_SDFF_PP0__841  (.L_HI(net841));
 sg13g2_tiehi \am_sdr0.cic1.count[5]$_SDFF_PP0__842  (.L_HI(net842));
 sg13g2_tiehi \am_sdr0.cic1.count[6]$_SDFF_PP0__843  (.L_HI(net843));
 sg13g2_tiehi \am_sdr0.cic1.count[7]$_SDFF_PP0__844  (.L_HI(net844));
 sg13g2_tiehi \am_sdr0.cic1.integ1[0]$_SDFF_PN0__845  (.L_HI(net845));
 sg13g2_tiehi \am_sdr0.cic1.integ1[10]$_SDFF_PN0__846  (.L_HI(net846));
 sg13g2_tiehi \am_sdr0.cic1.integ1[11]$_SDFF_PN0__847  (.L_HI(net847));
 sg13g2_tiehi \am_sdr0.cic1.integ1[12]$_SDFF_PN0__848  (.L_HI(net848));
 sg13g2_tiehi \am_sdr0.cic1.integ1[13]$_SDFF_PN0__849  (.L_HI(net849));
 sg13g2_tiehi \am_sdr0.cic1.integ1[14]$_SDFF_PN0__850  (.L_HI(net850));
 sg13g2_tiehi \am_sdr0.cic1.integ1[15]$_SDFF_PN0__851  (.L_HI(net851));
 sg13g2_tiehi \am_sdr0.cic1.integ1[16]$_SDFF_PN0__852  (.L_HI(net852));
 sg13g2_tiehi \am_sdr0.cic1.integ1[17]$_SDFF_PN0__853  (.L_HI(net853));
 sg13g2_tiehi \am_sdr0.cic1.integ1[18]$_SDFF_PN0__854  (.L_HI(net854));
 sg13g2_tiehi \am_sdr0.cic1.integ1[19]$_SDFF_PN0__855  (.L_HI(net855));
 sg13g2_tiehi \am_sdr0.cic1.integ1[1]$_SDFF_PN0__856  (.L_HI(net856));
 sg13g2_tiehi \am_sdr0.cic1.integ1[20]$_SDFF_PN0__857  (.L_HI(net857));
 sg13g2_tiehi \am_sdr0.cic1.integ1[21]$_SDFF_PN0__858  (.L_HI(net858));
 sg13g2_tiehi \am_sdr0.cic1.integ1[22]$_SDFF_PN0__859  (.L_HI(net859));
 sg13g2_tiehi \am_sdr0.cic1.integ1[23]$_SDFF_PN0__860  (.L_HI(net860));
 sg13g2_tiehi \am_sdr0.cic1.integ1[24]$_SDFF_PN0__861  (.L_HI(net861));
 sg13g2_tiehi \am_sdr0.cic1.integ1[25]$_SDFF_PN0__862  (.L_HI(net862));
 sg13g2_tiehi \am_sdr0.cic1.integ1[2]$_SDFF_PN0__863  (.L_HI(net863));
 sg13g2_tiehi \am_sdr0.cic1.integ1[3]$_SDFF_PN0__864  (.L_HI(net864));
 sg13g2_tiehi \am_sdr0.cic1.integ1[4]$_SDFF_PN0__865  (.L_HI(net865));
 sg13g2_tiehi \am_sdr0.cic1.integ1[5]$_SDFF_PN0__866  (.L_HI(net866));
 sg13g2_tiehi \am_sdr0.cic1.integ1[6]$_SDFF_PN0__867  (.L_HI(net867));
 sg13g2_tiehi \am_sdr0.cic1.integ1[7]$_SDFF_PN0__868  (.L_HI(net868));
 sg13g2_tiehi \am_sdr0.cic1.integ1[8]$_SDFF_PN0__869  (.L_HI(net869));
 sg13g2_tiehi \am_sdr0.cic1.integ1[9]$_SDFF_PN0__870  (.L_HI(net870));
 sg13g2_tiehi \am_sdr0.cic1.integ2[0]$_SDFF_PN0__871  (.L_HI(net871));
 sg13g2_tiehi \am_sdr0.cic1.integ2[10]$_SDFF_PN0__872  (.L_HI(net872));
 sg13g2_tiehi \am_sdr0.cic1.integ2[11]$_SDFF_PN0__873  (.L_HI(net873));
 sg13g2_tiehi \am_sdr0.cic1.integ2[12]$_SDFF_PN0__874  (.L_HI(net874));
 sg13g2_tiehi \am_sdr0.cic1.integ2[13]$_SDFF_PN0__875  (.L_HI(net875));
 sg13g2_tiehi \am_sdr0.cic1.integ2[14]$_SDFF_PN0__876  (.L_HI(net876));
 sg13g2_tiehi \am_sdr0.cic1.integ2[15]$_SDFF_PN0__877  (.L_HI(net877));
 sg13g2_tiehi \am_sdr0.cic1.integ2[16]$_SDFF_PN0__878  (.L_HI(net878));
 sg13g2_tiehi \am_sdr0.cic1.integ2[17]$_SDFF_PN0__879  (.L_HI(net879));
 sg13g2_tiehi \am_sdr0.cic1.integ2[18]$_SDFF_PN0__880  (.L_HI(net880));
 sg13g2_tiehi \am_sdr0.cic1.integ2[19]$_SDFF_PN0__881  (.L_HI(net881));
 sg13g2_tiehi \am_sdr0.cic1.integ2[1]$_SDFF_PN0__882  (.L_HI(net882));
 sg13g2_tiehi \am_sdr0.cic1.integ2[20]$_SDFF_PN0__883  (.L_HI(net883));
 sg13g2_tiehi \am_sdr0.cic1.integ2[21]$_SDFF_PN0__884  (.L_HI(net884));
 sg13g2_tiehi \am_sdr0.cic1.integ2[22]$_SDFF_PN0__885  (.L_HI(net885));
 sg13g2_tiehi \am_sdr0.cic1.integ2[2]$_SDFF_PN0__886  (.L_HI(net886));
 sg13g2_tiehi \am_sdr0.cic1.integ2[3]$_SDFF_PN0__887  (.L_HI(net887));
 sg13g2_tiehi \am_sdr0.cic1.integ2[4]$_SDFF_PN0__888  (.L_HI(net888));
 sg13g2_tiehi \am_sdr0.cic1.integ2[5]$_SDFF_PN0__889  (.L_HI(net889));
 sg13g2_tiehi \am_sdr0.cic1.integ2[6]$_SDFF_PN0__890  (.L_HI(net890));
 sg13g2_tiehi \am_sdr0.cic1.integ2[7]$_SDFF_PN0__891  (.L_HI(net891));
 sg13g2_tiehi \am_sdr0.cic1.integ2[8]$_SDFF_PN0__892  (.L_HI(net892));
 sg13g2_tiehi \am_sdr0.cic1.integ2[9]$_SDFF_PN0__893  (.L_HI(net893));
 sg13g2_tiehi \am_sdr0.cic1.integ3[0]$_SDFF_PN0__894  (.L_HI(net894));
 sg13g2_tiehi \am_sdr0.cic1.integ3[10]$_SDFF_PN0__895  (.L_HI(net895));
 sg13g2_tiehi \am_sdr0.cic1.integ3[11]$_SDFF_PN0__896  (.L_HI(net896));
 sg13g2_tiehi \am_sdr0.cic1.integ3[12]$_SDFF_PN0__897  (.L_HI(net897));
 sg13g2_tiehi \am_sdr0.cic1.integ3[13]$_SDFF_PN0__898  (.L_HI(net898));
 sg13g2_tiehi \am_sdr0.cic1.integ3[14]$_SDFF_PN0__899  (.L_HI(net899));
 sg13g2_tiehi \am_sdr0.cic1.integ3[15]$_SDFF_PN0__900  (.L_HI(net900));
 sg13g2_tiehi \am_sdr0.cic1.integ3[16]$_SDFF_PN0__901  (.L_HI(net901));
 sg13g2_tiehi \am_sdr0.cic1.integ3[17]$_SDFF_PN0__902  (.L_HI(net902));
 sg13g2_tiehi \am_sdr0.cic1.integ3[18]$_SDFF_PN0__903  (.L_HI(net903));
 sg13g2_tiehi \am_sdr0.cic1.integ3[19]$_SDFF_PN0__904  (.L_HI(net904));
 sg13g2_tiehi \am_sdr0.cic1.integ3[1]$_SDFF_PN0__905  (.L_HI(net905));
 sg13g2_tiehi \am_sdr0.cic1.integ3[2]$_SDFF_PN0__906  (.L_HI(net906));
 sg13g2_tiehi \am_sdr0.cic1.integ3[3]$_SDFF_PN0__907  (.L_HI(net907));
 sg13g2_tiehi \am_sdr0.cic1.integ3[4]$_SDFF_PN0__908  (.L_HI(net908));
 sg13g2_tiehi \am_sdr0.cic1.integ3[5]$_SDFF_PN0__909  (.L_HI(net909));
 sg13g2_tiehi \am_sdr0.cic1.integ3[6]$_SDFF_PN0__910  (.L_HI(net910));
 sg13g2_tiehi \am_sdr0.cic1.integ3[7]$_SDFF_PN0__911  (.L_HI(net911));
 sg13g2_tiehi \am_sdr0.cic1.integ3[8]$_SDFF_PN0__912  (.L_HI(net912));
 sg13g2_tiehi \am_sdr0.cic1.integ3[9]$_SDFF_PN0__913  (.L_HI(net913));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[0]$_DFFE_PP__914  (.L_HI(net914));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[10]$_DFFE_PP__915  (.L_HI(net915));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[11]$_DFFE_PP__916  (.L_HI(net916));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[12]$_DFFE_PP__917  (.L_HI(net917));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[13]$_DFFE_PP__918  (.L_HI(net918));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[14]$_DFFE_PP__919  (.L_HI(net919));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[15]$_DFFE_PP__920  (.L_HI(net920));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[16]$_DFFE_PP__921  (.L_HI(net921));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[17]$_DFFE_PP__922  (.L_HI(net922));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[18]$_DFFE_PP__923  (.L_HI(net923));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[19]$_DFFE_PP__924  (.L_HI(net924));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[1]$_DFFE_PP__925  (.L_HI(net925));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[2]$_DFFE_PP__926  (.L_HI(net926));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[3]$_DFFE_PP__927  (.L_HI(net927));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[4]$_DFFE_PP__928  (.L_HI(net928));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[5]$_DFFE_PP__929  (.L_HI(net929));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[6]$_DFFE_PP__930  (.L_HI(net930));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[7]$_DFFE_PP__931  (.L_HI(net931));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[8]$_DFFE_PP__932  (.L_HI(net932));
 sg13g2_tiehi \am_sdr0.cic1.integ_sample[9]$_DFFE_PP__933  (.L_HI(net933));
 sg13g2_tiehi \am_sdr0.cic1.out_tick$_SDFF_PN0__934  (.L_HI(net934));
 sg13g2_tiehi \am_sdr0.cic1.sample$_SDFF_PN0__935  (.L_HI(net935));
 sg13g2_tiehi \am_sdr0.cic1.x_out[10]$_SDFFE_PN0P__936  (.L_HI(net936));
 sg13g2_tiehi \am_sdr0.cic1.x_out[11]$_SDFFE_PN0P__937  (.L_HI(net937));
 sg13g2_tiehi \am_sdr0.cic1.x_out[12]$_SDFFE_PN0P__938  (.L_HI(net938));
 sg13g2_tiehi \am_sdr0.cic1.x_out[13]$_SDFFE_PN0P__939  (.L_HI(net939));
 sg13g2_tiehi \am_sdr0.cic1.x_out[14]$_SDFFE_PN0P__940  (.L_HI(net940));
 sg13g2_tiehi \am_sdr0.cic1.x_out[15]$_SDFFE_PN0P__941  (.L_HI(net941));
 sg13g2_tiehi \am_sdr0.cic1.x_out[8]$_SDFFE_PN0P__942  (.L_HI(net942));
 sg13g2_tiehi \am_sdr0.cic1.x_out[9]$_SDFFE_PN0P__943  (.L_HI(net943));
 sg13g2_tiehi \am_sdr0.cic2.comb1[0]$_SDFFE_PN0P__944  (.L_HI(net944));
 sg13g2_tiehi \am_sdr0.cic2.comb1[10]$_SDFFE_PN0P__945  (.L_HI(net945));
 sg13g2_tiehi \am_sdr0.cic2.comb1[11]$_SDFFE_PN0P__946  (.L_HI(net946));
 sg13g2_tiehi \am_sdr0.cic2.comb1[12]$_SDFFE_PN0P__947  (.L_HI(net947));
 sg13g2_tiehi \am_sdr0.cic2.comb1[13]$_SDFFE_PN0P__948  (.L_HI(net948));
 sg13g2_tiehi \am_sdr0.cic2.comb1[14]$_SDFFE_PN0P__949  (.L_HI(net949));
 sg13g2_tiehi \am_sdr0.cic2.comb1[15]$_SDFFE_PN0P__950  (.L_HI(net950));
 sg13g2_tiehi \am_sdr0.cic2.comb1[16]$_SDFFE_PN0P__951  (.L_HI(net951));
 sg13g2_tiehi \am_sdr0.cic2.comb1[17]$_SDFFE_PN0P__952  (.L_HI(net952));
 sg13g2_tiehi \am_sdr0.cic2.comb1[18]$_SDFFE_PN0P__953  (.L_HI(net953));
 sg13g2_tiehi \am_sdr0.cic2.comb1[19]$_SDFFE_PN0P__954  (.L_HI(net954));
 sg13g2_tiehi \am_sdr0.cic2.comb1[1]$_SDFFE_PN0P__955  (.L_HI(net955));
 sg13g2_tiehi \am_sdr0.cic2.comb1[2]$_SDFFE_PN0P__956  (.L_HI(net956));
 sg13g2_tiehi \am_sdr0.cic2.comb1[3]$_SDFFE_PN0P__957  (.L_HI(net957));
 sg13g2_tiehi \am_sdr0.cic2.comb1[4]$_SDFFE_PN0P__958  (.L_HI(net958));
 sg13g2_tiehi \am_sdr0.cic2.comb1[5]$_SDFFE_PN0P__959  (.L_HI(net959));
 sg13g2_tiehi \am_sdr0.cic2.comb1[6]$_SDFFE_PN0P__960  (.L_HI(net960));
 sg13g2_tiehi \am_sdr0.cic2.comb1[7]$_SDFFE_PN0P__961  (.L_HI(net961));
 sg13g2_tiehi \am_sdr0.cic2.comb1[8]$_SDFFE_PN0P__962  (.L_HI(net962));
 sg13g2_tiehi \am_sdr0.cic2.comb1[9]$_SDFFE_PN0P__963  (.L_HI(net963));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[0]$_SDFFE_PN0P__964  (.L_HI(net964));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[10]$_SDFFE_PN0P__965  (.L_HI(net965));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[11]$_SDFFE_PN0P__966  (.L_HI(net966));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[12]$_SDFFE_PN0P__967  (.L_HI(net967));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[13]$_SDFFE_PN0P__968  (.L_HI(net968));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[14]$_SDFFE_PN0P__969  (.L_HI(net969));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[15]$_SDFFE_PN0P__970  (.L_HI(net970));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[16]$_SDFFE_PN0P__971  (.L_HI(net971));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[17]$_SDFFE_PN0P__972  (.L_HI(net972));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[18]$_SDFFE_PN0P__973  (.L_HI(net973));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[19]$_SDFFE_PN0P__974  (.L_HI(net974));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[1]$_SDFFE_PN0P__975  (.L_HI(net975));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[2]$_SDFFE_PN0P__976  (.L_HI(net976));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[3]$_SDFFE_PN0P__977  (.L_HI(net977));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[4]$_SDFFE_PN0P__978  (.L_HI(net978));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[5]$_SDFFE_PN0P__979  (.L_HI(net979));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[6]$_SDFFE_PN0P__980  (.L_HI(net980));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[7]$_SDFFE_PN0P__981  (.L_HI(net981));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[8]$_SDFFE_PN0P__982  (.L_HI(net982));
 sg13g2_tiehi \am_sdr0.cic2.comb1_in_del[9]$_SDFFE_PN0P__983  (.L_HI(net983));
 sg13g2_tiehi \am_sdr0.cic2.comb2[0]$_SDFFE_PN0P__984  (.L_HI(net984));
 sg13g2_tiehi \am_sdr0.cic2.comb2[10]$_SDFFE_PN0P__985  (.L_HI(net985));
 sg13g2_tiehi \am_sdr0.cic2.comb2[11]$_SDFFE_PN0P__986  (.L_HI(net986));
 sg13g2_tiehi \am_sdr0.cic2.comb2[12]$_SDFFE_PN0P__987  (.L_HI(net987));
 sg13g2_tiehi \am_sdr0.cic2.comb2[13]$_SDFFE_PN0P__988  (.L_HI(net988));
 sg13g2_tiehi \am_sdr0.cic2.comb2[14]$_SDFFE_PN0P__989  (.L_HI(net989));
 sg13g2_tiehi \am_sdr0.cic2.comb2[15]$_SDFFE_PN0P__990  (.L_HI(net990));
 sg13g2_tiehi \am_sdr0.cic2.comb2[16]$_SDFFE_PN0P__991  (.L_HI(net991));
 sg13g2_tiehi \am_sdr0.cic2.comb2[17]$_SDFFE_PN0P__992  (.L_HI(net992));
 sg13g2_tiehi \am_sdr0.cic2.comb2[18]$_SDFFE_PN0P__993  (.L_HI(net993));
 sg13g2_tiehi \am_sdr0.cic2.comb2[19]$_SDFFE_PN0P__994  (.L_HI(net994));
 sg13g2_tiehi \am_sdr0.cic2.comb2[1]$_SDFFE_PN0P__995  (.L_HI(net995));
 sg13g2_tiehi \am_sdr0.cic2.comb2[2]$_SDFFE_PN0P__996  (.L_HI(net996));
 sg13g2_tiehi \am_sdr0.cic2.comb2[3]$_SDFFE_PN0P__997  (.L_HI(net997));
 sg13g2_tiehi \am_sdr0.cic2.comb2[4]$_SDFFE_PN0P__998  (.L_HI(net998));
 sg13g2_tiehi \am_sdr0.cic2.comb2[5]$_SDFFE_PN0P__999  (.L_HI(net999));
 sg13g2_tiehi \am_sdr0.cic2.comb2[6]$_SDFFE_PN0P__1000  (.L_HI(net1000));
 sg13g2_tiehi \am_sdr0.cic2.comb2[7]$_SDFFE_PN0P__1001  (.L_HI(net1001));
 sg13g2_tiehi \am_sdr0.cic2.comb2[8]$_SDFFE_PN0P__1002  (.L_HI(net1002));
 sg13g2_tiehi \am_sdr0.cic2.comb2[9]$_SDFFE_PN0P__1003  (.L_HI(net1003));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[0]$_SDFFE_PN0P__1004  (.L_HI(net1004));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[10]$_SDFFE_PN0P__1005  (.L_HI(net1005));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[11]$_SDFFE_PN0P__1006  (.L_HI(net1006));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[12]$_SDFFE_PN0P__1007  (.L_HI(net1007));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[13]$_SDFFE_PN0P__1008  (.L_HI(net1008));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[14]$_SDFFE_PN0P__1009  (.L_HI(net1009));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[15]$_SDFFE_PN0P__1010  (.L_HI(net1010));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[16]$_SDFFE_PN0P__1011  (.L_HI(net1011));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[17]$_SDFFE_PN0P__1012  (.L_HI(net1012));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[18]$_SDFFE_PN0P__1013  (.L_HI(net1013));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[19]$_SDFFE_PN0P__1014  (.L_HI(net1014));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[1]$_SDFFE_PN0P__1015  (.L_HI(net1015));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[2]$_SDFFE_PN0P__1016  (.L_HI(net1016));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[3]$_SDFFE_PN0P__1017  (.L_HI(net1017));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[4]$_SDFFE_PN0P__1018  (.L_HI(net1018));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[5]$_SDFFE_PN0P__1019  (.L_HI(net1019));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[6]$_SDFFE_PN0P__1020  (.L_HI(net1020));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[7]$_SDFFE_PN0P__1021  (.L_HI(net1021));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[8]$_SDFFE_PN0P__1022  (.L_HI(net1022));
 sg13g2_tiehi \am_sdr0.cic2.comb2_in_del[9]$_SDFFE_PN0P__1023  (.L_HI(net1023));
 sg13g2_tiehi \am_sdr0.cic2.comb3[12]$_SDFFE_PN0P__1024  (.L_HI(net1024));
 sg13g2_tiehi \am_sdr0.cic2.comb3[13]$_SDFFE_PN0P__1025  (.L_HI(net1025));
 sg13g2_tiehi \am_sdr0.cic2.comb3[14]$_SDFFE_PN0P__1026  (.L_HI(net1026));
 sg13g2_tiehi \am_sdr0.cic2.comb3[15]$_SDFFE_PN0P__1027  (.L_HI(net1027));
 sg13g2_tiehi \am_sdr0.cic2.comb3[16]$_SDFFE_PN0P__1028  (.L_HI(net1028));
 sg13g2_tiehi \am_sdr0.cic2.comb3[17]$_SDFFE_PN0P__1029  (.L_HI(net1029));
 sg13g2_tiehi \am_sdr0.cic2.comb3[18]$_SDFFE_PN0P__1030  (.L_HI(net1030));
 sg13g2_tiehi \am_sdr0.cic2.comb3[19]$_SDFFE_PN0P__1031  (.L_HI(net1031));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[0]$_SDFFE_PN0P__1032  (.L_HI(net1032));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[10]$_SDFFE_PN0P__1033  (.L_HI(net1033));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[11]$_SDFFE_PN0P__1034  (.L_HI(net1034));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[12]$_SDFFE_PN0P__1035  (.L_HI(net1035));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[13]$_SDFFE_PN0P__1036  (.L_HI(net1036));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[14]$_SDFFE_PN0P__1037  (.L_HI(net1037));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[15]$_SDFFE_PN0P__1038  (.L_HI(net1038));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[16]$_SDFFE_PN0P__1039  (.L_HI(net1039));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[17]$_SDFFE_PN0P__1040  (.L_HI(net1040));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[18]$_SDFFE_PN0P__1041  (.L_HI(net1041));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[19]$_SDFFE_PN0P__1042  (.L_HI(net1042));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[1]$_SDFFE_PN0P__1043  (.L_HI(net1043));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[2]$_SDFFE_PN0P__1044  (.L_HI(net1044));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[3]$_SDFFE_PN0P__1045  (.L_HI(net1045));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[4]$_SDFFE_PN0P__1046  (.L_HI(net1046));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[5]$_SDFFE_PN0P__1047  (.L_HI(net1047));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[6]$_SDFFE_PN0P__1048  (.L_HI(net1048));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[7]$_SDFFE_PN0P__1049  (.L_HI(net1049));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[8]$_SDFFE_PN0P__1050  (.L_HI(net1050));
 sg13g2_tiehi \am_sdr0.cic2.comb3_in_del[9]$_SDFFE_PN0P__1051  (.L_HI(net1051));
 sg13g2_tiehi \am_sdr0.cic2.count[0]$_SDFFE_PN0P__1052  (.L_HI(net1052));
 sg13g2_tiehi \am_sdr0.cic2.count[1]$_SDFFE_PN0P__1053  (.L_HI(net1053));
 sg13g2_tiehi \am_sdr0.cic2.count[2]$_SDFFE_PN0P__1054  (.L_HI(net1054));
 sg13g2_tiehi \am_sdr0.cic2.count[3]$_SDFFE_PN0P__1055  (.L_HI(net1055));
 sg13g2_tiehi \am_sdr0.cic2.count[4]$_SDFFE_PN0P__1056  (.L_HI(net1056));
 sg13g2_tiehi \am_sdr0.cic2.count[5]$_SDFFE_PN0P__1057  (.L_HI(net1057));
 sg13g2_tiehi \am_sdr0.cic2.count[6]$_SDFFE_PN0P__1058  (.L_HI(net1058));
 sg13g2_tiehi \am_sdr0.cic2.count[7]$_SDFFE_PN0P__1059  (.L_HI(net1059));
 sg13g2_tiehi \am_sdr0.cic2.integ1[0]$_SDFFE_PN0P__1060  (.L_HI(net1060));
 sg13g2_tiehi \am_sdr0.cic2.integ1[10]$_SDFFE_PN0P__1061  (.L_HI(net1061));
 sg13g2_tiehi \am_sdr0.cic2.integ1[11]$_SDFFE_PN0P__1062  (.L_HI(net1062));
 sg13g2_tiehi \am_sdr0.cic2.integ1[12]$_SDFFE_PN0P__1063  (.L_HI(net1063));
 sg13g2_tiehi \am_sdr0.cic2.integ1[13]$_SDFFE_PN0P__1064  (.L_HI(net1064));
 sg13g2_tiehi \am_sdr0.cic2.integ1[14]$_SDFFE_PN0P__1065  (.L_HI(net1065));
 sg13g2_tiehi \am_sdr0.cic2.integ1[15]$_SDFFE_PN0P__1066  (.L_HI(net1066));
 sg13g2_tiehi \am_sdr0.cic2.integ1[16]$_SDFFE_PN0P__1067  (.L_HI(net1067));
 sg13g2_tiehi \am_sdr0.cic2.integ1[17]$_SDFFE_PN0P__1068  (.L_HI(net1068));
 sg13g2_tiehi \am_sdr0.cic2.integ1[18]$_SDFFE_PN0P__1069  (.L_HI(net1069));
 sg13g2_tiehi \am_sdr0.cic2.integ1[19]$_SDFFE_PN0P__1070  (.L_HI(net1070));
 sg13g2_tiehi \am_sdr0.cic2.integ1[1]$_SDFFE_PN0P__1071  (.L_HI(net1071));
 sg13g2_tiehi \am_sdr0.cic2.integ1[20]$_SDFFE_PN0P__1072  (.L_HI(net1072));
 sg13g2_tiehi \am_sdr0.cic2.integ1[21]$_SDFFE_PN0P__1073  (.L_HI(net1073));
 sg13g2_tiehi \am_sdr0.cic2.integ1[22]$_SDFFE_PN0P__1074  (.L_HI(net1074));
 sg13g2_tiehi \am_sdr0.cic2.integ1[23]$_SDFFE_PN0P__1075  (.L_HI(net1075));
 sg13g2_tiehi \am_sdr0.cic2.integ1[24]$_SDFFE_PN0P__1076  (.L_HI(net1076));
 sg13g2_tiehi \am_sdr0.cic2.integ1[25]$_SDFFE_PN0P__1077  (.L_HI(net1077));
 sg13g2_tiehi \am_sdr0.cic2.integ1[2]$_SDFFE_PN0P__1078  (.L_HI(net1078));
 sg13g2_tiehi \am_sdr0.cic2.integ1[3]$_SDFFE_PN0P__1079  (.L_HI(net1079));
 sg13g2_tiehi \am_sdr0.cic2.integ1[4]$_SDFFE_PN0P__1080  (.L_HI(net1080));
 sg13g2_tiehi \am_sdr0.cic2.integ1[5]$_SDFFE_PN0P__1081  (.L_HI(net1081));
 sg13g2_tiehi \am_sdr0.cic2.integ1[6]$_SDFFE_PN0P__1082  (.L_HI(net1082));
 sg13g2_tiehi \am_sdr0.cic2.integ1[7]$_SDFFE_PN0P__1083  (.L_HI(net1083));
 sg13g2_tiehi \am_sdr0.cic2.integ1[8]$_SDFFE_PN0P__1084  (.L_HI(net1084));
 sg13g2_tiehi \am_sdr0.cic2.integ1[9]$_SDFFE_PN0P__1085  (.L_HI(net1085));
 sg13g2_tiehi \am_sdr0.cic2.integ2[0]$_SDFFE_PN0P__1086  (.L_HI(net1086));
 sg13g2_tiehi \am_sdr0.cic2.integ2[10]$_SDFFE_PN0P__1087  (.L_HI(net1087));
 sg13g2_tiehi \am_sdr0.cic2.integ2[11]$_SDFFE_PN0P__1088  (.L_HI(net1088));
 sg13g2_tiehi \am_sdr0.cic2.integ2[12]$_SDFFE_PN0P__1089  (.L_HI(net1089));
 sg13g2_tiehi \am_sdr0.cic2.integ2[13]$_SDFFE_PN0P__1090  (.L_HI(net1090));
 sg13g2_tiehi \am_sdr0.cic2.integ2[14]$_SDFFE_PN0P__1091  (.L_HI(net1091));
 sg13g2_tiehi \am_sdr0.cic2.integ2[15]$_SDFFE_PN0P__1092  (.L_HI(net1092));
 sg13g2_tiehi \am_sdr0.cic2.integ2[16]$_SDFFE_PN0P__1093  (.L_HI(net1093));
 sg13g2_tiehi \am_sdr0.cic2.integ2[17]$_SDFFE_PN0P__1094  (.L_HI(net1094));
 sg13g2_tiehi \am_sdr0.cic2.integ2[18]$_SDFFE_PN0P__1095  (.L_HI(net1095));
 sg13g2_tiehi \am_sdr0.cic2.integ2[19]$_SDFFE_PN0P__1096  (.L_HI(net1096));
 sg13g2_tiehi \am_sdr0.cic2.integ2[1]$_SDFFE_PN0P__1097  (.L_HI(net1097));
 sg13g2_tiehi \am_sdr0.cic2.integ2[20]$_SDFFE_PN0P__1098  (.L_HI(net1098));
 sg13g2_tiehi \am_sdr0.cic2.integ2[21]$_SDFFE_PN0P__1099  (.L_HI(net1099));
 sg13g2_tiehi \am_sdr0.cic2.integ2[22]$_SDFFE_PN0P__1100  (.L_HI(net1100));
 sg13g2_tiehi \am_sdr0.cic2.integ2[2]$_SDFFE_PN0P__1101  (.L_HI(net1101));
 sg13g2_tiehi \am_sdr0.cic2.integ2[3]$_SDFFE_PN0P__1102  (.L_HI(net1102));
 sg13g2_tiehi \am_sdr0.cic2.integ2[4]$_SDFFE_PN0P__1103  (.L_HI(net1103));
 sg13g2_tiehi \am_sdr0.cic2.integ2[5]$_SDFFE_PN0P__1104  (.L_HI(net1104));
 sg13g2_tiehi \am_sdr0.cic2.integ2[6]$_SDFFE_PN0P__1105  (.L_HI(net1105));
 sg13g2_tiehi \am_sdr0.cic2.integ2[7]$_SDFFE_PN0P__1106  (.L_HI(net1106));
 sg13g2_tiehi \am_sdr0.cic2.integ2[8]$_SDFFE_PN0P__1107  (.L_HI(net1107));
 sg13g2_tiehi \am_sdr0.cic2.integ2[9]$_SDFFE_PN0P__1108  (.L_HI(net1108));
 sg13g2_tiehi \am_sdr0.cic2.integ3[0]$_SDFFE_PN0P__1109  (.L_HI(net1109));
 sg13g2_tiehi \am_sdr0.cic2.integ3[10]$_SDFFE_PN0P__1110  (.L_HI(net1110));
 sg13g2_tiehi \am_sdr0.cic2.integ3[11]$_SDFFE_PN0P__1111  (.L_HI(net1111));
 sg13g2_tiehi \am_sdr0.cic2.integ3[12]$_SDFFE_PN0P__1112  (.L_HI(net1112));
 sg13g2_tiehi \am_sdr0.cic2.integ3[13]$_SDFFE_PN0P__1113  (.L_HI(net1113));
 sg13g2_tiehi \am_sdr0.cic2.integ3[14]$_SDFFE_PN0P__1114  (.L_HI(net1114));
 sg13g2_tiehi \am_sdr0.cic2.integ3[15]$_SDFFE_PN0P__1115  (.L_HI(net1115));
 sg13g2_tiehi \am_sdr0.cic2.integ3[16]$_SDFFE_PN0P__1116  (.L_HI(net1116));
 sg13g2_tiehi \am_sdr0.cic2.integ3[17]$_SDFFE_PN0P__1117  (.L_HI(net1117));
 sg13g2_tiehi \am_sdr0.cic2.integ3[18]$_SDFFE_PN0P__1118  (.L_HI(net1118));
 sg13g2_tiehi \am_sdr0.cic2.integ3[19]$_SDFFE_PN0P__1119  (.L_HI(net1119));
 sg13g2_tiehi \am_sdr0.cic2.integ3[1]$_SDFFE_PN0P__1120  (.L_HI(net1120));
 sg13g2_tiehi \am_sdr0.cic2.integ3[2]$_SDFFE_PN0P__1121  (.L_HI(net1121));
 sg13g2_tiehi \am_sdr0.cic2.integ3[3]$_SDFFE_PN0P__1122  (.L_HI(net1122));
 sg13g2_tiehi \am_sdr0.cic2.integ3[4]$_SDFFE_PN0P__1123  (.L_HI(net1123));
 sg13g2_tiehi \am_sdr0.cic2.integ3[5]$_SDFFE_PN0P__1124  (.L_HI(net1124));
 sg13g2_tiehi \am_sdr0.cic2.integ3[6]$_SDFFE_PN0P__1125  (.L_HI(net1125));
 sg13g2_tiehi \am_sdr0.cic2.integ3[7]$_SDFFE_PN0P__1126  (.L_HI(net1126));
 sg13g2_tiehi \am_sdr0.cic2.integ3[8]$_SDFFE_PN0P__1127  (.L_HI(net1127));
 sg13g2_tiehi \am_sdr0.cic2.integ3[9]$_SDFFE_PN0P__1128  (.L_HI(net1128));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[0]$_DFFE_PP__1129  (.L_HI(net1129));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[10]$_DFFE_PP__1130  (.L_HI(net1130));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[11]$_DFFE_PP__1131  (.L_HI(net1131));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[12]$_DFFE_PP__1132  (.L_HI(net1132));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[13]$_DFFE_PP__1133  (.L_HI(net1133));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[14]$_DFFE_PP__1134  (.L_HI(net1134));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[15]$_DFFE_PP__1135  (.L_HI(net1135));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[16]$_DFFE_PP__1136  (.L_HI(net1136));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[17]$_DFFE_PP__1137  (.L_HI(net1137));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[18]$_DFFE_PP__1138  (.L_HI(net1138));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[19]$_DFFE_PP__1139  (.L_HI(net1139));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[1]$_DFFE_PP__1140  (.L_HI(net1140));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[2]$_DFFE_PP__1141  (.L_HI(net1141));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[3]$_DFFE_PP__1142  (.L_HI(net1142));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[4]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[5]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[6]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[7]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[8]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \am_sdr0.cic2.integ_sample[9]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \am_sdr0.cic2.out_tick$_SDFF_PN0__1149  (.L_HI(net1149));
 sg13g2_tiehi \am_sdr0.cic2.sample$_SDFF_PN0__1150  (.L_HI(net1150));
 sg13g2_tiehi \am_sdr0.cic2.x_out[10]$_SDFFE_PN0P__1151  (.L_HI(net1151));
 sg13g2_tiehi \am_sdr0.cic2.x_out[11]$_SDFFE_PN0P__1152  (.L_HI(net1152));
 sg13g2_tiehi \am_sdr0.cic2.x_out[12]$_SDFFE_PN0P__1153  (.L_HI(net1153));
 sg13g2_tiehi \am_sdr0.cic2.x_out[13]$_SDFFE_PN0P__1154  (.L_HI(net1154));
 sg13g2_tiehi \am_sdr0.cic2.x_out[14]$_SDFFE_PN0P__1155  (.L_HI(net1155));
 sg13g2_tiehi \am_sdr0.cic2.x_out[15]$_SDFFE_PN0P__1156  (.L_HI(net1156));
 sg13g2_tiehi \am_sdr0.cic2.x_out[8]$_SDFFE_PN0P__1157  (.L_HI(net1157));
 sg13g2_tiehi \am_sdr0.cic2.x_out[9]$_SDFFE_PN0P__1158  (.L_HI(net1158));
 sg13g2_tiehi \am_sdr0.cic3.comb1[0]$_SDFFE_PN0P__1159  (.L_HI(net1159));
 sg13g2_tiehi \am_sdr0.cic3.comb1[10]$_SDFFE_PN0P__1160  (.L_HI(net1160));
 sg13g2_tiehi \am_sdr0.cic3.comb1[11]$_SDFFE_PN0P__1161  (.L_HI(net1161));
 sg13g2_tiehi \am_sdr0.cic3.comb1[12]$_SDFFE_PN0P__1162  (.L_HI(net1162));
 sg13g2_tiehi \am_sdr0.cic3.comb1[13]$_SDFFE_PN0P__1163  (.L_HI(net1163));
 sg13g2_tiehi \am_sdr0.cic3.comb1[14]$_SDFFE_PN0P__1164  (.L_HI(net1164));
 sg13g2_tiehi \am_sdr0.cic3.comb1[15]$_SDFFE_PN0P__1165  (.L_HI(net1165));
 sg13g2_tiehi \am_sdr0.cic3.comb1[16]$_SDFFE_PN0P__1166  (.L_HI(net1166));
 sg13g2_tiehi \am_sdr0.cic3.comb1[17]$_SDFFE_PN0P__1167  (.L_HI(net1167));
 sg13g2_tiehi \am_sdr0.cic3.comb1[18]$_SDFFE_PN0P__1168  (.L_HI(net1168));
 sg13g2_tiehi \am_sdr0.cic3.comb1[19]$_SDFFE_PN0P__1169  (.L_HI(net1169));
 sg13g2_tiehi \am_sdr0.cic3.comb1[1]$_SDFFE_PN0P__1170  (.L_HI(net1170));
 sg13g2_tiehi \am_sdr0.cic3.comb1[2]$_SDFFE_PN0P__1171  (.L_HI(net1171));
 sg13g2_tiehi \am_sdr0.cic3.comb1[3]$_SDFFE_PN0P__1172  (.L_HI(net1172));
 sg13g2_tiehi \am_sdr0.cic3.comb1[4]$_SDFFE_PN0P__1173  (.L_HI(net1173));
 sg13g2_tiehi \am_sdr0.cic3.comb1[5]$_SDFFE_PN0P__1174  (.L_HI(net1174));
 sg13g2_tiehi \am_sdr0.cic3.comb1[6]$_SDFFE_PN0P__1175  (.L_HI(net1175));
 sg13g2_tiehi \am_sdr0.cic3.comb1[7]$_SDFFE_PN0P__1176  (.L_HI(net1176));
 sg13g2_tiehi \am_sdr0.cic3.comb1[8]$_SDFFE_PN0P__1177  (.L_HI(net1177));
 sg13g2_tiehi \am_sdr0.cic3.comb1[9]$_SDFFE_PN0P__1178  (.L_HI(net1178));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[0]$_SDFFE_PN0P__1179  (.L_HI(net1179));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[10]$_SDFFE_PN0P__1180  (.L_HI(net1180));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[11]$_SDFFE_PN0P__1181  (.L_HI(net1181));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[12]$_SDFFE_PN0P__1182  (.L_HI(net1182));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[13]$_SDFFE_PN0P__1183  (.L_HI(net1183));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[14]$_SDFFE_PN0P__1184  (.L_HI(net1184));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[15]$_SDFFE_PN0P__1185  (.L_HI(net1185));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[16]$_SDFFE_PN0P__1186  (.L_HI(net1186));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[17]$_SDFFE_PN0P__1187  (.L_HI(net1187));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[18]$_SDFFE_PN0P__1188  (.L_HI(net1188));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[19]$_SDFFE_PN0P__1189  (.L_HI(net1189));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[1]$_SDFFE_PN0P__1190  (.L_HI(net1190));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[2]$_SDFFE_PN0P__1191  (.L_HI(net1191));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[3]$_SDFFE_PN0P__1192  (.L_HI(net1192));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[4]$_SDFFE_PN0P__1193  (.L_HI(net1193));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[5]$_SDFFE_PN0P__1194  (.L_HI(net1194));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[6]$_SDFFE_PN0P__1195  (.L_HI(net1195));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[7]$_SDFFE_PN0P__1196  (.L_HI(net1196));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[8]$_SDFFE_PN0P__1197  (.L_HI(net1197));
 sg13g2_tiehi \am_sdr0.cic3.comb1_in_del[9]$_SDFFE_PN0P__1198  (.L_HI(net1198));
 sg13g2_tiehi \am_sdr0.cic3.comb2[0]$_SDFFE_PN0P__1199  (.L_HI(net1199));
 sg13g2_tiehi \am_sdr0.cic3.comb2[10]$_SDFFE_PN0P__1200  (.L_HI(net1200));
 sg13g2_tiehi \am_sdr0.cic3.comb2[11]$_SDFFE_PN0P__1201  (.L_HI(net1201));
 sg13g2_tiehi \am_sdr0.cic3.comb2[12]$_SDFFE_PN0P__1202  (.L_HI(net1202));
 sg13g2_tiehi \am_sdr0.cic3.comb2[13]$_SDFFE_PN0P__1203  (.L_HI(net1203));
 sg13g2_tiehi \am_sdr0.cic3.comb2[14]$_SDFFE_PN0P__1204  (.L_HI(net1204));
 sg13g2_tiehi \am_sdr0.cic3.comb2[15]$_SDFFE_PN0P__1205  (.L_HI(net1205));
 sg13g2_tiehi \am_sdr0.cic3.comb2[16]$_SDFFE_PN0P__1206  (.L_HI(net1206));
 sg13g2_tiehi \am_sdr0.cic3.comb2[17]$_SDFFE_PN0P__1207  (.L_HI(net1207));
 sg13g2_tiehi \am_sdr0.cic3.comb2[18]$_SDFFE_PN0P__1208  (.L_HI(net1208));
 sg13g2_tiehi \am_sdr0.cic3.comb2[19]$_SDFFE_PN0P__1209  (.L_HI(net1209));
 sg13g2_tiehi \am_sdr0.cic3.comb2[1]$_SDFFE_PN0P__1210  (.L_HI(net1210));
 sg13g2_tiehi \am_sdr0.cic3.comb2[2]$_SDFFE_PN0P__1211  (.L_HI(net1211));
 sg13g2_tiehi \am_sdr0.cic3.comb2[3]$_SDFFE_PN0P__1212  (.L_HI(net1212));
 sg13g2_tiehi \am_sdr0.cic3.comb2[4]$_SDFFE_PN0P__1213  (.L_HI(net1213));
 sg13g2_tiehi \am_sdr0.cic3.comb2[5]$_SDFFE_PN0P__1214  (.L_HI(net1214));
 sg13g2_tiehi \am_sdr0.cic3.comb2[6]$_SDFFE_PN0P__1215  (.L_HI(net1215));
 sg13g2_tiehi \am_sdr0.cic3.comb2[7]$_SDFFE_PN0P__1216  (.L_HI(net1216));
 sg13g2_tiehi \am_sdr0.cic3.comb2[8]$_SDFFE_PN0P__1217  (.L_HI(net1217));
 sg13g2_tiehi \am_sdr0.cic3.comb2[9]$_SDFFE_PN0P__1218  (.L_HI(net1218));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[0]$_SDFFE_PN0P__1219  (.L_HI(net1219));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[10]$_SDFFE_PN0P__1220  (.L_HI(net1220));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[11]$_SDFFE_PN0P__1221  (.L_HI(net1221));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[12]$_SDFFE_PN0P__1222  (.L_HI(net1222));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[13]$_SDFFE_PN0P__1223  (.L_HI(net1223));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[14]$_SDFFE_PN0P__1224  (.L_HI(net1224));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[15]$_SDFFE_PN0P__1225  (.L_HI(net1225));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[16]$_SDFFE_PN0P__1226  (.L_HI(net1226));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[17]$_SDFFE_PN0P__1227  (.L_HI(net1227));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[18]$_SDFFE_PN0P__1228  (.L_HI(net1228));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[19]$_SDFFE_PN0P__1229  (.L_HI(net1229));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[1]$_SDFFE_PN0P__1230  (.L_HI(net1230));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[2]$_SDFFE_PN0P__1231  (.L_HI(net1231));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[3]$_SDFFE_PN0P__1232  (.L_HI(net1232));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[4]$_SDFFE_PN0P__1233  (.L_HI(net1233));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[5]$_SDFFE_PN0P__1234  (.L_HI(net1234));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[6]$_SDFFE_PN0P__1235  (.L_HI(net1235));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[7]$_SDFFE_PN0P__1236  (.L_HI(net1236));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[8]$_SDFFE_PN0P__1237  (.L_HI(net1237));
 sg13g2_tiehi \am_sdr0.cic3.comb2_in_del[9]$_SDFFE_PN0P__1238  (.L_HI(net1238));
 sg13g2_tiehi \am_sdr0.cic3.comb3[12]$_SDFFE_PN0P__1239  (.L_HI(net1239));
 sg13g2_tiehi \am_sdr0.cic3.comb3[13]$_SDFFE_PN0P__1240  (.L_HI(net1240));
 sg13g2_tiehi \am_sdr0.cic3.comb3[14]$_SDFFE_PN0P__1241  (.L_HI(net1241));
 sg13g2_tiehi \am_sdr0.cic3.comb3[15]$_SDFFE_PN0P__1242  (.L_HI(net1242));
 sg13g2_tiehi \am_sdr0.cic3.comb3[16]$_SDFFE_PN0P__1243  (.L_HI(net1243));
 sg13g2_tiehi \am_sdr0.cic3.comb3[17]$_SDFFE_PN0P__1244  (.L_HI(net1244));
 sg13g2_tiehi \am_sdr0.cic3.comb3[18]$_SDFFE_PN0P__1245  (.L_HI(net1245));
 sg13g2_tiehi \am_sdr0.cic3.comb3[19]$_SDFFE_PN0P__1246  (.L_HI(net1246));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[0]$_SDFFE_PN0P__1247  (.L_HI(net1247));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[10]$_SDFFE_PN0P__1248  (.L_HI(net1248));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[11]$_SDFFE_PN0P__1249  (.L_HI(net1249));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[12]$_SDFFE_PN0P__1250  (.L_HI(net1250));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[13]$_SDFFE_PN0P__1251  (.L_HI(net1251));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[14]$_SDFFE_PN0P__1252  (.L_HI(net1252));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[15]$_SDFFE_PN0P__1253  (.L_HI(net1253));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[16]$_SDFFE_PN0P__1254  (.L_HI(net1254));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[17]$_SDFFE_PN0P__1255  (.L_HI(net1255));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[18]$_SDFFE_PN0P__1256  (.L_HI(net1256));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[19]$_SDFFE_PN0P__1257  (.L_HI(net1257));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[1]$_SDFFE_PN0P__1258  (.L_HI(net1258));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[2]$_SDFFE_PN0P__1259  (.L_HI(net1259));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[3]$_SDFFE_PN0P__1260  (.L_HI(net1260));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[4]$_SDFFE_PN0P__1261  (.L_HI(net1261));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[5]$_SDFFE_PN0P__1262  (.L_HI(net1262));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[6]$_SDFFE_PN0P__1263  (.L_HI(net1263));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[7]$_SDFFE_PN0P__1264  (.L_HI(net1264));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[8]$_SDFFE_PN0P__1265  (.L_HI(net1265));
 sg13g2_tiehi \am_sdr0.cic3.comb3_in_del[9]$_SDFFE_PN0P__1266  (.L_HI(net1266));
 sg13g2_tiehi \am_sdr0.cic3.count[0]$_SDFFE_PN0P__1267  (.L_HI(net1267));
 sg13g2_tiehi \am_sdr0.cic3.count[1]$_SDFFE_PN0P__1268  (.L_HI(net1268));
 sg13g2_tiehi \am_sdr0.cic3.count[2]$_SDFFE_PN0P__1269  (.L_HI(net1269));
 sg13g2_tiehi \am_sdr0.cic3.count[3]$_SDFFE_PN0P__1270  (.L_HI(net1270));
 sg13g2_tiehi \am_sdr0.cic3.count[4]$_SDFFE_PN0P__1271  (.L_HI(net1271));
 sg13g2_tiehi \am_sdr0.cic3.count[5]$_SDFFE_PN0P__1272  (.L_HI(net1272));
 sg13g2_tiehi \am_sdr0.cic3.count[6]$_SDFFE_PN0P__1273  (.L_HI(net1273));
 sg13g2_tiehi \am_sdr0.cic3.count[7]$_SDFFE_PN0P__1274  (.L_HI(net1274));
 sg13g2_tiehi \am_sdr0.cic3.integ1[0]$_SDFFE_PN0P__1275  (.L_HI(net1275));
 sg13g2_tiehi \am_sdr0.cic3.integ1[10]$_SDFFE_PN0P__1276  (.L_HI(net1276));
 sg13g2_tiehi \am_sdr0.cic3.integ1[11]$_SDFFE_PN0P__1277  (.L_HI(net1277));
 sg13g2_tiehi \am_sdr0.cic3.integ1[12]$_SDFFE_PN0P__1278  (.L_HI(net1278));
 sg13g2_tiehi \am_sdr0.cic3.integ1[13]$_SDFFE_PN0P__1279  (.L_HI(net1279));
 sg13g2_tiehi \am_sdr0.cic3.integ1[14]$_SDFFE_PN0P__1280  (.L_HI(net1280));
 sg13g2_tiehi \am_sdr0.cic3.integ1[15]$_SDFFE_PN0P__1281  (.L_HI(net1281));
 sg13g2_tiehi \am_sdr0.cic3.integ1[16]$_SDFFE_PN0P__1282  (.L_HI(net1282));
 sg13g2_tiehi \am_sdr0.cic3.integ1[17]$_SDFFE_PN0P__1283  (.L_HI(net1283));
 sg13g2_tiehi \am_sdr0.cic3.integ1[18]$_SDFFE_PN0P__1284  (.L_HI(net1284));
 sg13g2_tiehi \am_sdr0.cic3.integ1[19]$_SDFFE_PN0P__1285  (.L_HI(net1285));
 sg13g2_tiehi \am_sdr0.cic3.integ1[1]$_SDFFE_PN0P__1286  (.L_HI(net1286));
 sg13g2_tiehi \am_sdr0.cic3.integ1[20]$_SDFFE_PN0P__1287  (.L_HI(net1287));
 sg13g2_tiehi \am_sdr0.cic3.integ1[21]$_SDFFE_PN0P__1288  (.L_HI(net1288));
 sg13g2_tiehi \am_sdr0.cic3.integ1[22]$_SDFFE_PN0P__1289  (.L_HI(net1289));
 sg13g2_tiehi \am_sdr0.cic3.integ1[23]$_SDFFE_PN0P__1290  (.L_HI(net1290));
 sg13g2_tiehi \am_sdr0.cic3.integ1[24]$_SDFFE_PN0P__1291  (.L_HI(net1291));
 sg13g2_tiehi \am_sdr0.cic3.integ1[25]$_SDFFE_PN0P__1292  (.L_HI(net1292));
 sg13g2_tiehi \am_sdr0.cic3.integ1[2]$_SDFFE_PN0P__1293  (.L_HI(net1293));
 sg13g2_tiehi \am_sdr0.cic3.integ1[3]$_SDFFE_PN0P__1294  (.L_HI(net1294));
 sg13g2_tiehi \am_sdr0.cic3.integ1[4]$_SDFFE_PN0P__1295  (.L_HI(net1295));
 sg13g2_tiehi \am_sdr0.cic3.integ1[5]$_SDFFE_PN0P__1296  (.L_HI(net1296));
 sg13g2_tiehi \am_sdr0.cic3.integ1[6]$_SDFFE_PN0P__1297  (.L_HI(net1297));
 sg13g2_tiehi \am_sdr0.cic3.integ1[7]$_SDFFE_PN0P__1298  (.L_HI(net1298));
 sg13g2_tiehi \am_sdr0.cic3.integ1[8]$_SDFFE_PN0P__1299  (.L_HI(net1299));
 sg13g2_tiehi \am_sdr0.cic3.integ1[9]$_SDFFE_PN0P__1300  (.L_HI(net1300));
 sg13g2_tiehi \am_sdr0.cic3.integ2[0]$_SDFFE_PN0P__1301  (.L_HI(net1301));
 sg13g2_tiehi \am_sdr0.cic3.integ2[10]$_SDFFE_PN0P__1302  (.L_HI(net1302));
 sg13g2_tiehi \am_sdr0.cic3.integ2[11]$_SDFFE_PN0P__1303  (.L_HI(net1303));
 sg13g2_tiehi \am_sdr0.cic3.integ2[12]$_SDFFE_PN0P__1304  (.L_HI(net1304));
 sg13g2_tiehi \am_sdr0.cic3.integ2[13]$_SDFFE_PN0P__1305  (.L_HI(net1305));
 sg13g2_tiehi \am_sdr0.cic3.integ2[14]$_SDFFE_PN0P__1306  (.L_HI(net1306));
 sg13g2_tiehi \am_sdr0.cic3.integ2[15]$_SDFFE_PN0P__1307  (.L_HI(net1307));
 sg13g2_tiehi \am_sdr0.cic3.integ2[16]$_SDFFE_PN0P__1308  (.L_HI(net1308));
 sg13g2_tiehi \am_sdr0.cic3.integ2[17]$_SDFFE_PN0P__1309  (.L_HI(net1309));
 sg13g2_tiehi \am_sdr0.cic3.integ2[18]$_SDFFE_PN0P__1310  (.L_HI(net1310));
 sg13g2_tiehi \am_sdr0.cic3.integ2[19]$_SDFFE_PN0P__1311  (.L_HI(net1311));
 sg13g2_tiehi \am_sdr0.cic3.integ2[1]$_SDFFE_PN0P__1312  (.L_HI(net1312));
 sg13g2_tiehi \am_sdr0.cic3.integ2[20]$_SDFFE_PN0P__1313  (.L_HI(net1313));
 sg13g2_tiehi \am_sdr0.cic3.integ2[21]$_SDFFE_PN0P__1314  (.L_HI(net1314));
 sg13g2_tiehi \am_sdr0.cic3.integ2[22]$_SDFFE_PN0P__1315  (.L_HI(net1315));
 sg13g2_tiehi \am_sdr0.cic3.integ2[2]$_SDFFE_PN0P__1316  (.L_HI(net1316));
 sg13g2_tiehi \am_sdr0.cic3.integ2[3]$_SDFFE_PN0P__1317  (.L_HI(net1317));
 sg13g2_tiehi \am_sdr0.cic3.integ2[4]$_SDFFE_PN0P__1318  (.L_HI(net1318));
 sg13g2_tiehi \am_sdr0.cic3.integ2[5]$_SDFFE_PN0P__1319  (.L_HI(net1319));
 sg13g2_tiehi \am_sdr0.cic3.integ2[6]$_SDFFE_PN0P__1320  (.L_HI(net1320));
 sg13g2_tiehi \am_sdr0.cic3.integ2[7]$_SDFFE_PN0P__1321  (.L_HI(net1321));
 sg13g2_tiehi \am_sdr0.cic3.integ2[8]$_SDFFE_PN0P__1322  (.L_HI(net1322));
 sg13g2_tiehi \am_sdr0.cic3.integ2[9]$_SDFFE_PN0P__1323  (.L_HI(net1323));
 sg13g2_tiehi \am_sdr0.cic3.integ3[0]$_SDFFE_PN0P__1324  (.L_HI(net1324));
 sg13g2_tiehi \am_sdr0.cic3.integ3[10]$_SDFFE_PN0P__1325  (.L_HI(net1325));
 sg13g2_tiehi \am_sdr0.cic3.integ3[11]$_SDFFE_PN0P__1326  (.L_HI(net1326));
 sg13g2_tiehi \am_sdr0.cic3.integ3[12]$_SDFFE_PN0P__1327  (.L_HI(net1327));
 sg13g2_tiehi \am_sdr0.cic3.integ3[13]$_SDFFE_PN0P__1328  (.L_HI(net1328));
 sg13g2_tiehi \am_sdr0.cic3.integ3[14]$_SDFFE_PN0P__1329  (.L_HI(net1329));
 sg13g2_tiehi \am_sdr0.cic3.integ3[15]$_SDFFE_PN0P__1330  (.L_HI(net1330));
 sg13g2_tiehi \am_sdr0.cic3.integ3[16]$_SDFFE_PN0P__1331  (.L_HI(net1331));
 sg13g2_tiehi \am_sdr0.cic3.integ3[17]$_SDFFE_PN0P__1332  (.L_HI(net1332));
 sg13g2_tiehi \am_sdr0.cic3.integ3[18]$_SDFFE_PN0P__1333  (.L_HI(net1333));
 sg13g2_tiehi \am_sdr0.cic3.integ3[19]$_SDFFE_PN0P__1334  (.L_HI(net1334));
 sg13g2_tiehi \am_sdr0.cic3.integ3[1]$_SDFFE_PN0P__1335  (.L_HI(net1335));
 sg13g2_tiehi \am_sdr0.cic3.integ3[2]$_SDFFE_PN0P__1336  (.L_HI(net1336));
 sg13g2_tiehi \am_sdr0.cic3.integ3[3]$_SDFFE_PN0P__1337  (.L_HI(net1337));
 sg13g2_tiehi \am_sdr0.cic3.integ3[4]$_SDFFE_PN0P__1338  (.L_HI(net1338));
 sg13g2_tiehi \am_sdr0.cic3.integ3[5]$_SDFFE_PN0P__1339  (.L_HI(net1339));
 sg13g2_tiehi \am_sdr0.cic3.integ3[6]$_SDFFE_PN0P__1340  (.L_HI(net1340));
 sg13g2_tiehi \am_sdr0.cic3.integ3[7]$_SDFFE_PN0P__1341  (.L_HI(net1341));
 sg13g2_tiehi \am_sdr0.cic3.integ3[8]$_SDFFE_PN0P__1342  (.L_HI(net1342));
 sg13g2_tiehi \am_sdr0.cic3.integ3[9]$_SDFFE_PN0P__1343  (.L_HI(net1343));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[0]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[10]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[11]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[12]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[13]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[14]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[15]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[16]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[17]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[18]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[19]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[1]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[2]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[3]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[4]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[5]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[6]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[7]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[8]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \am_sdr0.cic3.integ_sample[9]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \am_sdr0.cic3.sample$_SDFF_PN0__1364  (.L_HI(net1364));
 sg13g2_tiehi \am_sdr0.cic3.x_out[10]$_SDFFE_PN0P__1365  (.L_HI(net1365));
 sg13g2_tiehi \am_sdr0.cic3.x_out[11]$_SDFFE_PN0P__1366  (.L_HI(net1366));
 sg13g2_tiehi \am_sdr0.cic3.x_out[12]$_SDFFE_PN0P__1367  (.L_HI(net1367));
 sg13g2_tiehi \am_sdr0.cic3.x_out[13]$_SDFFE_PN0P__1368  (.L_HI(net1368));
 sg13g2_tiehi \am_sdr0.cic3.x_out[14]$_SDFFE_PN0P__1369  (.L_HI(net1369));
 sg13g2_tiehi \am_sdr0.cic3.x_out[15]$_SDFFE_PN0P__1370  (.L_HI(net1370));
 sg13g2_tiehi \am_sdr0.cic3.x_out[8]$_SDFFE_PN0P__1371  (.L_HI(net1371));
 sg13g2_tiehi \am_sdr0.cic3.x_out[9]$_SDFFE_PN0P__1372  (.L_HI(net1372));
 sg13g2_tiehi \am_sdr0.count[0]$_SDFF_PN0__1373  (.L_HI(net1373));
 sg13g2_tiehi \am_sdr0.count[1]$_SDFF_PN0__1374  (.L_HI(net1374));
 sg13g2_tiehi \am_sdr0.count[2]$_SDFF_PN0__1375  (.L_HI(net1375));
 sg13g2_tiehi \am_sdr0.count[3]$_SDFF_PN0__1376  (.L_HI(net1376));
 sg13g2_tiehi \am_sdr0.count[4]$_SDFF_PN0__1377  (.L_HI(net1377));
 sg13g2_tiehi \am_sdr0.count[5]$_SDFF_PN0__1378  (.L_HI(net1378));
 sg13g2_tiehi \am_sdr0.count[6]$_SDFF_PN0__1379  (.L_HI(net1379));
 sg13g2_tiehi \am_sdr0.count[7]$_SDFF_PN0__1380  (.L_HI(net1380));
 sg13g2_tiehi \am_sdr0.mix0.I_out[0]$_DFF_P__1381  (.L_HI(net1381));
 sg13g2_tiehi \am_sdr0.mix0.I_out[1]$_DFF_P__1382  (.L_HI(net1382));
 sg13g2_tiehi \am_sdr0.mix0.I_out[2]$_DFF_P__1383  (.L_HI(net1383));
 sg13g2_tiehi \am_sdr0.mix0.I_out[3]$_DFF_P__1384  (.L_HI(net1384));
 sg13g2_tiehi \am_sdr0.mix0.I_out[4]$_DFF_P__1385  (.L_HI(net1385));
 sg13g2_tiehi \am_sdr0.mix0.I_out[5]$_DFF_P__1386  (.L_HI(net1386));
 sg13g2_tiehi \am_sdr0.mix0.I_out[6]$_DFF_P__1387  (.L_HI(net1387));
 sg13g2_tiehi \am_sdr0.mix0.I_out[7]$_DFF_P__1388  (.L_HI(net1388));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[0]$_DFF_P__1389  (.L_HI(net1389));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[1]$_DFF_P__1390  (.L_HI(net1390));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[2]$_DFF_P__1391  (.L_HI(net1391));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[3]$_DFF_P__1392  (.L_HI(net1392));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[4]$_DFF_P__1393  (.L_HI(net1393));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[5]$_DFF_P__1394  (.L_HI(net1394));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[6]$_DFF_P__1395  (.L_HI(net1395));
 sg13g2_tiehi \am_sdr0.mix0.Q_out[7]$_DFF_P__1396  (.L_HI(net1396));
 sg13g2_tiehi \am_sdr0.mix0.RF_in_q$_SDFF_PN0__1397  (.L_HI(net1397));
 sg13g2_tiehi \am_sdr0.mix0.RF_in_qq$_SDFF_PN0__1398  (.L_HI(net1398));
 sg13g2_tiehi \am_sdr0.mix0.RF_out$_SDFF_PN0__1399  (.L_HI(net1399));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[0]$_SDFF_PN0__1400  (.L_HI(net1400));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[1]$_SDFF_PN0__1401  (.L_HI(net1401));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[2]$_SDFF_PN0__1402  (.L_HI(net1402));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[3]$_SDFF_PN0__1403  (.L_HI(net1403));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[4]$_SDFF_PN0__1404  (.L_HI(net1404));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[5]$_SDFF_PN0__1405  (.L_HI(net1405));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[6]$_SDFF_PN0__1406  (.L_HI(net1406));
 sg13g2_tiehi \am_sdr0.mix0.cos_q[7]$_SDFF_PN0__1407  (.L_HI(net1407));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[0]$_SDFF_PN0__1408  (.L_HI(net1408));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[1]$_SDFF_PN0__1409  (.L_HI(net1409));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[2]$_SDFF_PN0__1410  (.L_HI(net1410));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[3]$_SDFF_PN0__1411  (.L_HI(net1411));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[4]$_SDFF_PN0__1412  (.L_HI(net1412));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[5]$_SDFF_PN0__1413  (.L_HI(net1413));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[6]$_SDFF_PN0__1414  (.L_HI(net1414));
 sg13g2_tiehi \am_sdr0.mix0.sin_q[7]$_SDFF_PN0__1415  (.L_HI(net1415));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[0]$_DFF_P__1416  (.L_HI(net1416));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[1]$_DFF_P__1417  (.L_HI(net1417));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[2]$_DFF_P__1418  (.L_HI(net1418));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[3]$_DFF_P__1419  (.L_HI(net1419));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[4]$_DFF_P__1420  (.L_HI(net1420));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[5]$_DFF_P__1421  (.L_HI(net1421));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[6]$_DFF_P__1422  (.L_HI(net1422));
 sg13g2_tiehi \am_sdr0.nco0.cos0.data[7]$_DFF_P__1423  (.L_HI(net1423));
 sg13g2_tiehi \am_sdr0.nco0.phase[0]$_SDFF_PN0__1424  (.L_HI(net1424));
 sg13g2_tiehi \am_sdr0.nco0.phase[10]$_SDFF_PN0__1425  (.L_HI(net1425));
 sg13g2_tiehi \am_sdr0.nco0.phase[11]$_SDFF_PN0__1426  (.L_HI(net1426));
 sg13g2_tiehi \am_sdr0.nco0.phase[12]$_SDFF_PN0__1427  (.L_HI(net1427));
 sg13g2_tiehi \am_sdr0.nco0.phase[13]$_SDFF_PN0__1428  (.L_HI(net1428));
 sg13g2_tiehi \am_sdr0.nco0.phase[14]$_SDFF_PN0__1429  (.L_HI(net1429));
 sg13g2_tiehi \am_sdr0.nco0.phase[15]$_SDFF_PN0__1430  (.L_HI(net1430));
 sg13g2_tiehi \am_sdr0.nco0.phase[16]$_SDFF_PN0__1431  (.L_HI(net1431));
 sg13g2_tiehi \am_sdr0.nco0.phase[17]$_SDFF_PN0__1432  (.L_HI(net1432));
 sg13g2_tiehi \am_sdr0.nco0.phase[18]$_SDFF_PN0__1433  (.L_HI(net1433));
 sg13g2_tiehi \am_sdr0.nco0.phase[19]$_SDFF_PN0__1434  (.L_HI(net1434));
 sg13g2_tiehi \am_sdr0.nco0.phase[1]$_SDFF_PN0__1435  (.L_HI(net1435));
 sg13g2_tiehi \am_sdr0.nco0.phase[20]$_SDFF_PN0__1436  (.L_HI(net1436));
 sg13g2_tiehi \am_sdr0.nco0.phase[21]$_SDFF_PN0__1437  (.L_HI(net1437));
 sg13g2_tiehi \am_sdr0.nco0.phase[22]$_SDFF_PN0__1438  (.L_HI(net1438));
 sg13g2_tiehi \am_sdr0.nco0.phase[23]$_SDFF_PN0__1439  (.L_HI(net1439));
 sg13g2_tiehi \am_sdr0.nco0.phase[24]$_SDFF_PN0__1440  (.L_HI(net1440));
 sg13g2_tiehi \am_sdr0.nco0.phase[25]$_SDFF_PN0__1441  (.L_HI(net1441));
 sg13g2_tiehi \am_sdr0.nco0.phase[2]$_SDFF_PN0__1442  (.L_HI(net1442));
 sg13g2_tiehi \am_sdr0.nco0.phase[3]$_SDFF_PN0__1443  (.L_HI(net1443));
 sg13g2_tiehi \am_sdr0.nco0.phase[4]$_SDFF_PN0__1444  (.L_HI(net1444));
 sg13g2_tiehi \am_sdr0.nco0.phase[5]$_SDFF_PN0__1445  (.L_HI(net1445));
 sg13g2_tiehi \am_sdr0.nco0.phase[6]$_SDFF_PN0__1446  (.L_HI(net1446));
 sg13g2_tiehi \am_sdr0.nco0.phase[7]$_SDFF_PN0__1447  (.L_HI(net1447));
 sg13g2_tiehi \am_sdr0.nco0.phase[8]$_SDFF_PN0__1448  (.L_HI(net1448));
 sg13g2_tiehi \am_sdr0.nco0.phase[9]$_SDFF_PN0__1449  (.L_HI(net1449));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[0]$_DFF_P__1450  (.L_HI(net1450));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[1]$_DFF_P__1451  (.L_HI(net1451));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[2]$_DFF_P__1452  (.L_HI(net1452));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[3]$_DFF_P__1453  (.L_HI(net1453));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[4]$_DFF_P__1454  (.L_HI(net1454));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[5]$_DFF_P__1455  (.L_HI(net1455));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[6]$_DFF_P__1456  (.L_HI(net1456));
 sg13g2_tiehi \am_sdr0.nco0.sin0.data[7]$_SDFF_PN0__1457  (.L_HI(net1457));
 sg13g2_tiehi \am_sdr0.spi0.CS_q$_SDFF_PN0__1458  (.L_HI(net1458));
 sg13g2_tiehi \am_sdr0.spi0.CS_qq$_SDFF_PN0__1459  (.L_HI(net1459));
 sg13g2_tiehi \am_sdr0.spi0.CS_qqq$_SDFF_PN0__1460  (.L_HI(net1460));
 sg13g2_tiehi \am_sdr0.spi0.MOSI_q$_SDFF_PN0__1461  (.L_HI(net1461));
 sg13g2_tiehi \am_sdr0.spi0.MOSI_qq$_SDFF_PN0__1462  (.L_HI(net1462));
 sg13g2_tiehi \am_sdr0.spi0.SCK_q$_SDFF_PN0__1463  (.L_HI(net1463));
 sg13g2_tiehi \am_sdr0.spi0.SCK_qq$_SDFF_PN0__1464  (.L_HI(net1464));
 sg13g2_tiehi \am_sdr0.spi0.SCK_qqq$_SDFF_PN0__1465  (.L_HI(net1465));
 sg13g2_tiehi \am_sdr0.spi0.gain[0]$_SDFFE_PN0N__1466  (.L_HI(net1466));
 sg13g2_tiehi \am_sdr0.spi0.gain[1]$_SDFFE_PN1N__1467  (.L_HI(net1467));
 sg13g2_tiehi \am_sdr0.spi0.gain[2]$_SDFFE_PN0N__1468  (.L_HI(net1468));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[0]$_SDFFE_PN1N__1469  (.L_HI(net1469));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[10]$_SDFFE_PN0N__1470  (.L_HI(net1470));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[11]$_SDFFE_PN0N__1471  (.L_HI(net1471));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[12]$_SDFFE_PN1N__1472  (.L_HI(net1472));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[13]$_SDFFE_PN0N__1473  (.L_HI(net1473));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[14]$_SDFFE_PN0N__1474  (.L_HI(net1474));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[15]$_SDFFE_PN0N__1475  (.L_HI(net1475));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[16]$_SDFFE_PN1N__1476  (.L_HI(net1476));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[17]$_SDFFE_PN1N__1477  (.L_HI(net1477));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[18]$_SDFFE_PN0N__1478  (.L_HI(net1478));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[19]$_SDFFE_PN0N__1479  (.L_HI(net1479));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[1]$_SDFFE_PN1N__1480  (.L_HI(net1480));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[20]$_SDFFE_PN1N__1481  (.L_HI(net1481));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[21]$_SDFFE_PN0N__1482  (.L_HI(net1482));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[22]$_SDFFE_PN0N__1483  (.L_HI(net1483));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[23]$_SDFFE_PN0N__1484  (.L_HI(net1484));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[24]$_SDFFE_PN0N__1485  (.L_HI(net1485));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[25]$_SDFFE_PN0N__1486  (.L_HI(net1486));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[2]$_SDFFE_PN0N__1487  (.L_HI(net1487));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[3]$_SDFFE_PN1N__1488  (.L_HI(net1488));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[4]$_SDFFE_PN0N__1489  (.L_HI(net1489));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[5]$_SDFFE_PN1N__1490  (.L_HI(net1490));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[6]$_SDFFE_PN1N__1491  (.L_HI(net1491));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[7]$_SDFFE_PN1N__1492  (.L_HI(net1492));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[8]$_SDFFE_PN0N__1493  (.L_HI(net1493));
 sg13g2_tiehi \am_sdr0.spi0.phase_inc[9]$_SDFFE_PN1N__1494  (.L_HI(net1494));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[0]$_SDFFCE_PN0P__1495  (.L_HI(net1495));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[10]$_SDFFCE_PN0P__1496  (.L_HI(net1496));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[11]$_SDFFCE_PN0P__1497  (.L_HI(net1497));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[12]$_SDFFCE_PN0P__1498  (.L_HI(net1498));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[13]$_SDFFCE_PN0P__1499  (.L_HI(net1499));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[14]$_SDFFCE_PN0P__1500  (.L_HI(net1500));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[15]$_SDFFCE_PN0P__1501  (.L_HI(net1501));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[16]$_SDFFCE_PN0P__1502  (.L_HI(net1502));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[17]$_SDFFCE_PN0P__1503  (.L_HI(net1503));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[18]$_SDFFCE_PN0P__1504  (.L_HI(net1504));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[19]$_SDFFCE_PN0P__1505  (.L_HI(net1505));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[1]$_SDFFCE_PN0P__1506  (.L_HI(net1506));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[20]$_SDFFCE_PN0P__1507  (.L_HI(net1507));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[21]$_SDFFCE_PN0P__1508  (.L_HI(net1508));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[22]$_SDFFCE_PN0P__1509  (.L_HI(net1509));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[23]$_SDFFCE_PN0P__1510  (.L_HI(net1510));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[24]$_SDFFCE_PN0P__1511  (.L_HI(net1511));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[25]$_SDFFCE_PN0P__1512  (.L_HI(net1512));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[26]$_SDFFCE_PN0P__1513  (.L_HI(net1513));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[27]$_SDFFCE_PN0P__1514  (.L_HI(net1514));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[28]$_SDFFCE_PN0P__1515  (.L_HI(net1515));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[2]$_SDFFCE_PN0P__1516  (.L_HI(net1516));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[3]$_SDFFCE_PN0P__1517  (.L_HI(net1517));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[4]$_SDFFCE_PN0P__1518  (.L_HI(net1518));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[5]$_SDFFCE_PN0P__1519  (.L_HI(net1519));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[6]$_SDFFCE_PN0P__1520  (.L_HI(net1520));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[7]$_SDFFCE_PN0P__1521  (.L_HI(net1521));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[8]$_SDFFCE_PN0P__1522  (.L_HI(net1522));
 sg13g2_tiehi \am_sdr0.spi0.shift_reg[9]$_SDFFCE_PN0P__1523  (.L_HI(net1523));
 sg13g2_tiehi \am_sdr0.spi0.state[0]$_SDFFE_PN0P__1524  (.L_HI(net1524));
 sg13g2_tiehi \am_sdr0.spi0.state[1]$_SDFFE_PN0P__1525  (.L_HI(net1525));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_77_clk (.X(clknet_leaf_77_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_138_clk (.X(clknet_leaf_138_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_139_clk (.X(clknet_leaf_139_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_140_clk (.X(clknet_leaf_140_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_141_clk (.X(clknet_leaf_141_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_142_clk (.X(clknet_leaf_142_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_143_clk (.X(clknet_leaf_143_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_144_clk (.X(clknet_leaf_144_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_145_clk (.X(clknet_leaf_145_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_146_clk (.X(clknet_leaf_146_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkload10 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkload11 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkload12 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_145_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_146_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_135_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_29_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_36_clk));
 sg13g2_inv_1 clkload20 (.A(clknet_leaf_22_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_118_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_120_clk));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_125_clk));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_96_clk));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_110_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_107_clk));
 sg13g2_inv_1 clkload28 (.A(clknet_leaf_65_clk));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_94_clk));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_66_clk));
 sg13g2_inv_1 clkload31 (.A(clknet_leaf_92_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_89_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_01558_));
 sg13g2_antennanp ANTENNA_2 (.A(_01558_));
 sg13g2_antennanp ANTENNA_3 (.A(_01558_));
 sg13g2_antennanp ANTENNA_4 (.A(_01558_));
 sg13g2_antennanp ANTENNA_5 (.A(_04198_));
 sg13g2_antennanp ANTENNA_6 (.A(_04198_));
 sg13g2_antennanp ANTENNA_7 (.A(_04198_));
 sg13g2_antennanp ANTENNA_8 (.A(_04198_));
 sg13g2_antennanp ANTENNA_9 (.A(_05246_));
 sg13g2_antennanp ANTENNA_10 (.A(_05246_));
 sg13g2_antennanp ANTENNA_11 (.A(_05246_));
 sg13g2_antennanp ANTENNA_12 (.A(_07113_));
 sg13g2_antennanp ANTENNA_13 (.A(_07113_));
 sg13g2_antennanp ANTENNA_14 (.A(_07113_));
 sg13g2_antennanp ANTENNA_15 (.A(_07113_));
 sg13g2_antennanp ANTENNA_16 (.A(_07113_));
 sg13g2_antennanp ANTENNA_17 (.A(_07113_));
 sg13g2_antennanp ANTENNA_18 (.A(_07113_));
 sg13g2_antennanp ANTENNA_19 (.A(_07113_));
 sg13g2_antennanp ANTENNA_20 (.A(clk));
 sg13g2_antennanp ANTENNA_21 (.A(net191));
 sg13g2_antennanp ANTENNA_22 (.A(net191));
 sg13g2_antennanp ANTENNA_23 (.A(net191));
 sg13g2_antennanp ANTENNA_24 (.A(net191));
 sg13g2_antennanp ANTENNA_25 (.A(net191));
 sg13g2_antennanp ANTENNA_26 (.A(net191));
 sg13g2_antennanp ANTENNA_27 (.A(net191));
 sg13g2_antennanp ANTENNA_28 (.A(net191));
 sg13g2_antennanp ANTENNA_29 (.A(net210));
 sg13g2_antennanp ANTENNA_30 (.A(net210));
 sg13g2_antennanp ANTENNA_31 (.A(net210));
 sg13g2_antennanp ANTENNA_32 (.A(net210));
 sg13g2_antennanp ANTENNA_33 (.A(net210));
 sg13g2_antennanp ANTENNA_34 (.A(net210));
 sg13g2_antennanp ANTENNA_35 (.A(net210));
 sg13g2_antennanp ANTENNA_36 (.A(net210));
 sg13g2_antennanp ANTENNA_37 (.A(net210));
 sg13g2_antennanp ANTENNA_38 (.A(net297));
 sg13g2_antennanp ANTENNA_39 (.A(net297));
 sg13g2_antennanp ANTENNA_40 (.A(net297));
 sg13g2_antennanp ANTENNA_41 (.A(net297));
 sg13g2_antennanp ANTENNA_42 (.A(net297));
 sg13g2_antennanp ANTENNA_43 (.A(net297));
 sg13g2_antennanp ANTENNA_44 (.A(net297));
 sg13g2_antennanp ANTENNA_45 (.A(net297));
 sg13g2_antennanp ANTENNA_46 (.A(net297));
 sg13g2_antennanp ANTENNA_47 (.A(net297));
 sg13g2_antennanp ANTENNA_48 (.A(net297));
 sg13g2_antennanp ANTENNA_49 (.A(net297));
 sg13g2_antennanp ANTENNA_50 (.A(net297));
 sg13g2_antennanp ANTENNA_51 (.A(net297));
 sg13g2_antennanp ANTENNA_52 (.A(net297));
 sg13g2_antennanp ANTENNA_53 (.A(net297));
 sg13g2_antennanp ANTENNA_54 (.A(net297));
 sg13g2_antennanp ANTENNA_55 (.A(net297));
 sg13g2_antennanp ANTENNA_56 (.A(net297));
 sg13g2_antennanp ANTENNA_57 (.A(net297));
 sg13g2_antennanp ANTENNA_58 (.A(net297));
 sg13g2_antennanp ANTENNA_59 (.A(net297));
 sg13g2_antennanp ANTENNA_60 (.A(_01558_));
 sg13g2_antennanp ANTENNA_61 (.A(_01558_));
 sg13g2_antennanp ANTENNA_62 (.A(_01558_));
 sg13g2_antennanp ANTENNA_63 (.A(_01558_));
 sg13g2_antennanp ANTENNA_64 (.A(_04198_));
 sg13g2_antennanp ANTENNA_65 (.A(_04198_));
 sg13g2_antennanp ANTENNA_66 (.A(_04198_));
 sg13g2_antennanp ANTENNA_67 (.A(_04198_));
 sg13g2_antennanp ANTENNA_68 (.A(_05246_));
 sg13g2_antennanp ANTENNA_69 (.A(_05246_));
 sg13g2_antennanp ANTENNA_70 (.A(_05246_));
 sg13g2_antennanp ANTENNA_71 (.A(_07113_));
 sg13g2_antennanp ANTENNA_72 (.A(_07113_));
 sg13g2_antennanp ANTENNA_73 (.A(_07113_));
 sg13g2_antennanp ANTENNA_74 (.A(_07113_));
 sg13g2_antennanp ANTENNA_75 (.A(_07113_));
 sg13g2_antennanp ANTENNA_76 (.A(_07113_));
 sg13g2_antennanp ANTENNA_77 (.A(_07113_));
 sg13g2_antennanp ANTENNA_78 (.A(_07113_));
 sg13g2_antennanp ANTENNA_79 (.A(clk));
 sg13g2_antennanp ANTENNA_80 (.A(net210));
 sg13g2_antennanp ANTENNA_81 (.A(net210));
 sg13g2_antennanp ANTENNA_82 (.A(net210));
 sg13g2_antennanp ANTENNA_83 (.A(net210));
 sg13g2_antennanp ANTENNA_84 (.A(net210));
 sg13g2_antennanp ANTENNA_85 (.A(net210));
 sg13g2_antennanp ANTENNA_86 (.A(net210));
 sg13g2_antennanp ANTENNA_87 (.A(net210));
 sg13g2_antennanp ANTENNA_88 (.A(net210));
 sg13g2_antennanp ANTENNA_89 (.A(_01558_));
 sg13g2_antennanp ANTENNA_90 (.A(_01558_));
 sg13g2_antennanp ANTENNA_91 (.A(_01558_));
 sg13g2_antennanp ANTENNA_92 (.A(_01558_));
 sg13g2_antennanp ANTENNA_93 (.A(_04198_));
 sg13g2_antennanp ANTENNA_94 (.A(_04198_));
 sg13g2_antennanp ANTENNA_95 (.A(_04198_));
 sg13g2_antennanp ANTENNA_96 (.A(_04198_));
 sg13g2_antennanp ANTENNA_97 (.A(_05246_));
 sg13g2_antennanp ANTENNA_98 (.A(_05246_));
 sg13g2_antennanp ANTENNA_99 (.A(_05246_));
 sg13g2_antennanp ANTENNA_100 (.A(_07113_));
 sg13g2_antennanp ANTENNA_101 (.A(_07113_));
 sg13g2_antennanp ANTENNA_102 (.A(_07113_));
 sg13g2_antennanp ANTENNA_103 (.A(_07113_));
 sg13g2_antennanp ANTENNA_104 (.A(_07113_));
 sg13g2_antennanp ANTENNA_105 (.A(_07113_));
 sg13g2_antennanp ANTENNA_106 (.A(_07113_));
 sg13g2_antennanp ANTENNA_107 (.A(_07113_));
 sg13g2_antennanp ANTENNA_108 (.A(clk));
 sg13g2_antennanp ANTENNA_109 (.A(clk));
 sg13g2_antennanp ANTENNA_110 (.A(net210));
 sg13g2_antennanp ANTENNA_111 (.A(net210));
 sg13g2_antennanp ANTENNA_112 (.A(net210));
 sg13g2_antennanp ANTENNA_113 (.A(net210));
 sg13g2_antennanp ANTENNA_114 (.A(net210));
 sg13g2_antennanp ANTENNA_115 (.A(net210));
 sg13g2_antennanp ANTENNA_116 (.A(net210));
 sg13g2_antennanp ANTENNA_117 (.A(net210));
 sg13g2_antennanp ANTENNA_118 (.A(net210));
 sg13g2_antennanp ANTENNA_119 (.A(_01558_));
 sg13g2_antennanp ANTENNA_120 (.A(_01558_));
 sg13g2_antennanp ANTENNA_121 (.A(_01558_));
 sg13g2_antennanp ANTENNA_122 (.A(_05246_));
 sg13g2_antennanp ANTENNA_123 (.A(_05246_));
 sg13g2_antennanp ANTENNA_124 (.A(_05246_));
 sg13g2_antennanp ANTENNA_125 (.A(_07113_));
 sg13g2_antennanp ANTENNA_126 (.A(_07113_));
 sg13g2_antennanp ANTENNA_127 (.A(_07113_));
 sg13g2_antennanp ANTENNA_128 (.A(_07113_));
 sg13g2_antennanp ANTENNA_129 (.A(_07113_));
 sg13g2_antennanp ANTENNA_130 (.A(_07113_));
 sg13g2_antennanp ANTENNA_131 (.A(_07113_));
 sg13g2_antennanp ANTENNA_132 (.A(_07113_));
 sg13g2_antennanp ANTENNA_133 (.A(clk));
 sg13g2_antennanp ANTENNA_134 (.A(clk));
 sg13g2_antennanp ANTENNA_135 (.A(net210));
 sg13g2_antennanp ANTENNA_136 (.A(net210));
 sg13g2_antennanp ANTENNA_137 (.A(net210));
 sg13g2_antennanp ANTENNA_138 (.A(net210));
 sg13g2_antennanp ANTENNA_139 (.A(net210));
 sg13g2_antennanp ANTENNA_140 (.A(net210));
 sg13g2_antennanp ANTENNA_141 (.A(net210));
 sg13g2_antennanp ANTENNA_142 (.A(net210));
 sg13g2_antennanp ANTENNA_143 (.A(net210));
 sg13g2_antennanp ANTENNA_144 (.A(_01558_));
 sg13g2_antennanp ANTENNA_145 (.A(_01558_));
 sg13g2_antennanp ANTENNA_146 (.A(_01558_));
 sg13g2_antennanp ANTENNA_147 (.A(_05246_));
 sg13g2_antennanp ANTENNA_148 (.A(_05246_));
 sg13g2_antennanp ANTENNA_149 (.A(_05246_));
 sg13g2_antennanp ANTENNA_150 (.A(_07113_));
 sg13g2_antennanp ANTENNA_151 (.A(_07113_));
 sg13g2_antennanp ANTENNA_152 (.A(_07113_));
 sg13g2_antennanp ANTENNA_153 (.A(_07113_));
 sg13g2_antennanp ANTENNA_154 (.A(_07113_));
 sg13g2_antennanp ANTENNA_155 (.A(_07113_));
 sg13g2_antennanp ANTENNA_156 (.A(_07113_));
 sg13g2_antennanp ANTENNA_157 (.A(_07113_));
 sg13g2_antennanp ANTENNA_158 (.A(clk));
 sg13g2_antennanp ANTENNA_159 (.A(clk));
 sg13g2_antennanp ANTENNA_160 (.A(net210));
 sg13g2_antennanp ANTENNA_161 (.A(net210));
 sg13g2_antennanp ANTENNA_162 (.A(net210));
 sg13g2_antennanp ANTENNA_163 (.A(net210));
 sg13g2_antennanp ANTENNA_164 (.A(net210));
 sg13g2_antennanp ANTENNA_165 (.A(net210));
 sg13g2_antennanp ANTENNA_166 (.A(net210));
 sg13g2_antennanp ANTENNA_167 (.A(net210));
 sg13g2_antennanp ANTENNA_168 (.A(net210));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_fill_1 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_467 ();
 sg13g2_decap_4 FILLER_0_474 ();
 sg13g2_decap_8 FILLER_0_508 ();
 sg13g2_decap_8 FILLER_0_515 ();
 sg13g2_decap_8 FILLER_0_522 ();
 sg13g2_decap_8 FILLER_0_529 ();
 sg13g2_decap_8 FILLER_0_540 ();
 sg13g2_decap_8 FILLER_0_547 ();
 sg13g2_decap_8 FILLER_0_554 ();
 sg13g2_decap_8 FILLER_0_561 ();
 sg13g2_decap_8 FILLER_0_568 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_decap_8 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_589 ();
 sg13g2_decap_8 FILLER_0_596 ();
 sg13g2_decap_8 FILLER_0_603 ();
 sg13g2_decap_8 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_617 ();
 sg13g2_decap_8 FILLER_0_624 ();
 sg13g2_decap_8 FILLER_0_631 ();
 sg13g2_decap_4 FILLER_0_638 ();
 sg13g2_fill_2 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_decap_8 FILLER_0_663 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_8 FILLER_0_698 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_decap_8 FILLER_0_712 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_747 ();
 sg13g2_fill_2 FILLER_0_754 ();
 sg13g2_decap_8 FILLER_0_782 ();
 sg13g2_decap_8 FILLER_0_789 ();
 sg13g2_decap_8 FILLER_0_796 ();
 sg13g2_decap_8 FILLER_0_803 ();
 sg13g2_decap_8 FILLER_0_810 ();
 sg13g2_decap_8 FILLER_0_817 ();
 sg13g2_decap_8 FILLER_0_824 ();
 sg13g2_fill_2 FILLER_0_857 ();
 sg13g2_fill_1 FILLER_0_859 ();
 sg13g2_decap_8 FILLER_0_894 ();
 sg13g2_decap_8 FILLER_0_901 ();
 sg13g2_decap_8 FILLER_0_908 ();
 sg13g2_decap_8 FILLER_0_915 ();
 sg13g2_decap_8 FILLER_0_922 ();
 sg13g2_decap_8 FILLER_0_929 ();
 sg13g2_decap_8 FILLER_0_936 ();
 sg13g2_decap_4 FILLER_0_943 ();
 sg13g2_fill_2 FILLER_0_977 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_8 FILLER_0_999 ();
 sg13g2_decap_8 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1013 ();
 sg13g2_decap_8 FILLER_0_1020 ();
 sg13g2_decap_8 FILLER_0_1027 ();
 sg13g2_decap_8 FILLER_0_1034 ();
 sg13g2_decap_8 FILLER_0_1041 ();
 sg13g2_decap_8 FILLER_0_1048 ();
 sg13g2_decap_8 FILLER_0_1055 ();
 sg13g2_decap_8 FILLER_0_1062 ();
 sg13g2_decap_8 FILLER_0_1069 ();
 sg13g2_decap_8 FILLER_0_1076 ();
 sg13g2_decap_8 FILLER_0_1083 ();
 sg13g2_decap_8 FILLER_0_1090 ();
 sg13g2_decap_8 FILLER_0_1097 ();
 sg13g2_decap_8 FILLER_0_1104 ();
 sg13g2_decap_8 FILLER_0_1111 ();
 sg13g2_decap_8 FILLER_0_1118 ();
 sg13g2_decap_8 FILLER_0_1125 ();
 sg13g2_decap_8 FILLER_0_1132 ();
 sg13g2_decap_8 FILLER_0_1139 ();
 sg13g2_decap_8 FILLER_0_1146 ();
 sg13g2_decap_8 FILLER_0_1153 ();
 sg13g2_decap_8 FILLER_0_1160 ();
 sg13g2_decap_8 FILLER_0_1167 ();
 sg13g2_decap_8 FILLER_0_1174 ();
 sg13g2_decap_8 FILLER_0_1181 ();
 sg13g2_decap_8 FILLER_0_1188 ();
 sg13g2_decap_8 FILLER_0_1195 ();
 sg13g2_decap_8 FILLER_0_1202 ();
 sg13g2_decap_8 FILLER_0_1209 ();
 sg13g2_decap_8 FILLER_0_1216 ();
 sg13g2_decap_8 FILLER_0_1223 ();
 sg13g2_decap_8 FILLER_0_1230 ();
 sg13g2_decap_8 FILLER_0_1237 ();
 sg13g2_decap_8 FILLER_0_1244 ();
 sg13g2_decap_8 FILLER_0_1251 ();
 sg13g2_decap_8 FILLER_0_1258 ();
 sg13g2_decap_8 FILLER_0_1265 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_8 FILLER_0_1286 ();
 sg13g2_decap_8 FILLER_0_1293 ();
 sg13g2_decap_8 FILLER_0_1300 ();
 sg13g2_decap_8 FILLER_0_1307 ();
 sg13g2_decap_8 FILLER_0_1314 ();
 sg13g2_decap_4 FILLER_0_1321 ();
 sg13g2_fill_1 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_4 FILLER_1_238 ();
 sg13g2_fill_2 FILLER_1_242 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_fill_2 FILLER_1_297 ();
 sg13g2_fill_1 FILLER_1_299 ();
 sg13g2_decap_4 FILLER_1_309 ();
 sg13g2_fill_1 FILLER_1_313 ();
 sg13g2_fill_2 FILLER_1_335 ();
 sg13g2_fill_1 FILLER_1_346 ();
 sg13g2_fill_1 FILLER_1_351 ();
 sg13g2_fill_1 FILLER_1_356 ();
 sg13g2_fill_1 FILLER_1_361 ();
 sg13g2_fill_1 FILLER_1_380 ();
 sg13g2_fill_1 FILLER_1_398 ();
 sg13g2_fill_2 FILLER_1_403 ();
 sg13g2_fill_1 FILLER_1_434 ();
 sg13g2_fill_2 FILLER_1_440 ();
 sg13g2_fill_2 FILLER_1_447 ();
 sg13g2_fill_1 FILLER_1_474 ();
 sg13g2_fill_2 FILLER_1_501 ();
 sg13g2_decap_8 FILLER_1_555 ();
 sg13g2_decap_8 FILLER_1_562 ();
 sg13g2_decap_8 FILLER_1_569 ();
 sg13g2_decap_8 FILLER_1_576 ();
 sg13g2_decap_8 FILLER_1_583 ();
 sg13g2_decap_8 FILLER_1_590 ();
 sg13g2_fill_2 FILLER_1_597 ();
 sg13g2_fill_1 FILLER_1_599 ();
 sg13g2_decap_8 FILLER_1_604 ();
 sg13g2_fill_2 FILLER_1_611 ();
 sg13g2_fill_1 FILLER_1_613 ();
 sg13g2_fill_2 FILLER_1_619 ();
 sg13g2_fill_1 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_decap_8 FILLER_1_685 ();
 sg13g2_decap_8 FILLER_1_692 ();
 sg13g2_decap_8 FILLER_1_699 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_4 FILLER_1_720 ();
 sg13g2_fill_2 FILLER_1_724 ();
 sg13g2_decap_8 FILLER_1_731 ();
 sg13g2_fill_2 FILLER_1_738 ();
 sg13g2_fill_1 FILLER_1_740 ();
 sg13g2_fill_2 FILLER_1_753 ();
 sg13g2_fill_2 FILLER_1_759 ();
 sg13g2_fill_1 FILLER_1_769 ();
 sg13g2_decap_4 FILLER_1_774 ();
 sg13g2_fill_2 FILLER_1_778 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_4 FILLER_1_805 ();
 sg13g2_fill_2 FILLER_1_809 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_4 FILLER_1_826 ();
 sg13g2_fill_2 FILLER_1_830 ();
 sg13g2_fill_2 FILLER_1_841 ();
 sg13g2_fill_2 FILLER_1_847 ();
 sg13g2_fill_2 FILLER_1_859 ();
 sg13g2_fill_1 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_901 ();
 sg13g2_fill_2 FILLER_1_908 ();
 sg13g2_decap_8 FILLER_1_936 ();
 sg13g2_fill_2 FILLER_1_943 ();
 sg13g2_fill_1 FILLER_1_945 ();
 sg13g2_fill_2 FILLER_1_951 ();
 sg13g2_decap_4 FILLER_1_961 ();
 sg13g2_fill_2 FILLER_1_965 ();
 sg13g2_fill_2 FILLER_1_993 ();
 sg13g2_fill_1 FILLER_1_995 ();
 sg13g2_decap_8 FILLER_1_1026 ();
 sg13g2_decap_8 FILLER_1_1033 ();
 sg13g2_decap_4 FILLER_1_1040 ();
 sg13g2_fill_1 FILLER_1_1044 ();
 sg13g2_decap_8 FILLER_1_1049 ();
 sg13g2_decap_8 FILLER_1_1056 ();
 sg13g2_decap_8 FILLER_1_1063 ();
 sg13g2_decap_8 FILLER_1_1070 ();
 sg13g2_decap_8 FILLER_1_1077 ();
 sg13g2_decap_8 FILLER_1_1084 ();
 sg13g2_decap_8 FILLER_1_1091 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_decap_8 FILLER_1_1119 ();
 sg13g2_decap_8 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1133 ();
 sg13g2_decap_8 FILLER_1_1140 ();
 sg13g2_decap_8 FILLER_1_1147 ();
 sg13g2_decap_8 FILLER_1_1154 ();
 sg13g2_decap_8 FILLER_1_1161 ();
 sg13g2_decap_8 FILLER_1_1168 ();
 sg13g2_decap_8 FILLER_1_1175 ();
 sg13g2_decap_8 FILLER_1_1182 ();
 sg13g2_decap_8 FILLER_1_1189 ();
 sg13g2_decap_8 FILLER_1_1196 ();
 sg13g2_decap_8 FILLER_1_1203 ();
 sg13g2_decap_8 FILLER_1_1210 ();
 sg13g2_decap_8 FILLER_1_1217 ();
 sg13g2_decap_8 FILLER_1_1224 ();
 sg13g2_decap_8 FILLER_1_1231 ();
 sg13g2_decap_8 FILLER_1_1238 ();
 sg13g2_decap_8 FILLER_1_1245 ();
 sg13g2_decap_8 FILLER_1_1252 ();
 sg13g2_decap_8 FILLER_1_1259 ();
 sg13g2_decap_8 FILLER_1_1266 ();
 sg13g2_decap_8 FILLER_1_1273 ();
 sg13g2_decap_8 FILLER_1_1280 ();
 sg13g2_decap_8 FILLER_1_1287 ();
 sg13g2_decap_8 FILLER_1_1294 ();
 sg13g2_decap_8 FILLER_1_1301 ();
 sg13g2_decap_8 FILLER_1_1308 ();
 sg13g2_decap_8 FILLER_1_1315 ();
 sg13g2_decap_4 FILLER_1_1322 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_fill_2 FILLER_2_263 ();
 sg13g2_fill_2 FILLER_2_269 ();
 sg13g2_fill_1 FILLER_2_305 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_fill_1 FILLER_2_328 ();
 sg13g2_fill_2 FILLER_2_354 ();
 sg13g2_fill_1 FILLER_2_361 ();
 sg13g2_fill_2 FILLER_2_392 ();
 sg13g2_fill_2 FILLER_2_399 ();
 sg13g2_fill_1 FILLER_2_417 ();
 sg13g2_fill_2 FILLER_2_440 ();
 sg13g2_fill_1 FILLER_2_450 ();
 sg13g2_fill_1 FILLER_2_463 ();
 sg13g2_fill_1 FILLER_2_468 ();
 sg13g2_fill_1 FILLER_2_478 ();
 sg13g2_fill_1 FILLER_2_483 ();
 sg13g2_decap_4 FILLER_2_492 ();
 sg13g2_fill_1 FILLER_2_496 ();
 sg13g2_fill_1 FILLER_2_501 ();
 sg13g2_fill_2 FILLER_2_522 ();
 sg13g2_fill_1 FILLER_2_524 ();
 sg13g2_fill_2 FILLER_2_534 ();
 sg13g2_decap_4 FILLER_2_540 ();
 sg13g2_fill_2 FILLER_2_549 ();
 sg13g2_decap_8 FILLER_2_555 ();
 sg13g2_decap_4 FILLER_2_562 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_fill_1 FILLER_2_588 ();
 sg13g2_fill_2 FILLER_2_635 ();
 sg13g2_fill_1 FILLER_2_637 ();
 sg13g2_fill_1 FILLER_2_646 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_fill_2 FILLER_2_669 ();
 sg13g2_fill_1 FILLER_2_680 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_fill_2 FILLER_2_718 ();
 sg13g2_fill_1 FILLER_2_753 ();
 sg13g2_fill_1 FILLER_2_762 ();
 sg13g2_fill_1 FILLER_2_793 ();
 sg13g2_fill_2 FILLER_2_834 ();
 sg13g2_fill_1 FILLER_2_836 ();
 sg13g2_decap_4 FILLER_2_841 ();
 sg13g2_fill_1 FILLER_2_868 ();
 sg13g2_fill_1 FILLER_2_894 ();
 sg13g2_fill_2 FILLER_2_900 ();
 sg13g2_decap_4 FILLER_2_906 ();
 sg13g2_fill_2 FILLER_2_915 ();
 sg13g2_decap_4 FILLER_2_925 ();
 sg13g2_fill_2 FILLER_2_933 ();
 sg13g2_decap_4 FILLER_2_943 ();
 sg13g2_fill_1 FILLER_2_947 ();
 sg13g2_fill_2 FILLER_2_952 ();
 sg13g2_decap_4 FILLER_2_993 ();
 sg13g2_fill_1 FILLER_2_1002 ();
 sg13g2_fill_1 FILLER_2_1007 ();
 sg13g2_fill_1 FILLER_2_1013 ();
 sg13g2_fill_1 FILLER_2_1018 ();
 sg13g2_fill_2 FILLER_2_1023 ();
 sg13g2_fill_2 FILLER_2_1029 ();
 sg13g2_decap_8 FILLER_2_1061 ();
 sg13g2_decap_8 FILLER_2_1068 ();
 sg13g2_decap_8 FILLER_2_1075 ();
 sg13g2_decap_8 FILLER_2_1082 ();
 sg13g2_decap_8 FILLER_2_1089 ();
 sg13g2_decap_8 FILLER_2_1096 ();
 sg13g2_decap_8 FILLER_2_1103 ();
 sg13g2_decap_8 FILLER_2_1110 ();
 sg13g2_decap_8 FILLER_2_1117 ();
 sg13g2_decap_8 FILLER_2_1124 ();
 sg13g2_decap_8 FILLER_2_1131 ();
 sg13g2_decap_8 FILLER_2_1138 ();
 sg13g2_decap_8 FILLER_2_1145 ();
 sg13g2_decap_8 FILLER_2_1152 ();
 sg13g2_decap_8 FILLER_2_1159 ();
 sg13g2_decap_8 FILLER_2_1166 ();
 sg13g2_decap_8 FILLER_2_1173 ();
 sg13g2_decap_8 FILLER_2_1180 ();
 sg13g2_decap_8 FILLER_2_1187 ();
 sg13g2_decap_8 FILLER_2_1194 ();
 sg13g2_decap_8 FILLER_2_1201 ();
 sg13g2_decap_8 FILLER_2_1208 ();
 sg13g2_decap_8 FILLER_2_1215 ();
 sg13g2_decap_8 FILLER_2_1222 ();
 sg13g2_decap_8 FILLER_2_1229 ();
 sg13g2_decap_8 FILLER_2_1236 ();
 sg13g2_decap_8 FILLER_2_1243 ();
 sg13g2_decap_8 FILLER_2_1250 ();
 sg13g2_decap_8 FILLER_2_1257 ();
 sg13g2_decap_8 FILLER_2_1264 ();
 sg13g2_decap_8 FILLER_2_1271 ();
 sg13g2_decap_8 FILLER_2_1278 ();
 sg13g2_decap_8 FILLER_2_1285 ();
 sg13g2_decap_8 FILLER_2_1292 ();
 sg13g2_decap_8 FILLER_2_1299 ();
 sg13g2_decap_8 FILLER_2_1306 ();
 sg13g2_decap_8 FILLER_2_1313 ();
 sg13g2_decap_4 FILLER_2_1320 ();
 sg13g2_fill_2 FILLER_2_1324 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_4 FILLER_3_231 ();
 sg13g2_fill_2 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_decap_4 FILLER_3_315 ();
 sg13g2_fill_2 FILLER_3_319 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_decap_4 FILLER_3_354 ();
 sg13g2_fill_2 FILLER_3_358 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_377 ();
 sg13g2_fill_1 FILLER_3_418 ();
 sg13g2_fill_1 FILLER_3_461 ();
 sg13g2_fill_1 FILLER_3_466 ();
 sg13g2_fill_1 FILLER_3_472 ();
 sg13g2_fill_2 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_549 ();
 sg13g2_fill_1 FILLER_3_577 ();
 sg13g2_fill_1 FILLER_3_582 ();
 sg13g2_fill_1 FILLER_3_603 ();
 sg13g2_fill_2 FILLER_3_608 ();
 sg13g2_fill_1 FILLER_3_642 ();
 sg13g2_fill_2 FILLER_3_652 ();
 sg13g2_fill_1 FILLER_3_654 ();
 sg13g2_decap_4 FILLER_3_662 ();
 sg13g2_fill_1 FILLER_3_666 ();
 sg13g2_fill_1 FILLER_3_675 ();
 sg13g2_fill_1 FILLER_3_684 ();
 sg13g2_fill_2 FILLER_3_697 ();
 sg13g2_fill_2 FILLER_3_703 ();
 sg13g2_fill_1 FILLER_3_740 ();
 sg13g2_decap_8 FILLER_3_839 ();
 sg13g2_fill_2 FILLER_3_846 ();
 sg13g2_fill_1 FILLER_3_848 ();
 sg13g2_fill_1 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_860 ();
 sg13g2_decap_4 FILLER_3_878 ();
 sg13g2_fill_1 FILLER_3_882 ();
 sg13g2_fill_2 FILLER_3_887 ();
 sg13g2_fill_1 FILLER_3_905 ();
 sg13g2_fill_2 FILLER_3_941 ();
 sg13g2_decap_4 FILLER_3_952 ();
 sg13g2_fill_1 FILLER_3_960 ();
 sg13g2_fill_1 FILLER_3_992 ();
 sg13g2_fill_2 FILLER_3_1001 ();
 sg13g2_fill_2 FILLER_3_1007 ();
 sg13g2_fill_2 FILLER_3_1048 ();
 sg13g2_fill_1 FILLER_3_1060 ();
 sg13g2_decap_8 FILLER_3_1091 ();
 sg13g2_decap_8 FILLER_3_1098 ();
 sg13g2_decap_8 FILLER_3_1105 ();
 sg13g2_decap_8 FILLER_3_1112 ();
 sg13g2_decap_8 FILLER_3_1119 ();
 sg13g2_decap_8 FILLER_3_1126 ();
 sg13g2_decap_8 FILLER_3_1133 ();
 sg13g2_decap_8 FILLER_3_1140 ();
 sg13g2_decap_8 FILLER_3_1147 ();
 sg13g2_decap_8 FILLER_3_1154 ();
 sg13g2_decap_8 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1168 ();
 sg13g2_decap_8 FILLER_3_1175 ();
 sg13g2_decap_8 FILLER_3_1182 ();
 sg13g2_decap_8 FILLER_3_1189 ();
 sg13g2_decap_8 FILLER_3_1196 ();
 sg13g2_decap_8 FILLER_3_1203 ();
 sg13g2_decap_8 FILLER_3_1210 ();
 sg13g2_decap_8 FILLER_3_1217 ();
 sg13g2_decap_8 FILLER_3_1224 ();
 sg13g2_decap_8 FILLER_3_1231 ();
 sg13g2_decap_8 FILLER_3_1238 ();
 sg13g2_decap_8 FILLER_3_1245 ();
 sg13g2_decap_8 FILLER_3_1252 ();
 sg13g2_decap_8 FILLER_3_1259 ();
 sg13g2_decap_8 FILLER_3_1266 ();
 sg13g2_decap_8 FILLER_3_1273 ();
 sg13g2_decap_8 FILLER_3_1280 ();
 sg13g2_decap_8 FILLER_3_1287 ();
 sg13g2_decap_8 FILLER_3_1294 ();
 sg13g2_decap_8 FILLER_3_1301 ();
 sg13g2_decap_8 FILLER_3_1308 ();
 sg13g2_decap_8 FILLER_3_1315 ();
 sg13g2_decap_4 FILLER_3_1322 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_197 ();
 sg13g2_decap_8 FILLER_4_204 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_decap_8 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_fill_2 FILLER_4_232 ();
 sg13g2_fill_1 FILLER_4_274 ();
 sg13g2_fill_1 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_344 ();
 sg13g2_fill_2 FILLER_4_393 ();
 sg13g2_fill_1 FILLER_4_399 ();
 sg13g2_fill_1 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_fill_1 FILLER_4_441 ();
 sg13g2_fill_2 FILLER_4_458 ();
 sg13g2_fill_2 FILLER_4_495 ();
 sg13g2_fill_1 FILLER_4_497 ();
 sg13g2_fill_1 FILLER_4_528 ();
 sg13g2_fill_1 FILLER_4_534 ();
 sg13g2_fill_2 FILLER_4_538 ();
 sg13g2_fill_1 FILLER_4_546 ();
 sg13g2_fill_1 FILLER_4_551 ();
 sg13g2_fill_2 FILLER_4_557 ();
 sg13g2_fill_2 FILLER_4_563 ();
 sg13g2_fill_2 FILLER_4_599 ();
 sg13g2_fill_1 FILLER_4_612 ();
 sg13g2_fill_1 FILLER_4_621 ();
 sg13g2_fill_1 FILLER_4_625 ();
 sg13g2_fill_1 FILLER_4_637 ();
 sg13g2_fill_2 FILLER_4_656 ();
 sg13g2_fill_1 FILLER_4_668 ();
 sg13g2_fill_1 FILLER_4_673 ();
 sg13g2_fill_1 FILLER_4_678 ();
 sg13g2_fill_1 FILLER_4_687 ();
 sg13g2_fill_1 FILLER_4_714 ();
 sg13g2_fill_2 FILLER_4_719 ();
 sg13g2_decap_8 FILLER_4_733 ();
 sg13g2_fill_2 FILLER_4_748 ();
 sg13g2_fill_2 FILLER_4_787 ();
 sg13g2_fill_1 FILLER_4_793 ();
 sg13g2_fill_2 FILLER_4_797 ();
 sg13g2_fill_1 FILLER_4_803 ();
 sg13g2_fill_2 FILLER_4_814 ();
 sg13g2_decap_8 FILLER_4_820 ();
 sg13g2_fill_1 FILLER_4_827 ();
 sg13g2_fill_1 FILLER_4_833 ();
 sg13g2_fill_1 FILLER_4_839 ();
 sg13g2_fill_1 FILLER_4_844 ();
 sg13g2_fill_2 FILLER_4_849 ();
 sg13g2_fill_2 FILLER_4_855 ();
 sg13g2_fill_2 FILLER_4_865 ();
 sg13g2_decap_4 FILLER_4_907 ();
 sg13g2_decap_4 FILLER_4_916 ();
 sg13g2_fill_1 FILLER_4_925 ();
 sg13g2_fill_2 FILLER_4_930 ();
 sg13g2_fill_1 FILLER_4_932 ();
 sg13g2_fill_1 FILLER_4_979 ();
 sg13g2_decap_4 FILLER_4_994 ();
 sg13g2_fill_2 FILLER_4_998 ();
 sg13g2_fill_1 FILLER_4_1004 ();
 sg13g2_fill_1 FILLER_4_1010 ();
 sg13g2_fill_2 FILLER_4_1015 ();
 sg13g2_fill_1 FILLER_4_1017 ();
 sg13g2_fill_2 FILLER_4_1030 ();
 sg13g2_fill_1 FILLER_4_1032 ();
 sg13g2_fill_1 FILLER_4_1046 ();
 sg13g2_fill_1 FILLER_4_1071 ();
 sg13g2_decap_8 FILLER_4_1079 ();
 sg13g2_decap_8 FILLER_4_1086 ();
 sg13g2_decap_8 FILLER_4_1093 ();
 sg13g2_decap_8 FILLER_4_1100 ();
 sg13g2_decap_8 FILLER_4_1107 ();
 sg13g2_decap_8 FILLER_4_1114 ();
 sg13g2_decap_8 FILLER_4_1121 ();
 sg13g2_decap_8 FILLER_4_1128 ();
 sg13g2_decap_8 FILLER_4_1135 ();
 sg13g2_decap_8 FILLER_4_1142 ();
 sg13g2_decap_8 FILLER_4_1149 ();
 sg13g2_decap_8 FILLER_4_1156 ();
 sg13g2_decap_8 FILLER_4_1163 ();
 sg13g2_decap_8 FILLER_4_1170 ();
 sg13g2_decap_8 FILLER_4_1177 ();
 sg13g2_decap_8 FILLER_4_1184 ();
 sg13g2_decap_8 FILLER_4_1191 ();
 sg13g2_decap_8 FILLER_4_1198 ();
 sg13g2_decap_8 FILLER_4_1205 ();
 sg13g2_decap_8 FILLER_4_1212 ();
 sg13g2_decap_8 FILLER_4_1219 ();
 sg13g2_decap_8 FILLER_4_1226 ();
 sg13g2_decap_8 FILLER_4_1233 ();
 sg13g2_decap_8 FILLER_4_1240 ();
 sg13g2_decap_8 FILLER_4_1247 ();
 sg13g2_decap_8 FILLER_4_1254 ();
 sg13g2_decap_8 FILLER_4_1261 ();
 sg13g2_decap_8 FILLER_4_1268 ();
 sg13g2_decap_8 FILLER_4_1275 ();
 sg13g2_decap_8 FILLER_4_1282 ();
 sg13g2_decap_8 FILLER_4_1289 ();
 sg13g2_decap_8 FILLER_4_1296 ();
 sg13g2_decap_8 FILLER_4_1303 ();
 sg13g2_decap_8 FILLER_4_1310 ();
 sg13g2_decap_8 FILLER_4_1317 ();
 sg13g2_fill_2 FILLER_4_1324 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_226 ();
 sg13g2_fill_2 FILLER_5_233 ();
 sg13g2_fill_1 FILLER_5_235 ();
 sg13g2_fill_2 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_fill_1 FILLER_5_300 ();
 sg13g2_decap_4 FILLER_5_313 ();
 sg13g2_fill_2 FILLER_5_317 ();
 sg13g2_decap_4 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_fill_2 FILLER_5_348 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_fill_1 FILLER_5_441 ();
 sg13g2_fill_1 FILLER_5_446 ();
 sg13g2_fill_1 FILLER_5_455 ();
 sg13g2_fill_2 FILLER_5_459 ();
 sg13g2_fill_1 FILLER_5_465 ();
 sg13g2_fill_1 FILLER_5_471 ();
 sg13g2_fill_1 FILLER_5_476 ();
 sg13g2_fill_1 FILLER_5_503 ();
 sg13g2_fill_2 FILLER_5_518 ();
 sg13g2_fill_1 FILLER_5_520 ();
 sg13g2_decap_4 FILLER_5_533 ();
 sg13g2_fill_1 FILLER_5_577 ();
 sg13g2_decap_8 FILLER_5_582 ();
 sg13g2_fill_2 FILLER_5_595 ();
 sg13g2_fill_2 FILLER_5_635 ();
 sg13g2_fill_1 FILLER_5_642 ();
 sg13g2_fill_1 FILLER_5_647 ();
 sg13g2_fill_2 FILLER_5_673 ();
 sg13g2_fill_1 FILLER_5_687 ();
 sg13g2_fill_1 FILLER_5_692 ();
 sg13g2_fill_1 FILLER_5_722 ();
 sg13g2_fill_2 FILLER_5_749 ();
 sg13g2_fill_1 FILLER_5_773 ();
 sg13g2_fill_2 FILLER_5_860 ();
 sg13g2_fill_1 FILLER_5_862 ();
 sg13g2_fill_1 FILLER_5_891 ();
 sg13g2_fill_1 FILLER_5_896 ();
 sg13g2_fill_1 FILLER_5_900 ();
 sg13g2_fill_1 FILLER_5_909 ();
 sg13g2_decap_8 FILLER_5_953 ();
 sg13g2_fill_1 FILLER_5_960 ();
 sg13g2_fill_2 FILLER_5_964 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_fill_2 FILLER_5_977 ();
 sg13g2_decap_4 FILLER_5_996 ();
 sg13g2_fill_2 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1063 ();
 sg13g2_decap_8 FILLER_5_1070 ();
 sg13g2_decap_8 FILLER_5_1077 ();
 sg13g2_decap_8 FILLER_5_1084 ();
 sg13g2_decap_8 FILLER_5_1091 ();
 sg13g2_decap_8 FILLER_5_1098 ();
 sg13g2_decap_8 FILLER_5_1105 ();
 sg13g2_decap_8 FILLER_5_1112 ();
 sg13g2_decap_8 FILLER_5_1119 ();
 sg13g2_decap_8 FILLER_5_1126 ();
 sg13g2_decap_8 FILLER_5_1133 ();
 sg13g2_decap_8 FILLER_5_1140 ();
 sg13g2_decap_8 FILLER_5_1147 ();
 sg13g2_decap_8 FILLER_5_1154 ();
 sg13g2_decap_8 FILLER_5_1161 ();
 sg13g2_decap_8 FILLER_5_1168 ();
 sg13g2_decap_8 FILLER_5_1175 ();
 sg13g2_decap_8 FILLER_5_1182 ();
 sg13g2_decap_8 FILLER_5_1189 ();
 sg13g2_decap_8 FILLER_5_1196 ();
 sg13g2_decap_8 FILLER_5_1203 ();
 sg13g2_decap_8 FILLER_5_1210 ();
 sg13g2_decap_8 FILLER_5_1217 ();
 sg13g2_decap_8 FILLER_5_1224 ();
 sg13g2_decap_8 FILLER_5_1231 ();
 sg13g2_decap_8 FILLER_5_1238 ();
 sg13g2_decap_8 FILLER_5_1245 ();
 sg13g2_decap_8 FILLER_5_1252 ();
 sg13g2_decap_8 FILLER_5_1259 ();
 sg13g2_decap_8 FILLER_5_1266 ();
 sg13g2_decap_8 FILLER_5_1273 ();
 sg13g2_decap_8 FILLER_5_1280 ();
 sg13g2_decap_8 FILLER_5_1287 ();
 sg13g2_decap_8 FILLER_5_1294 ();
 sg13g2_decap_8 FILLER_5_1301 ();
 sg13g2_decap_8 FILLER_5_1308 ();
 sg13g2_decap_8 FILLER_5_1315 ();
 sg13g2_decap_4 FILLER_5_1322 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_161 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_decap_4 FILLER_6_190 ();
 sg13g2_decap_8 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_248 ();
 sg13g2_fill_1 FILLER_6_250 ();
 sg13g2_fill_1 FILLER_6_255 ();
 sg13g2_fill_1 FILLER_6_282 ();
 sg13g2_fill_1 FILLER_6_287 ();
 sg13g2_fill_2 FILLER_6_293 ();
 sg13g2_fill_1 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_fill_2 FILLER_6_335 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_fill_1 FILLER_6_384 ();
 sg13g2_fill_1 FILLER_6_390 ();
 sg13g2_fill_2 FILLER_6_395 ();
 sg13g2_fill_2 FILLER_6_402 ();
 sg13g2_fill_2 FILLER_6_408 ();
 sg13g2_fill_1 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_446 ();
 sg13g2_fill_1 FILLER_6_451 ();
 sg13g2_fill_1 FILLER_6_533 ();
 sg13g2_fill_1 FILLER_6_543 ();
 sg13g2_decap_4 FILLER_6_553 ();
 sg13g2_fill_2 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_563 ();
 sg13g2_fill_2 FILLER_6_570 ();
 sg13g2_fill_1 FILLER_6_572 ();
 sg13g2_decap_8 FILLER_6_577 ();
 sg13g2_decap_4 FILLER_6_584 ();
 sg13g2_fill_2 FILLER_6_588 ();
 sg13g2_fill_2 FILLER_6_618 ();
 sg13g2_fill_1 FILLER_6_620 ();
 sg13g2_decap_4 FILLER_6_659 ();
 sg13g2_fill_1 FILLER_6_667 ();
 sg13g2_fill_1 FILLER_6_672 ();
 sg13g2_fill_2 FILLER_6_678 ();
 sg13g2_fill_2 FILLER_6_684 ();
 sg13g2_fill_2 FILLER_6_689 ();
 sg13g2_fill_1 FILLER_6_713 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_733 ();
 sg13g2_decap_4 FILLER_6_740 ();
 sg13g2_fill_1 FILLER_6_744 ();
 sg13g2_decap_8 FILLER_6_750 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_4 FILLER_6_822 ();
 sg13g2_fill_2 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_863 ();
 sg13g2_fill_1 FILLER_6_883 ();
 sg13g2_fill_1 FILLER_6_892 ();
 sg13g2_fill_1 FILLER_6_901 ();
 sg13g2_fill_1 FILLER_6_907 ();
 sg13g2_fill_1 FILLER_6_911 ();
 sg13g2_fill_2 FILLER_6_920 ();
 sg13g2_decap_4 FILLER_6_942 ();
 sg13g2_fill_1 FILLER_6_983 ();
 sg13g2_decap_8 FILLER_6_1023 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_fill_2 FILLER_6_1037 ();
 sg13g2_fill_1 FILLER_6_1039 ();
 sg13g2_decap_4 FILLER_6_1052 ();
 sg13g2_fill_1 FILLER_6_1061 ();
 sg13g2_decap_8 FILLER_6_1073 ();
 sg13g2_decap_8 FILLER_6_1080 ();
 sg13g2_decap_8 FILLER_6_1087 ();
 sg13g2_decap_8 FILLER_6_1094 ();
 sg13g2_decap_8 FILLER_6_1101 ();
 sg13g2_decap_8 FILLER_6_1108 ();
 sg13g2_decap_8 FILLER_6_1115 ();
 sg13g2_decap_8 FILLER_6_1122 ();
 sg13g2_decap_8 FILLER_6_1129 ();
 sg13g2_decap_8 FILLER_6_1136 ();
 sg13g2_decap_8 FILLER_6_1143 ();
 sg13g2_decap_8 FILLER_6_1150 ();
 sg13g2_decap_8 FILLER_6_1157 ();
 sg13g2_decap_8 FILLER_6_1164 ();
 sg13g2_decap_8 FILLER_6_1171 ();
 sg13g2_decap_8 FILLER_6_1178 ();
 sg13g2_decap_8 FILLER_6_1185 ();
 sg13g2_decap_8 FILLER_6_1192 ();
 sg13g2_decap_8 FILLER_6_1199 ();
 sg13g2_decap_8 FILLER_6_1206 ();
 sg13g2_decap_8 FILLER_6_1213 ();
 sg13g2_decap_8 FILLER_6_1220 ();
 sg13g2_decap_8 FILLER_6_1227 ();
 sg13g2_decap_8 FILLER_6_1234 ();
 sg13g2_decap_8 FILLER_6_1241 ();
 sg13g2_decap_8 FILLER_6_1248 ();
 sg13g2_decap_8 FILLER_6_1255 ();
 sg13g2_decap_8 FILLER_6_1262 ();
 sg13g2_decap_8 FILLER_6_1269 ();
 sg13g2_decap_8 FILLER_6_1276 ();
 sg13g2_decap_8 FILLER_6_1283 ();
 sg13g2_decap_8 FILLER_6_1290 ();
 sg13g2_decap_8 FILLER_6_1297 ();
 sg13g2_decap_8 FILLER_6_1304 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1318 ();
 sg13g2_fill_1 FILLER_6_1325 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_4 FILLER_7_56 ();
 sg13g2_fill_1 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_208 ();
 sg13g2_fill_2 FILLER_7_222 ();
 sg13g2_fill_2 FILLER_7_310 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_326 ();
 sg13g2_decap_4 FILLER_7_332 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_decap_4 FILLER_7_341 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_fill_1 FILLER_7_352 ();
 sg13g2_fill_1 FILLER_7_357 ();
 sg13g2_fill_1 FILLER_7_363 ();
 sg13g2_fill_1 FILLER_7_390 ();
 sg13g2_fill_1 FILLER_7_417 ();
 sg13g2_fill_1 FILLER_7_449 ();
 sg13g2_fill_1 FILLER_7_453 ();
 sg13g2_fill_1 FILLER_7_458 ();
 sg13g2_fill_1 FILLER_7_464 ();
 sg13g2_fill_2 FILLER_7_504 ();
 sg13g2_fill_1 FILLER_7_519 ();
 sg13g2_fill_2 FILLER_7_528 ();
 sg13g2_fill_1 FILLER_7_535 ();
 sg13g2_fill_2 FILLER_7_597 ();
 sg13g2_decap_4 FILLER_7_604 ();
 sg13g2_fill_1 FILLER_7_608 ();
 sg13g2_decap_8 FILLER_7_613 ();
 sg13g2_decap_4 FILLER_7_620 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_decap_4 FILLER_7_629 ();
 sg13g2_fill_2 FILLER_7_633 ();
 sg13g2_fill_1 FILLER_7_639 ();
 sg13g2_fill_2 FILLER_7_645 ();
 sg13g2_fill_1 FILLER_7_655 ();
 sg13g2_fill_1 FILLER_7_682 ();
 sg13g2_fill_2 FILLER_7_698 ();
 sg13g2_fill_2 FILLER_7_711 ();
 sg13g2_fill_1 FILLER_7_713 ();
 sg13g2_fill_1 FILLER_7_756 ();
 sg13g2_fill_1 FILLER_7_778 ();
 sg13g2_fill_2 FILLER_7_844 ();
 sg13g2_decap_8 FILLER_7_850 ();
 sg13g2_fill_2 FILLER_7_857 ();
 sg13g2_fill_1 FILLER_7_862 ();
 sg13g2_fill_1 FILLER_7_868 ();
 sg13g2_fill_1 FILLER_7_873 ();
 sg13g2_fill_1 FILLER_7_881 ();
 sg13g2_fill_1 FILLER_7_885 ();
 sg13g2_fill_1 FILLER_7_890 ();
 sg13g2_fill_1 FILLER_7_895 ();
 sg13g2_fill_1 FILLER_7_904 ();
 sg13g2_fill_1 FILLER_7_910 ();
 sg13g2_fill_1 FILLER_7_915 ();
 sg13g2_fill_2 FILLER_7_920 ();
 sg13g2_fill_1 FILLER_7_922 ();
 sg13g2_fill_1 FILLER_7_954 ();
 sg13g2_fill_1 FILLER_7_959 ();
 sg13g2_fill_1 FILLER_7_972 ();
 sg13g2_fill_2 FILLER_7_977 ();
 sg13g2_fill_2 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_7_1085 ();
 sg13g2_decap_8 FILLER_7_1092 ();
 sg13g2_decap_8 FILLER_7_1099 ();
 sg13g2_decap_8 FILLER_7_1106 ();
 sg13g2_decap_8 FILLER_7_1113 ();
 sg13g2_decap_8 FILLER_7_1120 ();
 sg13g2_decap_8 FILLER_7_1127 ();
 sg13g2_decap_8 FILLER_7_1134 ();
 sg13g2_decap_8 FILLER_7_1141 ();
 sg13g2_decap_8 FILLER_7_1148 ();
 sg13g2_decap_8 FILLER_7_1155 ();
 sg13g2_decap_8 FILLER_7_1162 ();
 sg13g2_decap_8 FILLER_7_1169 ();
 sg13g2_decap_8 FILLER_7_1176 ();
 sg13g2_decap_8 FILLER_7_1183 ();
 sg13g2_decap_8 FILLER_7_1190 ();
 sg13g2_decap_8 FILLER_7_1197 ();
 sg13g2_decap_8 FILLER_7_1204 ();
 sg13g2_decap_8 FILLER_7_1211 ();
 sg13g2_decap_8 FILLER_7_1218 ();
 sg13g2_decap_8 FILLER_7_1225 ();
 sg13g2_decap_8 FILLER_7_1232 ();
 sg13g2_decap_8 FILLER_7_1239 ();
 sg13g2_decap_8 FILLER_7_1246 ();
 sg13g2_decap_8 FILLER_7_1253 ();
 sg13g2_decap_8 FILLER_7_1260 ();
 sg13g2_decap_8 FILLER_7_1267 ();
 sg13g2_decap_8 FILLER_7_1274 ();
 sg13g2_decap_8 FILLER_7_1281 ();
 sg13g2_decap_8 FILLER_7_1288 ();
 sg13g2_decap_8 FILLER_7_1295 ();
 sg13g2_decap_8 FILLER_7_1302 ();
 sg13g2_decap_8 FILLER_7_1309 ();
 sg13g2_decap_8 FILLER_7_1316 ();
 sg13g2_fill_2 FILLER_7_1323 ();
 sg13g2_fill_1 FILLER_7_1325 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_decap_4 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_140 ();
 sg13g2_fill_1 FILLER_8_159 ();
 sg13g2_fill_1 FILLER_8_172 ();
 sg13g2_fill_1 FILLER_8_177 ();
 sg13g2_fill_1 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_194 ();
 sg13g2_fill_2 FILLER_8_199 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_fill_2 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_1 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_294 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_410 ();
 sg13g2_decap_4 FILLER_8_446 ();
 sg13g2_fill_1 FILLER_8_450 ();
 sg13g2_fill_1 FILLER_8_474 ();
 sg13g2_fill_2 FILLER_8_501 ();
 sg13g2_fill_2 FILLER_8_508 ();
 sg13g2_fill_1 FILLER_8_545 ();
 sg13g2_fill_2 FILLER_8_577 ();
 sg13g2_fill_2 FILLER_8_605 ();
 sg13g2_fill_1 FILLER_8_607 ();
 sg13g2_decap_4 FILLER_8_612 ();
 sg13g2_fill_1 FILLER_8_689 ();
 sg13g2_fill_1 FILLER_8_715 ();
 sg13g2_fill_2 FILLER_8_744 ();
 sg13g2_decap_4 FILLER_8_786 ();
 sg13g2_decap_4 FILLER_8_794 ();
 sg13g2_decap_4 FILLER_8_812 ();
 sg13g2_fill_1 FILLER_8_824 ();
 sg13g2_fill_2 FILLER_8_866 ();
 sg13g2_fill_1 FILLER_8_868 ();
 sg13g2_fill_1 FILLER_8_911 ();
 sg13g2_fill_2 FILLER_8_951 ();
 sg13g2_fill_1 FILLER_8_958 ();
 sg13g2_fill_1 FILLER_8_1006 ();
 sg13g2_fill_2 FILLER_8_1012 ();
 sg13g2_fill_1 FILLER_8_1018 ();
 sg13g2_fill_2 FILLER_8_1023 ();
 sg13g2_fill_2 FILLER_8_1029 ();
 sg13g2_fill_1 FILLER_8_1048 ();
 sg13g2_fill_1 FILLER_8_1053 ();
 sg13g2_fill_1 FILLER_8_1061 ();
 sg13g2_decap_8 FILLER_8_1078 ();
 sg13g2_decap_8 FILLER_8_1085 ();
 sg13g2_decap_8 FILLER_8_1092 ();
 sg13g2_decap_8 FILLER_8_1099 ();
 sg13g2_decap_8 FILLER_8_1106 ();
 sg13g2_decap_8 FILLER_8_1113 ();
 sg13g2_decap_8 FILLER_8_1120 ();
 sg13g2_decap_8 FILLER_8_1127 ();
 sg13g2_decap_8 FILLER_8_1134 ();
 sg13g2_decap_8 FILLER_8_1141 ();
 sg13g2_decap_8 FILLER_8_1148 ();
 sg13g2_decap_8 FILLER_8_1155 ();
 sg13g2_decap_8 FILLER_8_1162 ();
 sg13g2_decap_8 FILLER_8_1169 ();
 sg13g2_decap_8 FILLER_8_1176 ();
 sg13g2_decap_8 FILLER_8_1183 ();
 sg13g2_decap_8 FILLER_8_1190 ();
 sg13g2_decap_8 FILLER_8_1197 ();
 sg13g2_decap_8 FILLER_8_1204 ();
 sg13g2_decap_8 FILLER_8_1211 ();
 sg13g2_decap_8 FILLER_8_1218 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_8 FILLER_8_1232 ();
 sg13g2_decap_8 FILLER_8_1239 ();
 sg13g2_decap_8 FILLER_8_1246 ();
 sg13g2_decap_8 FILLER_8_1253 ();
 sg13g2_decap_8 FILLER_8_1260 ();
 sg13g2_decap_8 FILLER_8_1267 ();
 sg13g2_decap_8 FILLER_8_1274 ();
 sg13g2_decap_8 FILLER_8_1281 ();
 sg13g2_decap_8 FILLER_8_1288 ();
 sg13g2_decap_8 FILLER_8_1295 ();
 sg13g2_decap_8 FILLER_8_1302 ();
 sg13g2_decap_8 FILLER_8_1309 ();
 sg13g2_decap_8 FILLER_8_1316 ();
 sg13g2_fill_2 FILLER_8_1323 ();
 sg13g2_fill_1 FILLER_8_1325 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_fill_1 FILLER_9_63 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_fill_1 FILLER_9_91 ();
 sg13g2_fill_2 FILLER_9_97 ();
 sg13g2_fill_1 FILLER_9_104 ();
 sg13g2_fill_1 FILLER_9_161 ();
 sg13g2_fill_1 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_197 ();
 sg13g2_fill_1 FILLER_9_205 ();
 sg13g2_fill_1 FILLER_9_210 ();
 sg13g2_fill_1 FILLER_9_216 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_fill_2 FILLER_9_240 ();
 sg13g2_fill_1 FILLER_9_322 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_342 ();
 sg13g2_fill_1 FILLER_9_356 ();
 sg13g2_fill_2 FILLER_9_422 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_9_434 ();
 sg13g2_fill_2 FILLER_9_439 ();
 sg13g2_fill_1 FILLER_9_454 ();
 sg13g2_fill_2 FILLER_9_468 ();
 sg13g2_fill_2 FILLER_9_492 ();
 sg13g2_fill_1 FILLER_9_499 ();
 sg13g2_fill_2 FILLER_9_519 ();
 sg13g2_fill_2 FILLER_9_529 ();
 sg13g2_fill_1 FILLER_9_531 ();
 sg13g2_fill_1 FILLER_9_542 ();
 sg13g2_fill_2 FILLER_9_551 ();
 sg13g2_fill_1 FILLER_9_553 ();
 sg13g2_decap_4 FILLER_9_629 ();
 sg13g2_fill_1 FILLER_9_633 ();
 sg13g2_fill_2 FILLER_9_638 ();
 sg13g2_fill_2 FILLER_9_649 ();
 sg13g2_decap_8 FILLER_9_663 ();
 sg13g2_fill_2 FILLER_9_670 ();
 sg13g2_fill_2 FILLER_9_676 ();
 sg13g2_fill_1 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_688 ();
 sg13g2_fill_2 FILLER_9_695 ();
 sg13g2_fill_2 FILLER_9_702 ();
 sg13g2_fill_2 FILLER_9_724 ();
 sg13g2_fill_2 FILLER_9_752 ();
 sg13g2_fill_1 FILLER_9_754 ();
 sg13g2_fill_1 FILLER_9_770 ();
 sg13g2_fill_2 FILLER_9_775 ();
 sg13g2_fill_2 FILLER_9_807 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_fill_2 FILLER_9_887 ();
 sg13g2_decap_4 FILLER_9_902 ();
 sg13g2_fill_1 FILLER_9_910 ();
 sg13g2_fill_2 FILLER_9_937 ();
 sg13g2_fill_1 FILLER_9_965 ();
 sg13g2_fill_2 FILLER_9_971 ();
 sg13g2_fill_1 FILLER_9_1032 ();
 sg13g2_fill_2 FILLER_9_1072 ();
 sg13g2_fill_1 FILLER_9_1074 ();
 sg13g2_decap_8 FILLER_9_1079 ();
 sg13g2_decap_8 FILLER_9_1086 ();
 sg13g2_decap_8 FILLER_9_1093 ();
 sg13g2_decap_8 FILLER_9_1100 ();
 sg13g2_decap_8 FILLER_9_1107 ();
 sg13g2_decap_8 FILLER_9_1114 ();
 sg13g2_decap_8 FILLER_9_1121 ();
 sg13g2_decap_8 FILLER_9_1128 ();
 sg13g2_decap_8 FILLER_9_1135 ();
 sg13g2_decap_8 FILLER_9_1142 ();
 sg13g2_decap_8 FILLER_9_1149 ();
 sg13g2_decap_8 FILLER_9_1156 ();
 sg13g2_decap_8 FILLER_9_1163 ();
 sg13g2_decap_8 FILLER_9_1170 ();
 sg13g2_decap_8 FILLER_9_1177 ();
 sg13g2_decap_8 FILLER_9_1184 ();
 sg13g2_decap_8 FILLER_9_1191 ();
 sg13g2_decap_8 FILLER_9_1198 ();
 sg13g2_decap_8 FILLER_9_1205 ();
 sg13g2_decap_8 FILLER_9_1212 ();
 sg13g2_decap_8 FILLER_9_1219 ();
 sg13g2_decap_8 FILLER_9_1226 ();
 sg13g2_decap_8 FILLER_9_1233 ();
 sg13g2_decap_8 FILLER_9_1240 ();
 sg13g2_decap_8 FILLER_9_1247 ();
 sg13g2_decap_8 FILLER_9_1254 ();
 sg13g2_decap_8 FILLER_9_1261 ();
 sg13g2_decap_8 FILLER_9_1268 ();
 sg13g2_decap_8 FILLER_9_1275 ();
 sg13g2_decap_8 FILLER_9_1282 ();
 sg13g2_decap_8 FILLER_9_1289 ();
 sg13g2_decap_8 FILLER_9_1296 ();
 sg13g2_decap_8 FILLER_9_1303 ();
 sg13g2_decap_8 FILLER_9_1310 ();
 sg13g2_decap_8 FILLER_9_1317 ();
 sg13g2_fill_2 FILLER_9_1324 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_56 ();
 sg13g2_fill_2 FILLER_10_60 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_76 ();
 sg13g2_fill_2 FILLER_10_95 ();
 sg13g2_fill_1 FILLER_10_114 ();
 sg13g2_fill_1 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_125 ();
 sg13g2_fill_2 FILLER_10_131 ();
 sg13g2_fill_1 FILLER_10_133 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_201 ();
 sg13g2_fill_2 FILLER_10_211 ();
 sg13g2_fill_2 FILLER_10_218 ();
 sg13g2_fill_2 FILLER_10_224 ();
 sg13g2_fill_2 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_271 ();
 sg13g2_fill_2 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_283 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_decap_4 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_2 FILLER_10_382 ();
 sg13g2_fill_1 FILLER_10_389 ();
 sg13g2_fill_1 FILLER_10_394 ();
 sg13g2_fill_2 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_405 ();
 sg13g2_fill_2 FILLER_10_411 ();
 sg13g2_fill_2 FILLER_10_421 ();
 sg13g2_fill_1 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_466 ();
 sg13g2_fill_1 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_572 ();
 sg13g2_fill_1 FILLER_10_581 ();
 sg13g2_fill_1 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_607 ();
 sg13g2_fill_1 FILLER_10_614 ();
 sg13g2_fill_1 FILLER_10_623 ();
 sg13g2_fill_2 FILLER_10_648 ();
 sg13g2_fill_1 FILLER_10_650 ();
 sg13g2_fill_2 FILLER_10_659 ();
 sg13g2_fill_1 FILLER_10_661 ();
 sg13g2_fill_1 FILLER_10_693 ();
 sg13g2_fill_2 FILLER_10_698 ();
 sg13g2_fill_2 FILLER_10_714 ();
 sg13g2_fill_2 FILLER_10_731 ();
 sg13g2_fill_1 FILLER_10_759 ();
 sg13g2_fill_2 FILLER_10_765 ();
 sg13g2_fill_1 FILLER_10_780 ();
 sg13g2_fill_1 FILLER_10_785 ();
 sg13g2_decap_4 FILLER_10_794 ();
 sg13g2_fill_1 FILLER_10_798 ();
 sg13g2_fill_2 FILLER_10_809 ();
 sg13g2_fill_1 FILLER_10_811 ();
 sg13g2_fill_2 FILLER_10_816 ();
 sg13g2_fill_1 FILLER_10_866 ();
 sg13g2_fill_1 FILLER_10_876 ();
 sg13g2_fill_1 FILLER_10_882 ();
 sg13g2_fill_1 FILLER_10_891 ();
 sg13g2_fill_2 FILLER_10_904 ();
 sg13g2_fill_2 FILLER_10_932 ();
 sg13g2_fill_1 FILLER_10_934 ();
 sg13g2_fill_2 FILLER_10_956 ();
 sg13g2_fill_1 FILLER_10_962 ();
 sg13g2_fill_2 FILLER_10_967 ();
 sg13g2_fill_1 FILLER_10_973 ();
 sg13g2_fill_2 FILLER_10_979 ();
 sg13g2_fill_2 FILLER_10_985 ();
 sg13g2_fill_1 FILLER_10_987 ();
 sg13g2_decap_8 FILLER_10_996 ();
 sg13g2_decap_8 FILLER_10_1003 ();
 sg13g2_fill_2 FILLER_10_1010 ();
 sg13g2_decap_4 FILLER_10_1020 ();
 sg13g2_fill_2 FILLER_10_1024 ();
 sg13g2_decap_8 FILLER_10_1077 ();
 sg13g2_decap_8 FILLER_10_1084 ();
 sg13g2_decap_8 FILLER_10_1091 ();
 sg13g2_decap_8 FILLER_10_1098 ();
 sg13g2_decap_8 FILLER_10_1105 ();
 sg13g2_decap_8 FILLER_10_1112 ();
 sg13g2_decap_8 FILLER_10_1119 ();
 sg13g2_decap_8 FILLER_10_1126 ();
 sg13g2_decap_8 FILLER_10_1133 ();
 sg13g2_decap_8 FILLER_10_1140 ();
 sg13g2_decap_8 FILLER_10_1147 ();
 sg13g2_decap_8 FILLER_10_1154 ();
 sg13g2_decap_8 FILLER_10_1161 ();
 sg13g2_decap_8 FILLER_10_1168 ();
 sg13g2_decap_8 FILLER_10_1175 ();
 sg13g2_decap_8 FILLER_10_1182 ();
 sg13g2_decap_8 FILLER_10_1189 ();
 sg13g2_decap_8 FILLER_10_1196 ();
 sg13g2_decap_8 FILLER_10_1203 ();
 sg13g2_decap_8 FILLER_10_1210 ();
 sg13g2_decap_8 FILLER_10_1217 ();
 sg13g2_decap_8 FILLER_10_1224 ();
 sg13g2_decap_8 FILLER_10_1231 ();
 sg13g2_decap_8 FILLER_10_1238 ();
 sg13g2_decap_8 FILLER_10_1245 ();
 sg13g2_decap_8 FILLER_10_1252 ();
 sg13g2_decap_8 FILLER_10_1259 ();
 sg13g2_decap_8 FILLER_10_1266 ();
 sg13g2_decap_8 FILLER_10_1273 ();
 sg13g2_decap_8 FILLER_10_1280 ();
 sg13g2_decap_8 FILLER_10_1287 ();
 sg13g2_decap_8 FILLER_10_1294 ();
 sg13g2_decap_8 FILLER_10_1301 ();
 sg13g2_decap_8 FILLER_10_1308 ();
 sg13g2_decap_8 FILLER_10_1315 ();
 sg13g2_decap_4 FILLER_10_1322 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_92 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_fill_1 FILLER_11_141 ();
 sg13g2_fill_2 FILLER_11_147 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_2 FILLER_11_205 ();
 sg13g2_fill_2 FILLER_11_230 ();
 sg13g2_decap_4 FILLER_11_240 ();
 sg13g2_fill_2 FILLER_11_294 ();
 sg13g2_decap_4 FILLER_11_325 ();
 sg13g2_fill_1 FILLER_11_329 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_fill_2 FILLER_11_353 ();
 sg13g2_fill_1 FILLER_11_355 ();
 sg13g2_decap_4 FILLER_11_360 ();
 sg13g2_fill_1 FILLER_11_364 ();
 sg13g2_fill_2 FILLER_11_369 ();
 sg13g2_fill_1 FILLER_11_401 ();
 sg13g2_fill_1 FILLER_11_451 ();
 sg13g2_fill_1 FILLER_11_482 ();
 sg13g2_fill_2 FILLER_11_492 ();
 sg13g2_fill_1 FILLER_11_494 ();
 sg13g2_fill_2 FILLER_11_511 ();
 sg13g2_fill_1 FILLER_11_518 ();
 sg13g2_fill_2 FILLER_11_524 ();
 sg13g2_fill_2 FILLER_11_535 ();
 sg13g2_fill_1 FILLER_11_537 ();
 sg13g2_fill_1 FILLER_11_572 ();
 sg13g2_fill_2 FILLER_11_586 ();
 sg13g2_fill_1 FILLER_11_588 ();
 sg13g2_fill_1 FILLER_11_622 ();
 sg13g2_fill_2 FILLER_11_640 ();
 sg13g2_decap_4 FILLER_11_654 ();
 sg13g2_fill_2 FILLER_11_658 ();
 sg13g2_fill_1 FILLER_11_672 ();
 sg13g2_fill_2 FILLER_11_703 ();
 sg13g2_fill_2 FILLER_11_743 ();
 sg13g2_fill_1 FILLER_11_749 ();
 sg13g2_fill_1 FILLER_11_755 ();
 sg13g2_fill_1 FILLER_11_760 ();
 sg13g2_fill_2 FILLER_11_766 ();
 sg13g2_fill_1 FILLER_11_773 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_fill_1 FILLER_11_844 ();
 sg13g2_fill_2 FILLER_11_850 ();
 sg13g2_decap_8 FILLER_11_856 ();
 sg13g2_fill_2 FILLER_11_932 ();
 sg13g2_fill_1 FILLER_11_960 ();
 sg13g2_fill_2 FILLER_11_991 ();
 sg13g2_fill_1 FILLER_11_993 ();
 sg13g2_fill_1 FILLER_11_998 ();
 sg13g2_fill_1 FILLER_11_1007 ();
 sg13g2_decap_8 FILLER_11_1072 ();
 sg13g2_decap_8 FILLER_11_1079 ();
 sg13g2_decap_8 FILLER_11_1086 ();
 sg13g2_decap_8 FILLER_11_1093 ();
 sg13g2_decap_8 FILLER_11_1100 ();
 sg13g2_decap_8 FILLER_11_1107 ();
 sg13g2_decap_8 FILLER_11_1114 ();
 sg13g2_decap_8 FILLER_11_1121 ();
 sg13g2_decap_8 FILLER_11_1128 ();
 sg13g2_decap_8 FILLER_11_1135 ();
 sg13g2_decap_8 FILLER_11_1142 ();
 sg13g2_decap_8 FILLER_11_1149 ();
 sg13g2_decap_8 FILLER_11_1156 ();
 sg13g2_decap_8 FILLER_11_1163 ();
 sg13g2_decap_8 FILLER_11_1170 ();
 sg13g2_decap_8 FILLER_11_1177 ();
 sg13g2_decap_8 FILLER_11_1184 ();
 sg13g2_decap_8 FILLER_11_1191 ();
 sg13g2_decap_8 FILLER_11_1198 ();
 sg13g2_decap_8 FILLER_11_1205 ();
 sg13g2_decap_8 FILLER_11_1212 ();
 sg13g2_decap_8 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1226 ();
 sg13g2_decap_8 FILLER_11_1233 ();
 sg13g2_decap_8 FILLER_11_1240 ();
 sg13g2_decap_8 FILLER_11_1247 ();
 sg13g2_decap_8 FILLER_11_1254 ();
 sg13g2_decap_8 FILLER_11_1261 ();
 sg13g2_decap_8 FILLER_11_1268 ();
 sg13g2_decap_8 FILLER_11_1275 ();
 sg13g2_decap_8 FILLER_11_1282 ();
 sg13g2_decap_8 FILLER_11_1289 ();
 sg13g2_decap_8 FILLER_11_1296 ();
 sg13g2_decap_8 FILLER_11_1303 ();
 sg13g2_decap_8 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1317 ();
 sg13g2_fill_2 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_56 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_162 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_decap_4 FILLER_12_247 ();
 sg13g2_decap_4 FILLER_12_255 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_268 ();
 sg13g2_decap_4 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_279 ();
 sg13g2_decap_4 FILLER_12_311 ();
 sg13g2_fill_2 FILLER_12_365 ();
 sg13g2_fill_1 FILLER_12_367 ();
 sg13g2_fill_2 FILLER_12_394 ();
 sg13g2_fill_1 FILLER_12_415 ();
 sg13g2_fill_1 FILLER_12_442 ();
 sg13g2_fill_1 FILLER_12_448 ();
 sg13g2_fill_1 FILLER_12_453 ();
 sg13g2_fill_1 FILLER_12_459 ();
 sg13g2_fill_1 FILLER_12_465 ();
 sg13g2_fill_2 FILLER_12_479 ();
 sg13g2_fill_1 FILLER_12_481 ();
 sg13g2_fill_1 FILLER_12_486 ();
 sg13g2_fill_2 FILLER_12_492 ();
 sg13g2_fill_2 FILLER_12_556 ();
 sg13g2_fill_2 FILLER_12_571 ();
 sg13g2_fill_1 FILLER_12_573 ();
 sg13g2_fill_1 FILLER_12_581 ();
 sg13g2_fill_1 FILLER_12_587 ();
 sg13g2_fill_1 FILLER_12_593 ();
 sg13g2_fill_2 FILLER_12_612 ();
 sg13g2_fill_2 FILLER_12_619 ();
 sg13g2_fill_2 FILLER_12_641 ();
 sg13g2_decap_4 FILLER_12_652 ();
 sg13g2_fill_2 FILLER_12_685 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_fill_2 FILLER_12_698 ();
 sg13g2_fill_1 FILLER_12_700 ();
 sg13g2_fill_2 FILLER_12_709 ();
 sg13g2_fill_2 FILLER_12_725 ();
 sg13g2_fill_1 FILLER_12_727 ();
 sg13g2_fill_1 FILLER_12_736 ();
 sg13g2_fill_1 FILLER_12_763 ();
 sg13g2_fill_1 FILLER_12_773 ();
 sg13g2_fill_1 FILLER_12_782 ();
 sg13g2_decap_4 FILLER_12_791 ();
 sg13g2_fill_2 FILLER_12_795 ();
 sg13g2_decap_4 FILLER_12_801 ();
 sg13g2_decap_4 FILLER_12_815 ();
 sg13g2_fill_1 FILLER_12_823 ();
 sg13g2_fill_2 FILLER_12_866 ();
 sg13g2_fill_2 FILLER_12_876 ();
 sg13g2_fill_2 FILLER_12_887 ();
 sg13g2_fill_2 FILLER_12_894 ();
 sg13g2_fill_2 FILLER_12_912 ();
 sg13g2_decap_4 FILLER_12_937 ();
 sg13g2_fill_2 FILLER_12_949 ();
 sg13g2_fill_1 FILLER_12_951 ();
 sg13g2_fill_1 FILLER_12_960 ();
 sg13g2_fill_1 FILLER_12_973 ();
 sg13g2_fill_1 FILLER_12_982 ();
 sg13g2_fill_2 FILLER_12_1041 ();
 sg13g2_fill_1 FILLER_12_1043 ();
 sg13g2_decap_8 FILLER_12_1075 ();
 sg13g2_decap_8 FILLER_12_1082 ();
 sg13g2_decap_8 FILLER_12_1089 ();
 sg13g2_decap_8 FILLER_12_1096 ();
 sg13g2_decap_8 FILLER_12_1103 ();
 sg13g2_decap_8 FILLER_12_1110 ();
 sg13g2_decap_8 FILLER_12_1117 ();
 sg13g2_decap_8 FILLER_12_1124 ();
 sg13g2_decap_8 FILLER_12_1131 ();
 sg13g2_decap_8 FILLER_12_1138 ();
 sg13g2_decap_8 FILLER_12_1145 ();
 sg13g2_decap_8 FILLER_12_1152 ();
 sg13g2_decap_8 FILLER_12_1159 ();
 sg13g2_decap_8 FILLER_12_1166 ();
 sg13g2_decap_8 FILLER_12_1173 ();
 sg13g2_decap_8 FILLER_12_1180 ();
 sg13g2_decap_8 FILLER_12_1187 ();
 sg13g2_decap_8 FILLER_12_1194 ();
 sg13g2_decap_8 FILLER_12_1201 ();
 sg13g2_decap_8 FILLER_12_1208 ();
 sg13g2_decap_8 FILLER_12_1215 ();
 sg13g2_decap_8 FILLER_12_1222 ();
 sg13g2_decap_8 FILLER_12_1229 ();
 sg13g2_decap_8 FILLER_12_1236 ();
 sg13g2_decap_8 FILLER_12_1243 ();
 sg13g2_decap_8 FILLER_12_1250 ();
 sg13g2_decap_8 FILLER_12_1257 ();
 sg13g2_decap_8 FILLER_12_1264 ();
 sg13g2_decap_8 FILLER_12_1271 ();
 sg13g2_decap_8 FILLER_12_1278 ();
 sg13g2_decap_8 FILLER_12_1285 ();
 sg13g2_decap_8 FILLER_12_1292 ();
 sg13g2_decap_8 FILLER_12_1299 ();
 sg13g2_decap_8 FILLER_12_1306 ();
 sg13g2_decap_8 FILLER_12_1313 ();
 sg13g2_decap_4 FILLER_12_1320 ();
 sg13g2_fill_2 FILLER_12_1324 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_80 ();
 sg13g2_decap_8 FILLER_13_86 ();
 sg13g2_decap_4 FILLER_13_93 ();
 sg13g2_fill_1 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_13_150 ();
 sg13g2_decap_8 FILLER_13_155 ();
 sg13g2_fill_2 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_232 ();
 sg13g2_fill_2 FILLER_13_237 ();
 sg13g2_decap_4 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_1 FILLER_13_309 ();
 sg13g2_fill_1 FILLER_13_323 ();
 sg13g2_fill_1 FILLER_13_329 ();
 sg13g2_fill_1 FILLER_13_335 ();
 sg13g2_fill_1 FILLER_13_342 ();
 sg13g2_decap_4 FILLER_13_347 ();
 sg13g2_fill_2 FILLER_13_361 ();
 sg13g2_fill_1 FILLER_13_367 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_400 ();
 sg13g2_fill_1 FILLER_13_421 ();
 sg13g2_decap_4 FILLER_13_440 ();
 sg13g2_decap_4 FILLER_13_452 ();
 sg13g2_fill_2 FILLER_13_456 ();
 sg13g2_fill_1 FILLER_13_462 ();
 sg13g2_fill_1 FILLER_13_467 ();
 sg13g2_fill_2 FILLER_13_494 ();
 sg13g2_fill_1 FILLER_13_496 ();
 sg13g2_fill_2 FILLER_13_506 ();
 sg13g2_fill_2 FILLER_13_526 ();
 sg13g2_fill_1 FILLER_13_528 ();
 sg13g2_fill_2 FILLER_13_546 ();
 sg13g2_fill_1 FILLER_13_583 ();
 sg13g2_fill_1 FILLER_13_587 ();
 sg13g2_fill_1 FILLER_13_596 ();
 sg13g2_fill_1 FILLER_13_613 ();
 sg13g2_fill_1 FILLER_13_620 ();
 sg13g2_fill_1 FILLER_13_654 ();
 sg13g2_fill_1 FILLER_13_677 ();
 sg13g2_fill_1 FILLER_13_686 ();
 sg13g2_fill_1 FILLER_13_762 ();
 sg13g2_fill_2 FILLER_13_780 ();
 sg13g2_fill_1 FILLER_13_877 ();
 sg13g2_fill_1 FILLER_13_916 ();
 sg13g2_fill_2 FILLER_13_948 ();
 sg13g2_fill_1 FILLER_13_950 ();
 sg13g2_fill_1 FILLER_13_996 ();
 sg13g2_fill_2 FILLER_13_1010 ();
 sg13g2_decap_4 FILLER_13_1049 ();
 sg13g2_decap_8 FILLER_13_1062 ();
 sg13g2_decap_8 FILLER_13_1069 ();
 sg13g2_decap_8 FILLER_13_1076 ();
 sg13g2_decap_8 FILLER_13_1083 ();
 sg13g2_decap_8 FILLER_13_1090 ();
 sg13g2_decap_8 FILLER_13_1097 ();
 sg13g2_decap_8 FILLER_13_1104 ();
 sg13g2_decap_8 FILLER_13_1111 ();
 sg13g2_decap_8 FILLER_13_1118 ();
 sg13g2_decap_8 FILLER_13_1125 ();
 sg13g2_decap_8 FILLER_13_1132 ();
 sg13g2_decap_8 FILLER_13_1139 ();
 sg13g2_decap_8 FILLER_13_1146 ();
 sg13g2_decap_8 FILLER_13_1153 ();
 sg13g2_decap_8 FILLER_13_1160 ();
 sg13g2_decap_8 FILLER_13_1167 ();
 sg13g2_decap_8 FILLER_13_1174 ();
 sg13g2_decap_8 FILLER_13_1181 ();
 sg13g2_decap_8 FILLER_13_1188 ();
 sg13g2_decap_8 FILLER_13_1195 ();
 sg13g2_decap_8 FILLER_13_1202 ();
 sg13g2_decap_8 FILLER_13_1209 ();
 sg13g2_decap_8 FILLER_13_1216 ();
 sg13g2_decap_8 FILLER_13_1223 ();
 sg13g2_decap_8 FILLER_13_1230 ();
 sg13g2_decap_8 FILLER_13_1237 ();
 sg13g2_decap_8 FILLER_13_1244 ();
 sg13g2_decap_8 FILLER_13_1251 ();
 sg13g2_decap_8 FILLER_13_1258 ();
 sg13g2_decap_8 FILLER_13_1265 ();
 sg13g2_decap_8 FILLER_13_1272 ();
 sg13g2_decap_8 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1286 ();
 sg13g2_decap_8 FILLER_13_1293 ();
 sg13g2_decap_8 FILLER_13_1300 ();
 sg13g2_decap_8 FILLER_13_1307 ();
 sg13g2_decap_8 FILLER_13_1314 ();
 sg13g2_decap_4 FILLER_13_1321 ();
 sg13g2_fill_1 FILLER_13_1325 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_4 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_128 ();
 sg13g2_fill_1 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_fill_2 FILLER_14_158 ();
 sg13g2_fill_1 FILLER_14_160 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_fill_1 FILLER_14_213 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_231 ();
 sg13g2_decap_4 FILLER_14_258 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_4 FILLER_14_345 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_fill_2 FILLER_14_363 ();
 sg13g2_fill_1 FILLER_14_430 ();
 sg13g2_fill_1 FILLER_14_436 ();
 sg13g2_fill_1 FILLER_14_445 ();
 sg13g2_fill_1 FILLER_14_477 ();
 sg13g2_fill_2 FILLER_14_483 ();
 sg13g2_fill_2 FILLER_14_511 ();
 sg13g2_fill_2 FILLER_14_564 ();
 sg13g2_decap_4 FILLER_14_570 ();
 sg13g2_fill_2 FILLER_14_579 ();
 sg13g2_fill_1 FILLER_14_601 ();
 sg13g2_decap_4 FILLER_14_607 ();
 sg13g2_fill_1 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_621 ();
 sg13g2_fill_1 FILLER_14_627 ();
 sg13g2_fill_1 FILLER_14_633 ();
 sg13g2_fill_2 FILLER_14_638 ();
 sg13g2_fill_1 FILLER_14_645 ();
 sg13g2_fill_2 FILLER_14_657 ();
 sg13g2_fill_1 FILLER_14_659 ();
 sg13g2_fill_2 FILLER_14_665 ();
 sg13g2_fill_1 FILLER_14_673 ();
 sg13g2_fill_1 FILLER_14_683 ();
 sg13g2_fill_2 FILLER_14_688 ();
 sg13g2_fill_1 FILLER_14_690 ();
 sg13g2_fill_2 FILLER_14_699 ();
 sg13g2_fill_1 FILLER_14_705 ();
 sg13g2_fill_2 FILLER_14_731 ();
 sg13g2_fill_1 FILLER_14_733 ();
 sg13g2_fill_2 FILLER_14_763 ();
 sg13g2_fill_2 FILLER_14_799 ();
 sg13g2_decap_4 FILLER_14_805 ();
 sg13g2_fill_1 FILLER_14_817 ();
 sg13g2_fill_1 FILLER_14_822 ();
 sg13g2_fill_1 FILLER_14_828 ();
 sg13g2_fill_1 FILLER_14_834 ();
 sg13g2_decap_4 FILLER_14_839 ();
 sg13g2_fill_2 FILLER_14_843 ();
 sg13g2_decap_4 FILLER_14_858 ();
 sg13g2_fill_1 FILLER_14_862 ();
 sg13g2_fill_2 FILLER_14_872 ();
 sg13g2_fill_1 FILLER_14_891 ();
 sg13g2_fill_1 FILLER_14_900 ();
 sg13g2_fill_1 FILLER_14_905 ();
 sg13g2_fill_2 FILLER_14_936 ();
 sg13g2_fill_2 FILLER_14_947 ();
 sg13g2_fill_1 FILLER_14_949 ();
 sg13g2_fill_2 FILLER_14_989 ();
 sg13g2_fill_1 FILLER_14_1011 ();
 sg13g2_fill_2 FILLER_14_1054 ();
 sg13g2_fill_1 FILLER_14_1056 ();
 sg13g2_decap_8 FILLER_14_1083 ();
 sg13g2_decap_8 FILLER_14_1090 ();
 sg13g2_decap_8 FILLER_14_1097 ();
 sg13g2_decap_8 FILLER_14_1104 ();
 sg13g2_decap_8 FILLER_14_1111 ();
 sg13g2_decap_8 FILLER_14_1118 ();
 sg13g2_decap_8 FILLER_14_1125 ();
 sg13g2_decap_8 FILLER_14_1132 ();
 sg13g2_decap_8 FILLER_14_1139 ();
 sg13g2_decap_8 FILLER_14_1146 ();
 sg13g2_decap_8 FILLER_14_1153 ();
 sg13g2_decap_8 FILLER_14_1160 ();
 sg13g2_decap_8 FILLER_14_1167 ();
 sg13g2_decap_8 FILLER_14_1174 ();
 sg13g2_decap_8 FILLER_14_1181 ();
 sg13g2_decap_8 FILLER_14_1188 ();
 sg13g2_decap_8 FILLER_14_1195 ();
 sg13g2_decap_8 FILLER_14_1202 ();
 sg13g2_decap_8 FILLER_14_1209 ();
 sg13g2_decap_8 FILLER_14_1216 ();
 sg13g2_decap_8 FILLER_14_1223 ();
 sg13g2_decap_8 FILLER_14_1230 ();
 sg13g2_decap_8 FILLER_14_1237 ();
 sg13g2_decap_8 FILLER_14_1244 ();
 sg13g2_decap_8 FILLER_14_1251 ();
 sg13g2_decap_8 FILLER_14_1258 ();
 sg13g2_decap_8 FILLER_14_1265 ();
 sg13g2_decap_8 FILLER_14_1272 ();
 sg13g2_decap_8 FILLER_14_1279 ();
 sg13g2_decap_8 FILLER_14_1286 ();
 sg13g2_decap_8 FILLER_14_1293 ();
 sg13g2_decap_8 FILLER_14_1300 ();
 sg13g2_decap_8 FILLER_14_1307 ();
 sg13g2_decap_8 FILLER_14_1314 ();
 sg13g2_decap_4 FILLER_14_1321 ();
 sg13g2_fill_1 FILLER_14_1325 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_2 FILLER_15_80 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_89 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_fill_2 FILLER_15_103 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_114 ();
 sg13g2_fill_1 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_145 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_1 FILLER_15_157 ();
 sg13g2_fill_2 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_174 ();
 sg13g2_fill_2 FILLER_15_180 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_1 FILLER_15_229 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_237 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_269 ();
 sg13g2_fill_2 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_284 ();
 sg13g2_fill_2 FILLER_15_323 ();
 sg13g2_fill_1 FILLER_15_347 ();
 sg13g2_fill_2 FILLER_15_374 ();
 sg13g2_fill_2 FILLER_15_411 ();
 sg13g2_fill_2 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_15_436 ();
 sg13g2_fill_2 FILLER_15_443 ();
 sg13g2_fill_1 FILLER_15_445 ();
 sg13g2_fill_1 FILLER_15_464 ();
 sg13g2_fill_2 FILLER_15_495 ();
 sg13g2_fill_2 FILLER_15_542 ();
 sg13g2_fill_2 FILLER_15_579 ();
 sg13g2_fill_2 FILLER_15_589 ();
 sg13g2_fill_2 FILLER_15_599 ();
 sg13g2_fill_1 FILLER_15_601 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_fill_1 FILLER_15_613 ();
 sg13g2_fill_2 FILLER_15_661 ();
 sg13g2_fill_1 FILLER_15_674 ();
 sg13g2_fill_2 FILLER_15_680 ();
 sg13g2_fill_2 FILLER_15_723 ();
 sg13g2_fill_1 FILLER_15_729 ();
 sg13g2_fill_2 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_752 ();
 sg13g2_fill_1 FILLER_15_759 ();
 sg13g2_fill_1 FILLER_15_820 ();
 sg13g2_fill_1 FILLER_15_851 ();
 sg13g2_fill_1 FILLER_15_887 ();
 sg13g2_fill_1 FILLER_15_892 ();
 sg13g2_fill_1 FILLER_15_898 ();
 sg13g2_fill_2 FILLER_15_907 ();
 sg13g2_fill_1 FILLER_15_940 ();
 sg13g2_fill_2 FILLER_15_954 ();
 sg13g2_fill_1 FILLER_15_982 ();
 sg13g2_fill_2 FILLER_15_1043 ();
 sg13g2_decap_4 FILLER_15_1076 ();
 sg13g2_fill_2 FILLER_15_1080 ();
 sg13g2_decap_8 FILLER_15_1090 ();
 sg13g2_decap_8 FILLER_15_1097 ();
 sg13g2_decap_8 FILLER_15_1104 ();
 sg13g2_decap_8 FILLER_15_1111 ();
 sg13g2_decap_8 FILLER_15_1118 ();
 sg13g2_decap_8 FILLER_15_1125 ();
 sg13g2_decap_8 FILLER_15_1132 ();
 sg13g2_decap_8 FILLER_15_1139 ();
 sg13g2_decap_8 FILLER_15_1146 ();
 sg13g2_decap_8 FILLER_15_1153 ();
 sg13g2_decap_8 FILLER_15_1160 ();
 sg13g2_decap_8 FILLER_15_1167 ();
 sg13g2_decap_8 FILLER_15_1174 ();
 sg13g2_decap_8 FILLER_15_1181 ();
 sg13g2_decap_8 FILLER_15_1188 ();
 sg13g2_decap_8 FILLER_15_1195 ();
 sg13g2_decap_8 FILLER_15_1202 ();
 sg13g2_decap_8 FILLER_15_1209 ();
 sg13g2_decap_8 FILLER_15_1216 ();
 sg13g2_decap_8 FILLER_15_1223 ();
 sg13g2_decap_8 FILLER_15_1230 ();
 sg13g2_decap_8 FILLER_15_1237 ();
 sg13g2_decap_8 FILLER_15_1244 ();
 sg13g2_decap_8 FILLER_15_1251 ();
 sg13g2_decap_8 FILLER_15_1258 ();
 sg13g2_decap_8 FILLER_15_1265 ();
 sg13g2_decap_8 FILLER_15_1272 ();
 sg13g2_decap_8 FILLER_15_1279 ();
 sg13g2_decap_8 FILLER_15_1286 ();
 sg13g2_decap_8 FILLER_15_1293 ();
 sg13g2_decap_8 FILLER_15_1300 ();
 sg13g2_decap_8 FILLER_15_1307 ();
 sg13g2_decap_8 FILLER_15_1314 ();
 sg13g2_decap_4 FILLER_15_1321 ();
 sg13g2_fill_1 FILLER_15_1325 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_4 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_53 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_124 ();
 sg13g2_fill_1 FILLER_16_130 ();
 sg13g2_fill_2 FILLER_16_136 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_294 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_decap_4 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_388 ();
 sg13g2_fill_1 FILLER_16_390 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_397 ();
 sg13g2_fill_2 FILLER_16_402 ();
 sg13g2_fill_1 FILLER_16_411 ();
 sg13g2_fill_2 FILLER_16_479 ();
 sg13g2_fill_2 FILLER_16_559 ();
 sg13g2_fill_1 FILLER_16_588 ();
 sg13g2_fill_2 FILLER_16_640 ();
 sg13g2_fill_2 FILLER_16_708 ();
 sg13g2_fill_1 FILLER_16_718 ();
 sg13g2_fill_2 FILLER_16_782 ();
 sg13g2_fill_2 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_820 ();
 sg13g2_fill_1 FILLER_16_827 ();
 sg13g2_fill_1 FILLER_16_859 ();
 sg13g2_fill_1 FILLER_16_924 ();
 sg13g2_fill_2 FILLER_16_964 ();
 sg13g2_fill_1 FILLER_16_983 ();
 sg13g2_fill_1 FILLER_16_989 ();
 sg13g2_fill_1 FILLER_16_995 ();
 sg13g2_fill_2 FILLER_16_1035 ();
 sg13g2_fill_1 FILLER_16_1037 ();
 sg13g2_decap_4 FILLER_16_1047 ();
 sg13g2_fill_2 FILLER_16_1068 ();
 sg13g2_fill_1 FILLER_16_1078 ();
 sg13g2_decap_8 FILLER_16_1105 ();
 sg13g2_decap_8 FILLER_16_1112 ();
 sg13g2_decap_8 FILLER_16_1119 ();
 sg13g2_decap_8 FILLER_16_1126 ();
 sg13g2_decap_8 FILLER_16_1133 ();
 sg13g2_decap_8 FILLER_16_1140 ();
 sg13g2_decap_8 FILLER_16_1147 ();
 sg13g2_decap_8 FILLER_16_1154 ();
 sg13g2_decap_8 FILLER_16_1161 ();
 sg13g2_decap_8 FILLER_16_1168 ();
 sg13g2_decap_8 FILLER_16_1175 ();
 sg13g2_decap_8 FILLER_16_1182 ();
 sg13g2_decap_8 FILLER_16_1189 ();
 sg13g2_decap_8 FILLER_16_1196 ();
 sg13g2_decap_8 FILLER_16_1203 ();
 sg13g2_decap_8 FILLER_16_1210 ();
 sg13g2_decap_8 FILLER_16_1217 ();
 sg13g2_decap_8 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1231 ();
 sg13g2_decap_8 FILLER_16_1238 ();
 sg13g2_decap_8 FILLER_16_1245 ();
 sg13g2_decap_8 FILLER_16_1252 ();
 sg13g2_decap_8 FILLER_16_1259 ();
 sg13g2_decap_8 FILLER_16_1266 ();
 sg13g2_decap_8 FILLER_16_1273 ();
 sg13g2_decap_8 FILLER_16_1280 ();
 sg13g2_decap_8 FILLER_16_1287 ();
 sg13g2_decap_8 FILLER_16_1294 ();
 sg13g2_decap_8 FILLER_16_1301 ();
 sg13g2_decap_8 FILLER_16_1308 ();
 sg13g2_decap_8 FILLER_16_1315 ();
 sg13g2_decap_4 FILLER_16_1322 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_56 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_17_78 ();
 sg13g2_decap_8 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_fill_2 FILLER_17_113 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_fill_2 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_fill_1 FILLER_17_415 ();
 sg13g2_fill_2 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_2 FILLER_17_477 ();
 sg13g2_fill_2 FILLER_17_501 ();
 sg13g2_fill_1 FILLER_17_529 ();
 sg13g2_fill_2 FILLER_17_548 ();
 sg13g2_fill_1 FILLER_17_550 ();
 sg13g2_fill_1 FILLER_17_577 ();
 sg13g2_fill_1 FILLER_17_595 ();
 sg13g2_fill_1 FILLER_17_604 ();
 sg13g2_fill_1 FILLER_17_609 ();
 sg13g2_fill_1 FILLER_17_615 ();
 sg13g2_fill_1 FILLER_17_624 ();
 sg13g2_decap_4 FILLER_17_649 ();
 sg13g2_fill_2 FILLER_17_661 ();
 sg13g2_fill_1 FILLER_17_663 ();
 sg13g2_decap_4 FILLER_17_669 ();
 sg13g2_fill_2 FILLER_17_673 ();
 sg13g2_fill_2 FILLER_17_687 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_fill_2 FILLER_17_708 ();
 sg13g2_fill_1 FILLER_17_710 ();
 sg13g2_fill_2 FILLER_17_750 ();
 sg13g2_fill_1 FILLER_17_752 ();
 sg13g2_fill_1 FILLER_17_758 ();
 sg13g2_fill_1 FILLER_17_763 ();
 sg13g2_fill_1 FILLER_17_796 ();
 sg13g2_fill_1 FILLER_17_841 ();
 sg13g2_fill_2 FILLER_17_859 ();
 sg13g2_fill_1 FILLER_17_881 ();
 sg13g2_fill_1 FILLER_17_931 ();
 sg13g2_fill_1 FILLER_17_945 ();
 sg13g2_fill_1 FILLER_17_950 ();
 sg13g2_fill_2 FILLER_17_972 ();
 sg13g2_fill_2 FILLER_17_979 ();
 sg13g2_fill_1 FILLER_17_981 ();
 sg13g2_fill_1 FILLER_17_991 ();
 sg13g2_fill_2 FILLER_17_1022 ();
 sg13g2_fill_2 FILLER_17_1028 ();
 sg13g2_decap_8 FILLER_17_1098 ();
 sg13g2_decap_8 FILLER_17_1105 ();
 sg13g2_decap_8 FILLER_17_1112 ();
 sg13g2_decap_8 FILLER_17_1119 ();
 sg13g2_decap_8 FILLER_17_1126 ();
 sg13g2_decap_8 FILLER_17_1133 ();
 sg13g2_decap_8 FILLER_17_1140 ();
 sg13g2_decap_8 FILLER_17_1147 ();
 sg13g2_decap_8 FILLER_17_1154 ();
 sg13g2_decap_8 FILLER_17_1161 ();
 sg13g2_decap_8 FILLER_17_1168 ();
 sg13g2_decap_8 FILLER_17_1175 ();
 sg13g2_decap_8 FILLER_17_1182 ();
 sg13g2_decap_8 FILLER_17_1189 ();
 sg13g2_decap_8 FILLER_17_1196 ();
 sg13g2_decap_8 FILLER_17_1203 ();
 sg13g2_decap_8 FILLER_17_1210 ();
 sg13g2_decap_8 FILLER_17_1217 ();
 sg13g2_decap_8 FILLER_17_1224 ();
 sg13g2_decap_8 FILLER_17_1231 ();
 sg13g2_decap_8 FILLER_17_1238 ();
 sg13g2_decap_8 FILLER_17_1245 ();
 sg13g2_decap_8 FILLER_17_1252 ();
 sg13g2_decap_8 FILLER_17_1259 ();
 sg13g2_decap_8 FILLER_17_1266 ();
 sg13g2_decap_8 FILLER_17_1273 ();
 sg13g2_decap_8 FILLER_17_1280 ();
 sg13g2_decap_8 FILLER_17_1287 ();
 sg13g2_decap_8 FILLER_17_1294 ();
 sg13g2_decap_8 FILLER_17_1301 ();
 sg13g2_decap_8 FILLER_17_1308 ();
 sg13g2_decap_8 FILLER_17_1315 ();
 sg13g2_decap_4 FILLER_17_1322 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_180 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_270 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_fill_2 FILLER_18_301 ();
 sg13g2_fill_2 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_fill_2 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_fill_1 FILLER_18_391 ();
 sg13g2_fill_2 FILLER_18_396 ();
 sg13g2_fill_2 FILLER_18_402 ();
 sg13g2_fill_1 FILLER_18_426 ();
 sg13g2_fill_2 FILLER_18_435 ();
 sg13g2_fill_2 FILLER_18_446 ();
 sg13g2_fill_1 FILLER_18_448 ();
 sg13g2_fill_2 FILLER_18_453 ();
 sg13g2_fill_2 FILLER_18_508 ();
 sg13g2_fill_2 FILLER_18_519 ();
 sg13g2_decap_8 FILLER_18_568 ();
 sg13g2_decap_4 FILLER_18_575 ();
 sg13g2_fill_2 FILLER_18_579 ();
 sg13g2_fill_1 FILLER_18_585 ();
 sg13g2_fill_2 FILLER_18_624 ();
 sg13g2_fill_1 FILLER_18_643 ();
 sg13g2_fill_2 FILLER_18_649 ();
 sg13g2_fill_1 FILLER_18_656 ();
 sg13g2_fill_2 FILLER_18_664 ();
 sg13g2_fill_1 FILLER_18_666 ();
 sg13g2_fill_1 FILLER_18_672 ();
 sg13g2_fill_1 FILLER_18_747 ();
 sg13g2_decap_8 FILLER_18_752 ();
 sg13g2_decap_4 FILLER_18_759 ();
 sg13g2_fill_1 FILLER_18_763 ();
 sg13g2_fill_2 FILLER_18_769 ();
 sg13g2_fill_1 FILLER_18_787 ();
 sg13g2_decap_4 FILLER_18_792 ();
 sg13g2_decap_4 FILLER_18_800 ();
 sg13g2_fill_1 FILLER_18_804 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_4 FILLER_18_830 ();
 sg13g2_fill_1 FILLER_18_850 ();
 sg13g2_fill_1 FILLER_18_869 ();
 sg13g2_fill_1 FILLER_18_874 ();
 sg13g2_fill_1 FILLER_18_880 ();
 sg13g2_fill_2 FILLER_18_903 ();
 sg13g2_fill_2 FILLER_18_914 ();
 sg13g2_decap_4 FILLER_18_955 ();
 sg13g2_fill_1 FILLER_18_974 ();
 sg13g2_fill_1 FILLER_18_988 ();
 sg13g2_fill_2 FILLER_18_994 ();
 sg13g2_fill_1 FILLER_18_996 ();
 sg13g2_fill_2 FILLER_18_1001 ();
 sg13g2_fill_1 FILLER_18_1003 ();
 sg13g2_fill_1 FILLER_18_1013 ();
 sg13g2_fill_1 FILLER_18_1044 ();
 sg13g2_fill_2 FILLER_18_1084 ();
 sg13g2_fill_2 FILLER_18_1095 ();
 sg13g2_decap_8 FILLER_18_1104 ();
 sg13g2_decap_8 FILLER_18_1111 ();
 sg13g2_decap_8 FILLER_18_1118 ();
 sg13g2_decap_8 FILLER_18_1125 ();
 sg13g2_decap_8 FILLER_18_1132 ();
 sg13g2_decap_8 FILLER_18_1139 ();
 sg13g2_decap_8 FILLER_18_1146 ();
 sg13g2_decap_8 FILLER_18_1153 ();
 sg13g2_decap_8 FILLER_18_1160 ();
 sg13g2_decap_8 FILLER_18_1167 ();
 sg13g2_decap_8 FILLER_18_1174 ();
 sg13g2_decap_8 FILLER_18_1181 ();
 sg13g2_decap_8 FILLER_18_1188 ();
 sg13g2_decap_8 FILLER_18_1195 ();
 sg13g2_decap_8 FILLER_18_1202 ();
 sg13g2_decap_8 FILLER_18_1209 ();
 sg13g2_decap_8 FILLER_18_1216 ();
 sg13g2_decap_8 FILLER_18_1223 ();
 sg13g2_decap_8 FILLER_18_1230 ();
 sg13g2_decap_8 FILLER_18_1237 ();
 sg13g2_decap_8 FILLER_18_1244 ();
 sg13g2_decap_8 FILLER_18_1251 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_8 FILLER_18_1265 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_8 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1286 ();
 sg13g2_decap_8 FILLER_18_1293 ();
 sg13g2_decap_8 FILLER_18_1300 ();
 sg13g2_decap_8 FILLER_18_1307 ();
 sg13g2_decap_8 FILLER_18_1314 ();
 sg13g2_decap_4 FILLER_18_1321 ();
 sg13g2_fill_1 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_110 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_fill_1 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_197 ();
 sg13g2_fill_2 FILLER_19_229 ();
 sg13g2_fill_2 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_416 ();
 sg13g2_fill_1 FILLER_19_418 ();
 sg13g2_fill_1 FILLER_19_428 ();
 sg13g2_fill_2 FILLER_19_434 ();
 sg13g2_fill_1 FILLER_19_444 ();
 sg13g2_fill_1 FILLER_19_454 ();
 sg13g2_fill_1 FILLER_19_496 ();
 sg13g2_fill_1 FILLER_19_502 ();
 sg13g2_fill_1 FILLER_19_508 ();
 sg13g2_fill_2 FILLER_19_520 ();
 sg13g2_fill_1 FILLER_19_526 ();
 sg13g2_fill_2 FILLER_19_532 ();
 sg13g2_fill_1 FILLER_19_538 ();
 sg13g2_fill_2 FILLER_19_543 ();
 sg13g2_fill_2 FILLER_19_549 ();
 sg13g2_decap_8 FILLER_19_590 ();
 sg13g2_fill_1 FILLER_19_605 ();
 sg13g2_fill_1 FILLER_19_614 ();
 sg13g2_fill_1 FILLER_19_625 ();
 sg13g2_fill_1 FILLER_19_649 ();
 sg13g2_fill_2 FILLER_19_673 ();
 sg13g2_fill_1 FILLER_19_675 ();
 sg13g2_decap_4 FILLER_19_733 ();
 sg13g2_fill_1 FILLER_19_737 ();
 sg13g2_fill_1 FILLER_19_870 ();
 sg13g2_fill_1 FILLER_19_881 ();
 sg13g2_fill_1 FILLER_19_890 ();
 sg13g2_fill_1 FILLER_19_921 ();
 sg13g2_fill_2 FILLER_19_982 ();
 sg13g2_fill_2 FILLER_19_996 ();
 sg13g2_fill_2 FILLER_19_1024 ();
 sg13g2_decap_4 FILLER_19_1030 ();
 sg13g2_fill_1 FILLER_19_1038 ();
 sg13g2_decap_4 FILLER_19_1053 ();
 sg13g2_fill_2 FILLER_19_1075 ();
 sg13g2_fill_1 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1112 ();
 sg13g2_decap_8 FILLER_19_1119 ();
 sg13g2_decap_8 FILLER_19_1126 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_decap_8 FILLER_19_1140 ();
 sg13g2_decap_8 FILLER_19_1147 ();
 sg13g2_decap_8 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1161 ();
 sg13g2_decap_8 FILLER_19_1168 ();
 sg13g2_decap_8 FILLER_19_1175 ();
 sg13g2_decap_8 FILLER_19_1182 ();
 sg13g2_decap_8 FILLER_19_1189 ();
 sg13g2_decap_8 FILLER_19_1196 ();
 sg13g2_decap_8 FILLER_19_1203 ();
 sg13g2_decap_8 FILLER_19_1210 ();
 sg13g2_decap_8 FILLER_19_1217 ();
 sg13g2_decap_8 FILLER_19_1224 ();
 sg13g2_decap_8 FILLER_19_1231 ();
 sg13g2_decap_8 FILLER_19_1238 ();
 sg13g2_decap_8 FILLER_19_1245 ();
 sg13g2_decap_8 FILLER_19_1252 ();
 sg13g2_decap_8 FILLER_19_1259 ();
 sg13g2_decap_8 FILLER_19_1266 ();
 sg13g2_decap_8 FILLER_19_1273 ();
 sg13g2_decap_8 FILLER_19_1280 ();
 sg13g2_decap_8 FILLER_19_1287 ();
 sg13g2_decap_8 FILLER_19_1294 ();
 sg13g2_decap_8 FILLER_19_1301 ();
 sg13g2_decap_8 FILLER_19_1308 ();
 sg13g2_decap_8 FILLER_19_1315 ();
 sg13g2_decap_4 FILLER_19_1322 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_42 ();
 sg13g2_fill_1 FILLER_20_46 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_100 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_204 ();
 sg13g2_fill_1 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_248 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_fill_2 FILLER_20_265 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_272 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_301 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_387 ();
 sg13g2_fill_2 FILLER_20_392 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_20_409 ();
 sg13g2_fill_1 FILLER_20_448 ();
 sg13g2_fill_1 FILLER_20_488 ();
 sg13g2_fill_1 FILLER_20_556 ();
 sg13g2_fill_2 FILLER_20_562 ();
 sg13g2_fill_2 FILLER_20_568 ();
 sg13g2_fill_2 FILLER_20_574 ();
 sg13g2_fill_2 FILLER_20_596 ();
 sg13g2_fill_2 FILLER_20_639 ();
 sg13g2_fill_1 FILLER_20_649 ();
 sg13g2_fill_1 FILLER_20_655 ();
 sg13g2_decap_4 FILLER_20_698 ();
 sg13g2_fill_2 FILLER_20_742 ();
 sg13g2_fill_1 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_761 ();
 sg13g2_decap_4 FILLER_20_797 ();
 sg13g2_fill_2 FILLER_20_806 ();
 sg13g2_fill_1 FILLER_20_808 ();
 sg13g2_decap_4 FILLER_20_813 ();
 sg13g2_fill_2 FILLER_20_827 ();
 sg13g2_fill_1 FILLER_20_829 ();
 sg13g2_fill_1 FILLER_20_860 ();
 sg13g2_decap_4 FILLER_20_945 ();
 sg13g2_fill_1 FILLER_20_949 ();
 sg13g2_fill_2 FILLER_20_970 ();
 sg13g2_fill_1 FILLER_20_979 ();
 sg13g2_decap_8 FILLER_20_985 ();
 sg13g2_decap_8 FILLER_20_992 ();
 sg13g2_decap_8 FILLER_20_999 ();
 sg13g2_fill_1 FILLER_20_1077 ();
 sg13g2_decap_8 FILLER_20_1094 ();
 sg13g2_decap_8 FILLER_20_1101 ();
 sg13g2_decap_8 FILLER_20_1108 ();
 sg13g2_decap_8 FILLER_20_1115 ();
 sg13g2_decap_8 FILLER_20_1122 ();
 sg13g2_decap_8 FILLER_20_1129 ();
 sg13g2_decap_8 FILLER_20_1136 ();
 sg13g2_decap_8 FILLER_20_1143 ();
 sg13g2_decap_8 FILLER_20_1150 ();
 sg13g2_decap_8 FILLER_20_1157 ();
 sg13g2_decap_8 FILLER_20_1164 ();
 sg13g2_decap_8 FILLER_20_1171 ();
 sg13g2_decap_8 FILLER_20_1178 ();
 sg13g2_decap_8 FILLER_20_1185 ();
 sg13g2_decap_8 FILLER_20_1192 ();
 sg13g2_decap_8 FILLER_20_1199 ();
 sg13g2_decap_8 FILLER_20_1206 ();
 sg13g2_decap_8 FILLER_20_1213 ();
 sg13g2_decap_8 FILLER_20_1220 ();
 sg13g2_decap_8 FILLER_20_1227 ();
 sg13g2_decap_8 FILLER_20_1234 ();
 sg13g2_decap_8 FILLER_20_1241 ();
 sg13g2_decap_8 FILLER_20_1248 ();
 sg13g2_decap_8 FILLER_20_1255 ();
 sg13g2_decap_8 FILLER_20_1262 ();
 sg13g2_decap_8 FILLER_20_1269 ();
 sg13g2_decap_8 FILLER_20_1276 ();
 sg13g2_decap_8 FILLER_20_1283 ();
 sg13g2_decap_8 FILLER_20_1290 ();
 sg13g2_decap_8 FILLER_20_1297 ();
 sg13g2_decap_8 FILLER_20_1304 ();
 sg13g2_decap_8 FILLER_20_1311 ();
 sg13g2_decap_8 FILLER_20_1318 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_39 ();
 sg13g2_decap_4 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_decap_4 FILLER_21_169 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_191 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_2 FILLER_21_204 ();
 sg13g2_fill_1 FILLER_21_206 ();
 sg13g2_fill_1 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_221 ();
 sg13g2_fill_1 FILLER_21_247 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_decap_4 FILLER_21_317 ();
 sg13g2_fill_1 FILLER_21_321 ();
 sg13g2_fill_2 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_364 ();
 sg13g2_fill_1 FILLER_21_369 ();
 sg13g2_fill_1 FILLER_21_375 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_21_414 ();
 sg13g2_decap_8 FILLER_21_435 ();
 sg13g2_fill_2 FILLER_21_446 ();
 sg13g2_fill_2 FILLER_21_453 ();
 sg13g2_fill_1 FILLER_21_455 ();
 sg13g2_fill_2 FILLER_21_461 ();
 sg13g2_fill_1 FILLER_21_463 ();
 sg13g2_fill_2 FILLER_21_468 ();
 sg13g2_fill_1 FILLER_21_491 ();
 sg13g2_fill_1 FILLER_21_496 ();
 sg13g2_fill_2 FILLER_21_519 ();
 sg13g2_fill_1 FILLER_21_521 ();
 sg13g2_fill_2 FILLER_21_526 ();
 sg13g2_fill_1 FILLER_21_528 ();
 sg13g2_fill_1 FILLER_21_611 ();
 sg13g2_fill_2 FILLER_21_624 ();
 sg13g2_fill_2 FILLER_21_649 ();
 sg13g2_fill_1 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_671 ();
 sg13g2_fill_1 FILLER_21_677 ();
 sg13g2_fill_1 FILLER_21_704 ();
 sg13g2_fill_2 FILLER_21_709 ();
 sg13g2_fill_2 FILLER_21_728 ();
 sg13g2_fill_1 FILLER_21_735 ();
 sg13g2_fill_2 FILLER_21_767 ();
 sg13g2_fill_1 FILLER_21_778 ();
 sg13g2_fill_2 FILLER_21_873 ();
 sg13g2_fill_1 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_884 ();
 sg13g2_fill_2 FILLER_21_890 ();
 sg13g2_fill_1 FILLER_21_917 ();
 sg13g2_decap_4 FILLER_21_935 ();
 sg13g2_fill_2 FILLER_21_939 ();
 sg13g2_decap_8 FILLER_21_945 ();
 sg13g2_fill_2 FILLER_21_952 ();
 sg13g2_fill_2 FILLER_21_962 ();
 sg13g2_fill_2 FILLER_21_982 ();
 sg13g2_fill_1 FILLER_21_996 ();
 sg13g2_fill_2 FILLER_21_1001 ();
 sg13g2_fill_1 FILLER_21_1008 ();
 sg13g2_fill_1 FILLER_21_1026 ();
 sg13g2_fill_1 FILLER_21_1076 ();
 sg13g2_fill_1 FILLER_21_1107 ();
 sg13g2_decap_8 FILLER_21_1112 ();
 sg13g2_decap_8 FILLER_21_1119 ();
 sg13g2_decap_8 FILLER_21_1126 ();
 sg13g2_decap_8 FILLER_21_1133 ();
 sg13g2_decap_8 FILLER_21_1140 ();
 sg13g2_decap_8 FILLER_21_1147 ();
 sg13g2_decap_8 FILLER_21_1154 ();
 sg13g2_decap_8 FILLER_21_1161 ();
 sg13g2_decap_8 FILLER_21_1168 ();
 sg13g2_decap_8 FILLER_21_1175 ();
 sg13g2_decap_8 FILLER_21_1182 ();
 sg13g2_decap_8 FILLER_21_1189 ();
 sg13g2_decap_8 FILLER_21_1196 ();
 sg13g2_decap_8 FILLER_21_1203 ();
 sg13g2_decap_8 FILLER_21_1210 ();
 sg13g2_decap_8 FILLER_21_1217 ();
 sg13g2_decap_8 FILLER_21_1224 ();
 sg13g2_decap_8 FILLER_21_1231 ();
 sg13g2_decap_8 FILLER_21_1238 ();
 sg13g2_decap_8 FILLER_21_1245 ();
 sg13g2_decap_8 FILLER_21_1252 ();
 sg13g2_decap_8 FILLER_21_1259 ();
 sg13g2_decap_8 FILLER_21_1266 ();
 sg13g2_decap_8 FILLER_21_1273 ();
 sg13g2_decap_8 FILLER_21_1280 ();
 sg13g2_decap_8 FILLER_21_1287 ();
 sg13g2_decap_8 FILLER_21_1294 ();
 sg13g2_decap_8 FILLER_21_1301 ();
 sg13g2_decap_8 FILLER_21_1308 ();
 sg13g2_decap_8 FILLER_21_1315 ();
 sg13g2_decap_4 FILLER_21_1322 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_fill_2 FILLER_22_144 ();
 sg13g2_decap_4 FILLER_22_150 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_decap_4 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_290 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_334 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_372 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_fill_2 FILLER_22_383 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_418 ();
 sg13g2_fill_2 FILLER_22_433 ();
 sg13g2_fill_2 FILLER_22_448 ();
 sg13g2_fill_1 FILLER_22_450 ();
 sg13g2_fill_2 FILLER_22_481 ();
 sg13g2_fill_2 FILLER_22_513 ();
 sg13g2_fill_1 FILLER_22_537 ();
 sg13g2_fill_2 FILLER_22_542 ();
 sg13g2_fill_2 FILLER_22_548 ();
 sg13g2_fill_2 FILLER_22_554 ();
 sg13g2_fill_1 FILLER_22_556 ();
 sg13g2_fill_2 FILLER_22_566 ();
 sg13g2_fill_2 FILLER_22_589 ();
 sg13g2_fill_1 FILLER_22_591 ();
 sg13g2_fill_1 FILLER_22_600 ();
 sg13g2_fill_1 FILLER_22_605 ();
 sg13g2_decap_8 FILLER_22_615 ();
 sg13g2_fill_2 FILLER_22_630 ();
 sg13g2_fill_1 FILLER_22_632 ();
 sg13g2_fill_1 FILLER_22_655 ();
 sg13g2_fill_2 FILLER_22_664 ();
 sg13g2_fill_1 FILLER_22_666 ();
 sg13g2_fill_2 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_685 ();
 sg13g2_fill_1 FILLER_22_687 ();
 sg13g2_decap_4 FILLER_22_692 ();
 sg13g2_fill_1 FILLER_22_696 ();
 sg13g2_fill_1 FILLER_22_710 ();
 sg13g2_fill_1 FILLER_22_787 ();
 sg13g2_decap_4 FILLER_22_792 ();
 sg13g2_fill_1 FILLER_22_796 ();
 sg13g2_fill_2 FILLER_22_801 ();
 sg13g2_fill_1 FILLER_22_813 ();
 sg13g2_decap_4 FILLER_22_818 ();
 sg13g2_fill_2 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_828 ();
 sg13g2_fill_1 FILLER_22_855 ();
 sg13g2_fill_2 FILLER_22_870 ();
 sg13g2_fill_1 FILLER_22_872 ();
 sg13g2_fill_1 FILLER_22_889 ();
 sg13g2_fill_1 FILLER_22_916 ();
 sg13g2_fill_1 FILLER_22_921 ();
 sg13g2_fill_1 FILLER_22_952 ();
 sg13g2_fill_1 FILLER_22_978 ();
 sg13g2_fill_2 FILLER_22_983 ();
 sg13g2_fill_1 FILLER_22_1086 ();
 sg13g2_fill_2 FILLER_22_1090 ();
 sg13g2_decap_8 FILLER_22_1096 ();
 sg13g2_decap_8 FILLER_22_1103 ();
 sg13g2_decap_8 FILLER_22_1110 ();
 sg13g2_decap_8 FILLER_22_1117 ();
 sg13g2_decap_8 FILLER_22_1124 ();
 sg13g2_decap_8 FILLER_22_1131 ();
 sg13g2_decap_8 FILLER_22_1138 ();
 sg13g2_decap_8 FILLER_22_1145 ();
 sg13g2_decap_8 FILLER_22_1152 ();
 sg13g2_decap_8 FILLER_22_1159 ();
 sg13g2_decap_8 FILLER_22_1166 ();
 sg13g2_decap_8 FILLER_22_1173 ();
 sg13g2_decap_8 FILLER_22_1180 ();
 sg13g2_decap_8 FILLER_22_1187 ();
 sg13g2_decap_8 FILLER_22_1194 ();
 sg13g2_decap_8 FILLER_22_1201 ();
 sg13g2_decap_8 FILLER_22_1208 ();
 sg13g2_decap_8 FILLER_22_1215 ();
 sg13g2_decap_8 FILLER_22_1222 ();
 sg13g2_decap_8 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1236 ();
 sg13g2_decap_8 FILLER_22_1243 ();
 sg13g2_decap_8 FILLER_22_1250 ();
 sg13g2_decap_8 FILLER_22_1257 ();
 sg13g2_decap_8 FILLER_22_1264 ();
 sg13g2_decap_8 FILLER_22_1271 ();
 sg13g2_decap_8 FILLER_22_1278 ();
 sg13g2_decap_8 FILLER_22_1285 ();
 sg13g2_decap_8 FILLER_22_1292 ();
 sg13g2_decap_8 FILLER_22_1299 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_decap_8 FILLER_22_1313 ();
 sg13g2_decap_4 FILLER_22_1320 ();
 sg13g2_fill_2 FILLER_22_1324 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_4 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_46 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_82 ();
 sg13g2_fill_1 FILLER_23_91 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_228 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_262 ();
 sg13g2_fill_2 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_1 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_335 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_fill_1 FILLER_23_345 ();
 sg13g2_fill_2 FILLER_23_373 ();
 sg13g2_fill_2 FILLER_23_378 ();
 sg13g2_fill_2 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_448 ();
 sg13g2_fill_1 FILLER_23_450 ();
 sg13g2_decap_4 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_471 ();
 sg13g2_fill_1 FILLER_23_478 ();
 sg13g2_fill_2 FILLER_23_483 ();
 sg13g2_fill_1 FILLER_23_485 ();
 sg13g2_fill_2 FILLER_23_498 ();
 sg13g2_fill_1 FILLER_23_517 ();
 sg13g2_fill_2 FILLER_23_522 ();
 sg13g2_fill_2 FILLER_23_555 ();
 sg13g2_fill_2 FILLER_23_583 ();
 sg13g2_fill_1 FILLER_23_642 ();
 sg13g2_fill_2 FILLER_23_668 ();
 sg13g2_fill_2 FILLER_23_674 ();
 sg13g2_fill_1 FILLER_23_676 ();
 sg13g2_fill_1 FILLER_23_703 ();
 sg13g2_fill_1 FILLER_23_709 ();
 sg13g2_fill_1 FILLER_23_715 ();
 sg13g2_fill_1 FILLER_23_724 ();
 sg13g2_fill_2 FILLER_23_785 ();
 sg13g2_fill_1 FILLER_23_880 ();
 sg13g2_fill_1 FILLER_23_907 ();
 sg13g2_fill_2 FILLER_23_913 ();
 sg13g2_fill_2 FILLER_23_919 ();
 sg13g2_decap_8 FILLER_23_925 ();
 sg13g2_fill_2 FILLER_23_936 ();
 sg13g2_fill_1 FILLER_23_965 ();
 sg13g2_fill_1 FILLER_23_992 ();
 sg13g2_fill_1 FILLER_23_1003 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_fill_1 FILLER_23_1020 ();
 sg13g2_fill_2 FILLER_23_1029 ();
 sg13g2_fill_1 FILLER_23_1031 ();
 sg13g2_decap_8 FILLER_23_1035 ();
 sg13g2_fill_2 FILLER_23_1042 ();
 sg13g2_decap_4 FILLER_23_1084 ();
 sg13g2_fill_1 FILLER_23_1088 ();
 sg13g2_decap_8 FILLER_23_1093 ();
 sg13g2_decap_8 FILLER_23_1100 ();
 sg13g2_decap_8 FILLER_23_1107 ();
 sg13g2_decap_8 FILLER_23_1114 ();
 sg13g2_decap_8 FILLER_23_1121 ();
 sg13g2_decap_8 FILLER_23_1128 ();
 sg13g2_decap_8 FILLER_23_1135 ();
 sg13g2_decap_8 FILLER_23_1142 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_decap_8 FILLER_23_1156 ();
 sg13g2_decap_8 FILLER_23_1163 ();
 sg13g2_decap_8 FILLER_23_1170 ();
 sg13g2_decap_8 FILLER_23_1177 ();
 sg13g2_decap_8 FILLER_23_1184 ();
 sg13g2_decap_8 FILLER_23_1191 ();
 sg13g2_decap_8 FILLER_23_1198 ();
 sg13g2_decap_8 FILLER_23_1205 ();
 sg13g2_decap_8 FILLER_23_1212 ();
 sg13g2_decap_8 FILLER_23_1219 ();
 sg13g2_decap_8 FILLER_23_1226 ();
 sg13g2_decap_8 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1240 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1261 ();
 sg13g2_decap_8 FILLER_23_1268 ();
 sg13g2_decap_8 FILLER_23_1275 ();
 sg13g2_decap_8 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_decap_8 FILLER_23_1296 ();
 sg13g2_decap_8 FILLER_23_1303 ();
 sg13g2_decap_8 FILLER_23_1310 ();
 sg13g2_decap_8 FILLER_23_1317 ();
 sg13g2_fill_2 FILLER_23_1324 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_44 ();
 sg13g2_decap_8 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_78 ();
 sg13g2_fill_2 FILLER_24_132 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_329 ();
 sg13g2_fill_1 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_394 ();
 sg13g2_fill_1 FILLER_24_400 ();
 sg13g2_fill_1 FILLER_24_406 ();
 sg13g2_decap_4 FILLER_24_444 ();
 sg13g2_fill_2 FILLER_24_458 ();
 sg13g2_fill_1 FILLER_24_460 ();
 sg13g2_fill_1 FILLER_24_495 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_fill_1 FILLER_24_547 ();
 sg13g2_fill_1 FILLER_24_552 ();
 sg13g2_fill_1 FILLER_24_557 ();
 sg13g2_fill_2 FILLER_24_606 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_fill_1 FILLER_24_618 ();
 sg13g2_fill_2 FILLER_24_627 ();
 sg13g2_fill_1 FILLER_24_633 ();
 sg13g2_fill_1 FILLER_24_639 ();
 sg13g2_fill_1 FILLER_24_645 ();
 sg13g2_fill_2 FILLER_24_651 ();
 sg13g2_fill_2 FILLER_24_657 ();
 sg13g2_fill_1 FILLER_24_693 ();
 sg13g2_fill_1 FILLER_24_702 ();
 sg13g2_fill_1 FILLER_24_730 ();
 sg13g2_fill_2 FILLER_24_735 ();
 sg13g2_fill_1 FILLER_24_763 ();
 sg13g2_fill_1 FILLER_24_779 ();
 sg13g2_fill_1 FILLER_24_797 ();
 sg13g2_decap_4 FILLER_24_802 ();
 sg13g2_fill_2 FILLER_24_806 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_4 FILLER_24_823 ();
 sg13g2_fill_2 FILLER_24_827 ();
 sg13g2_fill_1 FILLER_24_855 ();
 sg13g2_fill_1 FILLER_24_873 ();
 sg13g2_fill_1 FILLER_24_882 ();
 sg13g2_fill_2 FILLER_24_888 ();
 sg13g2_decap_4 FILLER_24_929 ();
 sg13g2_decap_4 FILLER_24_937 ();
 sg13g2_decap_4 FILLER_24_983 ();
 sg13g2_decap_8 FILLER_24_1035 ();
 sg13g2_fill_2 FILLER_24_1042 ();
 sg13g2_fill_1 FILLER_24_1044 ();
 sg13g2_fill_2 FILLER_24_1070 ();
 sg13g2_fill_1 FILLER_24_1080 ();
 sg13g2_fill_2 FILLER_24_1090 ();
 sg13g2_fill_1 FILLER_24_1092 ();
 sg13g2_decap_8 FILLER_24_1097 ();
 sg13g2_decap_8 FILLER_24_1104 ();
 sg13g2_decap_8 FILLER_24_1111 ();
 sg13g2_decap_8 FILLER_24_1118 ();
 sg13g2_decap_8 FILLER_24_1125 ();
 sg13g2_decap_8 FILLER_24_1132 ();
 sg13g2_decap_8 FILLER_24_1139 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1153 ();
 sg13g2_decap_8 FILLER_24_1160 ();
 sg13g2_decap_8 FILLER_24_1167 ();
 sg13g2_decap_8 FILLER_24_1174 ();
 sg13g2_decap_8 FILLER_24_1181 ();
 sg13g2_decap_8 FILLER_24_1188 ();
 sg13g2_decap_8 FILLER_24_1195 ();
 sg13g2_decap_8 FILLER_24_1202 ();
 sg13g2_decap_8 FILLER_24_1209 ();
 sg13g2_decap_8 FILLER_24_1216 ();
 sg13g2_decap_8 FILLER_24_1223 ();
 sg13g2_decap_8 FILLER_24_1230 ();
 sg13g2_decap_8 FILLER_24_1237 ();
 sg13g2_decap_8 FILLER_24_1244 ();
 sg13g2_decap_8 FILLER_24_1251 ();
 sg13g2_decap_8 FILLER_24_1258 ();
 sg13g2_decap_8 FILLER_24_1265 ();
 sg13g2_decap_8 FILLER_24_1272 ();
 sg13g2_decap_8 FILLER_24_1279 ();
 sg13g2_decap_8 FILLER_24_1286 ();
 sg13g2_decap_8 FILLER_24_1293 ();
 sg13g2_decap_8 FILLER_24_1300 ();
 sg13g2_decap_8 FILLER_24_1307 ();
 sg13g2_decap_8 FILLER_24_1314 ();
 sg13g2_decap_4 FILLER_24_1321 ();
 sg13g2_fill_1 FILLER_24_1325 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_4 FILLER_25_49 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_210 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_2 FILLER_25_263 ();
 sg13g2_fill_1 FILLER_25_269 ();
 sg13g2_fill_2 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_314 ();
 sg13g2_fill_1 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_395 ();
 sg13g2_fill_1 FILLER_25_468 ();
 sg13g2_decap_4 FILLER_25_472 ();
 sg13g2_fill_2 FILLER_25_561 ();
 sg13g2_fill_1 FILLER_25_563 ();
 sg13g2_fill_2 FILLER_25_568 ();
 sg13g2_fill_1 FILLER_25_570 ();
 sg13g2_fill_2 FILLER_25_639 ();
 sg13g2_fill_1 FILLER_25_648 ();
 sg13g2_fill_1 FILLER_25_654 ();
 sg13g2_fill_1 FILLER_25_661 ();
 sg13g2_fill_1 FILLER_25_667 ();
 sg13g2_fill_1 FILLER_25_676 ();
 sg13g2_fill_2 FILLER_25_704 ();
 sg13g2_fill_1 FILLER_25_710 ();
 sg13g2_fill_1 FILLER_25_717 ();
 sg13g2_fill_2 FILLER_25_722 ();
 sg13g2_fill_1 FILLER_25_730 ();
 sg13g2_fill_1 FILLER_25_739 ();
 sg13g2_fill_2 FILLER_25_747 ();
 sg13g2_fill_1 FILLER_25_749 ();
 sg13g2_fill_2 FILLER_25_773 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_1 FILLER_25_858 ();
 sg13g2_decap_4 FILLER_25_864 ();
 sg13g2_fill_1 FILLER_25_878 ();
 sg13g2_fill_2 FILLER_25_883 ();
 sg13g2_fill_1 FILLER_25_914 ();
 sg13g2_fill_2 FILLER_25_972 ();
 sg13g2_fill_2 FILLER_25_978 ();
 sg13g2_fill_1 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1057 ();
 sg13g2_fill_1 FILLER_25_1059 ();
 sg13g2_fill_2 FILLER_25_1064 ();
 sg13g2_fill_2 FILLER_25_1070 ();
 sg13g2_decap_4 FILLER_25_1077 ();
 sg13g2_fill_2 FILLER_25_1081 ();
 sg13g2_decap_8 FILLER_25_1109 ();
 sg13g2_decap_8 FILLER_25_1116 ();
 sg13g2_decap_8 FILLER_25_1123 ();
 sg13g2_decap_8 FILLER_25_1130 ();
 sg13g2_decap_8 FILLER_25_1137 ();
 sg13g2_decap_8 FILLER_25_1144 ();
 sg13g2_decap_8 FILLER_25_1151 ();
 sg13g2_decap_8 FILLER_25_1158 ();
 sg13g2_decap_8 FILLER_25_1165 ();
 sg13g2_decap_8 FILLER_25_1172 ();
 sg13g2_decap_8 FILLER_25_1179 ();
 sg13g2_decap_8 FILLER_25_1186 ();
 sg13g2_decap_8 FILLER_25_1193 ();
 sg13g2_decap_8 FILLER_25_1200 ();
 sg13g2_decap_8 FILLER_25_1207 ();
 sg13g2_decap_8 FILLER_25_1214 ();
 sg13g2_decap_8 FILLER_25_1221 ();
 sg13g2_decap_8 FILLER_25_1228 ();
 sg13g2_decap_8 FILLER_25_1235 ();
 sg13g2_decap_8 FILLER_25_1242 ();
 sg13g2_decap_8 FILLER_25_1249 ();
 sg13g2_decap_8 FILLER_25_1256 ();
 sg13g2_decap_8 FILLER_25_1263 ();
 sg13g2_decap_8 FILLER_25_1270 ();
 sg13g2_decap_8 FILLER_25_1277 ();
 sg13g2_decap_8 FILLER_25_1284 ();
 sg13g2_decap_8 FILLER_25_1291 ();
 sg13g2_decap_8 FILLER_25_1298 ();
 sg13g2_decap_8 FILLER_25_1305 ();
 sg13g2_decap_8 FILLER_25_1312 ();
 sg13g2_decap_8 FILLER_25_1319 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_fill_2 FILLER_26_86 ();
 sg13g2_decap_4 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_133 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_fill_2 FILLER_26_175 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_2 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_281 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_300 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_343 ();
 sg13g2_fill_2 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_394 ();
 sg13g2_fill_1 FILLER_26_426 ();
 sg13g2_fill_1 FILLER_26_455 ();
 sg13g2_fill_1 FILLER_26_460 ();
 sg13g2_fill_1 FILLER_26_473 ();
 sg13g2_fill_2 FILLER_26_513 ();
 sg13g2_fill_1 FILLER_26_515 ();
 sg13g2_fill_1 FILLER_26_521 ();
 sg13g2_decap_4 FILLER_26_534 ();
 sg13g2_fill_2 FILLER_26_538 ();
 sg13g2_fill_2 FILLER_26_544 ();
 sg13g2_fill_2 FILLER_26_572 ();
 sg13g2_fill_1 FILLER_26_578 ();
 sg13g2_fill_1 FILLER_26_583 ();
 sg13g2_fill_1 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_599 ();
 sg13g2_fill_2 FILLER_26_604 ();
 sg13g2_fill_1 FILLER_26_610 ();
 sg13g2_decap_4 FILLER_26_623 ();
 sg13g2_fill_2 FILLER_26_627 ();
 sg13g2_fill_1 FILLER_26_658 ();
 sg13g2_fill_2 FILLER_26_685 ();
 sg13g2_fill_2 FILLER_26_707 ();
 sg13g2_fill_1 FILLER_26_734 ();
 sg13g2_decap_4 FILLER_26_751 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_fill_2 FILLER_26_826 ();
 sg13g2_fill_1 FILLER_26_828 ();
 sg13g2_fill_1 FILLER_26_833 ();
 sg13g2_decap_4 FILLER_26_838 ();
 sg13g2_fill_2 FILLER_26_842 ();
 sg13g2_fill_2 FILLER_26_853 ();
 sg13g2_fill_1 FILLER_26_855 ();
 sg13g2_fill_2 FILLER_26_864 ();
 sg13g2_fill_2 FILLER_26_889 ();
 sg13g2_fill_2 FILLER_26_895 ();
 sg13g2_fill_2 FILLER_26_919 ();
 sg13g2_fill_1 FILLER_26_947 ();
 sg13g2_fill_1 FILLER_26_963 ();
 sg13g2_fill_2 FILLER_26_979 ();
 sg13g2_fill_1 FILLER_26_1010 ();
 sg13g2_fill_2 FILLER_26_1044 ();
 sg13g2_fill_1 FILLER_26_1059 ();
 sg13g2_decap_8 FILLER_26_1102 ();
 sg13g2_decap_8 FILLER_26_1109 ();
 sg13g2_decap_8 FILLER_26_1116 ();
 sg13g2_decap_8 FILLER_26_1123 ();
 sg13g2_decap_8 FILLER_26_1130 ();
 sg13g2_decap_8 FILLER_26_1137 ();
 sg13g2_decap_8 FILLER_26_1144 ();
 sg13g2_decap_8 FILLER_26_1151 ();
 sg13g2_decap_8 FILLER_26_1158 ();
 sg13g2_decap_8 FILLER_26_1165 ();
 sg13g2_decap_8 FILLER_26_1172 ();
 sg13g2_decap_8 FILLER_26_1179 ();
 sg13g2_decap_8 FILLER_26_1186 ();
 sg13g2_decap_8 FILLER_26_1193 ();
 sg13g2_decap_8 FILLER_26_1200 ();
 sg13g2_decap_8 FILLER_26_1207 ();
 sg13g2_decap_8 FILLER_26_1214 ();
 sg13g2_decap_8 FILLER_26_1221 ();
 sg13g2_decap_8 FILLER_26_1228 ();
 sg13g2_decap_8 FILLER_26_1235 ();
 sg13g2_decap_8 FILLER_26_1242 ();
 sg13g2_decap_8 FILLER_26_1249 ();
 sg13g2_decap_8 FILLER_26_1256 ();
 sg13g2_decap_8 FILLER_26_1263 ();
 sg13g2_decap_8 FILLER_26_1270 ();
 sg13g2_decap_8 FILLER_26_1277 ();
 sg13g2_decap_8 FILLER_26_1284 ();
 sg13g2_decap_8 FILLER_26_1291 ();
 sg13g2_decap_8 FILLER_26_1298 ();
 sg13g2_decap_8 FILLER_26_1305 ();
 sg13g2_decap_8 FILLER_26_1312 ();
 sg13g2_decap_8 FILLER_26_1319 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_188 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_211 ();
 sg13g2_decap_4 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_decap_4 FILLER_27_260 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_fill_2 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_330 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_1 FILLER_27_409 ();
 sg13g2_fill_1 FILLER_27_512 ();
 sg13g2_fill_2 FILLER_27_594 ();
 sg13g2_fill_1 FILLER_27_596 ();
 sg13g2_fill_2 FILLER_27_643 ();
 sg13g2_fill_2 FILLER_27_649 ();
 sg13g2_decap_4 FILLER_27_661 ();
 sg13g2_fill_2 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_671 ();
 sg13g2_decap_4 FILLER_27_678 ();
 sg13g2_fill_1 FILLER_27_682 ();
 sg13g2_fill_2 FILLER_27_687 ();
 sg13g2_fill_1 FILLER_27_689 ();
 sg13g2_fill_2 FILLER_27_791 ();
 sg13g2_fill_1 FILLER_27_832 ();
 sg13g2_fill_2 FILLER_27_863 ();
 sg13g2_fill_1 FILLER_27_878 ();
 sg13g2_fill_1 FILLER_27_893 ();
 sg13g2_fill_1 FILLER_27_963 ();
 sg13g2_fill_1 FILLER_27_977 ();
 sg13g2_fill_1 FILLER_27_982 ();
 sg13g2_fill_2 FILLER_27_988 ();
 sg13g2_decap_8 FILLER_27_1020 ();
 sg13g2_fill_1 FILLER_27_1027 ();
 sg13g2_fill_2 FILLER_27_1038 ();
 sg13g2_fill_1 FILLER_27_1045 ();
 sg13g2_decap_8 FILLER_27_1090 ();
 sg13g2_decap_8 FILLER_27_1097 ();
 sg13g2_decap_8 FILLER_27_1104 ();
 sg13g2_decap_8 FILLER_27_1111 ();
 sg13g2_decap_8 FILLER_27_1118 ();
 sg13g2_decap_8 FILLER_27_1125 ();
 sg13g2_decap_8 FILLER_27_1132 ();
 sg13g2_decap_8 FILLER_27_1139 ();
 sg13g2_decap_8 FILLER_27_1146 ();
 sg13g2_decap_8 FILLER_27_1153 ();
 sg13g2_decap_8 FILLER_27_1160 ();
 sg13g2_decap_8 FILLER_27_1167 ();
 sg13g2_decap_8 FILLER_27_1174 ();
 sg13g2_decap_8 FILLER_27_1181 ();
 sg13g2_decap_8 FILLER_27_1188 ();
 sg13g2_decap_8 FILLER_27_1195 ();
 sg13g2_decap_8 FILLER_27_1202 ();
 sg13g2_decap_8 FILLER_27_1209 ();
 sg13g2_decap_8 FILLER_27_1216 ();
 sg13g2_decap_8 FILLER_27_1223 ();
 sg13g2_decap_8 FILLER_27_1230 ();
 sg13g2_decap_8 FILLER_27_1237 ();
 sg13g2_decap_8 FILLER_27_1244 ();
 sg13g2_decap_8 FILLER_27_1251 ();
 sg13g2_decap_8 FILLER_27_1258 ();
 sg13g2_decap_8 FILLER_27_1265 ();
 sg13g2_decap_8 FILLER_27_1272 ();
 sg13g2_decap_8 FILLER_27_1279 ();
 sg13g2_decap_8 FILLER_27_1286 ();
 sg13g2_decap_8 FILLER_27_1293 ();
 sg13g2_decap_8 FILLER_27_1300 ();
 sg13g2_decap_8 FILLER_27_1307 ();
 sg13g2_decap_8 FILLER_27_1314 ();
 sg13g2_decap_4 FILLER_27_1321 ();
 sg13g2_fill_1 FILLER_27_1325 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_fill_1 FILLER_28_213 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_fill_2 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_2 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_345 ();
 sg13g2_fill_2 FILLER_28_354 ();
 sg13g2_fill_1 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_383 ();
 sg13g2_fill_2 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_433 ();
 sg13g2_fill_1 FILLER_28_442 ();
 sg13g2_decap_4 FILLER_28_471 ();
 sg13g2_fill_2 FILLER_28_530 ();
 sg13g2_fill_2 FILLER_28_541 ();
 sg13g2_fill_2 FILLER_28_590 ();
 sg13g2_fill_1 FILLER_28_608 ();
 sg13g2_fill_1 FILLER_28_639 ();
 sg13g2_fill_1 FILLER_28_678 ();
 sg13g2_fill_2 FILLER_28_683 ();
 sg13g2_fill_2 FILLER_28_695 ();
 sg13g2_fill_1 FILLER_28_697 ();
 sg13g2_fill_1 FILLER_28_716 ();
 sg13g2_fill_2 FILLER_28_721 ();
 sg13g2_fill_2 FILLER_28_728 ();
 sg13g2_fill_2 FILLER_28_734 ();
 sg13g2_fill_1 FILLER_28_736 ();
 sg13g2_fill_1 FILLER_28_741 ();
 sg13g2_fill_2 FILLER_28_747 ();
 sg13g2_fill_1 FILLER_28_749 ();
 sg13g2_fill_2 FILLER_28_773 ();
 sg13g2_fill_2 FILLER_28_809 ();
 sg13g2_decap_4 FILLER_28_841 ();
 sg13g2_fill_1 FILLER_28_845 ();
 sg13g2_decap_4 FILLER_28_850 ();
 sg13g2_fill_2 FILLER_28_867 ();
 sg13g2_fill_1 FILLER_28_900 ();
 sg13g2_fill_1 FILLER_28_906 ();
 sg13g2_fill_2 FILLER_28_936 ();
 sg13g2_fill_1 FILLER_28_942 ();
 sg13g2_fill_1 FILLER_28_948 ();
 sg13g2_fill_1 FILLER_28_965 ();
 sg13g2_fill_1 FILLER_28_979 ();
 sg13g2_fill_2 FILLER_28_1054 ();
 sg13g2_fill_1 FILLER_28_1056 ();
 sg13g2_fill_2 FILLER_28_1065 ();
 sg13g2_fill_1 FILLER_28_1067 ();
 sg13g2_decap_8 FILLER_28_1085 ();
 sg13g2_decap_8 FILLER_28_1092 ();
 sg13g2_decap_8 FILLER_28_1099 ();
 sg13g2_decap_8 FILLER_28_1106 ();
 sg13g2_decap_8 FILLER_28_1113 ();
 sg13g2_decap_8 FILLER_28_1120 ();
 sg13g2_decap_8 FILLER_28_1127 ();
 sg13g2_decap_8 FILLER_28_1134 ();
 sg13g2_decap_8 FILLER_28_1141 ();
 sg13g2_decap_8 FILLER_28_1148 ();
 sg13g2_decap_8 FILLER_28_1155 ();
 sg13g2_decap_8 FILLER_28_1162 ();
 sg13g2_decap_8 FILLER_28_1169 ();
 sg13g2_decap_8 FILLER_28_1176 ();
 sg13g2_decap_8 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1190 ();
 sg13g2_decap_8 FILLER_28_1197 ();
 sg13g2_decap_8 FILLER_28_1204 ();
 sg13g2_decap_8 FILLER_28_1211 ();
 sg13g2_decap_8 FILLER_28_1218 ();
 sg13g2_decap_8 FILLER_28_1225 ();
 sg13g2_decap_8 FILLER_28_1232 ();
 sg13g2_decap_8 FILLER_28_1239 ();
 sg13g2_decap_8 FILLER_28_1246 ();
 sg13g2_decap_8 FILLER_28_1253 ();
 sg13g2_decap_8 FILLER_28_1260 ();
 sg13g2_decap_8 FILLER_28_1267 ();
 sg13g2_decap_8 FILLER_28_1274 ();
 sg13g2_decap_8 FILLER_28_1281 ();
 sg13g2_decap_8 FILLER_28_1288 ();
 sg13g2_decap_8 FILLER_28_1295 ();
 sg13g2_decap_8 FILLER_28_1302 ();
 sg13g2_decap_8 FILLER_28_1309 ();
 sg13g2_decap_8 FILLER_28_1316 ();
 sg13g2_fill_2 FILLER_28_1323 ();
 sg13g2_fill_1 FILLER_28_1325 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_59 ();
 sg13g2_decap_8 FILLER_29_66 ();
 sg13g2_decap_4 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_112 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_fill_2 FILLER_29_193 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_339 ();
 sg13g2_fill_1 FILLER_29_419 ();
 sg13g2_fill_1 FILLER_29_437 ();
 sg13g2_fill_2 FILLER_29_446 ();
 sg13g2_fill_2 FILLER_29_457 ();
 sg13g2_fill_1 FILLER_29_459 ();
 sg13g2_fill_2 FILLER_29_464 ();
 sg13g2_fill_1 FILLER_29_475 ();
 sg13g2_fill_1 FILLER_29_481 ();
 sg13g2_fill_1 FILLER_29_499 ();
 sg13g2_decap_4 FILLER_29_547 ();
 sg13g2_fill_1 FILLER_29_551 ();
 sg13g2_decap_4 FILLER_29_681 ();
 sg13g2_fill_1 FILLER_29_685 ();
 sg13g2_fill_1 FILLER_29_778 ();
 sg13g2_fill_2 FILLER_29_796 ();
 sg13g2_fill_2 FILLER_29_811 ();
 sg13g2_fill_1 FILLER_29_865 ();
 sg13g2_fill_1 FILLER_29_889 ();
 sg13g2_fill_1 FILLER_29_963 ();
 sg13g2_fill_1 FILLER_29_975 ();
 sg13g2_fill_2 FILLER_29_1024 ();
 sg13g2_fill_1 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1031 ();
 sg13g2_fill_1 FILLER_29_1037 ();
 sg13g2_fill_2 FILLER_29_1056 ();
 sg13g2_fill_1 FILLER_29_1063 ();
 sg13g2_decap_8 FILLER_29_1094 ();
 sg13g2_decap_8 FILLER_29_1101 ();
 sg13g2_decap_8 FILLER_29_1108 ();
 sg13g2_decap_8 FILLER_29_1115 ();
 sg13g2_decap_8 FILLER_29_1122 ();
 sg13g2_decap_8 FILLER_29_1129 ();
 sg13g2_decap_8 FILLER_29_1136 ();
 sg13g2_decap_8 FILLER_29_1143 ();
 sg13g2_decap_8 FILLER_29_1150 ();
 sg13g2_decap_8 FILLER_29_1157 ();
 sg13g2_decap_8 FILLER_29_1164 ();
 sg13g2_decap_8 FILLER_29_1171 ();
 sg13g2_decap_8 FILLER_29_1178 ();
 sg13g2_decap_8 FILLER_29_1185 ();
 sg13g2_decap_8 FILLER_29_1192 ();
 sg13g2_decap_8 FILLER_29_1199 ();
 sg13g2_decap_8 FILLER_29_1206 ();
 sg13g2_decap_8 FILLER_29_1213 ();
 sg13g2_decap_8 FILLER_29_1220 ();
 sg13g2_decap_8 FILLER_29_1227 ();
 sg13g2_decap_8 FILLER_29_1234 ();
 sg13g2_decap_8 FILLER_29_1241 ();
 sg13g2_decap_8 FILLER_29_1248 ();
 sg13g2_decap_8 FILLER_29_1255 ();
 sg13g2_decap_8 FILLER_29_1262 ();
 sg13g2_decap_8 FILLER_29_1269 ();
 sg13g2_decap_8 FILLER_29_1276 ();
 sg13g2_decap_8 FILLER_29_1283 ();
 sg13g2_decap_8 FILLER_29_1290 ();
 sg13g2_decap_8 FILLER_29_1297 ();
 sg13g2_decap_8 FILLER_29_1304 ();
 sg13g2_decap_8 FILLER_29_1311 ();
 sg13g2_decap_8 FILLER_29_1318 ();
 sg13g2_fill_1 FILLER_29_1325 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_88 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_fill_2 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_111 ();
 sg13g2_fill_1 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_1 FILLER_30_155 ();
 sg13g2_fill_1 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_178 ();
 sg13g2_decap_4 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_386 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_fill_1 FILLER_30_433 ();
 sg13g2_fill_1 FILLER_30_439 ();
 sg13g2_fill_1 FILLER_30_474 ();
 sg13g2_fill_2 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_508 ();
 sg13g2_fill_2 FILLER_30_513 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_fill_2 FILLER_30_525 ();
 sg13g2_fill_1 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_558 ();
 sg13g2_fill_2 FILLER_30_603 ();
 sg13g2_fill_1 FILLER_30_605 ();
 sg13g2_fill_1 FILLER_30_610 ();
 sg13g2_decap_8 FILLER_30_641 ();
 sg13g2_fill_2 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_fill_2 FILLER_30_662 ();
 sg13g2_fill_1 FILLER_30_671 ();
 sg13g2_fill_2 FILLER_30_682 ();
 sg13g2_fill_1 FILLER_30_684 ();
 sg13g2_fill_1 FILLER_30_705 ();
 sg13g2_fill_1 FILLER_30_748 ();
 sg13g2_fill_1 FILLER_30_757 ();
 sg13g2_fill_1 FILLER_30_768 ();
 sg13g2_fill_2 FILLER_30_781 ();
 sg13g2_fill_2 FILLER_30_795 ();
 sg13g2_fill_1 FILLER_30_828 ();
 sg13g2_fill_1 FILLER_30_833 ();
 sg13g2_fill_1 FILLER_30_844 ();
 sg13g2_fill_1 FILLER_30_873 ();
 sg13g2_fill_2 FILLER_30_898 ();
 sg13g2_fill_2 FILLER_30_904 ();
 sg13g2_decap_4 FILLER_30_915 ();
 sg13g2_fill_1 FILLER_30_932 ();
 sg13g2_fill_2 FILLER_30_941 ();
 sg13g2_fill_2 FILLER_30_955 ();
 sg13g2_fill_1 FILLER_30_972 ();
 sg13g2_fill_2 FILLER_30_1020 ();
 sg13g2_fill_1 FILLER_30_1066 ();
 sg13g2_decap_8 FILLER_30_1097 ();
 sg13g2_decap_8 FILLER_30_1104 ();
 sg13g2_decap_8 FILLER_30_1111 ();
 sg13g2_decap_8 FILLER_30_1118 ();
 sg13g2_decap_8 FILLER_30_1125 ();
 sg13g2_decap_8 FILLER_30_1132 ();
 sg13g2_decap_8 FILLER_30_1139 ();
 sg13g2_decap_8 FILLER_30_1146 ();
 sg13g2_decap_8 FILLER_30_1153 ();
 sg13g2_decap_8 FILLER_30_1160 ();
 sg13g2_decap_8 FILLER_30_1167 ();
 sg13g2_decap_8 FILLER_30_1174 ();
 sg13g2_decap_8 FILLER_30_1181 ();
 sg13g2_decap_8 FILLER_30_1188 ();
 sg13g2_decap_8 FILLER_30_1195 ();
 sg13g2_decap_8 FILLER_30_1202 ();
 sg13g2_decap_8 FILLER_30_1209 ();
 sg13g2_decap_8 FILLER_30_1216 ();
 sg13g2_decap_8 FILLER_30_1223 ();
 sg13g2_decap_8 FILLER_30_1230 ();
 sg13g2_decap_8 FILLER_30_1237 ();
 sg13g2_decap_8 FILLER_30_1244 ();
 sg13g2_decap_8 FILLER_30_1251 ();
 sg13g2_decap_8 FILLER_30_1258 ();
 sg13g2_decap_8 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1272 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_decap_8 FILLER_30_1286 ();
 sg13g2_decap_8 FILLER_30_1293 ();
 sg13g2_decap_8 FILLER_30_1300 ();
 sg13g2_decap_8 FILLER_30_1307 ();
 sg13g2_decap_8 FILLER_30_1314 ();
 sg13g2_decap_4 FILLER_30_1321 ();
 sg13g2_fill_1 FILLER_30_1325 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_2 FILLER_31_141 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_fill_2 FILLER_31_463 ();
 sg13g2_decap_4 FILLER_31_469 ();
 sg13g2_fill_2 FILLER_31_473 ();
 sg13g2_fill_2 FILLER_31_480 ();
 sg13g2_fill_1 FILLER_31_538 ();
 sg13g2_fill_2 FILLER_31_599 ();
 sg13g2_fill_2 FILLER_31_605 ();
 sg13g2_fill_1 FILLER_31_607 ();
 sg13g2_fill_2 FILLER_31_627 ();
 sg13g2_fill_1 FILLER_31_689 ();
 sg13g2_fill_1 FILLER_31_704 ();
 sg13g2_fill_2 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_738 ();
 sg13g2_fill_2 FILLER_31_745 ();
 sg13g2_fill_2 FILLER_31_820 ();
 sg13g2_fill_2 FILLER_31_848 ();
 sg13g2_fill_2 FILLER_31_959 ();
 sg13g2_fill_1 FILLER_31_971 ();
 sg13g2_fill_2 FILLER_31_996 ();
 sg13g2_fill_1 FILLER_31_998 ();
 sg13g2_fill_2 FILLER_31_1054 ();
 sg13g2_fill_1 FILLER_31_1069 ();
 sg13g2_decap_8 FILLER_31_1087 ();
 sg13g2_decap_8 FILLER_31_1094 ();
 sg13g2_decap_8 FILLER_31_1101 ();
 sg13g2_decap_8 FILLER_31_1108 ();
 sg13g2_decap_8 FILLER_31_1115 ();
 sg13g2_decap_8 FILLER_31_1122 ();
 sg13g2_decap_8 FILLER_31_1129 ();
 sg13g2_decap_8 FILLER_31_1136 ();
 sg13g2_decap_8 FILLER_31_1143 ();
 sg13g2_decap_8 FILLER_31_1150 ();
 sg13g2_decap_8 FILLER_31_1157 ();
 sg13g2_decap_8 FILLER_31_1164 ();
 sg13g2_decap_8 FILLER_31_1171 ();
 sg13g2_decap_8 FILLER_31_1178 ();
 sg13g2_decap_8 FILLER_31_1185 ();
 sg13g2_decap_8 FILLER_31_1192 ();
 sg13g2_decap_8 FILLER_31_1199 ();
 sg13g2_decap_8 FILLER_31_1206 ();
 sg13g2_decap_8 FILLER_31_1213 ();
 sg13g2_decap_8 FILLER_31_1220 ();
 sg13g2_decap_8 FILLER_31_1227 ();
 sg13g2_decap_8 FILLER_31_1234 ();
 sg13g2_decap_8 FILLER_31_1241 ();
 sg13g2_decap_8 FILLER_31_1248 ();
 sg13g2_decap_8 FILLER_31_1255 ();
 sg13g2_decap_8 FILLER_31_1262 ();
 sg13g2_decap_8 FILLER_31_1269 ();
 sg13g2_decap_8 FILLER_31_1276 ();
 sg13g2_decap_8 FILLER_31_1283 ();
 sg13g2_decap_8 FILLER_31_1290 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_decap_8 FILLER_31_1311 ();
 sg13g2_decap_8 FILLER_31_1318 ();
 sg13g2_fill_1 FILLER_31_1325 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_112 ();
 sg13g2_decap_4 FILLER_32_118 ();
 sg13g2_fill_1 FILLER_32_122 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_194 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_decap_4 FILLER_32_217 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_fill_2 FILLER_32_245 ();
 sg13g2_fill_1 FILLER_32_253 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_271 ();
 sg13g2_fill_1 FILLER_32_278 ();
 sg13g2_fill_1 FILLER_32_354 ();
 sg13g2_fill_2 FILLER_32_385 ();
 sg13g2_fill_2 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_424 ();
 sg13g2_decap_4 FILLER_32_500 ();
 sg13g2_decap_4 FILLER_32_508 ();
 sg13g2_fill_1 FILLER_32_529 ();
 sg13g2_fill_1 FILLER_32_538 ();
 sg13g2_fill_2 FILLER_32_561 ();
 sg13g2_fill_1 FILLER_32_563 ();
 sg13g2_fill_2 FILLER_32_640 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_fill_1 FILLER_32_658 ();
 sg13g2_decap_4 FILLER_32_663 ();
 sg13g2_fill_1 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_676 ();
 sg13g2_fill_2 FILLER_32_681 ();
 sg13g2_fill_1 FILLER_32_687 ();
 sg13g2_fill_1 FILLER_32_721 ();
 sg13g2_fill_2 FILLER_32_774 ();
 sg13g2_fill_1 FILLER_32_787 ();
 sg13g2_fill_2 FILLER_32_798 ();
 sg13g2_fill_2 FILLER_32_883 ();
 sg13g2_fill_1 FILLER_32_913 ();
 sg13g2_fill_1 FILLER_32_922 ();
 sg13g2_fill_1 FILLER_32_954 ();
 sg13g2_fill_1 FILLER_32_980 ();
 sg13g2_fill_1 FILLER_32_1007 ();
 sg13g2_fill_1 FILLER_32_1012 ();
 sg13g2_fill_1 FILLER_32_1017 ();
 sg13g2_fill_1 FILLER_32_1023 ();
 sg13g2_fill_2 FILLER_32_1034 ();
 sg13g2_fill_1 FILLER_32_1036 ();
 sg13g2_fill_1 FILLER_32_1042 ();
 sg13g2_decap_8 FILLER_32_1098 ();
 sg13g2_decap_8 FILLER_32_1105 ();
 sg13g2_decap_8 FILLER_32_1112 ();
 sg13g2_decap_8 FILLER_32_1119 ();
 sg13g2_decap_8 FILLER_32_1126 ();
 sg13g2_decap_8 FILLER_32_1133 ();
 sg13g2_decap_8 FILLER_32_1140 ();
 sg13g2_decap_8 FILLER_32_1147 ();
 sg13g2_decap_8 FILLER_32_1154 ();
 sg13g2_decap_8 FILLER_32_1161 ();
 sg13g2_decap_8 FILLER_32_1168 ();
 sg13g2_decap_8 FILLER_32_1175 ();
 sg13g2_decap_8 FILLER_32_1182 ();
 sg13g2_decap_8 FILLER_32_1189 ();
 sg13g2_decap_8 FILLER_32_1196 ();
 sg13g2_decap_8 FILLER_32_1203 ();
 sg13g2_decap_8 FILLER_32_1210 ();
 sg13g2_decap_8 FILLER_32_1217 ();
 sg13g2_decap_8 FILLER_32_1224 ();
 sg13g2_decap_8 FILLER_32_1231 ();
 sg13g2_decap_8 FILLER_32_1238 ();
 sg13g2_decap_8 FILLER_32_1245 ();
 sg13g2_decap_8 FILLER_32_1252 ();
 sg13g2_decap_8 FILLER_32_1259 ();
 sg13g2_decap_8 FILLER_32_1266 ();
 sg13g2_decap_8 FILLER_32_1273 ();
 sg13g2_decap_8 FILLER_32_1280 ();
 sg13g2_decap_8 FILLER_32_1287 ();
 sg13g2_decap_8 FILLER_32_1294 ();
 sg13g2_decap_8 FILLER_32_1301 ();
 sg13g2_decap_8 FILLER_32_1308 ();
 sg13g2_decap_8 FILLER_32_1315 ();
 sg13g2_decap_4 FILLER_32_1322 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_132 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_260 ();
 sg13g2_decap_4 FILLER_33_292 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_decap_4 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_fill_2 FILLER_33_433 ();
 sg13g2_fill_2 FILLER_33_461 ();
 sg13g2_decap_4 FILLER_33_467 ();
 sg13g2_fill_1 FILLER_33_471 ();
 sg13g2_fill_2 FILLER_33_496 ();
 sg13g2_fill_1 FILLER_33_542 ();
 sg13g2_fill_2 FILLER_33_573 ();
 sg13g2_decap_4 FILLER_33_588 ();
 sg13g2_decap_4 FILLER_33_631 ();
 sg13g2_fill_2 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_657 ();
 sg13g2_decap_8 FILLER_33_696 ();
 sg13g2_fill_1 FILLER_33_703 ();
 sg13g2_fill_2 FILLER_33_747 ();
 sg13g2_fill_2 FILLER_33_793 ();
 sg13g2_fill_1 FILLER_33_795 ();
 sg13g2_decap_4 FILLER_33_830 ();
 sg13g2_fill_1 FILLER_33_838 ();
 sg13g2_fill_2 FILLER_33_848 ();
 sg13g2_fill_2 FILLER_33_887 ();
 sg13g2_fill_1 FILLER_33_889 ();
 sg13g2_fill_1 FILLER_33_916 ();
 sg13g2_fill_1 FILLER_33_922 ();
 sg13g2_fill_1 FILLER_33_957 ();
 sg13g2_fill_1 FILLER_33_963 ();
 sg13g2_fill_1 FILLER_33_970 ();
 sg13g2_fill_1 FILLER_33_976 ();
 sg13g2_fill_1 FILLER_33_981 ();
 sg13g2_fill_1 FILLER_33_1000 ();
 sg13g2_fill_1 FILLER_33_1006 ();
 sg13g2_fill_1 FILLER_33_1012 ();
 sg13g2_fill_2 FILLER_33_1030 ();
 sg13g2_fill_1 FILLER_33_1032 ();
 sg13g2_fill_2 FILLER_33_1049 ();
 sg13g2_decap_8 FILLER_33_1097 ();
 sg13g2_decap_8 FILLER_33_1104 ();
 sg13g2_decap_8 FILLER_33_1111 ();
 sg13g2_decap_8 FILLER_33_1118 ();
 sg13g2_decap_8 FILLER_33_1125 ();
 sg13g2_decap_8 FILLER_33_1132 ();
 sg13g2_decap_8 FILLER_33_1139 ();
 sg13g2_decap_8 FILLER_33_1146 ();
 sg13g2_decap_8 FILLER_33_1153 ();
 sg13g2_decap_8 FILLER_33_1160 ();
 sg13g2_decap_8 FILLER_33_1167 ();
 sg13g2_decap_8 FILLER_33_1174 ();
 sg13g2_decap_8 FILLER_33_1181 ();
 sg13g2_decap_8 FILLER_33_1188 ();
 sg13g2_decap_8 FILLER_33_1195 ();
 sg13g2_decap_8 FILLER_33_1202 ();
 sg13g2_decap_8 FILLER_33_1209 ();
 sg13g2_decap_8 FILLER_33_1216 ();
 sg13g2_decap_8 FILLER_33_1223 ();
 sg13g2_decap_8 FILLER_33_1230 ();
 sg13g2_decap_8 FILLER_33_1237 ();
 sg13g2_decap_8 FILLER_33_1244 ();
 sg13g2_decap_8 FILLER_33_1251 ();
 sg13g2_decap_8 FILLER_33_1258 ();
 sg13g2_decap_8 FILLER_33_1265 ();
 sg13g2_decap_8 FILLER_33_1272 ();
 sg13g2_decap_8 FILLER_33_1279 ();
 sg13g2_decap_8 FILLER_33_1286 ();
 sg13g2_decap_8 FILLER_33_1293 ();
 sg13g2_decap_8 FILLER_33_1300 ();
 sg13g2_decap_8 FILLER_33_1307 ();
 sg13g2_decap_8 FILLER_33_1314 ();
 sg13g2_decap_4 FILLER_33_1321 ();
 sg13g2_fill_1 FILLER_33_1325 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_66 ();
 sg13g2_decap_4 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_fill_2 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_164 ();
 sg13g2_fill_1 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_273 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_decap_4 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_307 ();
 sg13g2_fill_2 FILLER_34_369 ();
 sg13g2_fill_1 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_405 ();
 sg13g2_fill_2 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_fill_1 FILLER_34_457 ();
 sg13g2_fill_2 FILLER_34_496 ();
 sg13g2_fill_2 FILLER_34_521 ();
 sg13g2_decap_8 FILLER_34_536 ();
 sg13g2_decap_4 FILLER_34_543 ();
 sg13g2_fill_1 FILLER_34_547 ();
 sg13g2_fill_1 FILLER_34_574 ();
 sg13g2_fill_2 FILLER_34_601 ();
 sg13g2_fill_2 FILLER_34_624 ();
 sg13g2_fill_1 FILLER_34_631 ();
 sg13g2_fill_2 FILLER_34_636 ();
 sg13g2_fill_1 FILLER_34_650 ();
 sg13g2_fill_2 FILLER_34_670 ();
 sg13g2_decap_4 FILLER_34_711 ();
 sg13g2_fill_1 FILLER_34_719 ();
 sg13g2_fill_1 FILLER_34_728 ();
 sg13g2_decap_4 FILLER_34_733 ();
 sg13g2_fill_1 FILLER_34_737 ();
 sg13g2_fill_1 FILLER_34_742 ();
 sg13g2_fill_2 FILLER_34_762 ();
 sg13g2_fill_1 FILLER_34_790 ();
 sg13g2_fill_2 FILLER_34_796 ();
 sg13g2_fill_1 FILLER_34_802 ();
 sg13g2_fill_2 FILLER_34_807 ();
 sg13g2_fill_1 FILLER_34_835 ();
 sg13g2_fill_1 FILLER_34_840 ();
 sg13g2_fill_2 FILLER_34_872 ();
 sg13g2_fill_1 FILLER_34_905 ();
 sg13g2_fill_2 FILLER_34_945 ();
 sg13g2_fill_1 FILLER_34_1085 ();
 sg13g2_decap_8 FILLER_34_1095 ();
 sg13g2_decap_8 FILLER_34_1102 ();
 sg13g2_decap_8 FILLER_34_1109 ();
 sg13g2_decap_8 FILLER_34_1116 ();
 sg13g2_decap_8 FILLER_34_1123 ();
 sg13g2_decap_8 FILLER_34_1130 ();
 sg13g2_decap_8 FILLER_34_1137 ();
 sg13g2_decap_8 FILLER_34_1144 ();
 sg13g2_decap_8 FILLER_34_1151 ();
 sg13g2_decap_8 FILLER_34_1158 ();
 sg13g2_decap_8 FILLER_34_1165 ();
 sg13g2_decap_8 FILLER_34_1172 ();
 sg13g2_decap_8 FILLER_34_1179 ();
 sg13g2_decap_8 FILLER_34_1186 ();
 sg13g2_decap_8 FILLER_34_1193 ();
 sg13g2_decap_8 FILLER_34_1200 ();
 sg13g2_decap_8 FILLER_34_1207 ();
 sg13g2_decap_8 FILLER_34_1214 ();
 sg13g2_decap_8 FILLER_34_1221 ();
 sg13g2_decap_8 FILLER_34_1228 ();
 sg13g2_decap_8 FILLER_34_1235 ();
 sg13g2_decap_8 FILLER_34_1242 ();
 sg13g2_decap_8 FILLER_34_1249 ();
 sg13g2_decap_8 FILLER_34_1256 ();
 sg13g2_decap_8 FILLER_34_1263 ();
 sg13g2_decap_8 FILLER_34_1270 ();
 sg13g2_decap_8 FILLER_34_1277 ();
 sg13g2_decap_8 FILLER_34_1284 ();
 sg13g2_decap_8 FILLER_34_1291 ();
 sg13g2_decap_8 FILLER_34_1298 ();
 sg13g2_decap_8 FILLER_34_1305 ();
 sg13g2_decap_8 FILLER_34_1312 ();
 sg13g2_decap_8 FILLER_34_1319 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_4 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_2 FILLER_35_190 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_202 ();
 sg13g2_fill_1 FILLER_35_211 ();
 sg13g2_decap_4 FILLER_35_216 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_283 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_decap_4 FILLER_35_342 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_357 ();
 sg13g2_fill_1 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_403 ();
 sg13g2_fill_1 FILLER_35_439 ();
 sg13g2_fill_2 FILLER_35_465 ();
 sg13g2_fill_1 FILLER_35_472 ();
 sg13g2_fill_1 FILLER_35_477 ();
 sg13g2_fill_1 FILLER_35_483 ();
 sg13g2_fill_1 FILLER_35_489 ();
 sg13g2_fill_1 FILLER_35_495 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_fill_1 FILLER_35_509 ();
 sg13g2_fill_2 FILLER_35_515 ();
 sg13g2_fill_1 FILLER_35_530 ();
 sg13g2_fill_2 FILLER_35_539 ();
 sg13g2_fill_2 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_552 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_fill_1 FILLER_35_559 ();
 sg13g2_fill_2 FILLER_35_564 ();
 sg13g2_fill_2 FILLER_35_570 ();
 sg13g2_fill_2 FILLER_35_576 ();
 sg13g2_fill_1 FILLER_35_586 ();
 sg13g2_fill_1 FILLER_35_592 ();
 sg13g2_fill_2 FILLER_35_609 ();
 sg13g2_fill_1 FILLER_35_611 ();
 sg13g2_fill_1 FILLER_35_655 ();
 sg13g2_decap_4 FILLER_35_687 ();
 sg13g2_fill_1 FILLER_35_763 ();
 sg13g2_fill_2 FILLER_35_788 ();
 sg13g2_fill_2 FILLER_35_814 ();
 sg13g2_fill_1 FILLER_35_816 ();
 sg13g2_decap_4 FILLER_35_822 ();
 sg13g2_fill_2 FILLER_35_859 ();
 sg13g2_fill_1 FILLER_35_886 ();
 sg13g2_decap_4 FILLER_35_911 ();
 sg13g2_fill_2 FILLER_35_915 ();
 sg13g2_decap_8 FILLER_35_921 ();
 sg13g2_fill_1 FILLER_35_928 ();
 sg13g2_fill_1 FILLER_35_942 ();
 sg13g2_fill_1 FILLER_35_958 ();
 sg13g2_fill_2 FILLER_35_964 ();
 sg13g2_fill_2 FILLER_35_971 ();
 sg13g2_fill_1 FILLER_35_973 ();
 sg13g2_fill_1 FILLER_35_978 ();
 sg13g2_fill_2 FILLER_35_984 ();
 sg13g2_fill_1 FILLER_35_986 ();
 sg13g2_fill_1 FILLER_35_991 ();
 sg13g2_fill_1 FILLER_35_997 ();
 sg13g2_fill_1 FILLER_35_1002 ();
 sg13g2_fill_2 FILLER_35_1007 ();
 sg13g2_fill_2 FILLER_35_1045 ();
 sg13g2_fill_1 FILLER_35_1055 ();
 sg13g2_fill_1 FILLER_35_1065 ();
 sg13g2_fill_1 FILLER_35_1070 ();
 sg13g2_decap_8 FILLER_35_1080 ();
 sg13g2_decap_8 FILLER_35_1087 ();
 sg13g2_decap_8 FILLER_35_1094 ();
 sg13g2_decap_8 FILLER_35_1101 ();
 sg13g2_decap_8 FILLER_35_1108 ();
 sg13g2_decap_8 FILLER_35_1115 ();
 sg13g2_decap_8 FILLER_35_1122 ();
 sg13g2_decap_8 FILLER_35_1129 ();
 sg13g2_decap_8 FILLER_35_1136 ();
 sg13g2_decap_8 FILLER_35_1143 ();
 sg13g2_decap_8 FILLER_35_1150 ();
 sg13g2_decap_8 FILLER_35_1157 ();
 sg13g2_decap_8 FILLER_35_1164 ();
 sg13g2_decap_8 FILLER_35_1171 ();
 sg13g2_decap_8 FILLER_35_1178 ();
 sg13g2_decap_8 FILLER_35_1185 ();
 sg13g2_decap_8 FILLER_35_1192 ();
 sg13g2_decap_8 FILLER_35_1199 ();
 sg13g2_decap_8 FILLER_35_1206 ();
 sg13g2_decap_8 FILLER_35_1213 ();
 sg13g2_decap_8 FILLER_35_1220 ();
 sg13g2_decap_8 FILLER_35_1227 ();
 sg13g2_decap_8 FILLER_35_1234 ();
 sg13g2_decap_8 FILLER_35_1241 ();
 sg13g2_decap_8 FILLER_35_1248 ();
 sg13g2_decap_8 FILLER_35_1255 ();
 sg13g2_decap_8 FILLER_35_1262 ();
 sg13g2_decap_8 FILLER_35_1269 ();
 sg13g2_decap_8 FILLER_35_1276 ();
 sg13g2_decap_8 FILLER_35_1283 ();
 sg13g2_decap_8 FILLER_35_1290 ();
 sg13g2_decap_8 FILLER_35_1297 ();
 sg13g2_decap_8 FILLER_35_1304 ();
 sg13g2_decap_8 FILLER_35_1311 ();
 sg13g2_decap_8 FILLER_35_1318 ();
 sg13g2_fill_1 FILLER_35_1325 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_fill_2 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_decap_4 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_257 ();
 sg13g2_fill_2 FILLER_36_264 ();
 sg13g2_fill_1 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_295 ();
 sg13g2_fill_2 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_358 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_fill_2 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_fill_2 FILLER_36_418 ();
 sg13g2_fill_1 FILLER_36_420 ();
 sg13g2_fill_2 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_427 ();
 sg13g2_decap_4 FILLER_36_471 ();
 sg13g2_fill_2 FILLER_36_479 ();
 sg13g2_decap_4 FILLER_36_503 ();
 sg13g2_fill_2 FILLER_36_520 ();
 sg13g2_fill_1 FILLER_36_522 ();
 sg13g2_fill_1 FILLER_36_544 ();
 sg13g2_fill_1 FILLER_36_575 ();
 sg13g2_fill_2 FILLER_36_581 ();
 sg13g2_fill_2 FILLER_36_609 ();
 sg13g2_fill_2 FILLER_36_614 ();
 sg13g2_fill_2 FILLER_36_624 ();
 sg13g2_fill_1 FILLER_36_626 ();
 sg13g2_fill_2 FILLER_36_632 ();
 sg13g2_fill_1 FILLER_36_634 ();
 sg13g2_fill_2 FILLER_36_660 ();
 sg13g2_fill_1 FILLER_36_662 ();
 sg13g2_fill_1 FILLER_36_705 ();
 sg13g2_fill_1 FILLER_36_729 ();
 sg13g2_fill_1 FILLER_36_747 ();
 sg13g2_fill_1 FILLER_36_753 ();
 sg13g2_fill_1 FILLER_36_764 ();
 sg13g2_fill_1 FILLER_36_796 ();
 sg13g2_fill_2 FILLER_36_853 ();
 sg13g2_fill_1 FILLER_36_855 ();
 sg13g2_fill_2 FILLER_36_907 ();
 sg13g2_fill_2 FILLER_36_948 ();
 sg13g2_fill_1 FILLER_36_950 ();
 sg13g2_fill_2 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1095 ();
 sg13g2_decap_4 FILLER_36_1102 ();
 sg13g2_fill_1 FILLER_36_1106 ();
 sg13g2_decap_8 FILLER_36_1112 ();
 sg13g2_decap_8 FILLER_36_1119 ();
 sg13g2_decap_8 FILLER_36_1126 ();
 sg13g2_decap_8 FILLER_36_1133 ();
 sg13g2_decap_8 FILLER_36_1140 ();
 sg13g2_decap_8 FILLER_36_1147 ();
 sg13g2_decap_8 FILLER_36_1154 ();
 sg13g2_decap_8 FILLER_36_1161 ();
 sg13g2_decap_8 FILLER_36_1168 ();
 sg13g2_decap_8 FILLER_36_1175 ();
 sg13g2_decap_8 FILLER_36_1182 ();
 sg13g2_decap_8 FILLER_36_1189 ();
 sg13g2_decap_8 FILLER_36_1196 ();
 sg13g2_decap_8 FILLER_36_1203 ();
 sg13g2_decap_8 FILLER_36_1210 ();
 sg13g2_decap_8 FILLER_36_1217 ();
 sg13g2_decap_8 FILLER_36_1224 ();
 sg13g2_decap_8 FILLER_36_1231 ();
 sg13g2_decap_8 FILLER_36_1238 ();
 sg13g2_decap_8 FILLER_36_1245 ();
 sg13g2_decap_8 FILLER_36_1252 ();
 sg13g2_decap_8 FILLER_36_1259 ();
 sg13g2_decap_8 FILLER_36_1266 ();
 sg13g2_decap_8 FILLER_36_1273 ();
 sg13g2_decap_8 FILLER_36_1280 ();
 sg13g2_decap_8 FILLER_36_1287 ();
 sg13g2_decap_8 FILLER_36_1294 ();
 sg13g2_decap_8 FILLER_36_1301 ();
 sg13g2_decap_8 FILLER_36_1308 ();
 sg13g2_decap_8 FILLER_36_1315 ();
 sg13g2_decap_4 FILLER_36_1322 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_4 FILLER_37_63 ();
 sg13g2_fill_1 FILLER_37_67 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_194 ();
 sg13g2_fill_1 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_282 ();
 sg13g2_fill_2 FILLER_37_295 ();
 sg13g2_fill_2 FILLER_37_319 ();
 sg13g2_fill_1 FILLER_37_321 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_fill_1 FILLER_37_415 ();
 sg13g2_fill_1 FILLER_37_420 ();
 sg13g2_fill_2 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_37_431 ();
 sg13g2_fill_2 FILLER_37_488 ();
 sg13g2_fill_1 FILLER_37_502 ();
 sg13g2_fill_2 FILLER_37_511 ();
 sg13g2_fill_1 FILLER_37_518 ();
 sg13g2_fill_2 FILLER_37_523 ();
 sg13g2_fill_1 FILLER_37_529 ();
 sg13g2_fill_2 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_585 ();
 sg13g2_fill_2 FILLER_37_590 ();
 sg13g2_decap_4 FILLER_37_596 ();
 sg13g2_fill_1 FILLER_37_600 ();
 sg13g2_fill_2 FILLER_37_605 ();
 sg13g2_fill_1 FILLER_37_612 ();
 sg13g2_fill_2 FILLER_37_633 ();
 sg13g2_fill_1 FILLER_37_635 ();
 sg13g2_fill_2 FILLER_37_640 ();
 sg13g2_fill_2 FILLER_37_694 ();
 sg13g2_fill_1 FILLER_37_696 ();
 sg13g2_decap_8 FILLER_37_780 ();
 sg13g2_fill_1 FILLER_37_787 ();
 sg13g2_fill_2 FILLER_37_801 ();
 sg13g2_fill_1 FILLER_37_803 ();
 sg13g2_decap_4 FILLER_37_808 ();
 sg13g2_fill_1 FILLER_37_812 ();
 sg13g2_decap_4 FILLER_37_825 ();
 sg13g2_fill_2 FILLER_37_833 ();
 sg13g2_fill_2 FILLER_37_853 ();
 sg13g2_fill_2 FILLER_37_879 ();
 sg13g2_fill_1 FILLER_37_881 ();
 sg13g2_decap_8 FILLER_37_894 ();
 sg13g2_fill_2 FILLER_37_901 ();
 sg13g2_fill_1 FILLER_37_903 ();
 sg13g2_decap_4 FILLER_37_916 ();
 sg13g2_decap_4 FILLER_37_924 ();
 sg13g2_fill_1 FILLER_37_933 ();
 sg13g2_fill_2 FILLER_37_968 ();
 sg13g2_decap_4 FILLER_37_1008 ();
 sg13g2_fill_2 FILLER_37_1020 ();
 sg13g2_fill_1 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1036 ();
 sg13g2_fill_2 FILLER_37_1058 ();
 sg13g2_fill_2 FILLER_37_1064 ();
 sg13g2_fill_1 FILLER_37_1066 ();
 sg13g2_fill_2 FILLER_37_1071 ();
 sg13g2_fill_1 FILLER_37_1073 ();
 sg13g2_fill_1 FILLER_37_1079 ();
 sg13g2_decap_8 FILLER_37_1084 ();
 sg13g2_fill_2 FILLER_37_1091 ();
 sg13g2_fill_1 FILLER_37_1093 ();
 sg13g2_decap_4 FILLER_37_1105 ();
 sg13g2_decap_8 FILLER_37_1113 ();
 sg13g2_decap_8 FILLER_37_1120 ();
 sg13g2_decap_8 FILLER_37_1127 ();
 sg13g2_decap_8 FILLER_37_1134 ();
 sg13g2_decap_8 FILLER_37_1141 ();
 sg13g2_decap_8 FILLER_37_1148 ();
 sg13g2_decap_8 FILLER_37_1155 ();
 sg13g2_decap_8 FILLER_37_1162 ();
 sg13g2_decap_8 FILLER_37_1169 ();
 sg13g2_decap_8 FILLER_37_1176 ();
 sg13g2_decap_8 FILLER_37_1183 ();
 sg13g2_decap_8 FILLER_37_1190 ();
 sg13g2_decap_8 FILLER_37_1197 ();
 sg13g2_decap_8 FILLER_37_1204 ();
 sg13g2_decap_8 FILLER_37_1211 ();
 sg13g2_decap_8 FILLER_37_1218 ();
 sg13g2_decap_8 FILLER_37_1225 ();
 sg13g2_decap_8 FILLER_37_1232 ();
 sg13g2_decap_8 FILLER_37_1239 ();
 sg13g2_decap_8 FILLER_37_1246 ();
 sg13g2_decap_8 FILLER_37_1253 ();
 sg13g2_decap_8 FILLER_37_1260 ();
 sg13g2_decap_8 FILLER_37_1267 ();
 sg13g2_decap_8 FILLER_37_1274 ();
 sg13g2_decap_8 FILLER_37_1281 ();
 sg13g2_decap_8 FILLER_37_1288 ();
 sg13g2_decap_8 FILLER_37_1295 ();
 sg13g2_decap_8 FILLER_37_1302 ();
 sg13g2_decap_8 FILLER_37_1309 ();
 sg13g2_decap_8 FILLER_37_1316 ();
 sg13g2_fill_2 FILLER_37_1323 ();
 sg13g2_fill_1 FILLER_37_1325 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_1 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_168 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_2 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_fill_2 FILLER_38_300 ();
 sg13g2_decap_4 FILLER_38_307 ();
 sg13g2_decap_4 FILLER_38_315 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_2 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_2 FILLER_38_404 ();
 sg13g2_decap_8 FILLER_38_466 ();
 sg13g2_fill_1 FILLER_38_477 ();
 sg13g2_fill_1 FILLER_38_483 ();
 sg13g2_fill_2 FILLER_38_498 ();
 sg13g2_fill_2 FILLER_38_539 ();
 sg13g2_fill_1 FILLER_38_541 ();
 sg13g2_fill_2 FILLER_38_559 ();
 sg13g2_fill_2 FILLER_38_565 ();
 sg13g2_fill_1 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_572 ();
 sg13g2_fill_1 FILLER_38_574 ();
 sg13g2_fill_1 FILLER_38_579 ();
 sg13g2_fill_1 FILLER_38_606 ();
 sg13g2_fill_1 FILLER_38_628 ();
 sg13g2_fill_1 FILLER_38_633 ();
 sg13g2_fill_2 FILLER_38_643 ();
 sg13g2_fill_1 FILLER_38_654 ();
 sg13g2_fill_1 FILLER_38_664 ();
 sg13g2_fill_1 FILLER_38_674 ();
 sg13g2_fill_1 FILLER_38_706 ();
 sg13g2_fill_2 FILLER_38_715 ();
 sg13g2_fill_1 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_729 ();
 sg13g2_fill_1 FILLER_38_784 ();
 sg13g2_fill_1 FILLER_38_807 ();
 sg13g2_fill_2 FILLER_38_813 ();
 sg13g2_fill_1 FILLER_38_823 ();
 sg13g2_fill_2 FILLER_38_828 ();
 sg13g2_fill_1 FILLER_38_856 ();
 sg13g2_fill_1 FILLER_38_860 ();
 sg13g2_fill_1 FILLER_38_871 ();
 sg13g2_fill_2 FILLER_38_891 ();
 sg13g2_fill_1 FILLER_38_893 ();
 sg13g2_fill_1 FILLER_38_904 ();
 sg13g2_decap_8 FILLER_38_913 ();
 sg13g2_decap_4 FILLER_38_920 ();
 sg13g2_decap_8 FILLER_38_927 ();
 sg13g2_fill_1 FILLER_38_942 ();
 sg13g2_fill_1 FILLER_38_947 ();
 sg13g2_fill_1 FILLER_38_978 ();
 sg13g2_fill_1 FILLER_38_983 ();
 sg13g2_fill_1 FILLER_38_988 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_fill_2 FILLER_38_1013 ();
 sg13g2_fill_2 FILLER_38_1031 ();
 sg13g2_fill_2 FILLER_38_1041 ();
 sg13g2_fill_2 FILLER_38_1069 ();
 sg13g2_decap_8 FILLER_38_1097 ();
 sg13g2_decap_8 FILLER_38_1104 ();
 sg13g2_decap_8 FILLER_38_1111 ();
 sg13g2_decap_8 FILLER_38_1118 ();
 sg13g2_decap_8 FILLER_38_1125 ();
 sg13g2_decap_8 FILLER_38_1132 ();
 sg13g2_decap_8 FILLER_38_1139 ();
 sg13g2_decap_8 FILLER_38_1146 ();
 sg13g2_decap_8 FILLER_38_1153 ();
 sg13g2_decap_8 FILLER_38_1160 ();
 sg13g2_decap_8 FILLER_38_1167 ();
 sg13g2_decap_8 FILLER_38_1174 ();
 sg13g2_decap_8 FILLER_38_1181 ();
 sg13g2_decap_8 FILLER_38_1188 ();
 sg13g2_decap_8 FILLER_38_1195 ();
 sg13g2_decap_8 FILLER_38_1202 ();
 sg13g2_decap_8 FILLER_38_1209 ();
 sg13g2_decap_8 FILLER_38_1216 ();
 sg13g2_decap_8 FILLER_38_1223 ();
 sg13g2_decap_8 FILLER_38_1230 ();
 sg13g2_decap_8 FILLER_38_1237 ();
 sg13g2_decap_8 FILLER_38_1244 ();
 sg13g2_decap_8 FILLER_38_1251 ();
 sg13g2_decap_8 FILLER_38_1258 ();
 sg13g2_decap_8 FILLER_38_1265 ();
 sg13g2_decap_8 FILLER_38_1272 ();
 sg13g2_decap_8 FILLER_38_1279 ();
 sg13g2_decap_8 FILLER_38_1286 ();
 sg13g2_decap_8 FILLER_38_1293 ();
 sg13g2_decap_8 FILLER_38_1300 ();
 sg13g2_decap_8 FILLER_38_1307 ();
 sg13g2_decap_8 FILLER_38_1314 ();
 sg13g2_decap_4 FILLER_38_1321 ();
 sg13g2_fill_1 FILLER_38_1325 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_42 ();
 sg13g2_fill_2 FILLER_39_51 ();
 sg13g2_fill_1 FILLER_39_57 ();
 sg13g2_fill_1 FILLER_39_141 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_4 FILLER_39_175 ();
 sg13g2_fill_1 FILLER_39_179 ();
 sg13g2_fill_2 FILLER_39_230 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_fill_1 FILLER_39_299 ();
 sg13g2_fill_2 FILLER_39_304 ();
 sg13g2_fill_1 FILLER_39_306 ();
 sg13g2_fill_1 FILLER_39_318 ();
 sg13g2_decap_4 FILLER_39_371 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_fill_2 FILLER_39_381 ();
 sg13g2_fill_1 FILLER_39_413 ();
 sg13g2_decap_4 FILLER_39_426 ();
 sg13g2_fill_1 FILLER_39_451 ();
 sg13g2_fill_2 FILLER_39_508 ();
 sg13g2_fill_1 FILLER_39_510 ();
 sg13g2_fill_2 FILLER_39_515 ();
 sg13g2_fill_1 FILLER_39_517 ();
 sg13g2_decap_4 FILLER_39_522 ();
 sg13g2_fill_1 FILLER_39_541 ();
 sg13g2_fill_2 FILLER_39_545 ();
 sg13g2_fill_1 FILLER_39_547 ();
 sg13g2_fill_1 FILLER_39_578 ();
 sg13g2_fill_2 FILLER_39_583 ();
 sg13g2_fill_1 FILLER_39_585 ();
 sg13g2_fill_1 FILLER_39_590 ();
 sg13g2_fill_1 FILLER_39_604 ();
 sg13g2_fill_2 FILLER_39_678 ();
 sg13g2_fill_1 FILLER_39_689 ();
 sg13g2_fill_1 FILLER_39_720 ();
 sg13g2_fill_1 FILLER_39_735 ();
 sg13g2_fill_2 FILLER_39_762 ();
 sg13g2_fill_1 FILLER_39_764 ();
 sg13g2_fill_2 FILLER_39_769 ();
 sg13g2_decap_8 FILLER_39_775 ();
 sg13g2_decap_4 FILLER_39_799 ();
 sg13g2_fill_2 FILLER_39_803 ();
 sg13g2_fill_1 FILLER_39_835 ();
 sg13g2_fill_1 FILLER_39_907 ();
 sg13g2_fill_1 FILLER_39_918 ();
 sg13g2_fill_2 FILLER_39_927 ();
 sg13g2_fill_2 FILLER_39_953 ();
 sg13g2_decap_8 FILLER_39_963 ();
 sg13g2_fill_2 FILLER_39_970 ();
 sg13g2_fill_1 FILLER_39_972 ();
 sg13g2_fill_2 FILLER_39_978 ();
 sg13g2_fill_1 FILLER_39_1006 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_fill_1 FILLER_39_1075 ();
 sg13g2_fill_2 FILLER_39_1080 ();
 sg13g2_fill_1 FILLER_39_1086 ();
 sg13g2_decap_8 FILLER_39_1095 ();
 sg13g2_decap_8 FILLER_39_1102 ();
 sg13g2_decap_8 FILLER_39_1109 ();
 sg13g2_decap_8 FILLER_39_1116 ();
 sg13g2_decap_8 FILLER_39_1123 ();
 sg13g2_decap_4 FILLER_39_1130 ();
 sg13g2_fill_2 FILLER_39_1134 ();
 sg13g2_fill_2 FILLER_39_1141 ();
 sg13g2_decap_8 FILLER_39_1147 ();
 sg13g2_fill_2 FILLER_39_1154 ();
 sg13g2_decap_8 FILLER_39_1186 ();
 sg13g2_decap_8 FILLER_39_1193 ();
 sg13g2_decap_8 FILLER_39_1200 ();
 sg13g2_decap_8 FILLER_39_1207 ();
 sg13g2_decap_8 FILLER_39_1214 ();
 sg13g2_decap_8 FILLER_39_1221 ();
 sg13g2_decap_8 FILLER_39_1228 ();
 sg13g2_decap_8 FILLER_39_1235 ();
 sg13g2_decap_8 FILLER_39_1242 ();
 sg13g2_decap_8 FILLER_39_1249 ();
 sg13g2_decap_8 FILLER_39_1256 ();
 sg13g2_decap_8 FILLER_39_1263 ();
 sg13g2_decap_8 FILLER_39_1270 ();
 sg13g2_decap_8 FILLER_39_1277 ();
 sg13g2_decap_8 FILLER_39_1284 ();
 sg13g2_decap_8 FILLER_39_1291 ();
 sg13g2_decap_8 FILLER_39_1298 ();
 sg13g2_decap_8 FILLER_39_1305 ();
 sg13g2_decap_8 FILLER_39_1312 ();
 sg13g2_decap_8 FILLER_39_1319 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_fill_2 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_129 ();
 sg13g2_fill_1 FILLER_40_146 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_fill_1 FILLER_40_215 ();
 sg13g2_decap_4 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_255 ();
 sg13g2_fill_2 FILLER_40_264 ();
 sg13g2_decap_4 FILLER_40_296 ();
 sg13g2_fill_2 FILLER_40_331 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_348 ();
 sg13g2_fill_2 FILLER_40_354 ();
 sg13g2_fill_1 FILLER_40_386 ();
 sg13g2_fill_2 FILLER_40_405 ();
 sg13g2_fill_1 FILLER_40_457 ();
 sg13g2_fill_2 FILLER_40_466 ();
 sg13g2_decap_4 FILLER_40_472 ();
 sg13g2_fill_2 FILLER_40_476 ();
 sg13g2_fill_1 FILLER_40_482 ();
 sg13g2_fill_1 FILLER_40_487 ();
 sg13g2_fill_2 FILLER_40_491 ();
 sg13g2_fill_1 FILLER_40_497 ();
 sg13g2_fill_1 FILLER_40_528 ();
 sg13g2_fill_1 FILLER_40_542 ();
 sg13g2_fill_1 FILLER_40_577 ();
 sg13g2_fill_1 FILLER_40_668 ();
 sg13g2_fill_2 FILLER_40_673 ();
 sg13g2_decap_4 FILLER_40_679 ();
 sg13g2_fill_1 FILLER_40_683 ();
 sg13g2_fill_2 FILLER_40_692 ();
 sg13g2_fill_2 FILLER_40_700 ();
 sg13g2_fill_1 FILLER_40_715 ();
 sg13g2_fill_2 FILLER_40_754 ();
 sg13g2_fill_2 FILLER_40_803 ();
 sg13g2_fill_1 FILLER_40_812 ();
 sg13g2_fill_2 FILLER_40_821 ();
 sg13g2_fill_2 FILLER_40_827 ();
 sg13g2_fill_2 FILLER_40_833 ();
 sg13g2_decap_4 FILLER_40_847 ();
 sg13g2_fill_1 FILLER_40_851 ();
 sg13g2_fill_1 FILLER_40_856 ();
 sg13g2_fill_2 FILLER_40_895 ();
 sg13g2_fill_1 FILLER_40_909 ();
 sg13g2_fill_2 FILLER_40_923 ();
 sg13g2_fill_1 FILLER_40_933 ();
 sg13g2_fill_2 FILLER_40_946 ();
 sg13g2_decap_4 FILLER_40_979 ();
 sg13g2_fill_2 FILLER_40_995 ();
 sg13g2_fill_1 FILLER_40_1001 ();
 sg13g2_fill_2 FILLER_40_1007 ();
 sg13g2_fill_1 FILLER_40_1009 ();
 sg13g2_decap_4 FILLER_40_1014 ();
 sg13g2_decap_4 FILLER_40_1043 ();
 sg13g2_fill_2 FILLER_40_1047 ();
 sg13g2_decap_4 FILLER_40_1061 ();
 sg13g2_fill_2 FILLER_40_1065 ();
 sg13g2_fill_2 FILLER_40_1111 ();
 sg13g2_fill_2 FILLER_40_1117 ();
 sg13g2_decap_4 FILLER_40_1123 ();
 sg13g2_fill_1 FILLER_40_1161 ();
 sg13g2_fill_1 FILLER_40_1166 ();
 sg13g2_fill_1 FILLER_40_1171 ();
 sg13g2_decap_8 FILLER_40_1207 ();
 sg13g2_decap_8 FILLER_40_1214 ();
 sg13g2_decap_8 FILLER_40_1221 ();
 sg13g2_decap_8 FILLER_40_1228 ();
 sg13g2_decap_8 FILLER_40_1235 ();
 sg13g2_decap_8 FILLER_40_1242 ();
 sg13g2_decap_8 FILLER_40_1249 ();
 sg13g2_decap_8 FILLER_40_1256 ();
 sg13g2_decap_8 FILLER_40_1263 ();
 sg13g2_decap_8 FILLER_40_1270 ();
 sg13g2_decap_8 FILLER_40_1277 ();
 sg13g2_decap_8 FILLER_40_1284 ();
 sg13g2_decap_8 FILLER_40_1291 ();
 sg13g2_decap_8 FILLER_40_1298 ();
 sg13g2_decap_8 FILLER_40_1305 ();
 sg13g2_decap_8 FILLER_40_1312 ();
 sg13g2_decap_8 FILLER_40_1319 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_23 ();
 sg13g2_fill_1 FILLER_41_90 ();
 sg13g2_fill_2 FILLER_41_125 ();
 sg13g2_decap_8 FILLER_41_188 ();
 sg13g2_decap_4 FILLER_41_195 ();
 sg13g2_decap_8 FILLER_41_215 ();
 sg13g2_decap_4 FILLER_41_226 ();
 sg13g2_fill_1 FILLER_41_230 ();
 sg13g2_fill_2 FILLER_41_235 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_262 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_1 FILLER_41_276 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_fill_1 FILLER_41_285 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_fill_2 FILLER_41_312 ();
 sg13g2_fill_2 FILLER_41_365 ();
 sg13g2_fill_1 FILLER_41_371 ();
 sg13g2_fill_2 FILLER_41_401 ();
 sg13g2_decap_8 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_41_457 ();
 sg13g2_fill_2 FILLER_41_494 ();
 sg13g2_fill_1 FILLER_41_505 ();
 sg13g2_fill_2 FILLER_41_510 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_fill_1 FILLER_41_522 ();
 sg13g2_fill_1 FILLER_41_535 ();
 sg13g2_decap_4 FILLER_41_562 ();
 sg13g2_fill_1 FILLER_41_588 ();
 sg13g2_fill_2 FILLER_41_593 ();
 sg13g2_decap_4 FILLER_41_598 ();
 sg13g2_fill_1 FILLER_41_602 ();
 sg13g2_fill_2 FILLER_41_624 ();
 sg13g2_fill_1 FILLER_41_637 ();
 sg13g2_decap_4 FILLER_41_707 ();
 sg13g2_fill_1 FILLER_41_747 ();
 sg13g2_fill_2 FILLER_41_752 ();
 sg13g2_fill_1 FILLER_41_754 ();
 sg13g2_fill_2 FILLER_41_760 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_fill_2 FILLER_41_779 ();
 sg13g2_fill_1 FILLER_41_781 ();
 sg13g2_fill_2 FILLER_41_810 ();
 sg13g2_decap_4 FILLER_41_816 ();
 sg13g2_fill_2 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_856 ();
 sg13g2_fill_2 FILLER_41_865 ();
 sg13g2_fill_1 FILLER_41_867 ();
 sg13g2_fill_2 FILLER_41_880 ();
 sg13g2_fill_1 FILLER_41_892 ();
 sg13g2_fill_2 FILLER_41_942 ();
 sg13g2_fill_1 FILLER_41_944 ();
 sg13g2_fill_2 FILLER_41_980 ();
 sg13g2_fill_1 FILLER_41_1025 ();
 sg13g2_fill_1 FILLER_41_1034 ();
 sg13g2_fill_1 FILLER_41_1043 ();
 sg13g2_fill_2 FILLER_41_1070 ();
 sg13g2_fill_2 FILLER_41_1082 ();
 sg13g2_fill_2 FILLER_41_1110 ();
 sg13g2_fill_1 FILLER_41_1112 ();
 sg13g2_fill_1 FILLER_41_1143 ();
 sg13g2_decap_4 FILLER_41_1148 ();
 sg13g2_fill_1 FILLER_41_1171 ();
 sg13g2_fill_2 FILLER_41_1192 ();
 sg13g2_decap_8 FILLER_41_1202 ();
 sg13g2_decap_8 FILLER_41_1209 ();
 sg13g2_decap_8 FILLER_41_1216 ();
 sg13g2_decap_8 FILLER_41_1223 ();
 sg13g2_decap_8 FILLER_41_1230 ();
 sg13g2_decap_8 FILLER_41_1237 ();
 sg13g2_decap_8 FILLER_41_1244 ();
 sg13g2_decap_8 FILLER_41_1251 ();
 sg13g2_decap_8 FILLER_41_1258 ();
 sg13g2_decap_8 FILLER_41_1265 ();
 sg13g2_decap_8 FILLER_41_1272 ();
 sg13g2_decap_8 FILLER_41_1279 ();
 sg13g2_decap_8 FILLER_41_1286 ();
 sg13g2_decap_8 FILLER_41_1293 ();
 sg13g2_decap_8 FILLER_41_1300 ();
 sg13g2_decap_8 FILLER_41_1307 ();
 sg13g2_decap_8 FILLER_41_1314 ();
 sg13g2_decap_4 FILLER_41_1321 ();
 sg13g2_fill_1 FILLER_41_1325 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_4 FILLER_42_28 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_1 FILLER_42_64 ();
 sg13g2_decap_4 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_137 ();
 sg13g2_fill_1 FILLER_42_148 ();
 sg13g2_fill_2 FILLER_42_161 ();
 sg13g2_fill_1 FILLER_42_197 ();
 sg13g2_decap_8 FILLER_42_212 ();
 sg13g2_decap_8 FILLER_42_223 ();
 sg13g2_decap_4 FILLER_42_230 ();
 sg13g2_fill_2 FILLER_42_234 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_294 ();
 sg13g2_decap_4 FILLER_42_307 ();
 sg13g2_fill_1 FILLER_42_311 ();
 sg13g2_fill_2 FILLER_42_332 ();
 sg13g2_fill_1 FILLER_42_334 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_decap_8 FILLER_42_344 ();
 sg13g2_decap_4 FILLER_42_351 ();
 sg13g2_decap_4 FILLER_42_367 ();
 sg13g2_decap_4 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_4 FILLER_42_391 ();
 sg13g2_fill_1 FILLER_42_398 ();
 sg13g2_fill_2 FILLER_42_405 ();
 sg13g2_fill_1 FILLER_42_407 ();
 sg13g2_fill_1 FILLER_42_424 ();
 sg13g2_decap_8 FILLER_42_429 ();
 sg13g2_decap_4 FILLER_42_476 ();
 sg13g2_fill_2 FILLER_42_510 ();
 sg13g2_decap_4 FILLER_42_539 ();
 sg13g2_fill_1 FILLER_42_543 ();
 sg13g2_fill_1 FILLER_42_552 ();
 sg13g2_fill_2 FILLER_42_557 ();
 sg13g2_fill_2 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_597 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_fill_1 FILLER_42_610 ();
 sg13g2_fill_2 FILLER_42_615 ();
 sg13g2_fill_2 FILLER_42_652 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_fill_2 FILLER_42_669 ();
 sg13g2_fill_1 FILLER_42_676 ();
 sg13g2_fill_1 FILLER_42_681 ();
 sg13g2_fill_1 FILLER_42_685 ();
 sg13g2_fill_2 FILLER_42_690 ();
 sg13g2_fill_2 FILLER_42_702 ();
 sg13g2_fill_1 FILLER_42_704 ();
 sg13g2_fill_2 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_829 ();
 sg13g2_fill_2 FILLER_42_836 ();
 sg13g2_decap_4 FILLER_42_849 ();
 sg13g2_fill_1 FILLER_42_892 ();
 sg13g2_fill_1 FILLER_42_897 ();
 sg13g2_fill_1 FILLER_42_910 ();
 sg13g2_fill_2 FILLER_42_916 ();
 sg13g2_decap_4 FILLER_42_922 ();
 sg13g2_fill_2 FILLER_42_950 ();
 sg13g2_decap_4 FILLER_42_956 ();
 sg13g2_fill_2 FILLER_42_996 ();
 sg13g2_fill_2 FILLER_42_1006 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_fill_2 FILLER_42_1070 ();
 sg13g2_fill_1 FILLER_42_1108 ();
 sg13g2_decap_4 FILLER_42_1114 ();
 sg13g2_fill_2 FILLER_42_1118 ();
 sg13g2_fill_1 FILLER_42_1124 ();
 sg13g2_fill_1 FILLER_42_1130 ();
 sg13g2_fill_1 FILLER_42_1136 ();
 sg13g2_fill_1 FILLER_42_1141 ();
 sg13g2_fill_2 FILLER_42_1145 ();
 sg13g2_fill_2 FILLER_42_1150 ();
 sg13g2_decap_8 FILLER_42_1206 ();
 sg13g2_decap_8 FILLER_42_1213 ();
 sg13g2_decap_8 FILLER_42_1220 ();
 sg13g2_decap_8 FILLER_42_1227 ();
 sg13g2_decap_8 FILLER_42_1234 ();
 sg13g2_decap_8 FILLER_42_1241 ();
 sg13g2_decap_8 FILLER_42_1248 ();
 sg13g2_decap_8 FILLER_42_1255 ();
 sg13g2_decap_8 FILLER_42_1262 ();
 sg13g2_decap_8 FILLER_42_1269 ();
 sg13g2_decap_8 FILLER_42_1276 ();
 sg13g2_decap_8 FILLER_42_1283 ();
 sg13g2_decap_8 FILLER_42_1290 ();
 sg13g2_decap_8 FILLER_42_1297 ();
 sg13g2_decap_8 FILLER_42_1304 ();
 sg13g2_decap_8 FILLER_42_1311 ();
 sg13g2_decap_8 FILLER_42_1318 ();
 sg13g2_fill_1 FILLER_42_1325 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_4 FILLER_43_35 ();
 sg13g2_fill_2 FILLER_43_39 ();
 sg13g2_fill_2 FILLER_43_71 ();
 sg13g2_fill_1 FILLER_43_160 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_decap_4 FILLER_43_238 ();
 sg13g2_fill_2 FILLER_43_242 ();
 sg13g2_fill_1 FILLER_43_300 ();
 sg13g2_fill_2 FILLER_43_305 ();
 sg13g2_fill_2 FILLER_43_311 ();
 sg13g2_fill_1 FILLER_43_313 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_fill_2 FILLER_43_362 ();
 sg13g2_fill_2 FILLER_43_420 ();
 sg13g2_fill_1 FILLER_43_422 ();
 sg13g2_fill_2 FILLER_43_431 ();
 sg13g2_fill_2 FILLER_43_454 ();
 sg13g2_fill_1 FILLER_43_456 ();
 sg13g2_fill_2 FILLER_43_461 ();
 sg13g2_fill_2 FILLER_43_468 ();
 sg13g2_fill_2 FILLER_43_475 ();
 sg13g2_fill_1 FILLER_43_477 ();
 sg13g2_fill_1 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_493 ();
 sg13g2_fill_1 FILLER_43_524 ();
 sg13g2_fill_2 FILLER_43_533 ();
 sg13g2_fill_2 FILLER_43_543 ();
 sg13g2_decap_4 FILLER_43_579 ();
 sg13g2_fill_1 FILLER_43_583 ();
 sg13g2_fill_2 FILLER_43_624 ();
 sg13g2_fill_1 FILLER_43_635 ();
 sg13g2_decap_8 FILLER_43_701 ();
 sg13g2_fill_1 FILLER_43_718 ();
 sg13g2_fill_1 FILLER_43_723 ();
 sg13g2_fill_1 FILLER_43_729 ();
 sg13g2_fill_2 FILLER_43_735 ();
 sg13g2_fill_1 FILLER_43_741 ();
 sg13g2_decap_4 FILLER_43_747 ();
 sg13g2_fill_1 FILLER_43_751 ();
 sg13g2_fill_2 FILLER_43_761 ();
 sg13g2_fill_2 FILLER_43_768 ();
 sg13g2_fill_1 FILLER_43_770 ();
 sg13g2_fill_2 FILLER_43_818 ();
 sg13g2_fill_1 FILLER_43_862 ();
 sg13g2_fill_2 FILLER_43_875 ();
 sg13g2_fill_1 FILLER_43_903 ();
 sg13g2_fill_1 FILLER_43_912 ();
 sg13g2_fill_2 FILLER_43_918 ();
 sg13g2_fill_2 FILLER_43_924 ();
 sg13g2_decap_4 FILLER_43_934 ();
 sg13g2_fill_1 FILLER_43_938 ();
 sg13g2_fill_1 FILLER_43_973 ();
 sg13g2_fill_2 FILLER_43_986 ();
 sg13g2_fill_1 FILLER_43_1017 ();
 sg13g2_fill_2 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_43_1028 ();
 sg13g2_decap_4 FILLER_43_1035 ();
 sg13g2_fill_2 FILLER_43_1039 ();
 sg13g2_fill_2 FILLER_43_1045 ();
 sg13g2_fill_2 FILLER_43_1096 ();
 sg13g2_fill_2 FILLER_43_1115 ();
 sg13g2_decap_4 FILLER_43_1148 ();
 sg13g2_fill_2 FILLER_43_1171 ();
 sg13g2_fill_1 FILLER_43_1173 ();
 sg13g2_fill_1 FILLER_43_1190 ();
 sg13g2_decap_8 FILLER_43_1207 ();
 sg13g2_decap_8 FILLER_43_1214 ();
 sg13g2_decap_8 FILLER_43_1221 ();
 sg13g2_decap_8 FILLER_43_1228 ();
 sg13g2_decap_8 FILLER_43_1235 ();
 sg13g2_decap_8 FILLER_43_1242 ();
 sg13g2_decap_8 FILLER_43_1249 ();
 sg13g2_decap_8 FILLER_43_1256 ();
 sg13g2_decap_8 FILLER_43_1263 ();
 sg13g2_decap_8 FILLER_43_1270 ();
 sg13g2_decap_8 FILLER_43_1277 ();
 sg13g2_decap_8 FILLER_43_1284 ();
 sg13g2_decap_8 FILLER_43_1291 ();
 sg13g2_decap_8 FILLER_43_1298 ();
 sg13g2_decap_8 FILLER_43_1305 ();
 sg13g2_decap_8 FILLER_43_1312 ();
 sg13g2_decap_8 FILLER_43_1319 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_44 ();
 sg13g2_fill_1 FILLER_44_92 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_106 ();
 sg13g2_fill_2 FILLER_44_112 ();
 sg13g2_fill_2 FILLER_44_119 ();
 sg13g2_fill_2 FILLER_44_125 ();
 sg13g2_fill_1 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_149 ();
 sg13g2_fill_1 FILLER_44_156 ();
 sg13g2_decap_4 FILLER_44_170 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_fill_2 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_201 ();
 sg13g2_fill_2 FILLER_44_206 ();
 sg13g2_fill_2 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_214 ();
 sg13g2_decap_4 FILLER_44_219 ();
 sg13g2_fill_2 FILLER_44_270 ();
 sg13g2_fill_2 FILLER_44_319 ();
 sg13g2_fill_1 FILLER_44_321 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_fill_1 FILLER_44_398 ();
 sg13g2_fill_1 FILLER_44_409 ();
 sg13g2_fill_1 FILLER_44_415 ();
 sg13g2_fill_2 FILLER_44_435 ();
 sg13g2_fill_1 FILLER_44_437 ();
 sg13g2_fill_1 FILLER_44_464 ();
 sg13g2_fill_2 FILLER_44_495 ();
 sg13g2_fill_1 FILLER_44_505 ();
 sg13g2_fill_2 FILLER_44_510 ();
 sg13g2_fill_2 FILLER_44_535 ();
 sg13g2_fill_1 FILLER_44_537 ();
 sg13g2_fill_2 FILLER_44_565 ();
 sg13g2_fill_1 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_572 ();
 sg13g2_fill_1 FILLER_44_608 ();
 sg13g2_fill_2 FILLER_44_617 ();
 sg13g2_fill_2 FILLER_44_624 ();
 sg13g2_fill_2 FILLER_44_652 ();
 sg13g2_fill_1 FILLER_44_654 ();
 sg13g2_fill_2 FILLER_44_660 ();
 sg13g2_fill_1 FILLER_44_662 ();
 sg13g2_decap_8 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_692 ();
 sg13g2_decap_8 FILLER_44_698 ();
 sg13g2_fill_1 FILLER_44_713 ();
 sg13g2_fill_1 FILLER_44_721 ();
 sg13g2_fill_1 FILLER_44_735 ();
 sg13g2_fill_2 FILLER_44_740 ();
 sg13g2_fill_1 FILLER_44_791 ();
 sg13g2_decap_4 FILLER_44_796 ();
 sg13g2_fill_2 FILLER_44_808 ();
 sg13g2_fill_1 FILLER_44_810 ();
 sg13g2_fill_1 FILLER_44_828 ();
 sg13g2_fill_2 FILLER_44_843 ();
 sg13g2_fill_2 FILLER_44_855 ();
 sg13g2_fill_1 FILLER_44_865 ();
 sg13g2_fill_1 FILLER_44_870 ();
 sg13g2_fill_1 FILLER_44_901 ();
 sg13g2_fill_2 FILLER_44_914 ();
 sg13g2_fill_1 FILLER_44_942 ();
 sg13g2_fill_2 FILLER_44_950 ();
 sg13g2_fill_2 FILLER_44_999 ();
 sg13g2_fill_1 FILLER_44_1009 ();
 sg13g2_fill_1 FILLER_44_1015 ();
 sg13g2_decap_8 FILLER_44_1058 ();
 sg13g2_fill_1 FILLER_44_1091 ();
 sg13g2_fill_2 FILLER_44_1135 ();
 sg13g2_fill_1 FILLER_44_1137 ();
 sg13g2_decap_4 FILLER_44_1147 ();
 sg13g2_fill_2 FILLER_44_1156 ();
 sg13g2_fill_2 FILLER_44_1171 ();
 sg13g2_decap_4 FILLER_44_1177 ();
 sg13g2_fill_1 FILLER_44_1181 ();
 sg13g2_fill_1 FILLER_44_1195 ();
 sg13g2_decap_8 FILLER_44_1204 ();
 sg13g2_decap_8 FILLER_44_1211 ();
 sg13g2_decap_8 FILLER_44_1218 ();
 sg13g2_decap_8 FILLER_44_1225 ();
 sg13g2_decap_8 FILLER_44_1232 ();
 sg13g2_decap_8 FILLER_44_1239 ();
 sg13g2_decap_8 FILLER_44_1246 ();
 sg13g2_decap_8 FILLER_44_1253 ();
 sg13g2_decap_8 FILLER_44_1260 ();
 sg13g2_decap_8 FILLER_44_1267 ();
 sg13g2_decap_8 FILLER_44_1274 ();
 sg13g2_decap_8 FILLER_44_1281 ();
 sg13g2_decap_8 FILLER_44_1288 ();
 sg13g2_decap_8 FILLER_44_1295 ();
 sg13g2_decap_8 FILLER_44_1302 ();
 sg13g2_decap_8 FILLER_44_1309 ();
 sg13g2_decap_8 FILLER_44_1316 ();
 sg13g2_fill_2 FILLER_44_1323 ();
 sg13g2_fill_1 FILLER_44_1325 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_39 ();
 sg13g2_decap_4 FILLER_45_46 ();
 sg13g2_fill_1 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_100 ();
 sg13g2_fill_1 FILLER_45_128 ();
 sg13g2_fill_1 FILLER_45_134 ();
 sg13g2_fill_1 FILLER_45_161 ();
 sg13g2_fill_2 FILLER_45_193 ();
 sg13g2_fill_1 FILLER_45_195 ();
 sg13g2_fill_2 FILLER_45_242 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_1 FILLER_45_254 ();
 sg13g2_fill_2 FILLER_45_259 ();
 sg13g2_fill_1 FILLER_45_269 ();
 sg13g2_fill_1 FILLER_45_296 ();
 sg13g2_fill_1 FILLER_45_302 ();
 sg13g2_decap_4 FILLER_45_313 ();
 sg13g2_fill_2 FILLER_45_317 ();
 sg13g2_fill_1 FILLER_45_331 ();
 sg13g2_fill_2 FILLER_45_351 ();
 sg13g2_decap_4 FILLER_45_374 ();
 sg13g2_fill_2 FILLER_45_390 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_fill_1 FILLER_45_435 ();
 sg13g2_fill_2 FILLER_45_475 ();
 sg13g2_fill_1 FILLER_45_477 ();
 sg13g2_fill_1 FILLER_45_482 ();
 sg13g2_fill_2 FILLER_45_487 ();
 sg13g2_fill_1 FILLER_45_494 ();
 sg13g2_fill_2 FILLER_45_501 ();
 sg13g2_fill_2 FILLER_45_509 ();
 sg13g2_fill_2 FILLER_45_515 ();
 sg13g2_fill_1 FILLER_45_517 ();
 sg13g2_fill_2 FILLER_45_544 ();
 sg13g2_fill_2 FILLER_45_576 ();
 sg13g2_fill_1 FILLER_45_578 ();
 sg13g2_fill_2 FILLER_45_588 ();
 sg13g2_fill_1 FILLER_45_590 ();
 sg13g2_fill_1 FILLER_45_596 ();
 sg13g2_fill_1 FILLER_45_602 ();
 sg13g2_fill_1 FILLER_45_607 ();
 sg13g2_fill_1 FILLER_45_612 ();
 sg13g2_decap_4 FILLER_45_617 ();
 sg13g2_fill_1 FILLER_45_621 ();
 sg13g2_fill_1 FILLER_45_628 ();
 sg13g2_fill_1 FILLER_45_732 ();
 sg13g2_fill_1 FILLER_45_738 ();
 sg13g2_fill_1 FILLER_45_747 ();
 sg13g2_fill_1 FILLER_45_796 ();
 sg13g2_fill_1 FILLER_45_801 ();
 sg13g2_decap_4 FILLER_45_814 ();
 sg13g2_fill_2 FILLER_45_818 ();
 sg13g2_fill_2 FILLER_45_854 ();
 sg13g2_fill_1 FILLER_45_860 ();
 sg13g2_fill_2 FILLER_45_873 ();
 sg13g2_fill_1 FILLER_45_888 ();
 sg13g2_fill_2 FILLER_45_893 ();
 sg13g2_fill_1 FILLER_45_910 ();
 sg13g2_fill_2 FILLER_45_965 ();
 sg13g2_fill_1 FILLER_45_971 ();
 sg13g2_fill_2 FILLER_45_1002 ();
 sg13g2_fill_1 FILLER_45_1004 ();
 sg13g2_fill_2 FILLER_45_1013 ();
 sg13g2_decap_4 FILLER_45_1035 ();
 sg13g2_fill_2 FILLER_45_1039 ();
 sg13g2_fill_1 FILLER_45_1076 ();
 sg13g2_decap_8 FILLER_45_1112 ();
 sg13g2_decap_8 FILLER_45_1119 ();
 sg13g2_fill_2 FILLER_45_1126 ();
 sg13g2_fill_1 FILLER_45_1128 ();
 sg13g2_fill_1 FILLER_45_1147 ();
 sg13g2_fill_2 FILLER_45_1152 ();
 sg13g2_fill_2 FILLER_45_1166 ();
 sg13g2_decap_8 FILLER_45_1203 ();
 sg13g2_decap_8 FILLER_45_1210 ();
 sg13g2_decap_8 FILLER_45_1217 ();
 sg13g2_decap_8 FILLER_45_1224 ();
 sg13g2_decap_8 FILLER_45_1231 ();
 sg13g2_decap_8 FILLER_45_1238 ();
 sg13g2_decap_8 FILLER_45_1245 ();
 sg13g2_decap_8 FILLER_45_1252 ();
 sg13g2_decap_8 FILLER_45_1259 ();
 sg13g2_decap_8 FILLER_45_1266 ();
 sg13g2_decap_8 FILLER_45_1273 ();
 sg13g2_decap_8 FILLER_45_1280 ();
 sg13g2_decap_8 FILLER_45_1287 ();
 sg13g2_decap_8 FILLER_45_1294 ();
 sg13g2_decap_8 FILLER_45_1301 ();
 sg13g2_decap_8 FILLER_45_1308 ();
 sg13g2_decap_8 FILLER_45_1315 ();
 sg13g2_decap_4 FILLER_45_1322 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_fill_2 FILLER_46_58 ();
 sg13g2_fill_1 FILLER_46_60 ();
 sg13g2_fill_2 FILLER_46_89 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_2 FILLER_46_103 ();
 sg13g2_fill_1 FILLER_46_109 ();
 sg13g2_fill_1 FILLER_46_145 ();
 sg13g2_fill_2 FILLER_46_180 ();
 sg13g2_fill_2 FILLER_46_207 ();
 sg13g2_fill_2 FILLER_46_213 ();
 sg13g2_fill_1 FILLER_46_215 ();
 sg13g2_fill_1 FILLER_46_220 ();
 sg13g2_fill_2 FILLER_46_225 ();
 sg13g2_fill_1 FILLER_46_227 ();
 sg13g2_decap_4 FILLER_46_245 ();
 sg13g2_fill_1 FILLER_46_249 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_fill_2 FILLER_46_320 ();
 sg13g2_fill_1 FILLER_46_353 ();
 sg13g2_fill_1 FILLER_46_361 ();
 sg13g2_fill_2 FILLER_46_369 ();
 sg13g2_fill_1 FILLER_46_389 ();
 sg13g2_decap_4 FILLER_46_394 ();
 sg13g2_fill_2 FILLER_46_403 ();
 sg13g2_fill_1 FILLER_46_409 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_fill_1 FILLER_46_442 ();
 sg13g2_fill_2 FILLER_46_460 ();
 sg13g2_fill_2 FILLER_46_466 ();
 sg13g2_fill_1 FILLER_46_472 ();
 sg13g2_decap_4 FILLER_46_477 ();
 sg13g2_fill_2 FILLER_46_529 ();
 sg13g2_fill_1 FILLER_46_535 ();
 sg13g2_fill_1 FILLER_46_544 ();
 sg13g2_fill_1 FILLER_46_550 ();
 sg13g2_fill_1 FILLER_46_635 ();
 sg13g2_fill_1 FILLER_46_645 ();
 sg13g2_fill_2 FILLER_46_650 ();
 sg13g2_decap_4 FILLER_46_656 ();
 sg13g2_fill_2 FILLER_46_660 ();
 sg13g2_decap_4 FILLER_46_678 ();
 sg13g2_fill_1 FILLER_46_687 ();
 sg13g2_fill_1 FILLER_46_696 ();
 sg13g2_fill_1 FILLER_46_701 ();
 sg13g2_fill_1 FILLER_46_707 ();
 sg13g2_decap_4 FILLER_46_761 ();
 sg13g2_fill_1 FILLER_46_765 ();
 sg13g2_fill_2 FILLER_46_865 ();
 sg13g2_fill_1 FILLER_46_867 ();
 sg13g2_fill_1 FILLER_46_910 ();
 sg13g2_decap_4 FILLER_46_979 ();
 sg13g2_fill_1 FILLER_46_983 ();
 sg13g2_fill_2 FILLER_46_1017 ();
 sg13g2_fill_2 FILLER_46_1049 ();
 sg13g2_fill_2 FILLER_46_1077 ();
 sg13g2_fill_1 FILLER_46_1079 ();
 sg13g2_fill_2 FILLER_46_1085 ();
 sg13g2_fill_1 FILLER_46_1087 ();
 sg13g2_fill_2 FILLER_46_1092 ();
 sg13g2_fill_1 FILLER_46_1094 ();
 sg13g2_fill_1 FILLER_46_1160 ();
 sg13g2_fill_1 FILLER_46_1169 ();
 sg13g2_fill_2 FILLER_46_1182 ();
 sg13g2_decap_8 FILLER_46_1196 ();
 sg13g2_decap_8 FILLER_46_1203 ();
 sg13g2_decap_8 FILLER_46_1210 ();
 sg13g2_decap_8 FILLER_46_1217 ();
 sg13g2_decap_8 FILLER_46_1224 ();
 sg13g2_decap_8 FILLER_46_1231 ();
 sg13g2_decap_8 FILLER_46_1238 ();
 sg13g2_decap_8 FILLER_46_1245 ();
 sg13g2_decap_8 FILLER_46_1252 ();
 sg13g2_decap_8 FILLER_46_1259 ();
 sg13g2_decap_8 FILLER_46_1266 ();
 sg13g2_decap_8 FILLER_46_1273 ();
 sg13g2_decap_8 FILLER_46_1280 ();
 sg13g2_decap_8 FILLER_46_1287 ();
 sg13g2_decap_8 FILLER_46_1294 ();
 sg13g2_decap_8 FILLER_46_1301 ();
 sg13g2_decap_8 FILLER_46_1308 ();
 sg13g2_decap_8 FILLER_46_1315 ();
 sg13g2_decap_4 FILLER_46_1322 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_fill_2 FILLER_47_76 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_97 ();
 sg13g2_fill_1 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_113 ();
 sg13g2_fill_2 FILLER_47_118 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_fill_2 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_263 ();
 sg13g2_decap_8 FILLER_47_269 ();
 sg13g2_fill_2 FILLER_47_276 ();
 sg13g2_fill_1 FILLER_47_282 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_fill_1 FILLER_47_356 ();
 sg13g2_fill_2 FILLER_47_366 ();
 sg13g2_fill_2 FILLER_47_377 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_decap_4 FILLER_47_451 ();
 sg13g2_decap_4 FILLER_47_485 ();
 sg13g2_fill_2 FILLER_47_525 ();
 sg13g2_fill_1 FILLER_47_527 ();
 sg13g2_fill_2 FILLER_47_567 ();
 sg13g2_fill_1 FILLER_47_573 ();
 sg13g2_fill_1 FILLER_47_578 ();
 sg13g2_fill_2 FILLER_47_583 ();
 sg13g2_fill_1 FILLER_47_585 ();
 sg13g2_fill_1 FILLER_47_599 ();
 sg13g2_fill_2 FILLER_47_638 ();
 sg13g2_fill_1 FILLER_47_640 ();
 sg13g2_fill_1 FILLER_47_650 ();
 sg13g2_fill_2 FILLER_47_681 ();
 sg13g2_fill_1 FILLER_47_744 ();
 sg13g2_fill_1 FILLER_47_776 ();
 sg13g2_decap_8 FILLER_47_815 ();
 sg13g2_fill_2 FILLER_47_822 ();
 sg13g2_fill_1 FILLER_47_824 ();
 sg13g2_fill_1 FILLER_47_839 ();
 sg13g2_fill_2 FILLER_47_884 ();
 sg13g2_fill_2 FILLER_47_890 ();
 sg13g2_fill_2 FILLER_47_897 ();
 sg13g2_fill_2 FILLER_47_903 ();
 sg13g2_fill_2 FILLER_47_914 ();
 sg13g2_fill_1 FILLER_47_916 ();
 sg13g2_fill_2 FILLER_47_931 ();
 sg13g2_fill_1 FILLER_47_957 ();
 sg13g2_fill_1 FILLER_47_989 ();
 sg13g2_fill_2 FILLER_47_1008 ();
 sg13g2_fill_2 FILLER_47_1031 ();
 sg13g2_fill_1 FILLER_47_1033 ();
 sg13g2_fill_2 FILLER_47_1039 ();
 sg13g2_fill_1 FILLER_47_1041 ();
 sg13g2_fill_1 FILLER_47_1052 ();
 sg13g2_fill_1 FILLER_47_1057 ();
 sg13g2_fill_2 FILLER_47_1066 ();
 sg13g2_fill_1 FILLER_47_1068 ();
 sg13g2_fill_2 FILLER_47_1103 ();
 sg13g2_fill_2 FILLER_47_1121 ();
 sg13g2_fill_1 FILLER_47_1127 ();
 sg13g2_fill_2 FILLER_47_1202 ();
 sg13g2_fill_1 FILLER_47_1204 ();
 sg13g2_fill_1 FILLER_47_1209 ();
 sg13g2_decap_8 FILLER_47_1223 ();
 sg13g2_decap_8 FILLER_47_1230 ();
 sg13g2_decap_8 FILLER_47_1237 ();
 sg13g2_decap_8 FILLER_47_1244 ();
 sg13g2_decap_8 FILLER_47_1251 ();
 sg13g2_decap_8 FILLER_47_1258 ();
 sg13g2_decap_8 FILLER_47_1265 ();
 sg13g2_decap_8 FILLER_47_1272 ();
 sg13g2_decap_8 FILLER_47_1279 ();
 sg13g2_decap_8 FILLER_47_1286 ();
 sg13g2_decap_8 FILLER_47_1293 ();
 sg13g2_decap_8 FILLER_47_1300 ();
 sg13g2_decap_8 FILLER_47_1307 ();
 sg13g2_decap_8 FILLER_47_1314 ();
 sg13g2_decap_4 FILLER_47_1321 ();
 sg13g2_fill_1 FILLER_47_1325 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_fill_2 FILLER_48_64 ();
 sg13g2_fill_1 FILLER_48_71 ();
 sg13g2_fill_1 FILLER_48_76 ();
 sg13g2_fill_2 FILLER_48_86 ();
 sg13g2_fill_1 FILLER_48_88 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_fill_2 FILLER_48_219 ();
 sg13g2_fill_2 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_227 ();
 sg13g2_fill_2 FILLER_48_233 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_2 FILLER_48_241 ();
 sg13g2_fill_2 FILLER_48_262 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_decap_4 FILLER_48_322 ();
 sg13g2_fill_1 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_331 ();
 sg13g2_fill_2 FILLER_48_338 ();
 sg13g2_fill_1 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_407 ();
 sg13g2_fill_1 FILLER_48_423 ();
 sg13g2_fill_1 FILLER_48_431 ();
 sg13g2_decap_4 FILLER_48_440 ();
 sg13g2_fill_2 FILLER_48_448 ();
 sg13g2_fill_1 FILLER_48_450 ();
 sg13g2_fill_2 FILLER_48_455 ();
 sg13g2_fill_1 FILLER_48_496 ();
 sg13g2_fill_1 FILLER_48_519 ();
 sg13g2_decap_8 FILLER_48_533 ();
 sg13g2_decap_4 FILLER_48_540 ();
 sg13g2_fill_1 FILLER_48_544 ();
 sg13g2_fill_2 FILLER_48_677 ();
 sg13g2_fill_1 FILLER_48_708 ();
 sg13g2_fill_2 FILLER_48_726 ();
 sg13g2_fill_1 FILLER_48_732 ();
 sg13g2_fill_1 FILLER_48_777 ();
 sg13g2_fill_1 FILLER_48_787 ();
 sg13g2_decap_4 FILLER_48_814 ();
 sg13g2_fill_2 FILLER_48_818 ();
 sg13g2_fill_2 FILLER_48_829 ();
 sg13g2_fill_1 FILLER_48_831 ();
 sg13g2_fill_2 FILLER_48_854 ();
 sg13g2_fill_1 FILLER_48_865 ();
 sg13g2_fill_2 FILLER_48_917 ();
 sg13g2_fill_1 FILLER_48_924 ();
 sg13g2_fill_2 FILLER_48_949 ();
 sg13g2_fill_2 FILLER_48_972 ();
 sg13g2_fill_2 FILLER_48_979 ();
 sg13g2_fill_1 FILLER_48_981 ();
 sg13g2_fill_2 FILLER_48_1039 ();
 sg13g2_fill_1 FILLER_48_1084 ();
 sg13g2_fill_1 FILLER_48_1089 ();
 sg13g2_decap_4 FILLER_48_1099 ();
 sg13g2_fill_1 FILLER_48_1116 ();
 sg13g2_fill_2 FILLER_48_1121 ();
 sg13g2_fill_1 FILLER_48_1123 ();
 sg13g2_fill_2 FILLER_48_1139 ();
 sg13g2_fill_2 FILLER_48_1146 ();
 sg13g2_fill_1 FILLER_48_1148 ();
 sg13g2_fill_1 FILLER_48_1154 ();
 sg13g2_fill_2 FILLER_48_1160 ();
 sg13g2_fill_1 FILLER_48_1162 ();
 sg13g2_fill_2 FILLER_48_1190 ();
 sg13g2_fill_2 FILLER_48_1196 ();
 sg13g2_decap_8 FILLER_48_1237 ();
 sg13g2_decap_8 FILLER_48_1244 ();
 sg13g2_decap_8 FILLER_48_1251 ();
 sg13g2_decap_8 FILLER_48_1258 ();
 sg13g2_decap_8 FILLER_48_1265 ();
 sg13g2_decap_8 FILLER_48_1272 ();
 sg13g2_decap_8 FILLER_48_1279 ();
 sg13g2_decap_8 FILLER_48_1286 ();
 sg13g2_decap_8 FILLER_48_1293 ();
 sg13g2_decap_8 FILLER_48_1300 ();
 sg13g2_decap_8 FILLER_48_1307 ();
 sg13g2_decap_8 FILLER_48_1314 ();
 sg13g2_decap_4 FILLER_48_1321 ();
 sg13g2_fill_1 FILLER_48_1325 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_139 ();
 sg13g2_fill_2 FILLER_49_203 ();
 sg13g2_fill_1 FILLER_49_259 ();
 sg13g2_fill_1 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_317 ();
 sg13g2_fill_2 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_383 ();
 sg13g2_decap_8 FILLER_49_418 ();
 sg13g2_fill_1 FILLER_49_425 ();
 sg13g2_fill_2 FILLER_49_465 ();
 sg13g2_fill_1 FILLER_49_467 ();
 sg13g2_fill_2 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_474 ();
 sg13g2_fill_2 FILLER_49_484 ();
 sg13g2_fill_1 FILLER_49_486 ();
 sg13g2_fill_1 FILLER_49_491 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_fill_1 FILLER_49_540 ();
 sg13g2_fill_1 FILLER_49_571 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_fill_1 FILLER_49_591 ();
 sg13g2_fill_1 FILLER_49_596 ();
 sg13g2_decap_4 FILLER_49_601 ();
 sg13g2_fill_1 FILLER_49_644 ();
 sg13g2_decap_4 FILLER_49_662 ();
 sg13g2_fill_2 FILLER_49_666 ();
 sg13g2_decap_4 FILLER_49_672 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_fill_1 FILLER_49_709 ();
 sg13g2_fill_2 FILLER_49_750 ();
 sg13g2_fill_1 FILLER_49_787 ();
 sg13g2_fill_1 FILLER_49_792 ();
 sg13g2_fill_2 FILLER_49_819 ();
 sg13g2_fill_2 FILLER_49_825 ();
 sg13g2_fill_1 FILLER_49_833 ();
 sg13g2_fill_1 FILLER_49_849 ();
 sg13g2_fill_1 FILLER_49_858 ();
 sg13g2_fill_2 FILLER_49_894 ();
 sg13g2_decap_4 FILLER_49_899 ();
 sg13g2_fill_1 FILLER_49_903 ();
 sg13g2_fill_1 FILLER_49_936 ();
 sg13g2_fill_2 FILLER_49_941 ();
 sg13g2_fill_1 FILLER_49_947 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_fill_2 FILLER_49_980 ();
 sg13g2_fill_2 FILLER_49_986 ();
 sg13g2_fill_2 FILLER_49_1017 ();
 sg13g2_fill_1 FILLER_49_1019 ();
 sg13g2_fill_2 FILLER_49_1174 ();
 sg13g2_decap_4 FILLER_49_1181 ();
 sg13g2_decap_8 FILLER_49_1246 ();
 sg13g2_decap_8 FILLER_49_1253 ();
 sg13g2_decap_8 FILLER_49_1260 ();
 sg13g2_decap_8 FILLER_49_1267 ();
 sg13g2_decap_8 FILLER_49_1274 ();
 sg13g2_decap_8 FILLER_49_1281 ();
 sg13g2_decap_8 FILLER_49_1288 ();
 sg13g2_decap_8 FILLER_49_1295 ();
 sg13g2_decap_8 FILLER_49_1302 ();
 sg13g2_decap_8 FILLER_49_1309 ();
 sg13g2_decap_8 FILLER_49_1316 ();
 sg13g2_fill_2 FILLER_49_1323 ();
 sg13g2_fill_1 FILLER_49_1325 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_4 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_46 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_fill_2 FILLER_50_73 ();
 sg13g2_fill_1 FILLER_50_75 ();
 sg13g2_fill_1 FILLER_50_85 ();
 sg13g2_fill_2 FILLER_50_90 ();
 sg13g2_fill_2 FILLER_50_102 ();
 sg13g2_fill_1 FILLER_50_130 ();
 sg13g2_fill_2 FILLER_50_144 ();
 sg13g2_fill_2 FILLER_50_178 ();
 sg13g2_fill_1 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_232 ();
 sg13g2_fill_1 FILLER_50_275 ();
 sg13g2_fill_1 FILLER_50_288 ();
 sg13g2_fill_2 FILLER_50_297 ();
 sg13g2_fill_1 FILLER_50_303 ();
 sg13g2_decap_4 FILLER_50_350 ();
 sg13g2_fill_2 FILLER_50_371 ();
 sg13g2_fill_1 FILLER_50_399 ();
 sg13g2_fill_2 FILLER_50_428 ();
 sg13g2_fill_1 FILLER_50_430 ();
 sg13g2_fill_1 FILLER_50_444 ();
 sg13g2_decap_4 FILLER_50_449 ();
 sg13g2_fill_2 FILLER_50_453 ();
 sg13g2_decap_4 FILLER_50_459 ();
 sg13g2_decap_4 FILLER_50_510 ();
 sg13g2_fill_1 FILLER_50_527 ();
 sg13g2_fill_1 FILLER_50_541 ();
 sg13g2_decap_8 FILLER_50_546 ();
 sg13g2_fill_1 FILLER_50_553 ();
 sg13g2_fill_1 FILLER_50_558 ();
 sg13g2_fill_2 FILLER_50_563 ();
 sg13g2_fill_1 FILLER_50_612 ();
 sg13g2_fill_1 FILLER_50_624 ();
 sg13g2_fill_1 FILLER_50_630 ();
 sg13g2_fill_2 FILLER_50_647 ();
 sg13g2_fill_2 FILLER_50_719 ();
 sg13g2_fill_2 FILLER_50_725 ();
 sg13g2_fill_2 FILLER_50_736 ();
 sg13g2_fill_2 FILLER_50_758 ();
 sg13g2_fill_1 FILLER_50_760 ();
 sg13g2_fill_2 FILLER_50_787 ();
 sg13g2_fill_2 FILLER_50_819 ();
 sg13g2_fill_1 FILLER_50_826 ();
 sg13g2_fill_2 FILLER_50_886 ();
 sg13g2_fill_1 FILLER_50_918 ();
 sg13g2_fill_2 FILLER_50_971 ();
 sg13g2_fill_2 FILLER_50_977 ();
 sg13g2_fill_1 FILLER_50_979 ();
 sg13g2_fill_1 FILLER_50_997 ();
 sg13g2_fill_1 FILLER_50_1003 ();
 sg13g2_fill_1 FILLER_50_1008 ();
 sg13g2_fill_2 FILLER_50_1046 ();
 sg13g2_fill_2 FILLER_50_1053 ();
 sg13g2_decap_4 FILLER_50_1068 ();
 sg13g2_decap_4 FILLER_50_1076 ();
 sg13g2_fill_2 FILLER_50_1084 ();
 sg13g2_fill_1 FILLER_50_1086 ();
 sg13g2_fill_1 FILLER_50_1099 ();
 sg13g2_fill_1 FILLER_50_1105 ();
 sg13g2_fill_1 FILLER_50_1165 ();
 sg13g2_fill_2 FILLER_50_1170 ();
 sg13g2_fill_2 FILLER_50_1236 ();
 sg13g2_fill_1 FILLER_50_1238 ();
 sg13g2_decap_4 FILLER_50_1244 ();
 sg13g2_decap_8 FILLER_50_1252 ();
 sg13g2_decap_8 FILLER_50_1259 ();
 sg13g2_decap_8 FILLER_50_1266 ();
 sg13g2_decap_8 FILLER_50_1273 ();
 sg13g2_decap_8 FILLER_50_1280 ();
 sg13g2_decap_8 FILLER_50_1287 ();
 sg13g2_decap_8 FILLER_50_1294 ();
 sg13g2_decap_8 FILLER_50_1301 ();
 sg13g2_decap_8 FILLER_50_1308 ();
 sg13g2_decap_8 FILLER_50_1315 ();
 sg13g2_decap_4 FILLER_50_1322 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_4 FILLER_51_42 ();
 sg13g2_fill_2 FILLER_51_46 ();
 sg13g2_fill_1 FILLER_51_61 ();
 sg13g2_fill_1 FILLER_51_68 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_2 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_133 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_fill_1 FILLER_51_208 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_fill_1 FILLER_51_234 ();
 sg13g2_fill_2 FILLER_51_240 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_2 FILLER_51_278 ();
 sg13g2_fill_1 FILLER_51_284 ();
 sg13g2_fill_1 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_295 ();
 sg13g2_fill_1 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_311 ();
 sg13g2_decap_4 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_325 ();
 sg13g2_decap_4 FILLER_51_331 ();
 sg13g2_fill_2 FILLER_51_352 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_367 ();
 sg13g2_fill_1 FILLER_51_369 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_437 ();
 sg13g2_fill_1 FILLER_51_464 ();
 sg13g2_fill_1 FILLER_51_469 ();
 sg13g2_fill_2 FILLER_51_474 ();
 sg13g2_fill_1 FILLER_51_485 ();
 sg13g2_fill_1 FILLER_51_495 ();
 sg13g2_fill_1 FILLER_51_501 ();
 sg13g2_decap_4 FILLER_51_526 ();
 sg13g2_fill_1 FILLER_51_530 ();
 sg13g2_fill_1 FILLER_51_604 ();
 sg13g2_fill_1 FILLER_51_608 ();
 sg13g2_fill_2 FILLER_51_650 ();
 sg13g2_fill_1 FILLER_51_660 ();
 sg13g2_fill_1 FILLER_51_665 ();
 sg13g2_fill_1 FILLER_51_670 ();
 sg13g2_decap_4 FILLER_51_711 ();
 sg13g2_fill_2 FILLER_51_715 ();
 sg13g2_fill_2 FILLER_51_721 ();
 sg13g2_fill_1 FILLER_51_723 ();
 sg13g2_fill_1 FILLER_51_747 ();
 sg13g2_fill_1 FILLER_51_753 ();
 sg13g2_fill_2 FILLER_51_797 ();
 sg13g2_fill_1 FILLER_51_849 ();
 sg13g2_fill_2 FILLER_51_867 ();
 sg13g2_fill_2 FILLER_51_873 ();
 sg13g2_decap_4 FILLER_51_905 ();
 sg13g2_fill_2 FILLER_51_909 ();
 sg13g2_fill_2 FILLER_51_920 ();
 sg13g2_fill_1 FILLER_51_922 ();
 sg13g2_fill_2 FILLER_51_958 ();
 sg13g2_decap_4 FILLER_51_995 ();
 sg13g2_fill_2 FILLER_51_1029 ();
 sg13g2_fill_2 FILLER_51_1061 ();
 sg13g2_fill_2 FILLER_51_1067 ();
 sg13g2_fill_1 FILLER_51_1069 ();
 sg13g2_decap_4 FILLER_51_1087 ();
 sg13g2_fill_2 FILLER_51_1091 ();
 sg13g2_fill_2 FILLER_51_1153 ();
 sg13g2_fill_1 FILLER_51_1159 ();
 sg13g2_fill_2 FILLER_51_1164 ();
 sg13g2_fill_1 FILLER_51_1170 ();
 sg13g2_fill_2 FILLER_51_1176 ();
 sg13g2_fill_2 FILLER_51_1191 ();
 sg13g2_fill_1 FILLER_51_1197 ();
 sg13g2_fill_2 FILLER_51_1237 ();
 sg13g2_decap_8 FILLER_51_1270 ();
 sg13g2_decap_8 FILLER_51_1277 ();
 sg13g2_decap_8 FILLER_51_1284 ();
 sg13g2_decap_8 FILLER_51_1291 ();
 sg13g2_decap_8 FILLER_51_1298 ();
 sg13g2_decap_8 FILLER_51_1305 ();
 sg13g2_decap_8 FILLER_51_1312 ();
 sg13g2_decap_8 FILLER_51_1319 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_33 ();
 sg13g2_decap_4 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_137 ();
 sg13g2_decap_8 FILLER_52_213 ();
 sg13g2_fill_2 FILLER_52_220 ();
 sg13g2_fill_1 FILLER_52_299 ();
 sg13g2_fill_1 FILLER_52_308 ();
 sg13g2_fill_2 FILLER_52_344 ();
 sg13g2_fill_1 FILLER_52_380 ();
 sg13g2_decap_4 FILLER_52_385 ();
 sg13g2_fill_1 FILLER_52_389 ();
 sg13g2_fill_2 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_453 ();
 sg13g2_fill_2 FILLER_52_460 ();
 sg13g2_fill_1 FILLER_52_462 ();
 sg13g2_fill_1 FILLER_52_493 ();
 sg13g2_fill_1 FILLER_52_502 ();
 sg13g2_fill_1 FILLER_52_539 ();
 sg13g2_fill_2 FILLER_52_592 ();
 sg13g2_fill_1 FILLER_52_612 ();
 sg13g2_fill_1 FILLER_52_617 ();
 sg13g2_fill_1 FILLER_52_622 ();
 sg13g2_fill_1 FILLER_52_636 ();
 sg13g2_fill_1 FILLER_52_642 ();
 sg13g2_fill_1 FILLER_52_647 ();
 sg13g2_fill_1 FILLER_52_661 ();
 sg13g2_fill_1 FILLER_52_672 ();
 sg13g2_fill_1 FILLER_52_699 ();
 sg13g2_fill_1 FILLER_52_752 ();
 sg13g2_fill_2 FILLER_52_756 ();
 sg13g2_fill_2 FILLER_52_767 ();
 sg13g2_decap_4 FILLER_52_773 ();
 sg13g2_fill_2 FILLER_52_777 ();
 sg13g2_decap_4 FILLER_52_818 ();
 sg13g2_fill_1 FILLER_52_871 ();
 sg13g2_fill_2 FILLER_52_880 ();
 sg13g2_fill_1 FILLER_52_913 ();
 sg13g2_fill_1 FILLER_52_918 ();
 sg13g2_fill_1 FILLER_52_923 ();
 sg13g2_fill_2 FILLER_52_928 ();
 sg13g2_fill_1 FILLER_52_942 ();
 sg13g2_fill_2 FILLER_52_998 ();
 sg13g2_fill_2 FILLER_52_1005 ();
 sg13g2_fill_2 FILLER_52_1011 ();
 sg13g2_decap_4 FILLER_52_1048 ();
 sg13g2_fill_2 FILLER_52_1103 ();
 sg13g2_decap_4 FILLER_52_1118 ();
 sg13g2_fill_1 FILLER_52_1137 ();
 sg13g2_fill_2 FILLER_52_1146 ();
 sg13g2_fill_1 FILLER_52_1148 ();
 sg13g2_fill_2 FILLER_52_1196 ();
 sg13g2_fill_1 FILLER_52_1198 ();
 sg13g2_fill_1 FILLER_52_1203 ();
 sg13g2_fill_2 FILLER_52_1224 ();
 sg13g2_fill_1 FILLER_52_1226 ();
 sg13g2_decap_8 FILLER_52_1270 ();
 sg13g2_decap_8 FILLER_52_1277 ();
 sg13g2_decap_8 FILLER_52_1284 ();
 sg13g2_decap_8 FILLER_52_1291 ();
 sg13g2_decap_8 FILLER_52_1298 ();
 sg13g2_decap_8 FILLER_52_1305 ();
 sg13g2_decap_8 FILLER_52_1312 ();
 sg13g2_decap_8 FILLER_52_1319 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_fill_2 FILLER_53_49 ();
 sg13g2_fill_1 FILLER_53_51 ();
 sg13g2_fill_2 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_84 ();
 sg13g2_decap_4 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_115 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_fill_1 FILLER_53_188 ();
 sg13g2_fill_2 FILLER_53_197 ();
 sg13g2_fill_2 FILLER_53_237 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_294 ();
 sg13g2_fill_1 FILLER_53_299 ();
 sg13g2_fill_1 FILLER_53_307 ();
 sg13g2_fill_1 FILLER_53_418 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_decap_4 FILLER_53_432 ();
 sg13g2_fill_2 FILLER_53_476 ();
 sg13g2_fill_1 FILLER_53_483 ();
 sg13g2_fill_1 FILLER_53_510 ();
 sg13g2_fill_1 FILLER_53_516 ();
 sg13g2_fill_2 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_570 ();
 sg13g2_fill_2 FILLER_53_632 ();
 sg13g2_fill_1 FILLER_53_634 ();
 sg13g2_fill_2 FILLER_53_654 ();
 sg13g2_fill_1 FILLER_53_672 ();
 sg13g2_fill_1 FILLER_53_678 ();
 sg13g2_decap_8 FILLER_53_683 ();
 sg13g2_decap_4 FILLER_53_690 ();
 sg13g2_fill_1 FILLER_53_703 ();
 sg13g2_fill_1 FILLER_53_708 ();
 sg13g2_fill_1 FILLER_53_713 ();
 sg13g2_fill_2 FILLER_53_722 ();
 sg13g2_fill_2 FILLER_53_727 ();
 sg13g2_fill_1 FILLER_53_732 ();
 sg13g2_fill_1 FILLER_53_741 ();
 sg13g2_fill_1 FILLER_53_746 ();
 sg13g2_decap_8 FILLER_53_785 ();
 sg13g2_fill_1 FILLER_53_792 ();
 sg13g2_decap_8 FILLER_53_797 ();
 sg13g2_decap_8 FILLER_53_804 ();
 sg13g2_fill_2 FILLER_53_811 ();
 sg13g2_fill_2 FILLER_53_821 ();
 sg13g2_fill_2 FILLER_53_832 ();
 sg13g2_fill_2 FILLER_53_902 ();
 sg13g2_decap_4 FILLER_53_908 ();
 sg13g2_fill_2 FILLER_53_947 ();
 sg13g2_fill_2 FILLER_53_966 ();
 sg13g2_decap_8 FILLER_53_972 ();
 sg13g2_fill_2 FILLER_53_979 ();
 sg13g2_fill_1 FILLER_53_981 ();
 sg13g2_fill_2 FILLER_53_1044 ();
 sg13g2_fill_1 FILLER_53_1080 ();
 sg13g2_fill_1 FILLER_53_1094 ();
 sg13g2_fill_2 FILLER_53_1103 ();
 sg13g2_fill_1 FILLER_53_1105 ();
 sg13g2_fill_2 FILLER_53_1147 ();
 sg13g2_fill_1 FILLER_53_1153 ();
 sg13g2_fill_1 FILLER_53_1158 ();
 sg13g2_fill_1 FILLER_53_1164 ();
 sg13g2_fill_2 FILLER_53_1169 ();
 sg13g2_fill_1 FILLER_53_1171 ();
 sg13g2_fill_2 FILLER_53_1181 ();
 sg13g2_fill_1 FILLER_53_1188 ();
 sg13g2_fill_1 FILLER_53_1215 ();
 sg13g2_fill_1 FILLER_53_1242 ();
 sg13g2_decap_8 FILLER_53_1256 ();
 sg13g2_fill_1 FILLER_53_1263 ();
 sg13g2_decap_8 FILLER_53_1268 ();
 sg13g2_decap_8 FILLER_53_1275 ();
 sg13g2_decap_8 FILLER_53_1282 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_8 FILLER_53_1303 ();
 sg13g2_decap_8 FILLER_53_1310 ();
 sg13g2_decap_8 FILLER_53_1317 ();
 sg13g2_fill_2 FILLER_53_1324 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_fill_1 FILLER_54_49 ();
 sg13g2_decap_4 FILLER_54_58 ();
 sg13g2_fill_2 FILLER_54_62 ();
 sg13g2_fill_1 FILLER_54_72 ();
 sg13g2_fill_2 FILLER_54_105 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_fill_2 FILLER_54_116 ();
 sg13g2_fill_1 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_fill_2 FILLER_54_243 ();
 sg13g2_fill_1 FILLER_54_279 ();
 sg13g2_fill_2 FILLER_54_285 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_302 ();
 sg13g2_fill_1 FILLER_54_311 ();
 sg13g2_fill_2 FILLER_54_317 ();
 sg13g2_fill_1 FILLER_54_341 ();
 sg13g2_fill_2 FILLER_54_361 ();
 sg13g2_fill_1 FILLER_54_363 ();
 sg13g2_decap_4 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_381 ();
 sg13g2_fill_1 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_402 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_1 FILLER_54_451 ();
 sg13g2_fill_2 FILLER_54_477 ();
 sg13g2_fill_2 FILLER_54_484 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_fill_1 FILLER_54_492 ();
 sg13g2_fill_2 FILLER_54_498 ();
 sg13g2_fill_2 FILLER_54_522 ();
 sg13g2_fill_2 FILLER_54_542 ();
 sg13g2_fill_2 FILLER_54_576 ();
 sg13g2_fill_2 FILLER_54_587 ();
 sg13g2_fill_2 FILLER_54_593 ();
 sg13g2_fill_1 FILLER_54_595 ();
 sg13g2_fill_1 FILLER_54_600 ();
 sg13g2_fill_2 FILLER_54_605 ();
 sg13g2_fill_1 FILLER_54_612 ();
 sg13g2_fill_2 FILLER_54_617 ();
 sg13g2_fill_1 FILLER_54_619 ();
 sg13g2_fill_1 FILLER_54_631 ();
 sg13g2_fill_2 FILLER_54_636 ();
 sg13g2_fill_1 FILLER_54_638 ();
 sg13g2_fill_1 FILLER_54_652 ();
 sg13g2_fill_1 FILLER_54_665 ();
 sg13g2_decap_8 FILLER_54_670 ();
 sg13g2_fill_2 FILLER_54_677 ();
 sg13g2_fill_2 FILLER_54_745 ();
 sg13g2_fill_1 FILLER_54_747 ();
 sg13g2_fill_2 FILLER_54_761 ();
 sg13g2_fill_1 FILLER_54_767 ();
 sg13g2_fill_1 FILLER_54_794 ();
 sg13g2_fill_1 FILLER_54_799 ();
 sg13g2_fill_1 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_820 ();
 sg13g2_fill_1 FILLER_54_832 ();
 sg13g2_fill_2 FILLER_54_901 ();
 sg13g2_fill_2 FILLER_54_932 ();
 sg13g2_fill_2 FILLER_54_940 ();
 sg13g2_fill_1 FILLER_54_980 ();
 sg13g2_fill_2 FILLER_54_988 ();
 sg13g2_fill_2 FILLER_54_1028 ();
 sg13g2_decap_4 FILLER_54_1048 ();
 sg13g2_fill_2 FILLER_54_1056 ();
 sg13g2_fill_1 FILLER_54_1058 ();
 sg13g2_decap_4 FILLER_54_1063 ();
 sg13g2_fill_2 FILLER_54_1067 ();
 sg13g2_fill_2 FILLER_54_1080 ();
 sg13g2_fill_1 FILLER_54_1092 ();
 sg13g2_fill_1 FILLER_54_1096 ();
 sg13g2_fill_1 FILLER_54_1102 ();
 sg13g2_fill_2 FILLER_54_1111 ();
 sg13g2_fill_2 FILLER_54_1139 ();
 sg13g2_fill_2 FILLER_54_1145 ();
 sg13g2_fill_1 FILLER_54_1147 ();
 sg13g2_fill_1 FILLER_54_1152 ();
 sg13g2_fill_2 FILLER_54_1226 ();
 sg13g2_fill_1 FILLER_54_1228 ();
 sg13g2_fill_2 FILLER_54_1261 ();
 sg13g2_fill_1 FILLER_54_1263 ();
 sg13g2_decap_8 FILLER_54_1268 ();
 sg13g2_decap_8 FILLER_54_1275 ();
 sg13g2_decap_8 FILLER_54_1282 ();
 sg13g2_decap_8 FILLER_54_1289 ();
 sg13g2_decap_8 FILLER_54_1296 ();
 sg13g2_decap_8 FILLER_54_1303 ();
 sg13g2_decap_8 FILLER_54_1310 ();
 sg13g2_decap_8 FILLER_54_1317 ();
 sg13g2_fill_2 FILLER_54_1324 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_4 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_60 ();
 sg13g2_fill_2 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_110 ();
 sg13g2_decap_8 FILLER_55_115 ();
 sg13g2_fill_2 FILLER_55_122 ();
 sg13g2_fill_1 FILLER_55_124 ();
 sg13g2_fill_2 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_178 ();
 sg13g2_fill_1 FILLER_55_180 ();
 sg13g2_fill_2 FILLER_55_185 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_206 ();
 sg13g2_fill_1 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_274 ();
 sg13g2_fill_1 FILLER_55_280 ();
 sg13g2_fill_1 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_315 ();
 sg13g2_fill_1 FILLER_55_326 ();
 sg13g2_fill_1 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_55_447 ();
 sg13g2_fill_2 FILLER_55_474 ();
 sg13g2_fill_1 FILLER_55_511 ();
 sg13g2_fill_1 FILLER_55_541 ();
 sg13g2_fill_1 FILLER_55_547 ();
 sg13g2_fill_1 FILLER_55_574 ();
 sg13g2_fill_1 FILLER_55_606 ();
 sg13g2_fill_2 FILLER_55_614 ();
 sg13g2_fill_1 FILLER_55_616 ();
 sg13g2_fill_2 FILLER_55_697 ();
 sg13g2_fill_1 FILLER_55_699 ();
 sg13g2_fill_2 FILLER_55_715 ();
 sg13g2_fill_1 FILLER_55_717 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_decap_8 FILLER_55_752 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_4 FILLER_55_777 ();
 sg13g2_fill_1 FILLER_55_781 ();
 sg13g2_fill_1 FILLER_55_808 ();
 sg13g2_fill_1 FILLER_55_826 ();
 sg13g2_fill_2 FILLER_55_842 ();
 sg13g2_fill_1 FILLER_55_876 ();
 sg13g2_fill_2 FILLER_55_881 ();
 sg13g2_fill_1 FILLER_55_939 ();
 sg13g2_fill_2 FILLER_55_944 ();
 sg13g2_fill_2 FILLER_55_972 ();
 sg13g2_decap_4 FILLER_55_995 ();
 sg13g2_fill_1 FILLER_55_999 ();
 sg13g2_fill_2 FILLER_55_1012 ();
 sg13g2_fill_1 FILLER_55_1018 ();
 sg13g2_fill_2 FILLER_55_1036 ();
 sg13g2_fill_2 FILLER_55_1041 ();
 sg13g2_fill_1 FILLER_55_1043 ();
 sg13g2_fill_1 FILLER_55_1074 ();
 sg13g2_fill_1 FILLER_55_1080 ();
 sg13g2_fill_2 FILLER_55_1085 ();
 sg13g2_fill_2 FILLER_55_1092 ();
 sg13g2_fill_1 FILLER_55_1102 ();
 sg13g2_fill_1 FILLER_55_1129 ();
 sg13g2_fill_1 FILLER_55_1156 ();
 sg13g2_fill_1 FILLER_55_1162 ();
 sg13g2_fill_2 FILLER_55_1167 ();
 sg13g2_fill_2 FILLER_55_1211 ();
 sg13g2_fill_1 FILLER_55_1213 ();
 sg13g2_fill_1 FILLER_55_1248 ();
 sg13g2_decap_8 FILLER_55_1274 ();
 sg13g2_decap_8 FILLER_55_1281 ();
 sg13g2_decap_8 FILLER_55_1288 ();
 sg13g2_decap_8 FILLER_55_1295 ();
 sg13g2_decap_8 FILLER_55_1302 ();
 sg13g2_decap_8 FILLER_55_1309 ();
 sg13g2_decap_8 FILLER_55_1316 ();
 sg13g2_fill_2 FILLER_55_1323 ();
 sg13g2_fill_1 FILLER_55_1325 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_58 ();
 sg13g2_fill_1 FILLER_56_71 ();
 sg13g2_fill_1 FILLER_56_77 ();
 sg13g2_fill_2 FILLER_56_83 ();
 sg13g2_fill_2 FILLER_56_142 ();
 sg13g2_fill_1 FILLER_56_144 ();
 sg13g2_fill_2 FILLER_56_150 ();
 sg13g2_fill_1 FILLER_56_152 ();
 sg13g2_fill_1 FILLER_56_157 ();
 sg13g2_fill_1 FILLER_56_236 ();
 sg13g2_fill_2 FILLER_56_250 ();
 sg13g2_fill_1 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_257 ();
 sg13g2_fill_1 FILLER_56_302 ();
 sg13g2_fill_1 FILLER_56_308 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_347 ();
 sg13g2_fill_2 FILLER_56_354 ();
 sg13g2_fill_1 FILLER_56_356 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_fill_2 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_fill_2 FILLER_56_392 ();
 sg13g2_fill_2 FILLER_56_411 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_decap_4 FILLER_56_419 ();
 sg13g2_fill_1 FILLER_56_423 ();
 sg13g2_decap_8 FILLER_56_428 ();
 sg13g2_decap_4 FILLER_56_435 ();
 sg13g2_fill_1 FILLER_56_439 ();
 sg13g2_fill_2 FILLER_56_450 ();
 sg13g2_fill_1 FILLER_56_478 ();
 sg13g2_fill_1 FILLER_56_483 ();
 sg13g2_fill_1 FILLER_56_488 ();
 sg13g2_fill_2 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_499 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_fill_2 FILLER_56_530 ();
 sg13g2_fill_2 FILLER_56_536 ();
 sg13g2_fill_2 FILLER_56_577 ();
 sg13g2_fill_1 FILLER_56_579 ();
 sg13g2_fill_2 FILLER_56_585 ();
 sg13g2_fill_1 FILLER_56_587 ();
 sg13g2_fill_2 FILLER_56_596 ();
 sg13g2_fill_1 FILLER_56_598 ();
 sg13g2_fill_2 FILLER_56_627 ();
 sg13g2_fill_2 FILLER_56_637 ();
 sg13g2_fill_1 FILLER_56_639 ();
 sg13g2_decap_8 FILLER_56_644 ();
 sg13g2_fill_1 FILLER_56_651 ();
 sg13g2_decap_4 FILLER_56_656 ();
 sg13g2_fill_2 FILLER_56_704 ();
 sg13g2_fill_1 FILLER_56_721 ();
 sg13g2_fill_1 FILLER_56_726 ();
 sg13g2_fill_1 FILLER_56_732 ();
 sg13g2_fill_1 FILLER_56_745 ();
 sg13g2_fill_1 FILLER_56_777 ();
 sg13g2_fill_1 FILLER_56_786 ();
 sg13g2_fill_2 FILLER_56_799 ();
 sg13g2_fill_1 FILLER_56_801 ();
 sg13g2_fill_1 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_862 ();
 sg13g2_fill_1 FILLER_56_864 ();
 sg13g2_fill_2 FILLER_56_869 ();
 sg13g2_fill_2 FILLER_56_877 ();
 sg13g2_fill_1 FILLER_56_879 ();
 sg13g2_decap_4 FILLER_56_885 ();
 sg13g2_fill_1 FILLER_56_889 ();
 sg13g2_fill_1 FILLER_56_894 ();
 sg13g2_decap_8 FILLER_56_900 ();
 sg13g2_fill_2 FILLER_56_916 ();
 sg13g2_fill_1 FILLER_56_922 ();
 sg13g2_fill_2 FILLER_56_951 ();
 sg13g2_fill_1 FILLER_56_961 ();
 sg13g2_decap_8 FILLER_56_966 ();
 sg13g2_decap_4 FILLER_56_973 ();
 sg13g2_fill_1 FILLER_56_977 ();
 sg13g2_fill_2 FILLER_56_983 ();
 sg13g2_fill_1 FILLER_56_998 ();
 sg13g2_fill_1 FILLER_56_1045 ();
 sg13g2_fill_2 FILLER_56_1055 ();
 sg13g2_fill_1 FILLER_56_1057 ();
 sg13g2_fill_1 FILLER_56_1090 ();
 sg13g2_fill_1 FILLER_56_1099 ();
 sg13g2_decap_4 FILLER_56_1107 ();
 sg13g2_decap_4 FILLER_56_1115 ();
 sg13g2_fill_2 FILLER_56_1119 ();
 sg13g2_fill_2 FILLER_56_1162 ();
 sg13g2_fill_1 FILLER_56_1164 ();
 sg13g2_fill_1 FILLER_56_1174 ();
 sg13g2_fill_2 FILLER_56_1227 ();
 sg13g2_fill_1 FILLER_56_1238 ();
 sg13g2_fill_1 FILLER_56_1247 ();
 sg13g2_fill_1 FILLER_56_1256 ();
 sg13g2_fill_1 FILLER_56_1262 ();
 sg13g2_fill_1 FILLER_56_1268 ();
 sg13g2_decap_8 FILLER_56_1273 ();
 sg13g2_decap_8 FILLER_56_1280 ();
 sg13g2_decap_8 FILLER_56_1287 ();
 sg13g2_decap_8 FILLER_56_1294 ();
 sg13g2_decap_8 FILLER_56_1301 ();
 sg13g2_decap_8 FILLER_56_1308 ();
 sg13g2_decap_8 FILLER_56_1315 ();
 sg13g2_decap_4 FILLER_56_1322 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_fill_2 FILLER_57_42 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_decap_4 FILLER_57_49 ();
 sg13g2_fill_2 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_87 ();
 sg13g2_fill_2 FILLER_57_105 ();
 sg13g2_fill_2 FILLER_57_126 ();
 sg13g2_fill_1 FILLER_57_128 ();
 sg13g2_decap_4 FILLER_57_172 ();
 sg13g2_decap_4 FILLER_57_180 ();
 sg13g2_fill_2 FILLER_57_184 ();
 sg13g2_fill_2 FILLER_57_190 ();
 sg13g2_fill_1 FILLER_57_192 ();
 sg13g2_fill_1 FILLER_57_257 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_fill_2 FILLER_57_272 ();
 sg13g2_fill_1 FILLER_57_282 ();
 sg13g2_fill_2 FILLER_57_288 ();
 sg13g2_fill_2 FILLER_57_294 ();
 sg13g2_fill_2 FILLER_57_325 ();
 sg13g2_fill_1 FILLER_57_327 ();
 sg13g2_fill_1 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_367 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_2 FILLER_57_403 ();
 sg13g2_fill_1 FILLER_57_413 ();
 sg13g2_fill_2 FILLER_57_418 ();
 sg13g2_fill_2 FILLER_57_446 ();
 sg13g2_fill_1 FILLER_57_448 ();
 sg13g2_fill_2 FILLER_57_484 ();
 sg13g2_fill_1 FILLER_57_490 ();
 sg13g2_fill_2 FILLER_57_499 ();
 sg13g2_decap_4 FILLER_57_514 ();
 sg13g2_fill_1 FILLER_57_523 ();
 sg13g2_fill_1 FILLER_57_539 ();
 sg13g2_decap_8 FILLER_57_544 ();
 sg13g2_fill_2 FILLER_57_551 ();
 sg13g2_fill_1 FILLER_57_553 ();
 sg13g2_decap_4 FILLER_57_558 ();
 sg13g2_fill_1 FILLER_57_562 ();
 sg13g2_fill_1 FILLER_57_567 ();
 sg13g2_fill_1 FILLER_57_572 ();
 sg13g2_fill_2 FILLER_57_599 ();
 sg13g2_fill_2 FILLER_57_605 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_2 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_676 ();
 sg13g2_fill_1 FILLER_57_690 ();
 sg13g2_fill_1 FILLER_57_836 ();
 sg13g2_fill_2 FILLER_57_883 ();
 sg13g2_fill_2 FILLER_57_906 ();
 sg13g2_fill_2 FILLER_57_928 ();
 sg13g2_decap_8 FILLER_57_1005 ();
 sg13g2_decap_4 FILLER_57_1012 ();
 sg13g2_fill_1 FILLER_57_1171 ();
 sg13g2_fill_1 FILLER_57_1202 ();
 sg13g2_fill_2 FILLER_57_1207 ();
 sg13g2_fill_1 FILLER_57_1217 ();
 sg13g2_fill_2 FILLER_57_1239 ();
 sg13g2_decap_8 FILLER_57_1288 ();
 sg13g2_decap_8 FILLER_57_1295 ();
 sg13g2_decap_8 FILLER_57_1302 ();
 sg13g2_decap_8 FILLER_57_1309 ();
 sg13g2_decap_8 FILLER_57_1316 ();
 sg13g2_fill_2 FILLER_57_1323 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_fill_2 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_37 ();
 sg13g2_fill_1 FILLER_58_82 ();
 sg13g2_fill_1 FILLER_58_145 ();
 sg13g2_fill_1 FILLER_58_185 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_1 FILLER_58_211 ();
 sg13g2_fill_1 FILLER_58_216 ();
 sg13g2_fill_1 FILLER_58_221 ();
 sg13g2_fill_1 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_246 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_decap_8 FILLER_58_278 ();
 sg13g2_decap_8 FILLER_58_285 ();
 sg13g2_fill_2 FILLER_58_292 ();
 sg13g2_fill_1 FILLER_58_294 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_fill_2 FILLER_58_329 ();
 sg13g2_fill_1 FILLER_58_331 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_2 FILLER_58_354 ();
 sg13g2_fill_1 FILLER_58_356 ();
 sg13g2_decap_4 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_413 ();
 sg13g2_fill_1 FILLER_58_415 ();
 sg13g2_fill_2 FILLER_58_450 ();
 sg13g2_fill_1 FILLER_58_468 ();
 sg13g2_fill_1 FILLER_58_473 ();
 sg13g2_fill_2 FILLER_58_478 ();
 sg13g2_fill_1 FILLER_58_480 ();
 sg13g2_fill_1 FILLER_58_486 ();
 sg13g2_fill_2 FILLER_58_513 ();
 sg13g2_fill_1 FILLER_58_515 ();
 sg13g2_fill_2 FILLER_58_519 ();
 sg13g2_fill_1 FILLER_58_521 ();
 sg13g2_fill_2 FILLER_58_533 ();
 sg13g2_fill_2 FILLER_58_574 ();
 sg13g2_fill_2 FILLER_58_605 ();
 sg13g2_fill_1 FILLER_58_607 ();
 sg13g2_fill_1 FILLER_58_625 ();
 sg13g2_decap_4 FILLER_58_635 ();
 sg13g2_fill_1 FILLER_58_639 ();
 sg13g2_fill_2 FILLER_58_680 ();
 sg13g2_fill_1 FILLER_58_694 ();
 sg13g2_fill_1 FILLER_58_707 ();
 sg13g2_decap_4 FILLER_58_717 ();
 sg13g2_fill_1 FILLER_58_734 ();
 sg13g2_fill_2 FILLER_58_739 ();
 sg13g2_fill_2 FILLER_58_752 ();
 sg13g2_decap_4 FILLER_58_758 ();
 sg13g2_fill_2 FILLER_58_774 ();
 sg13g2_fill_2 FILLER_58_797 ();
 sg13g2_fill_1 FILLER_58_841 ();
 sg13g2_decap_8 FILLER_58_858 ();
 sg13g2_decap_4 FILLER_58_865 ();
 sg13g2_fill_2 FILLER_58_874 ();
 sg13g2_fill_1 FILLER_58_891 ();
 sg13g2_fill_1 FILLER_58_902 ();
 sg13g2_fill_2 FILLER_58_947 ();
 sg13g2_fill_1 FILLER_58_996 ();
 sg13g2_decap_8 FILLER_58_1036 ();
 sg13g2_decap_4 FILLER_58_1043 ();
 sg13g2_fill_1 FILLER_58_1047 ();
 sg13g2_fill_1 FILLER_58_1060 ();
 sg13g2_fill_1 FILLER_58_1092 ();
 sg13g2_fill_1 FILLER_58_1097 ();
 sg13g2_fill_1 FILLER_58_1103 ();
 sg13g2_fill_1 FILLER_58_1108 ();
 sg13g2_fill_1 FILLER_58_1114 ();
 sg13g2_fill_2 FILLER_58_1147 ();
 sg13g2_decap_4 FILLER_58_1208 ();
 sg13g2_fill_1 FILLER_58_1212 ();
 sg13g2_fill_2 FILLER_58_1248 ();
 sg13g2_fill_1 FILLER_58_1254 ();
 sg13g2_decap_8 FILLER_58_1266 ();
 sg13g2_decap_8 FILLER_58_1273 ();
 sg13g2_decap_8 FILLER_58_1280 ();
 sg13g2_decap_8 FILLER_58_1287 ();
 sg13g2_decap_8 FILLER_58_1294 ();
 sg13g2_decap_8 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1308 ();
 sg13g2_decap_8 FILLER_58_1315 ();
 sg13g2_decap_4 FILLER_58_1322 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_4 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_50 ();
 sg13g2_decap_4 FILLER_59_62 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_97 ();
 sg13g2_fill_2 FILLER_59_111 ();
 sg13g2_fill_1 FILLER_59_125 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_141 ();
 sg13g2_fill_2 FILLER_59_155 ();
 sg13g2_fill_2 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_224 ();
 sg13g2_fill_2 FILLER_59_256 ();
 sg13g2_fill_1 FILLER_59_258 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_357 ();
 sg13g2_fill_1 FILLER_59_389 ();
 sg13g2_fill_2 FILLER_59_400 ();
 sg13g2_fill_1 FILLER_59_411 ();
 sg13g2_fill_2 FILLER_59_476 ();
 sg13g2_fill_1 FILLER_59_478 ();
 sg13g2_fill_1 FILLER_59_518 ();
 sg13g2_decap_8 FILLER_59_540 ();
 sg13g2_fill_2 FILLER_59_547 ();
 sg13g2_fill_1 FILLER_59_553 ();
 sg13g2_fill_1 FILLER_59_559 ();
 sg13g2_fill_1 FILLER_59_591 ();
 sg13g2_fill_1 FILLER_59_630 ();
 sg13g2_fill_1 FILLER_59_635 ();
 sg13g2_fill_1 FILLER_59_640 ();
 sg13g2_fill_1 FILLER_59_649 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_fill_2 FILLER_59_677 ();
 sg13g2_fill_1 FILLER_59_679 ();
 sg13g2_fill_1 FILLER_59_695 ();
 sg13g2_fill_2 FILLER_59_710 ();
 sg13g2_decap_4 FILLER_59_721 ();
 sg13g2_fill_2 FILLER_59_725 ();
 sg13g2_decap_4 FILLER_59_753 ();
 sg13g2_fill_1 FILLER_59_757 ();
 sg13g2_fill_2 FILLER_59_790 ();
 sg13g2_fill_1 FILLER_59_818 ();
 sg13g2_fill_2 FILLER_59_844 ();
 sg13g2_fill_1 FILLER_59_880 ();
 sg13g2_fill_1 FILLER_59_933 ();
 sg13g2_fill_2 FILLER_59_938 ();
 sg13g2_fill_2 FILLER_59_948 ();
 sg13g2_fill_1 FILLER_59_950 ();
 sg13g2_fill_2 FILLER_59_955 ();
 sg13g2_fill_1 FILLER_59_957 ();
 sg13g2_fill_2 FILLER_59_962 ();
 sg13g2_fill_1 FILLER_59_964 ();
 sg13g2_fill_2 FILLER_59_974 ();
 sg13g2_fill_1 FILLER_59_976 ();
 sg13g2_fill_2 FILLER_59_995 ();
 sg13g2_fill_1 FILLER_59_1007 ();
 sg13g2_decap_4 FILLER_59_1027 ();
 sg13g2_fill_2 FILLER_59_1061 ();
 sg13g2_fill_2 FILLER_59_1094 ();
 sg13g2_fill_1 FILLER_59_1126 ();
 sg13g2_fill_1 FILLER_59_1131 ();
 sg13g2_fill_1 FILLER_59_1137 ();
 sg13g2_fill_2 FILLER_59_1146 ();
 sg13g2_fill_1 FILLER_59_1148 ();
 sg13g2_fill_2 FILLER_59_1156 ();
 sg13g2_fill_2 FILLER_59_1162 ();
 sg13g2_fill_1 FILLER_59_1195 ();
 sg13g2_fill_2 FILLER_59_1227 ();
 sg13g2_fill_1 FILLER_59_1237 ();
 sg13g2_fill_1 FILLER_59_1247 ();
 sg13g2_fill_1 FILLER_59_1274 ();
 sg13g2_decap_8 FILLER_59_1279 ();
 sg13g2_decap_8 FILLER_59_1286 ();
 sg13g2_decap_8 FILLER_59_1293 ();
 sg13g2_decap_8 FILLER_59_1300 ();
 sg13g2_decap_8 FILLER_59_1307 ();
 sg13g2_decap_8 FILLER_59_1314 ();
 sg13g2_decap_4 FILLER_59_1321 ();
 sg13g2_fill_1 FILLER_59_1325 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_4 FILLER_60_35 ();
 sg13g2_fill_1 FILLER_60_72 ();
 sg13g2_fill_1 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_197 ();
 sg13g2_decap_4 FILLER_60_202 ();
 sg13g2_fill_1 FILLER_60_206 ();
 sg13g2_fill_2 FILLER_60_211 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_2 FILLER_60_223 ();
 sg13g2_fill_2 FILLER_60_233 ();
 sg13g2_fill_2 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_241 ();
 sg13g2_fill_1 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_298 ();
 sg13g2_fill_2 FILLER_60_303 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_fill_1 FILLER_60_345 ();
 sg13g2_fill_1 FILLER_60_372 ();
 sg13g2_fill_2 FILLER_60_378 ();
 sg13g2_fill_2 FILLER_60_390 ();
 sg13g2_fill_1 FILLER_60_392 ();
 sg13g2_fill_2 FILLER_60_510 ();
 sg13g2_fill_1 FILLER_60_512 ();
 sg13g2_decap_4 FILLER_60_533 ();
 sg13g2_fill_2 FILLER_60_537 ();
 sg13g2_fill_1 FILLER_60_547 ();
 sg13g2_fill_2 FILLER_60_566 ();
 sg13g2_fill_2 FILLER_60_573 ();
 sg13g2_fill_1 FILLER_60_604 ();
 sg13g2_fill_2 FILLER_60_631 ();
 sg13g2_fill_2 FILLER_60_786 ();
 sg13g2_fill_1 FILLER_60_860 ();
 sg13g2_fill_1 FILLER_60_871 ();
 sg13g2_fill_1 FILLER_60_913 ();
 sg13g2_fill_1 FILLER_60_918 ();
 sg13g2_fill_1 FILLER_60_931 ();
 sg13g2_fill_1 FILLER_60_1004 ();
 sg13g2_fill_1 FILLER_60_1041 ();
 sg13g2_fill_1 FILLER_60_1051 ();
 sg13g2_fill_1 FILLER_60_1104 ();
 sg13g2_fill_1 FILLER_60_1113 ();
 sg13g2_fill_1 FILLER_60_1119 ();
 sg13g2_fill_1 FILLER_60_1146 ();
 sg13g2_fill_1 FILLER_60_1152 ();
 sg13g2_fill_1 FILLER_60_1158 ();
 sg13g2_fill_1 FILLER_60_1163 ();
 sg13g2_fill_2 FILLER_60_1168 ();
 sg13g2_fill_2 FILLER_60_1174 ();
 sg13g2_fill_2 FILLER_60_1180 ();
 sg13g2_fill_2 FILLER_60_1187 ();
 sg13g2_fill_2 FILLER_60_1193 ();
 sg13g2_fill_2 FILLER_60_1204 ();
 sg13g2_fill_1 FILLER_60_1206 ();
 sg13g2_fill_1 FILLER_60_1229 ();
 sg13g2_fill_1 FILLER_60_1254 ();
 sg13g2_decap_8 FILLER_60_1286 ();
 sg13g2_decap_8 FILLER_60_1293 ();
 sg13g2_decap_8 FILLER_60_1300 ();
 sg13g2_decap_8 FILLER_60_1307 ();
 sg13g2_decap_8 FILLER_60_1314 ();
 sg13g2_decap_4 FILLER_60_1321 ();
 sg13g2_fill_1 FILLER_60_1325 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_fill_1 FILLER_61_78 ();
 sg13g2_fill_2 FILLER_61_84 ();
 sg13g2_fill_1 FILLER_61_94 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_2 FILLER_61_150 ();
 sg13g2_fill_2 FILLER_61_220 ();
 sg13g2_fill_1 FILLER_61_253 ();
 sg13g2_fill_2 FILLER_61_274 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_fill_1 FILLER_61_323 ();
 sg13g2_fill_2 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_339 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_fill_2 FILLER_61_353 ();
 sg13g2_fill_1 FILLER_61_355 ();
 sg13g2_fill_2 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_362 ();
 sg13g2_fill_1 FILLER_61_417 ();
 sg13g2_fill_2 FILLER_61_444 ();
 sg13g2_fill_1 FILLER_61_446 ();
 sg13g2_fill_2 FILLER_61_477 ();
 sg13g2_fill_2 FILLER_61_483 ();
 sg13g2_fill_1 FILLER_61_490 ();
 sg13g2_fill_1 FILLER_61_495 ();
 sg13g2_fill_2 FILLER_61_504 ();
 sg13g2_fill_1 FILLER_61_506 ();
 sg13g2_fill_2 FILLER_61_545 ();
 sg13g2_fill_1 FILLER_61_552 ();
 sg13g2_fill_2 FILLER_61_610 ();
 sg13g2_fill_2 FILLER_61_616 ();
 sg13g2_fill_1 FILLER_61_618 ();
 sg13g2_fill_1 FILLER_61_645 ();
 sg13g2_fill_2 FILLER_61_654 ();
 sg13g2_fill_1 FILLER_61_656 ();
 sg13g2_fill_2 FILLER_61_665 ();
 sg13g2_fill_1 FILLER_61_667 ();
 sg13g2_fill_2 FILLER_61_672 ();
 sg13g2_fill_1 FILLER_61_674 ();
 sg13g2_decap_8 FILLER_61_679 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_fill_1 FILLER_61_691 ();
 sg13g2_fill_2 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_702 ();
 sg13g2_fill_1 FILLER_61_707 ();
 sg13g2_fill_1 FILLER_61_712 ();
 sg13g2_fill_1 FILLER_61_717 ();
 sg13g2_fill_1 FILLER_61_726 ();
 sg13g2_fill_1 FILLER_61_735 ();
 sg13g2_fill_2 FILLER_61_744 ();
 sg13g2_fill_1 FILLER_61_751 ();
 sg13g2_fill_2 FILLER_61_782 ();
 sg13g2_fill_2 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_fill_2 FILLER_61_826 ();
 sg13g2_fill_1 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_842 ();
 sg13g2_fill_2 FILLER_61_849 ();
 sg13g2_fill_1 FILLER_61_851 ();
 sg13g2_fill_2 FILLER_61_865 ();
 sg13g2_fill_2 FILLER_61_875 ();
 sg13g2_fill_1 FILLER_61_901 ();
 sg13g2_fill_1 FILLER_61_907 ();
 sg13g2_decap_4 FILLER_61_955 ();
 sg13g2_fill_1 FILLER_61_963 ();
 sg13g2_fill_1 FILLER_61_968 ();
 sg13g2_fill_1 FILLER_61_974 ();
 sg13g2_fill_1 FILLER_61_979 ();
 sg13g2_fill_1 FILLER_61_984 ();
 sg13g2_fill_1 FILLER_61_989 ();
 sg13g2_fill_1 FILLER_61_995 ();
 sg13g2_fill_1 FILLER_61_1026 ();
 sg13g2_fill_2 FILLER_61_1031 ();
 sg13g2_fill_2 FILLER_61_1070 ();
 sg13g2_fill_2 FILLER_61_1100 ();
 sg13g2_fill_2 FILLER_61_1144 ();
 sg13g2_fill_1 FILLER_61_1155 ();
 sg13g2_fill_2 FILLER_61_1190 ();
 sg13g2_fill_2 FILLER_61_1218 ();
 sg13g2_fill_2 FILLER_61_1232 ();
 sg13g2_fill_1 FILLER_61_1234 ();
 sg13g2_fill_2 FILLER_61_1244 ();
 sg13g2_decap_4 FILLER_61_1250 ();
 sg13g2_fill_1 FILLER_61_1254 ();
 sg13g2_fill_2 FILLER_61_1263 ();
 sg13g2_fill_1 FILLER_61_1270 ();
 sg13g2_decap_8 FILLER_61_1275 ();
 sg13g2_fill_1 FILLER_61_1282 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_8 FILLER_61_1294 ();
 sg13g2_decap_8 FILLER_61_1301 ();
 sg13g2_decap_8 FILLER_61_1308 ();
 sg13g2_decap_8 FILLER_61_1315 ();
 sg13g2_decap_4 FILLER_61_1322 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_4 FILLER_62_21 ();
 sg13g2_fill_2 FILLER_62_55 ();
 sg13g2_fill_1 FILLER_62_79 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_fill_1 FILLER_62_95 ();
 sg13g2_fill_1 FILLER_62_141 ();
 sg13g2_fill_2 FILLER_62_146 ();
 sg13g2_fill_2 FILLER_62_163 ();
 sg13g2_fill_2 FILLER_62_172 ();
 sg13g2_fill_1 FILLER_62_182 ();
 sg13g2_fill_1 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_259 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_1 FILLER_62_270 ();
 sg13g2_fill_1 FILLER_62_276 ();
 sg13g2_fill_1 FILLER_62_297 ();
 sg13g2_decap_4 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_310 ();
 sg13g2_fill_1 FILLER_62_312 ();
 sg13g2_fill_1 FILLER_62_359 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_1 FILLER_62_427 ();
 sg13g2_fill_2 FILLER_62_582 ();
 sg13g2_fill_2 FILLER_62_588 ();
 sg13g2_fill_1 FILLER_62_590 ();
 sg13g2_decap_4 FILLER_62_595 ();
 sg13g2_fill_1 FILLER_62_599 ();
 sg13g2_fill_2 FILLER_62_605 ();
 sg13g2_decap_4 FILLER_62_615 ();
 sg13g2_fill_2 FILLER_62_619 ();
 sg13g2_fill_2 FILLER_62_625 ();
 sg13g2_fill_1 FILLER_62_627 ();
 sg13g2_fill_1 FILLER_62_753 ();
 sg13g2_fill_2 FILLER_62_768 ();
 sg13g2_fill_2 FILLER_62_775 ();
 sg13g2_fill_2 FILLER_62_841 ();
 sg13g2_fill_1 FILLER_62_847 ();
 sg13g2_fill_2 FILLER_62_853 ();
 sg13g2_fill_2 FILLER_62_864 ();
 sg13g2_fill_2 FILLER_62_915 ();
 sg13g2_fill_1 FILLER_62_917 ();
 sg13g2_fill_2 FILLER_62_922 ();
 sg13g2_fill_1 FILLER_62_929 ();
 sg13g2_fill_1 FILLER_62_934 ();
 sg13g2_fill_2 FILLER_62_943 ();
 sg13g2_decap_4 FILLER_62_997 ();
 sg13g2_fill_2 FILLER_62_1001 ();
 sg13g2_decap_4 FILLER_62_1007 ();
 sg13g2_fill_1 FILLER_62_1011 ();
 sg13g2_fill_1 FILLER_62_1064 ();
 sg13g2_fill_1 FILLER_62_1073 ();
 sg13g2_fill_1 FILLER_62_1079 ();
 sg13g2_fill_1 FILLER_62_1085 ();
 sg13g2_fill_1 FILLER_62_1094 ();
 sg13g2_fill_1 FILLER_62_1103 ();
 sg13g2_fill_2 FILLER_62_1161 ();
 sg13g2_fill_1 FILLER_62_1190 ();
 sg13g2_fill_2 FILLER_62_1204 ();
 sg13g2_fill_2 FILLER_62_1219 ();
 sg13g2_fill_2 FILLER_62_1226 ();
 sg13g2_fill_1 FILLER_62_1228 ();
 sg13g2_fill_2 FILLER_62_1233 ();
 sg13g2_fill_1 FILLER_62_1235 ();
 sg13g2_decap_8 FILLER_62_1288 ();
 sg13g2_decap_8 FILLER_62_1295 ();
 sg13g2_decap_8 FILLER_62_1302 ();
 sg13g2_decap_8 FILLER_62_1309 ();
 sg13g2_decap_8 FILLER_62_1316 ();
 sg13g2_fill_2 FILLER_62_1323 ();
 sg13g2_fill_1 FILLER_62_1325 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_28 ();
 sg13g2_fill_1 FILLER_63_30 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_71 ();
 sg13g2_fill_2 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_119 ();
 sg13g2_fill_1 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_228 ();
 sg13g2_fill_1 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_239 ();
 sg13g2_fill_1 FILLER_63_245 ();
 sg13g2_fill_2 FILLER_63_299 ();
 sg13g2_fill_1 FILLER_63_301 ();
 sg13g2_fill_2 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_339 ();
 sg13g2_fill_2 FILLER_63_346 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_fill_1 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_363 ();
 sg13g2_fill_1 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_63_396 ();
 sg13g2_fill_1 FILLER_63_400 ();
 sg13g2_fill_1 FILLER_63_411 ();
 sg13g2_fill_1 FILLER_63_442 ();
 sg13g2_fill_1 FILLER_63_469 ();
 sg13g2_fill_1 FILLER_63_514 ();
 sg13g2_fill_2 FILLER_63_519 ();
 sg13g2_fill_1 FILLER_63_521 ();
 sg13g2_fill_2 FILLER_63_526 ();
 sg13g2_fill_1 FILLER_63_528 ();
 sg13g2_fill_2 FILLER_63_557 ();
 sg13g2_fill_2 FILLER_63_567 ();
 sg13g2_fill_2 FILLER_63_603 ();
 sg13g2_fill_1 FILLER_63_605 ();
 sg13g2_fill_2 FILLER_63_632 ();
 sg13g2_decap_4 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_655 ();
 sg13g2_fill_1 FILLER_63_657 ();
 sg13g2_fill_1 FILLER_63_668 ();
 sg13g2_fill_2 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_683 ();
 sg13g2_fill_1 FILLER_63_685 ();
 sg13g2_decap_4 FILLER_63_695 ();
 sg13g2_fill_1 FILLER_63_699 ();
 sg13g2_decap_4 FILLER_63_704 ();
 sg13g2_fill_1 FILLER_63_708 ();
 sg13g2_fill_1 FILLER_63_713 ();
 sg13g2_fill_2 FILLER_63_726 ();
 sg13g2_fill_1 FILLER_63_728 ();
 sg13g2_fill_2 FILLER_63_755 ();
 sg13g2_fill_1 FILLER_63_761 ();
 sg13g2_fill_2 FILLER_63_822 ();
 sg13g2_fill_1 FILLER_63_824 ();
 sg13g2_decap_4 FILLER_63_851 ();
 sg13g2_fill_2 FILLER_63_980 ();
 sg13g2_fill_1 FILLER_63_982 ();
 sg13g2_fill_2 FILLER_63_986 ();
 sg13g2_fill_1 FILLER_63_988 ();
 sg13g2_fill_2 FILLER_63_1032 ();
 sg13g2_fill_2 FILLER_63_1052 ();
 sg13g2_fill_1 FILLER_63_1095 ();
 sg13g2_fill_1 FILLER_63_1109 ();
 sg13g2_fill_1 FILLER_63_1185 ();
 sg13g2_fill_1 FILLER_63_1194 ();
 sg13g2_fill_2 FILLER_63_1200 ();
 sg13g2_fill_2 FILLER_63_1206 ();
 sg13g2_fill_2 FILLER_63_1212 ();
 sg13g2_fill_1 FILLER_63_1214 ();
 sg13g2_fill_2 FILLER_63_1242 ();
 sg13g2_fill_1 FILLER_63_1244 ();
 sg13g2_fill_2 FILLER_63_1249 ();
 sg13g2_fill_1 FILLER_63_1251 ();
 sg13g2_fill_2 FILLER_63_1257 ();
 sg13g2_fill_1 FILLER_63_1259 ();
 sg13g2_fill_2 FILLER_63_1264 ();
 sg13g2_decap_8 FILLER_63_1278 ();
 sg13g2_decap_8 FILLER_63_1285 ();
 sg13g2_decap_8 FILLER_63_1292 ();
 sg13g2_decap_8 FILLER_63_1299 ();
 sg13g2_decap_8 FILLER_63_1306 ();
 sg13g2_decap_8 FILLER_63_1313 ();
 sg13g2_decap_4 FILLER_63_1320 ();
 sg13g2_fill_2 FILLER_63_1324 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_56 ();
 sg13g2_fill_1 FILLER_64_65 ();
 sg13g2_fill_1 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_146 ();
 sg13g2_fill_1 FILLER_64_196 ();
 sg13g2_fill_2 FILLER_64_223 ();
 sg13g2_fill_1 FILLER_64_230 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_263 ();
 sg13g2_decap_4 FILLER_64_270 ();
 sg13g2_fill_2 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_286 ();
 sg13g2_fill_2 FILLER_64_292 ();
 sg13g2_decap_4 FILLER_64_298 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_457 ();
 sg13g2_fill_2 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_497 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_fill_2 FILLER_64_526 ();
 sg13g2_decap_4 FILLER_64_536 ();
 sg13g2_fill_1 FILLER_64_606 ();
 sg13g2_fill_2 FILLER_64_618 ();
 sg13g2_fill_1 FILLER_64_649 ();
 sg13g2_fill_1 FILLER_64_656 ();
 sg13g2_fill_1 FILLER_64_720 ();
 sg13g2_fill_1 FILLER_64_777 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_4 FILLER_64_828 ();
 sg13g2_fill_2 FILLER_64_832 ();
 sg13g2_decap_4 FILLER_64_838 ();
 sg13g2_fill_1 FILLER_64_854 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_1 FILLER_64_867 ();
 sg13g2_fill_1 FILLER_64_897 ();
 sg13g2_fill_1 FILLER_64_903 ();
 sg13g2_fill_2 FILLER_64_923 ();
 sg13g2_fill_1 FILLER_64_933 ();
 sg13g2_fill_1 FILLER_64_942 ();
 sg13g2_fill_1 FILLER_64_989 ();
 sg13g2_fill_1 FILLER_64_1052 ();
 sg13g2_fill_1 FILLER_64_1069 ();
 sg13g2_fill_1 FILLER_64_1074 ();
 sg13g2_decap_4 FILLER_64_1079 ();
 sg13g2_fill_2 FILLER_64_1083 ();
 sg13g2_fill_2 FILLER_64_1089 ();
 sg13g2_fill_1 FILLER_64_1095 ();
 sg13g2_fill_1 FILLER_64_1126 ();
 sg13g2_fill_1 FILLER_64_1132 ();
 sg13g2_fill_1 FILLER_64_1149 ();
 sg13g2_fill_1 FILLER_64_1221 ();
 sg13g2_decap_8 FILLER_64_1286 ();
 sg13g2_decap_8 FILLER_64_1293 ();
 sg13g2_decap_8 FILLER_64_1300 ();
 sg13g2_decap_8 FILLER_64_1307 ();
 sg13g2_decap_8 FILLER_64_1314 ();
 sg13g2_decap_4 FILLER_64_1321 ();
 sg13g2_fill_1 FILLER_64_1325 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_fill_2 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_37 ();
 sg13g2_fill_2 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_48 ();
 sg13g2_fill_1 FILLER_65_96 ();
 sg13g2_fill_2 FILLER_65_101 ();
 sg13g2_fill_1 FILLER_65_108 ();
 sg13g2_fill_2 FILLER_65_113 ();
 sg13g2_fill_2 FILLER_65_228 ();
 sg13g2_decap_4 FILLER_65_273 ();
 sg13g2_fill_1 FILLER_65_277 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_fill_1 FILLER_65_300 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_400 ();
 sg13g2_fill_1 FILLER_65_420 ();
 sg13g2_fill_2 FILLER_65_496 ();
 sg13g2_fill_1 FILLER_65_503 ();
 sg13g2_fill_1 FILLER_65_542 ();
 sg13g2_fill_2 FILLER_65_548 ();
 sg13g2_fill_1 FILLER_65_550 ();
 sg13g2_fill_2 FILLER_65_586 ();
 sg13g2_fill_2 FILLER_65_638 ();
 sg13g2_fill_1 FILLER_65_666 ();
 sg13g2_fill_2 FILLER_65_670 ();
 sg13g2_fill_1 FILLER_65_676 ();
 sg13g2_fill_2 FILLER_65_681 ();
 sg13g2_decap_4 FILLER_65_688 ();
 sg13g2_fill_2 FILLER_65_692 ();
 sg13g2_decap_8 FILLER_65_702 ();
 sg13g2_fill_1 FILLER_65_709 ();
 sg13g2_fill_1 FILLER_65_736 ();
 sg13g2_fill_1 FILLER_65_741 ();
 sg13g2_fill_1 FILLER_65_747 ();
 sg13g2_fill_1 FILLER_65_755 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_fill_1 FILLER_65_788 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_798 ();
 sg13g2_fill_2 FILLER_65_803 ();
 sg13g2_fill_1 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_861 ();
 sg13g2_fill_2 FILLER_65_893 ();
 sg13g2_fill_2 FILLER_65_908 ();
 sg13g2_fill_1 FILLER_65_956 ();
 sg13g2_fill_1 FILLER_65_998 ();
 sg13g2_fill_2 FILLER_65_1009 ();
 sg13g2_fill_1 FILLER_65_1026 ();
 sg13g2_fill_2 FILLER_65_1031 ();
 sg13g2_fill_2 FILLER_65_1041 ();
 sg13g2_fill_1 FILLER_65_1061 ();
 sg13g2_fill_1 FILLER_65_1190 ();
 sg13g2_fill_1 FILLER_65_1199 ();
 sg13g2_fill_1 FILLER_65_1213 ();
 sg13g2_fill_1 FILLER_65_1249 ();
 sg13g2_fill_1 FILLER_65_1258 ();
 sg13g2_decap_8 FILLER_65_1285 ();
 sg13g2_decap_8 FILLER_65_1292 ();
 sg13g2_decap_8 FILLER_65_1299 ();
 sg13g2_decap_8 FILLER_65_1306 ();
 sg13g2_decap_8 FILLER_65_1313 ();
 sg13g2_decap_4 FILLER_65_1320 ();
 sg13g2_fill_2 FILLER_65_1324 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_4 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_41 ();
 sg13g2_fill_1 FILLER_66_50 ();
 sg13g2_fill_2 FILLER_66_59 ();
 sg13g2_fill_1 FILLER_66_74 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_1 FILLER_66_227 ();
 sg13g2_fill_2 FILLER_66_237 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_1 FILLER_66_336 ();
 sg13g2_fill_1 FILLER_66_380 ();
 sg13g2_fill_1 FILLER_66_413 ();
 sg13g2_fill_1 FILLER_66_418 ();
 sg13g2_fill_2 FILLER_66_464 ();
 sg13g2_fill_1 FILLER_66_469 ();
 sg13g2_fill_2 FILLER_66_475 ();
 sg13g2_fill_2 FILLER_66_498 ();
 sg13g2_fill_1 FILLER_66_500 ();
 sg13g2_fill_2 FILLER_66_527 ();
 sg13g2_fill_1 FILLER_66_529 ();
 sg13g2_fill_2 FILLER_66_538 ();
 sg13g2_fill_1 FILLER_66_569 ();
 sg13g2_fill_2 FILLER_66_607 ();
 sg13g2_fill_2 FILLER_66_613 ();
 sg13g2_fill_1 FILLER_66_615 ();
 sg13g2_fill_1 FILLER_66_642 ();
 sg13g2_fill_2 FILLER_66_647 ();
 sg13g2_fill_1 FILLER_66_649 ();
 sg13g2_fill_1 FILLER_66_657 ();
 sg13g2_fill_1 FILLER_66_682 ();
 sg13g2_fill_1 FILLER_66_690 ();
 sg13g2_fill_1 FILLER_66_695 ();
 sg13g2_fill_1 FILLER_66_706 ();
 sg13g2_fill_1 FILLER_66_712 ();
 sg13g2_fill_2 FILLER_66_724 ();
 sg13g2_fill_1 FILLER_66_726 ();
 sg13g2_fill_2 FILLER_66_731 ();
 sg13g2_fill_1 FILLER_66_749 ();
 sg13g2_fill_1 FILLER_66_754 ();
 sg13g2_decap_8 FILLER_66_759 ();
 sg13g2_fill_2 FILLER_66_766 ();
 sg13g2_fill_2 FILLER_66_772 ();
 sg13g2_fill_2 FILLER_66_782 ();
 sg13g2_fill_1 FILLER_66_818 ();
 sg13g2_fill_1 FILLER_66_875 ();
 sg13g2_fill_1 FILLER_66_902 ();
 sg13g2_fill_2 FILLER_66_937 ();
 sg13g2_fill_1 FILLER_66_972 ();
 sg13g2_fill_1 FILLER_66_1019 ();
 sg13g2_fill_2 FILLER_66_1024 ();
 sg13g2_fill_1 FILLER_66_1031 ();
 sg13g2_fill_1 FILLER_66_1036 ();
 sg13g2_fill_1 FILLER_66_1041 ();
 sg13g2_fill_1 FILLER_66_1060 ();
 sg13g2_fill_1 FILLER_66_1091 ();
 sg13g2_fill_1 FILLER_66_1113 ();
 sg13g2_fill_2 FILLER_66_1132 ();
 sg13g2_fill_1 FILLER_66_1146 ();
 sg13g2_fill_1 FILLER_66_1159 ();
 sg13g2_fill_2 FILLER_66_1169 ();
 sg13g2_fill_1 FILLER_66_1201 ();
 sg13g2_fill_1 FILLER_66_1273 ();
 sg13g2_fill_2 FILLER_66_1278 ();
 sg13g2_decap_8 FILLER_66_1288 ();
 sg13g2_decap_8 FILLER_66_1295 ();
 sg13g2_decap_8 FILLER_66_1302 ();
 sg13g2_decap_8 FILLER_66_1309 ();
 sg13g2_decap_8 FILLER_66_1316 ();
 sg13g2_fill_2 FILLER_66_1323 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_23 ();
 sg13g2_fill_1 FILLER_67_50 ();
 sg13g2_fill_1 FILLER_67_68 ();
 sg13g2_fill_2 FILLER_67_79 ();
 sg13g2_fill_2 FILLER_67_150 ();
 sg13g2_fill_2 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_281 ();
 sg13g2_fill_1 FILLER_67_295 ();
 sg13g2_fill_2 FILLER_67_307 ();
 sg13g2_fill_2 FILLER_67_361 ();
 sg13g2_fill_2 FILLER_67_367 ();
 sg13g2_fill_1 FILLER_67_375 ();
 sg13g2_fill_1 FILLER_67_380 ();
 sg13g2_fill_1 FILLER_67_387 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_1 FILLER_67_420 ();
 sg13g2_fill_1 FILLER_67_432 ();
 sg13g2_fill_1 FILLER_67_437 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_501 ();
 sg13g2_fill_2 FILLER_67_549 ();
 sg13g2_fill_2 FILLER_67_555 ();
 sg13g2_fill_1 FILLER_67_583 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_fill_1 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_600 ();
 sg13g2_fill_1 FILLER_67_607 ();
 sg13g2_fill_2 FILLER_67_612 ();
 sg13g2_fill_2 FILLER_67_619 ();
 sg13g2_fill_1 FILLER_67_621 ();
 sg13g2_fill_1 FILLER_67_673 ();
 sg13g2_fill_1 FILLER_67_695 ();
 sg13g2_decap_4 FILLER_67_720 ();
 sg13g2_fill_1 FILLER_67_743 ();
 sg13g2_fill_1 FILLER_67_749 ();
 sg13g2_fill_1 FILLER_67_759 ();
 sg13g2_fill_1 FILLER_67_769 ();
 sg13g2_fill_1 FILLER_67_775 ();
 sg13g2_fill_1 FILLER_67_781 ();
 sg13g2_fill_1 FILLER_67_791 ();
 sg13g2_fill_1 FILLER_67_797 ();
 sg13g2_fill_1 FILLER_67_811 ();
 sg13g2_fill_1 FILLER_67_816 ();
 sg13g2_fill_2 FILLER_67_847 ();
 sg13g2_fill_2 FILLER_67_854 ();
 sg13g2_fill_1 FILLER_67_861 ();
 sg13g2_fill_1 FILLER_67_867 ();
 sg13g2_fill_1 FILLER_67_874 ();
 sg13g2_fill_1 FILLER_67_879 ();
 sg13g2_fill_1 FILLER_67_884 ();
 sg13g2_fill_2 FILLER_67_898 ();
 sg13g2_fill_2 FILLER_67_904 ();
 sg13g2_fill_2 FILLER_67_919 ();
 sg13g2_fill_2 FILLER_67_1134 ();
 sg13g2_fill_2 FILLER_67_1178 ();
 sg13g2_fill_1 FILLER_67_1196 ();
 sg13g2_fill_1 FILLER_67_1209 ();
 sg13g2_fill_1 FILLER_67_1222 ();
 sg13g2_fill_2 FILLER_67_1227 ();
 sg13g2_fill_2 FILLER_67_1233 ();
 sg13g2_fill_1 FILLER_67_1240 ();
 sg13g2_fill_2 FILLER_67_1249 ();
 sg13g2_fill_1 FILLER_67_1273 ();
 sg13g2_fill_1 FILLER_67_1278 ();
 sg13g2_fill_1 FILLER_67_1283 ();
 sg13g2_decap_8 FILLER_67_1294 ();
 sg13g2_decap_8 FILLER_67_1301 ();
 sg13g2_decap_8 FILLER_67_1308 ();
 sg13g2_decap_8 FILLER_67_1315 ();
 sg13g2_decap_4 FILLER_67_1322 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_fill_1 FILLER_68_35 ();
 sg13g2_decap_4 FILLER_68_40 ();
 sg13g2_fill_2 FILLER_68_44 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_1 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_233 ();
 sg13g2_fill_1 FILLER_68_335 ();
 sg13g2_fill_1 FILLER_68_450 ();
 sg13g2_fill_1 FILLER_68_454 ();
 sg13g2_fill_1 FILLER_68_465 ();
 sg13g2_fill_1 FILLER_68_470 ();
 sg13g2_fill_1 FILLER_68_476 ();
 sg13g2_fill_1 FILLER_68_503 ();
 sg13g2_fill_2 FILLER_68_508 ();
 sg13g2_decap_4 FILLER_68_515 ();
 sg13g2_decap_4 FILLER_68_523 ();
 sg13g2_fill_2 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_571 ();
 sg13g2_decap_8 FILLER_68_650 ();
 sg13g2_decap_4 FILLER_68_657 ();
 sg13g2_decap_8 FILLER_68_669 ();
 sg13g2_fill_2 FILLER_68_680 ();
 sg13g2_fill_1 FILLER_68_732 ();
 sg13g2_fill_1 FILLER_68_764 ();
 sg13g2_fill_1 FILLER_68_787 ();
 sg13g2_fill_2 FILLER_68_796 ();
 sg13g2_fill_1 FILLER_68_798 ();
 sg13g2_fill_2 FILLER_68_817 ();
 sg13g2_fill_1 FILLER_68_837 ();
 sg13g2_fill_2 FILLER_68_852 ();
 sg13g2_fill_2 FILLER_68_901 ();
 sg13g2_fill_2 FILLER_68_916 ();
 sg13g2_fill_2 FILLER_68_945 ();
 sg13g2_fill_2 FILLER_68_960 ();
 sg13g2_fill_1 FILLER_68_972 ();
 sg13g2_fill_2 FILLER_68_982 ();
 sg13g2_fill_1 FILLER_68_989 ();
 sg13g2_fill_1 FILLER_68_1017 ();
 sg13g2_fill_1 FILLER_68_1031 ();
 sg13g2_fill_2 FILLER_68_1066 ();
 sg13g2_fill_2 FILLER_68_1087 ();
 sg13g2_fill_2 FILLER_68_1105 ();
 sg13g2_fill_1 FILLER_68_1111 ();
 sg13g2_fill_1 FILLER_68_1159 ();
 sg13g2_fill_2 FILLER_68_1173 ();
 sg13g2_fill_2 FILLER_68_1194 ();
 sg13g2_fill_2 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1289 ();
 sg13g2_decap_8 FILLER_68_1296 ();
 sg13g2_decap_8 FILLER_68_1303 ();
 sg13g2_decap_8 FILLER_68_1310 ();
 sg13g2_decap_8 FILLER_68_1317 ();
 sg13g2_fill_2 FILLER_68_1324 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_4 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_25 ();
 sg13g2_fill_1 FILLER_69_57 ();
 sg13g2_fill_2 FILLER_69_89 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_1 FILLER_69_125 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_fill_1 FILLER_69_162 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_fill_2 FILLER_69_222 ();
 sg13g2_fill_2 FILLER_69_270 ();
 sg13g2_fill_2 FILLER_69_276 ();
 sg13g2_decap_4 FILLER_69_311 ();
 sg13g2_fill_1 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_346 ();
 sg13g2_fill_2 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_379 ();
 sg13g2_fill_2 FILLER_69_389 ();
 sg13g2_fill_1 FILLER_69_434 ();
 sg13g2_fill_2 FILLER_69_462 ();
 sg13g2_fill_1 FILLER_69_499 ();
 sg13g2_fill_1 FILLER_69_525 ();
 sg13g2_fill_2 FILLER_69_541 ();
 sg13g2_fill_1 FILLER_69_543 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_fill_1 FILLER_69_554 ();
 sg13g2_fill_1 FILLER_69_560 ();
 sg13g2_fill_1 FILLER_69_599 ();
 sg13g2_decap_4 FILLER_69_619 ();
 sg13g2_fill_1 FILLER_69_623 ();
 sg13g2_fill_2 FILLER_69_629 ();
 sg13g2_decap_8 FILLER_69_646 ();
 sg13g2_fill_2 FILLER_69_653 ();
 sg13g2_fill_1 FILLER_69_655 ();
 sg13g2_fill_2 FILLER_69_696 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_decap_4 FILLER_69_719 ();
 sg13g2_fill_2 FILLER_69_739 ();
 sg13g2_decap_4 FILLER_69_753 ();
 sg13g2_fill_1 FILLER_69_761 ();
 sg13g2_fill_1 FILLER_69_767 ();
 sg13g2_fill_2 FILLER_69_772 ();
 sg13g2_fill_2 FILLER_69_779 ();
 sg13g2_decap_4 FILLER_69_856 ();
 sg13g2_fill_1 FILLER_69_874 ();
 sg13g2_fill_2 FILLER_69_888 ();
 sg13g2_fill_2 FILLER_69_920 ();
 sg13g2_fill_2 FILLER_69_1000 ();
 sg13g2_fill_1 FILLER_69_1041 ();
 sg13g2_fill_2 FILLER_69_1047 ();
 sg13g2_fill_1 FILLER_69_1049 ();
 sg13g2_fill_2 FILLER_69_1103 ();
 sg13g2_fill_1 FILLER_69_1105 ();
 sg13g2_fill_2 FILLER_69_1233 ();
 sg13g2_fill_1 FILLER_69_1251 ();
 sg13g2_fill_2 FILLER_69_1270 ();
 sg13g2_fill_1 FILLER_69_1272 ();
 sg13g2_decap_4 FILLER_69_1277 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_8 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_69_1318 ();
 sg13g2_fill_1 FILLER_69_1325 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_4 FILLER_70_28 ();
 sg13g2_fill_2 FILLER_70_32 ();
 sg13g2_fill_1 FILLER_70_64 ();
 sg13g2_fill_1 FILLER_70_73 ();
 sg13g2_fill_1 FILLER_70_111 ();
 sg13g2_fill_2 FILLER_70_148 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_2 FILLER_70_204 ();
 sg13g2_fill_1 FILLER_70_219 ();
 sg13g2_fill_2 FILLER_70_224 ();
 sg13g2_fill_2 FILLER_70_238 ();
 sg13g2_fill_1 FILLER_70_275 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_2 FILLER_70_293 ();
 sg13g2_fill_1 FILLER_70_299 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_decap_4 FILLER_70_319 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_70_375 ();
 sg13g2_fill_1 FILLER_70_402 ();
 sg13g2_fill_1 FILLER_70_472 ();
 sg13g2_fill_2 FILLER_70_495 ();
 sg13g2_fill_1 FILLER_70_502 ();
 sg13g2_fill_1 FILLER_70_513 ();
 sg13g2_fill_1 FILLER_70_528 ();
 sg13g2_fill_2 FILLER_70_577 ();
 sg13g2_fill_1 FILLER_70_579 ();
 sg13g2_fill_1 FILLER_70_585 ();
 sg13g2_fill_1 FILLER_70_612 ();
 sg13g2_fill_1 FILLER_70_618 ();
 sg13g2_fill_1 FILLER_70_624 ();
 sg13g2_fill_2 FILLER_70_629 ();
 sg13g2_fill_2 FILLER_70_635 ();
 sg13g2_fill_2 FILLER_70_642 ();
 sg13g2_decap_8 FILLER_70_682 ();
 sg13g2_fill_2 FILLER_70_739 ();
 sg13g2_fill_1 FILLER_70_749 ();
 sg13g2_fill_1 FILLER_70_758 ();
 sg13g2_fill_1 FILLER_70_777 ();
 sg13g2_fill_1 FILLER_70_787 ();
 sg13g2_fill_1 FILLER_70_793 ();
 sg13g2_fill_2 FILLER_70_803 ();
 sg13g2_fill_2 FILLER_70_814 ();
 sg13g2_fill_2 FILLER_70_821 ();
 sg13g2_fill_2 FILLER_70_858 ();
 sg13g2_fill_2 FILLER_70_870 ();
 sg13g2_fill_2 FILLER_70_908 ();
 sg13g2_fill_1 FILLER_70_910 ();
 sg13g2_fill_2 FILLER_70_915 ();
 sg13g2_fill_1 FILLER_70_922 ();
 sg13g2_fill_1 FILLER_70_967 ();
 sg13g2_fill_1 FILLER_70_977 ();
 sg13g2_fill_2 FILLER_70_986 ();
 sg13g2_fill_1 FILLER_70_996 ();
 sg13g2_fill_1 FILLER_70_1032 ();
 sg13g2_decap_4 FILLER_70_1086 ();
 sg13g2_fill_1 FILLER_70_1090 ();
 sg13g2_fill_1 FILLER_70_1105 ();
 sg13g2_fill_1 FILLER_70_1137 ();
 sg13g2_fill_1 FILLER_70_1146 ();
 sg13g2_fill_1 FILLER_70_1215 ();
 sg13g2_fill_2 FILLER_70_1220 ();
 sg13g2_fill_1 FILLER_70_1222 ();
 sg13g2_fill_1 FILLER_70_1232 ();
 sg13g2_fill_2 FILLER_70_1258 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_8 FILLER_70_1298 ();
 sg13g2_decap_8 FILLER_70_1305 ();
 sg13g2_decap_8 FILLER_70_1312 ();
 sg13g2_decap_8 FILLER_70_1319 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_fill_1 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_47 ();
 sg13g2_decap_4 FILLER_71_54 ();
 sg13g2_fill_2 FILLER_71_58 ();
 sg13g2_fill_2 FILLER_71_75 ();
 sg13g2_fill_1 FILLER_71_81 ();
 sg13g2_fill_1 FILLER_71_86 ();
 sg13g2_fill_1 FILLER_71_98 ();
 sg13g2_fill_2 FILLER_71_130 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_1 FILLER_71_185 ();
 sg13g2_fill_1 FILLER_71_217 ();
 sg13g2_fill_1 FILLER_71_244 ();
 sg13g2_fill_2 FILLER_71_254 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_286 ();
 sg13g2_fill_1 FILLER_71_293 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_2 FILLER_71_356 ();
 sg13g2_fill_2 FILLER_71_363 ();
 sg13g2_fill_2 FILLER_71_369 ();
 sg13g2_fill_2 FILLER_71_380 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_397 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_456 ();
 sg13g2_fill_1 FILLER_71_487 ();
 sg13g2_fill_2 FILLER_71_510 ();
 sg13g2_fill_1 FILLER_71_512 ();
 sg13g2_fill_1 FILLER_71_530 ();
 sg13g2_fill_1 FILLER_71_557 ();
 sg13g2_fill_1 FILLER_71_596 ();
 sg13g2_fill_1 FILLER_71_601 ();
 sg13g2_fill_2 FILLER_71_641 ();
 sg13g2_fill_1 FILLER_71_663 ();
 sg13g2_decap_8 FILLER_71_684 ();
 sg13g2_fill_1 FILLER_71_701 ();
 sg13g2_fill_1 FILLER_71_706 ();
 sg13g2_fill_1 FILLER_71_710 ();
 sg13g2_fill_1 FILLER_71_720 ();
 sg13g2_fill_2 FILLER_71_747 ();
 sg13g2_fill_1 FILLER_71_749 ();
 sg13g2_fill_2 FILLER_71_781 ();
 sg13g2_fill_2 FILLER_71_837 ();
 sg13g2_fill_2 FILLER_71_946 ();
 sg13g2_decap_4 FILLER_71_983 ();
 sg13g2_fill_1 FILLER_71_992 ();
 sg13g2_fill_1 FILLER_71_1002 ();
 sg13g2_fill_2 FILLER_71_1008 ();
 sg13g2_fill_2 FILLER_71_1014 ();
 sg13g2_decap_4 FILLER_71_1020 ();
 sg13g2_fill_2 FILLER_71_1024 ();
 sg13g2_fill_2 FILLER_71_1070 ();
 sg13g2_fill_1 FILLER_71_1072 ();
 sg13g2_decap_4 FILLER_71_1099 ();
 sg13g2_fill_2 FILLER_71_1129 ();
 sg13g2_fill_2 FILLER_71_1186 ();
 sg13g2_fill_1 FILLER_71_1218 ();
 sg13g2_fill_1 FILLER_71_1258 ();
 sg13g2_fill_1 FILLER_71_1263 ();
 sg13g2_fill_1 FILLER_71_1268 ();
 sg13g2_fill_2 FILLER_71_1273 ();
 sg13g2_decap_8 FILLER_71_1290 ();
 sg13g2_decap_8 FILLER_71_1297 ();
 sg13g2_decap_8 FILLER_71_1304 ();
 sg13g2_decap_8 FILLER_71_1311 ();
 sg13g2_decap_8 FILLER_71_1318 ();
 sg13g2_fill_1 FILLER_71_1325 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_4 FILLER_72_56 ();
 sg13g2_fill_1 FILLER_72_60 ();
 sg13g2_fill_1 FILLER_72_174 ();
 sg13g2_fill_1 FILLER_72_180 ();
 sg13g2_fill_2 FILLER_72_193 ();
 sg13g2_fill_1 FILLER_72_219 ();
 sg13g2_fill_1 FILLER_72_229 ();
 sg13g2_fill_1 FILLER_72_256 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_325 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_340 ();
 sg13g2_fill_1 FILLER_72_393 ();
 sg13g2_fill_1 FILLER_72_452 ();
 sg13g2_fill_1 FILLER_72_457 ();
 sg13g2_fill_1 FILLER_72_489 ();
 sg13g2_fill_2 FILLER_72_530 ();
 sg13g2_fill_1 FILLER_72_532 ();
 sg13g2_fill_1 FILLER_72_541 ();
 sg13g2_fill_2 FILLER_72_568 ();
 sg13g2_fill_2 FILLER_72_575 ();
 sg13g2_fill_2 FILLER_72_617 ();
 sg13g2_fill_1 FILLER_72_624 ();
 sg13g2_fill_2 FILLER_72_629 ();
 sg13g2_fill_2 FILLER_72_636 ();
 sg13g2_fill_1 FILLER_72_638 ();
 sg13g2_fill_2 FILLER_72_669 ();
 sg13g2_fill_1 FILLER_72_680 ();
 sg13g2_fill_1 FILLER_72_697 ();
 sg13g2_fill_1 FILLER_72_703 ();
 sg13g2_fill_2 FILLER_72_708 ();
 sg13g2_fill_1 FILLER_72_715 ();
 sg13g2_fill_1 FILLER_72_720 ();
 sg13g2_fill_1 FILLER_72_725 ();
 sg13g2_fill_2 FILLER_72_730 ();
 sg13g2_fill_1 FILLER_72_785 ();
 sg13g2_fill_2 FILLER_72_795 ();
 sg13g2_fill_1 FILLER_72_806 ();
 sg13g2_fill_1 FILLER_72_845 ();
 sg13g2_fill_1 FILLER_72_852 ();
 sg13g2_fill_2 FILLER_72_915 ();
 sg13g2_fill_1 FILLER_72_917 ();
 sg13g2_fill_1 FILLER_72_923 ();
 sg13g2_fill_2 FILLER_72_929 ();
 sg13g2_fill_1 FILLER_72_931 ();
 sg13g2_fill_2 FILLER_72_1001 ();
 sg13g2_fill_1 FILLER_72_1007 ();
 sg13g2_fill_2 FILLER_72_1044 ();
 sg13g2_fill_1 FILLER_72_1056 ();
 sg13g2_fill_2 FILLER_72_1077 ();
 sg13g2_fill_2 FILLER_72_1095 ();
 sg13g2_fill_1 FILLER_72_1107 ();
 sg13g2_fill_1 FILLER_72_1113 ();
 sg13g2_fill_2 FILLER_72_1158 ();
 sg13g2_fill_1 FILLER_72_1164 ();
 sg13g2_fill_1 FILLER_72_1174 ();
 sg13g2_fill_1 FILLER_72_1201 ();
 sg13g2_decap_8 FILLER_72_1285 ();
 sg13g2_decap_8 FILLER_72_1292 ();
 sg13g2_decap_8 FILLER_72_1299 ();
 sg13g2_decap_8 FILLER_72_1306 ();
 sg13g2_decap_8 FILLER_72_1313 ();
 sg13g2_decap_4 FILLER_72_1320 ();
 sg13g2_fill_2 FILLER_72_1324 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_4 FILLER_73_49 ();
 sg13g2_fill_2 FILLER_73_53 ();
 sg13g2_fill_2 FILLER_73_95 ();
 sg13g2_fill_1 FILLER_73_122 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_fill_2 FILLER_73_142 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_1 FILLER_73_160 ();
 sg13g2_fill_1 FILLER_73_173 ();
 sg13g2_fill_2 FILLER_73_223 ();
 sg13g2_fill_1 FILLER_73_229 ();
 sg13g2_fill_2 FILLER_73_247 ();
 sg13g2_fill_1 FILLER_73_253 ();
 sg13g2_fill_1 FILLER_73_259 ();
 sg13g2_fill_1 FILLER_73_295 ();
 sg13g2_fill_1 FILLER_73_299 ();
 sg13g2_fill_1 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_331 ();
 sg13g2_fill_1 FILLER_73_337 ();
 sg13g2_fill_1 FILLER_73_343 ();
 sg13g2_fill_2 FILLER_73_349 ();
 sg13g2_fill_1 FILLER_73_369 ();
 sg13g2_fill_2 FILLER_73_379 ();
 sg13g2_fill_1 FILLER_73_390 ();
 sg13g2_fill_1 FILLER_73_395 ();
 sg13g2_fill_1 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_405 ();
 sg13g2_fill_2 FILLER_73_424 ();
 sg13g2_fill_2 FILLER_73_463 ();
 sg13g2_fill_1 FILLER_73_492 ();
 sg13g2_fill_2 FILLER_73_534 ();
 sg13g2_fill_1 FILLER_73_541 ();
 sg13g2_fill_1 FILLER_73_547 ();
 sg13g2_fill_2 FILLER_73_552 ();
 sg13g2_fill_1 FILLER_73_559 ();
 sg13g2_fill_2 FILLER_73_565 ();
 sg13g2_fill_2 FILLER_73_571 ();
 sg13g2_fill_1 FILLER_73_573 ();
 sg13g2_fill_2 FILLER_73_620 ();
 sg13g2_fill_1 FILLER_73_648 ();
 sg13g2_decap_4 FILLER_73_666 ();
 sg13g2_fill_2 FILLER_73_670 ();
 sg13g2_fill_2 FILLER_73_697 ();
 sg13g2_fill_1 FILLER_73_712 ();
 sg13g2_decap_8 FILLER_73_743 ();
 sg13g2_decap_4 FILLER_73_750 ();
 sg13g2_fill_1 FILLER_73_754 ();
 sg13g2_fill_2 FILLER_73_789 ();
 sg13g2_fill_1 FILLER_73_791 ();
 sg13g2_fill_1 FILLER_73_796 ();
 sg13g2_fill_2 FILLER_73_815 ();
 sg13g2_fill_2 FILLER_73_840 ();
 sg13g2_fill_1 FILLER_73_917 ();
 sg13g2_fill_2 FILLER_73_923 ();
 sg13g2_fill_1 FILLER_73_925 ();
 sg13g2_decap_8 FILLER_73_956 ();
 sg13g2_decap_4 FILLER_73_963 ();
 sg13g2_fill_1 FILLER_73_967 ();
 sg13g2_decap_4 FILLER_73_982 ();
 sg13g2_decap_4 FILLER_73_991 ();
 sg13g2_decap_8 FILLER_73_1037 ();
 sg13g2_fill_2 FILLER_73_1044 ();
 sg13g2_fill_1 FILLER_73_1046 ();
 sg13g2_fill_2 FILLER_73_1073 ();
 sg13g2_fill_1 FILLER_73_1083 ();
 sg13g2_decap_4 FILLER_73_1146 ();
 sg13g2_fill_2 FILLER_73_1150 ();
 sg13g2_fill_2 FILLER_73_1156 ();
 sg13g2_fill_1 FILLER_73_1196 ();
 sg13g2_fill_2 FILLER_73_1215 ();
 sg13g2_fill_2 FILLER_73_1222 ();
 sg13g2_decap_8 FILLER_73_1277 ();
 sg13g2_decap_8 FILLER_73_1284 ();
 sg13g2_decap_8 FILLER_73_1291 ();
 sg13g2_decap_8 FILLER_73_1298 ();
 sg13g2_decap_8 FILLER_73_1305 ();
 sg13g2_decap_8 FILLER_73_1312 ();
 sg13g2_decap_8 FILLER_73_1319 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_56 ();
 sg13g2_fill_1 FILLER_74_58 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_4 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_87 ();
 sg13g2_fill_1 FILLER_74_91 ();
 sg13g2_fill_2 FILLER_74_122 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_2 FILLER_74_236 ();
 sg13g2_fill_2 FILLER_74_264 ();
 sg13g2_fill_1 FILLER_74_276 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_fill_2 FILLER_74_296 ();
 sg13g2_fill_1 FILLER_74_298 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_fill_1 FILLER_74_314 ();
 sg13g2_fill_1 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_325 ();
 sg13g2_fill_2 FILLER_74_352 ();
 sg13g2_fill_2 FILLER_74_380 ();
 sg13g2_fill_2 FILLER_74_387 ();
 sg13g2_fill_1 FILLER_74_441 ();
 sg13g2_fill_1 FILLER_74_454 ();
 sg13g2_fill_1 FILLER_74_481 ();
 sg13g2_fill_2 FILLER_74_605 ();
 sg13g2_fill_1 FILLER_74_612 ();
 sg13g2_fill_1 FILLER_74_618 ();
 sg13g2_fill_1 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_629 ();
 sg13g2_decap_8 FILLER_74_634 ();
 sg13g2_decap_8 FILLER_74_641 ();
 sg13g2_fill_2 FILLER_74_670 ();
 sg13g2_fill_2 FILLER_74_690 ();
 sg13g2_fill_1 FILLER_74_696 ();
 sg13g2_fill_2 FILLER_74_702 ();
 sg13g2_fill_1 FILLER_74_708 ();
 sg13g2_fill_2 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_fill_1 FILLER_74_727 ();
 sg13g2_fill_2 FILLER_74_763 ();
 sg13g2_fill_1 FILLER_74_765 ();
 sg13g2_fill_2 FILLER_74_792 ();
 sg13g2_fill_2 FILLER_74_820 ();
 sg13g2_decap_4 FILLER_74_830 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_fill_1 FILLER_74_878 ();
 sg13g2_fill_2 FILLER_74_893 ();
 sg13g2_decap_4 FILLER_74_923 ();
 sg13g2_decap_4 FILLER_74_949 ();
 sg13g2_fill_2 FILLER_74_1005 ();
 sg13g2_fill_1 FILLER_74_1007 ();
 sg13g2_decap_4 FILLER_74_1047 ();
 sg13g2_decap_4 FILLER_74_1059 ();
 sg13g2_fill_2 FILLER_74_1063 ();
 sg13g2_fill_2 FILLER_74_1070 ();
 sg13g2_fill_1 FILLER_74_1085 ();
 sg13g2_fill_2 FILLER_74_1129 ();
 sg13g2_decap_8 FILLER_74_1139 ();
 sg13g2_decap_4 FILLER_74_1146 ();
 sg13g2_decap_4 FILLER_74_1154 ();
 sg13g2_fill_2 FILLER_74_1174 ();
 sg13g2_fill_1 FILLER_74_1228 ();
 sg13g2_fill_2 FILLER_74_1246 ();
 sg13g2_decap_8 FILLER_74_1274 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_decap_8 FILLER_74_1288 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_8 FILLER_74_1309 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_fill_2 FILLER_74_1323 ();
 sg13g2_fill_1 FILLER_74_1325 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_fill_2 FILLER_75_124 ();
 sg13g2_fill_1 FILLER_75_147 ();
 sg13g2_fill_1 FILLER_75_178 ();
 sg13g2_fill_2 FILLER_75_198 ();
 sg13g2_fill_1 FILLER_75_204 ();
 sg13g2_fill_2 FILLER_75_276 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_308 ();
 sg13g2_fill_2 FILLER_75_313 ();
 sg13g2_decap_4 FILLER_75_330 ();
 sg13g2_fill_2 FILLER_75_348 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_2 FILLER_75_399 ();
 sg13g2_fill_1 FILLER_75_405 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_fill_1 FILLER_75_417 ();
 sg13g2_fill_1 FILLER_75_426 ();
 sg13g2_fill_1 FILLER_75_431 ();
 sg13g2_fill_2 FILLER_75_445 ();
 sg13g2_fill_2 FILLER_75_451 ();
 sg13g2_fill_1 FILLER_75_458 ();
 sg13g2_fill_1 FILLER_75_467 ();
 sg13g2_fill_1 FILLER_75_477 ();
 sg13g2_fill_2 FILLER_75_491 ();
 sg13g2_fill_1 FILLER_75_497 ();
 sg13g2_fill_1 FILLER_75_523 ();
 sg13g2_fill_2 FILLER_75_544 ();
 sg13g2_fill_2 FILLER_75_611 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_decap_4 FILLER_75_699 ();
 sg13g2_fill_2 FILLER_75_707 ();
 sg13g2_fill_1 FILLER_75_709 ();
 sg13g2_fill_2 FILLER_75_719 ();
 sg13g2_fill_1 FILLER_75_721 ();
 sg13g2_fill_1 FILLER_75_727 ();
 sg13g2_fill_1 FILLER_75_732 ();
 sg13g2_fill_1 FILLER_75_738 ();
 sg13g2_fill_2 FILLER_75_744 ();
 sg13g2_fill_2 FILLER_75_750 ();
 sg13g2_fill_1 FILLER_75_752 ();
 sg13g2_decap_4 FILLER_75_765 ();
 sg13g2_fill_1 FILLER_75_769 ();
 sg13g2_fill_1 FILLER_75_773 ();
 sg13g2_fill_1 FILLER_75_778 ();
 sg13g2_fill_1 FILLER_75_789 ();
 sg13g2_fill_2 FILLER_75_794 ();
 sg13g2_fill_2 FILLER_75_800 ();
 sg13g2_fill_2 FILLER_75_806 ();
 sg13g2_fill_2 FILLER_75_821 ();
 sg13g2_fill_1 FILLER_75_823 ();
 sg13g2_fill_1 FILLER_75_859 ();
 sg13g2_fill_2 FILLER_75_867 ();
 sg13g2_decap_4 FILLER_75_877 ();
 sg13g2_fill_1 FILLER_75_894 ();
 sg13g2_fill_1 FILLER_75_900 ();
 sg13g2_decap_8 FILLER_75_941 ();
 sg13g2_decap_8 FILLER_75_948 ();
 sg13g2_fill_2 FILLER_75_955 ();
 sg13g2_decap_8 FILLER_75_961 ();
 sg13g2_fill_2 FILLER_75_968 ();
 sg13g2_fill_1 FILLER_75_970 ();
 sg13g2_decap_4 FILLER_75_975 ();
 sg13g2_fill_1 FILLER_75_1030 ();
 sg13g2_fill_1 FILLER_75_1041 ();
 sg13g2_fill_1 FILLER_75_1094 ();
 sg13g2_fill_1 FILLER_75_1099 ();
 sg13g2_decap_4 FILLER_75_1108 ();
 sg13g2_decap_4 FILLER_75_1120 ();
 sg13g2_fill_2 FILLER_75_1140 ();
 sg13g2_fill_1 FILLER_75_1187 ();
 sg13g2_fill_1 FILLER_75_1193 ();
 sg13g2_fill_2 FILLER_75_1203 ();
 sg13g2_fill_1 FILLER_75_1205 ();
 sg13g2_fill_1 FILLER_75_1229 ();
 sg13g2_decap_8 FILLER_75_1261 ();
 sg13g2_decap_8 FILLER_75_1268 ();
 sg13g2_decap_8 FILLER_75_1275 ();
 sg13g2_decap_8 FILLER_75_1282 ();
 sg13g2_decap_8 FILLER_75_1289 ();
 sg13g2_decap_8 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1303 ();
 sg13g2_decap_8 FILLER_75_1310 ();
 sg13g2_decap_8 FILLER_75_1317 ();
 sg13g2_fill_2 FILLER_75_1324 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_fill_1 FILLER_76_84 ();
 sg13g2_fill_1 FILLER_76_90 ();
 sg13g2_fill_1 FILLER_76_117 ();
 sg13g2_fill_1 FILLER_76_126 ();
 sg13g2_fill_1 FILLER_76_135 ();
 sg13g2_fill_2 FILLER_76_146 ();
 sg13g2_fill_2 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_255 ();
 sg13g2_decap_4 FILLER_76_262 ();
 sg13g2_decap_4 FILLER_76_284 ();
 sg13g2_fill_2 FILLER_76_288 ();
 sg13g2_fill_1 FILLER_76_338 ();
 sg13g2_fill_1 FILLER_76_343 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_380 ();
 sg13g2_fill_1 FILLER_76_391 ();
 sg13g2_fill_2 FILLER_76_396 ();
 sg13g2_fill_2 FILLER_76_402 ();
 sg13g2_fill_1 FILLER_76_543 ();
 sg13g2_fill_1 FILLER_76_551 ();
 sg13g2_fill_1 FILLER_76_557 ();
 sg13g2_fill_1 FILLER_76_562 ();
 sg13g2_fill_1 FILLER_76_568 ();
 sg13g2_fill_1 FILLER_76_599 ();
 sg13g2_fill_1 FILLER_76_605 ();
 sg13g2_fill_2 FILLER_76_610 ();
 sg13g2_fill_1 FILLER_76_638 ();
 sg13g2_decap_8 FILLER_76_643 ();
 sg13g2_decap_8 FILLER_76_666 ();
 sg13g2_decap_8 FILLER_76_673 ();
 sg13g2_fill_2 FILLER_76_683 ();
 sg13g2_fill_1 FILLER_76_685 ();
 sg13g2_fill_2 FILLER_76_709 ();
 sg13g2_fill_2 FILLER_76_786 ();
 sg13g2_fill_1 FILLER_76_802 ();
 sg13g2_fill_2 FILLER_76_808 ();
 sg13g2_fill_2 FILLER_76_814 ();
 sg13g2_fill_2 FILLER_76_869 ();
 sg13g2_fill_1 FILLER_76_903 ();
 sg13g2_decap_8 FILLER_76_943 ();
 sg13g2_decap_8 FILLER_76_950 ();
 sg13g2_decap_8 FILLER_76_957 ();
 sg13g2_decap_8 FILLER_76_964 ();
 sg13g2_decap_8 FILLER_76_971 ();
 sg13g2_decap_4 FILLER_76_978 ();
 sg13g2_fill_2 FILLER_76_982 ();
 sg13g2_decap_8 FILLER_76_992 ();
 sg13g2_fill_2 FILLER_76_1004 ();
 sg13g2_fill_1 FILLER_76_1006 ();
 sg13g2_fill_1 FILLER_76_1038 ();
 sg13g2_fill_2 FILLER_76_1052 ();
 sg13g2_fill_1 FILLER_76_1054 ();
 sg13g2_fill_2 FILLER_76_1065 ();
 sg13g2_fill_1 FILLER_76_1075 ();
 sg13g2_fill_1 FILLER_76_1081 ();
 sg13g2_fill_2 FILLER_76_1092 ();
 sg13g2_fill_1 FILLER_76_1094 ();
 sg13g2_fill_1 FILLER_76_1100 ();
 sg13g2_fill_2 FILLER_76_1118 ();
 sg13g2_fill_2 FILLER_76_1150 ();
 sg13g2_fill_1 FILLER_76_1179 ();
 sg13g2_fill_1 FILLER_76_1185 ();
 sg13g2_fill_1 FILLER_76_1194 ();
 sg13g2_fill_1 FILLER_76_1200 ();
 sg13g2_fill_1 FILLER_76_1209 ();
 sg13g2_fill_1 FILLER_76_1222 ();
 sg13g2_decap_8 FILLER_76_1274 ();
 sg13g2_decap_8 FILLER_76_1281 ();
 sg13g2_decap_8 FILLER_76_1288 ();
 sg13g2_decap_8 FILLER_76_1295 ();
 sg13g2_decap_8 FILLER_76_1302 ();
 sg13g2_decap_8 FILLER_76_1309 ();
 sg13g2_decap_8 FILLER_76_1316 ();
 sg13g2_fill_2 FILLER_76_1323 ();
 sg13g2_fill_1 FILLER_76_1325 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_104 ();
 sg13g2_fill_1 FILLER_77_106 ();
 sg13g2_fill_2 FILLER_77_111 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_fill_2 FILLER_77_134 ();
 sg13g2_fill_2 FILLER_77_144 ();
 sg13g2_fill_2 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_171 ();
 sg13g2_fill_2 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_190 ();
 sg13g2_fill_1 FILLER_77_195 ();
 sg13g2_fill_2 FILLER_77_201 ();
 sg13g2_fill_1 FILLER_77_207 ();
 sg13g2_fill_2 FILLER_77_213 ();
 sg13g2_fill_1 FILLER_77_219 ();
 sg13g2_fill_2 FILLER_77_225 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_fill_1 FILLER_77_290 ();
 sg13g2_fill_1 FILLER_77_296 ();
 sg13g2_fill_1 FILLER_77_305 ();
 sg13g2_fill_1 FILLER_77_309 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_fill_1 FILLER_77_340 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_352 ();
 sg13g2_fill_2 FILLER_77_379 ();
 sg13g2_fill_2 FILLER_77_436 ();
 sg13g2_fill_1 FILLER_77_438 ();
 sg13g2_fill_2 FILLER_77_455 ();
 sg13g2_fill_1 FILLER_77_471 ();
 sg13g2_fill_2 FILLER_77_477 ();
 sg13g2_fill_2 FILLER_77_483 ();
 sg13g2_fill_2 FILLER_77_497 ();
 sg13g2_decap_4 FILLER_77_504 ();
 sg13g2_fill_2 FILLER_77_512 ();
 sg13g2_fill_1 FILLER_77_519 ();
 sg13g2_fill_1 FILLER_77_572 ();
 sg13g2_fill_1 FILLER_77_595 ();
 sg13g2_fill_1 FILLER_77_622 ();
 sg13g2_fill_1 FILLER_77_654 ();
 sg13g2_decap_4 FILLER_77_686 ();
 sg13g2_fill_1 FILLER_77_751 ();
 sg13g2_fill_2 FILLER_77_778 ();
 sg13g2_decap_4 FILLER_77_800 ();
 sg13g2_fill_2 FILLER_77_804 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_fill_2 FILLER_77_845 ();
 sg13g2_fill_1 FILLER_77_847 ();
 sg13g2_fill_1 FILLER_77_857 ();
 sg13g2_fill_2 FILLER_77_862 ();
 sg13g2_fill_1 FILLER_77_864 ();
 sg13g2_fill_2 FILLER_77_878 ();
 sg13g2_fill_1 FILLER_77_887 ();
 sg13g2_fill_1 FILLER_77_893 ();
 sg13g2_fill_1 FILLER_77_898 ();
 sg13g2_decap_8 FILLER_77_929 ();
 sg13g2_decap_8 FILLER_77_936 ();
 sg13g2_decap_8 FILLER_77_943 ();
 sg13g2_decap_8 FILLER_77_950 ();
 sg13g2_decap_8 FILLER_77_957 ();
 sg13g2_decap_8 FILLER_77_964 ();
 sg13g2_decap_8 FILLER_77_971 ();
 sg13g2_decap_8 FILLER_77_978 ();
 sg13g2_decap_8 FILLER_77_985 ();
 sg13g2_decap_8 FILLER_77_992 ();
 sg13g2_decap_4 FILLER_77_999 ();
 sg13g2_fill_1 FILLER_77_1003 ();
 sg13g2_decap_8 FILLER_77_1034 ();
 sg13g2_decap_8 FILLER_77_1041 ();
 sg13g2_decap_8 FILLER_77_1048 ();
 sg13g2_fill_1 FILLER_77_1055 ();
 sg13g2_fill_1 FILLER_77_1103 ();
 sg13g2_decap_8 FILLER_77_1109 ();
 sg13g2_fill_1 FILLER_77_1169 ();
 sg13g2_fill_2 FILLER_77_1200 ();
 sg13g2_decap_8 FILLER_77_1234 ();
 sg13g2_decap_8 FILLER_77_1241 ();
 sg13g2_fill_2 FILLER_77_1248 ();
 sg13g2_fill_1 FILLER_77_1250 ();
 sg13g2_decap_8 FILLER_77_1255 ();
 sg13g2_decap_8 FILLER_77_1262 ();
 sg13g2_decap_8 FILLER_77_1269 ();
 sg13g2_decap_8 FILLER_77_1276 ();
 sg13g2_decap_8 FILLER_77_1283 ();
 sg13g2_decap_8 FILLER_77_1290 ();
 sg13g2_decap_8 FILLER_77_1297 ();
 sg13g2_decap_8 FILLER_77_1304 ();
 sg13g2_decap_8 FILLER_77_1311 ();
 sg13g2_decap_8 FILLER_77_1318 ();
 sg13g2_fill_1 FILLER_77_1325 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_fill_2 FILLER_78_145 ();
 sg13g2_fill_1 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_240 ();
 sg13g2_fill_2 FILLER_78_246 ();
 sg13g2_fill_1 FILLER_78_278 ();
 sg13g2_fill_1 FILLER_78_287 ();
 sg13g2_fill_1 FILLER_78_292 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_fill_2 FILLER_78_302 ();
 sg13g2_fill_1 FILLER_78_309 ();
 sg13g2_fill_2 FILLER_78_314 ();
 sg13g2_fill_1 FILLER_78_371 ();
 sg13g2_fill_2 FILLER_78_381 ();
 sg13g2_fill_1 FILLER_78_383 ();
 sg13g2_fill_1 FILLER_78_401 ();
 sg13g2_decap_4 FILLER_78_445 ();
 sg13g2_fill_1 FILLER_78_462 ();
 sg13g2_fill_2 FILLER_78_493 ();
 sg13g2_fill_2 FILLER_78_521 ();
 sg13g2_fill_1 FILLER_78_523 ();
 sg13g2_decap_8 FILLER_78_538 ();
 sg13g2_fill_1 FILLER_78_605 ();
 sg13g2_fill_1 FILLER_78_616 ();
 sg13g2_fill_1 FILLER_78_621 ();
 sg13g2_fill_1 FILLER_78_627 ();
 sg13g2_fill_2 FILLER_78_633 ();
 sg13g2_fill_2 FILLER_78_640 ();
 sg13g2_fill_2 FILLER_78_647 ();
 sg13g2_fill_1 FILLER_78_661 ();
 sg13g2_fill_1 FILLER_78_667 ();
 sg13g2_fill_2 FILLER_78_673 ();
 sg13g2_fill_2 FILLER_78_707 ();
 sg13g2_fill_1 FILLER_78_714 ();
 sg13g2_decap_4 FILLER_78_760 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_fill_1 FILLER_78_776 ();
 sg13g2_fill_1 FILLER_78_816 ();
 sg13g2_fill_2 FILLER_78_829 ();
 sg13g2_fill_1 FILLER_78_856 ();
 sg13g2_fill_1 FILLER_78_880 ();
 sg13g2_decap_8 FILLER_78_925 ();
 sg13g2_decap_8 FILLER_78_932 ();
 sg13g2_decap_8 FILLER_78_939 ();
 sg13g2_decap_8 FILLER_78_946 ();
 sg13g2_decap_8 FILLER_78_953 ();
 sg13g2_decap_8 FILLER_78_960 ();
 sg13g2_decap_8 FILLER_78_967 ();
 sg13g2_decap_8 FILLER_78_974 ();
 sg13g2_decap_8 FILLER_78_981 ();
 sg13g2_decap_8 FILLER_78_988 ();
 sg13g2_decap_8 FILLER_78_995 ();
 sg13g2_decap_8 FILLER_78_1002 ();
 sg13g2_decap_4 FILLER_78_1009 ();
 sg13g2_decap_8 FILLER_78_1017 ();
 sg13g2_decap_8 FILLER_78_1024 ();
 sg13g2_decap_8 FILLER_78_1031 ();
 sg13g2_decap_8 FILLER_78_1038 ();
 sg13g2_decap_8 FILLER_78_1045 ();
 sg13g2_decap_8 FILLER_78_1052 ();
 sg13g2_fill_2 FILLER_78_1059 ();
 sg13g2_decap_8 FILLER_78_1065 ();
 sg13g2_decap_8 FILLER_78_1072 ();
 sg13g2_decap_8 FILLER_78_1079 ();
 sg13g2_fill_1 FILLER_78_1091 ();
 sg13g2_fill_2 FILLER_78_1109 ();
 sg13g2_fill_1 FILLER_78_1128 ();
 sg13g2_fill_1 FILLER_78_1133 ();
 sg13g2_fill_1 FILLER_78_1138 ();
 sg13g2_fill_1 FILLER_78_1143 ();
 sg13g2_fill_1 FILLER_78_1149 ();
 sg13g2_decap_4 FILLER_78_1196 ();
 sg13g2_fill_1 FILLER_78_1200 ();
 sg13g2_fill_1 FILLER_78_1210 ();
 sg13g2_decap_8 FILLER_78_1232 ();
 sg13g2_decap_8 FILLER_78_1239 ();
 sg13g2_decap_8 FILLER_78_1246 ();
 sg13g2_decap_8 FILLER_78_1253 ();
 sg13g2_decap_8 FILLER_78_1260 ();
 sg13g2_decap_8 FILLER_78_1267 ();
 sg13g2_decap_8 FILLER_78_1274 ();
 sg13g2_decap_8 FILLER_78_1281 ();
 sg13g2_decap_8 FILLER_78_1288 ();
 sg13g2_decap_8 FILLER_78_1295 ();
 sg13g2_decap_8 FILLER_78_1302 ();
 sg13g2_decap_8 FILLER_78_1309 ();
 sg13g2_decap_8 FILLER_78_1316 ();
 sg13g2_fill_2 FILLER_78_1323 ();
 sg13g2_fill_1 FILLER_78_1325 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_decap_4 FILLER_79_131 ();
 sg13g2_fill_2 FILLER_79_135 ();
 sg13g2_decap_8 FILLER_79_141 ();
 sg13g2_decap_4 FILLER_79_148 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_2 FILLER_79_161 ();
 sg13g2_fill_1 FILLER_79_167 ();
 sg13g2_decap_8 FILLER_79_198 ();
 sg13g2_decap_8 FILLER_79_205 ();
 sg13g2_decap_8 FILLER_79_212 ();
 sg13g2_decap_8 FILLER_79_219 ();
 sg13g2_decap_8 FILLER_79_230 ();
 sg13g2_decap_8 FILLER_79_237 ();
 sg13g2_decap_4 FILLER_79_244 ();
 sg13g2_decap_4 FILLER_79_274 ();
 sg13g2_fill_2 FILLER_79_320 ();
 sg13g2_fill_1 FILLER_79_326 ();
 sg13g2_fill_1 FILLER_79_336 ();
 sg13g2_fill_1 FILLER_79_341 ();
 sg13g2_fill_2 FILLER_79_346 ();
 sg13g2_fill_2 FILLER_79_374 ();
 sg13g2_fill_2 FILLER_79_402 ();
 sg13g2_fill_1 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_431 ();
 sg13g2_fill_2 FILLER_79_457 ();
 sg13g2_fill_2 FILLER_79_481 ();
 sg13g2_fill_1 FILLER_79_483 ();
 sg13g2_fill_1 FILLER_79_491 ();
 sg13g2_decap_4 FILLER_79_517 ();
 sg13g2_fill_1 FILLER_79_521 ();
 sg13g2_fill_2 FILLER_79_544 ();
 sg13g2_fill_1 FILLER_79_546 ();
 sg13g2_decap_4 FILLER_79_551 ();
 sg13g2_fill_2 FILLER_79_555 ();
 sg13g2_decap_8 FILLER_79_561 ();
 sg13g2_fill_2 FILLER_79_571 ();
 sg13g2_fill_1 FILLER_79_573 ();
 sg13g2_fill_2 FILLER_79_583 ();
 sg13g2_decap_8 FILLER_79_594 ();
 sg13g2_fill_1 FILLER_79_601 ();
 sg13g2_fill_1 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_642 ();
 sg13g2_decap_8 FILLER_79_649 ();
 sg13g2_decap_4 FILLER_79_656 ();
 sg13g2_fill_1 FILLER_79_660 ();
 sg13g2_fill_2 FILLER_79_687 ();
 sg13g2_fill_1 FILLER_79_689 ();
 sg13g2_decap_4 FILLER_79_737 ();
 sg13g2_fill_1 FILLER_79_750 ();
 sg13g2_decap_8 FILLER_79_765 ();
 sg13g2_fill_2 FILLER_79_785 ();
 sg13g2_fill_2 FILLER_79_816 ();
 sg13g2_fill_1 FILLER_79_818 ();
 sg13g2_decap_4 FILLER_79_823 ();
 sg13g2_fill_2 FILLER_79_832 ();
 sg13g2_fill_1 FILLER_79_834 ();
 sg13g2_fill_2 FILLER_79_845 ();
 sg13g2_fill_1 FILLER_79_847 ();
 sg13g2_decap_4 FILLER_79_860 ();
 sg13g2_fill_2 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_901 ();
 sg13g2_decap_8 FILLER_79_908 ();
 sg13g2_decap_8 FILLER_79_915 ();
 sg13g2_decap_8 FILLER_79_922 ();
 sg13g2_decap_8 FILLER_79_929 ();
 sg13g2_decap_8 FILLER_79_936 ();
 sg13g2_decap_8 FILLER_79_943 ();
 sg13g2_decap_8 FILLER_79_950 ();
 sg13g2_decap_8 FILLER_79_957 ();
 sg13g2_decap_8 FILLER_79_964 ();
 sg13g2_decap_8 FILLER_79_971 ();
 sg13g2_decap_8 FILLER_79_978 ();
 sg13g2_decap_8 FILLER_79_985 ();
 sg13g2_decap_8 FILLER_79_992 ();
 sg13g2_decap_8 FILLER_79_999 ();
 sg13g2_decap_8 FILLER_79_1006 ();
 sg13g2_decap_8 FILLER_79_1013 ();
 sg13g2_decap_8 FILLER_79_1020 ();
 sg13g2_decap_8 FILLER_79_1027 ();
 sg13g2_decap_8 FILLER_79_1034 ();
 sg13g2_decap_8 FILLER_79_1041 ();
 sg13g2_decap_8 FILLER_79_1048 ();
 sg13g2_decap_8 FILLER_79_1055 ();
 sg13g2_decap_8 FILLER_79_1062 ();
 sg13g2_decap_8 FILLER_79_1069 ();
 sg13g2_decap_4 FILLER_79_1076 ();
 sg13g2_fill_1 FILLER_79_1080 ();
 sg13g2_fill_1 FILLER_79_1107 ();
 sg13g2_fill_1 FILLER_79_1113 ();
 sg13g2_fill_1 FILLER_79_1145 ();
 sg13g2_fill_2 FILLER_79_1172 ();
 sg13g2_fill_2 FILLER_79_1186 ();
 sg13g2_fill_1 FILLER_79_1188 ();
 sg13g2_fill_2 FILLER_79_1194 ();
 sg13g2_decap_8 FILLER_79_1226 ();
 sg13g2_decap_8 FILLER_79_1233 ();
 sg13g2_decap_8 FILLER_79_1240 ();
 sg13g2_decap_8 FILLER_79_1247 ();
 sg13g2_decap_8 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1261 ();
 sg13g2_decap_8 FILLER_79_1268 ();
 sg13g2_decap_8 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1282 ();
 sg13g2_decap_8 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1296 ();
 sg13g2_decap_8 FILLER_79_1303 ();
 sg13g2_decap_8 FILLER_79_1310 ();
 sg13g2_decap_8 FILLER_79_1317 ();
 sg13g2_fill_2 FILLER_79_1324 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_decap_8 FILLER_80_249 ();
 sg13g2_fill_2 FILLER_80_264 ();
 sg13g2_decap_8 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_297 ();
 sg13g2_fill_1 FILLER_80_347 ();
 sg13g2_fill_1 FILLER_80_385 ();
 sg13g2_fill_2 FILLER_80_390 ();
 sg13g2_decap_4 FILLER_80_396 ();
 sg13g2_fill_2 FILLER_80_438 ();
 sg13g2_fill_2 FILLER_80_449 ();
 sg13g2_fill_2 FILLER_80_485 ();
 sg13g2_fill_2 FILLER_80_492 ();
 sg13g2_fill_1 FILLER_80_498 ();
 sg13g2_fill_2 FILLER_80_533 ();
 sg13g2_decap_8 FILLER_80_561 ();
 sg13g2_decap_8 FILLER_80_568 ();
 sg13g2_decap_8 FILLER_80_575 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_610 ();
 sg13g2_fill_1 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_622 ();
 sg13g2_decap_8 FILLER_80_629 ();
 sg13g2_decap_8 FILLER_80_636 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_8 FILLER_80_650 ();
 sg13g2_decap_8 FILLER_80_657 ();
 sg13g2_fill_2 FILLER_80_664 ();
 sg13g2_fill_1 FILLER_80_666 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_8 FILLER_80_678 ();
 sg13g2_fill_2 FILLER_80_685 ();
 sg13g2_fill_1 FILLER_80_687 ();
 sg13g2_fill_1 FILLER_80_692 ();
 sg13g2_fill_2 FILLER_80_719 ();
 sg13g2_decap_4 FILLER_80_747 ();
 sg13g2_fill_2 FILLER_80_789 ();
 sg13g2_fill_1 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_4 FILLER_80_839 ();
 sg13g2_decap_8 FILLER_80_853 ();
 sg13g2_decap_8 FILLER_80_860 ();
 sg13g2_decap_8 FILLER_80_867 ();
 sg13g2_fill_1 FILLER_80_874 ();
 sg13g2_decap_8 FILLER_80_879 ();
 sg13g2_decap_8 FILLER_80_886 ();
 sg13g2_decap_8 FILLER_80_893 ();
 sg13g2_decap_8 FILLER_80_900 ();
 sg13g2_decap_8 FILLER_80_907 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_949 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_977 ();
 sg13g2_decap_8 FILLER_80_984 ();
 sg13g2_decap_8 FILLER_80_991 ();
 sg13g2_decap_8 FILLER_80_998 ();
 sg13g2_decap_8 FILLER_80_1005 ();
 sg13g2_decap_8 FILLER_80_1012 ();
 sg13g2_decap_8 FILLER_80_1019 ();
 sg13g2_decap_8 FILLER_80_1026 ();
 sg13g2_decap_8 FILLER_80_1033 ();
 sg13g2_decap_8 FILLER_80_1040 ();
 sg13g2_decap_8 FILLER_80_1047 ();
 sg13g2_decap_8 FILLER_80_1054 ();
 sg13g2_decap_8 FILLER_80_1061 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_decap_8 FILLER_80_1075 ();
 sg13g2_decap_4 FILLER_80_1082 ();
 sg13g2_fill_1 FILLER_80_1086 ();
 sg13g2_decap_4 FILLER_80_1091 ();
 sg13g2_fill_1 FILLER_80_1095 ();
 sg13g2_decap_8 FILLER_80_1130 ();
 sg13g2_fill_2 FILLER_80_1137 ();
 sg13g2_fill_1 FILLER_80_1139 ();
 sg13g2_decap_4 FILLER_80_1144 ();
 sg13g2_fill_1 FILLER_80_1148 ();
 sg13g2_decap_4 FILLER_80_1157 ();
 sg13g2_fill_1 FILLER_80_1161 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_fill_2 FILLER_80_1181 ();
 sg13g2_decap_8 FILLER_80_1213 ();
 sg13g2_decap_8 FILLER_80_1220 ();
 sg13g2_decap_8 FILLER_80_1227 ();
 sg13g2_decap_8 FILLER_80_1234 ();
 sg13g2_decap_8 FILLER_80_1241 ();
 sg13g2_decap_8 FILLER_80_1248 ();
 sg13g2_decap_8 FILLER_80_1255 ();
 sg13g2_decap_8 FILLER_80_1262 ();
 sg13g2_decap_8 FILLER_80_1269 ();
 sg13g2_decap_8 FILLER_80_1276 ();
 sg13g2_decap_8 FILLER_80_1283 ();
 sg13g2_decap_8 FILLER_80_1290 ();
 sg13g2_decap_8 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1304 ();
 sg13g2_decap_8 FILLER_80_1311 ();
 sg13g2_decap_8 FILLER_80_1318 ();
 sg13g2_fill_1 FILLER_80_1325 ();
endmodule
