module tt_um_a1k0n_demo (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire _4704_;
 wire _4705_;
 wire _4706_;
 wire _4707_;
 wire _4708_;
 wire _4709_;
 wire _4710_;
 wire _4711_;
 wire _4712_;
 wire _4713_;
 wire _4714_;
 wire _4715_;
 wire _4716_;
 wire _4717_;
 wire _4718_;
 wire _4719_;
 wire _4720_;
 wire _4721_;
 wire _4722_;
 wire _4723_;
 wire _4724_;
 wire _4725_;
 wire _4726_;
 wire _4727_;
 wire _4728_;
 wire _4729_;
 wire _4730_;
 wire _4731_;
 wire _4732_;
 wire _4733_;
 wire _4734_;
 wire _4735_;
 wire _4736_;
 wire _4737_;
 wire _4738_;
 wire _4739_;
 wire _4740_;
 wire _4741_;
 wire _4742_;
 wire _4743_;
 wire _4744_;
 wire _4745_;
 wire _4746_;
 wire _4747_;
 wire _4748_;
 wire _4749_;
 wire _4750_;
 wire _4751_;
 wire _4752_;
 wire _4753_;
 wire _4754_;
 wire _4755_;
 wire _4756_;
 wire _4757_;
 wire _4758_;
 wire _4759_;
 wire _4760_;
 wire _4761_;
 wire _4762_;
 wire _4763_;
 wire _4764_;
 wire _4765_;
 wire _4766_;
 wire _4767_;
 wire _4768_;
 wire _4769_;
 wire _4770_;
 wire clknet_leaf_0_clk;
 wire net167;
 wire audio;
 wire hsync;
 wire \vgademo.a_cos[0] ;
 wire \vgademo.a_cos[10] ;
 wire \vgademo.a_cos[11] ;
 wire \vgademo.a_cos[12] ;
 wire \vgademo.a_cos[13] ;
 wire \vgademo.a_cos[14] ;
 wire \vgademo.a_cos[1] ;
 wire \vgademo.a_cos[2] ;
 wire \vgademo.a_cos[3] ;
 wire \vgademo.a_cos[4] ;
 wire \vgademo.a_cos[5] ;
 wire \vgademo.a_cos[6] ;
 wire \vgademo.a_cos[7] ;
 wire \vgademo.a_cos[8] ;
 wire \vgademo.a_cos[9] ;
 wire \vgademo.a_scrolly[10] ;
 wire \vgademo.a_scrolly[11] ;
 wire \vgademo.a_scrolly[12] ;
 wire \vgademo.a_scrolly[13] ;
 wire \vgademo.a_scrolly[3] ;
 wire \vgademo.a_scrolly[4] ;
 wire \vgademo.a_scrolly[5] ;
 wire \vgademo.a_scrolly[6] ;
 wire \vgademo.a_scrolly[7] ;
 wire \vgademo.a_scrolly[8] ;
 wire \vgademo.a_scrolly[9] ;
 wire \vgademo.a_sin[0] ;
 wire \vgademo.a_sin[10] ;
 wire \vgademo.a_sin[11] ;
 wire \vgademo.a_sin[12] ;
 wire \vgademo.a_sin[13] ;
 wire \vgademo.a_sin[14] ;
 wire \vgademo.a_sin[1] ;
 wire \vgademo.a_sin[2] ;
 wire \vgademo.a_sin[3] ;
 wire \vgademo.a_sin[4] ;
 wire \vgademo.a_sin[5] ;
 wire \vgademo.a_sin[6] ;
 wire \vgademo.a_sin[7] ;
 wire \vgademo.a_sin[8] ;
 wire \vgademo.a_sin[9] ;
 wire \vgademo.audio_beat_out[0] ;
 wire \vgademo.audio_beat_out[1] ;
 wire \vgademo.audio_beat_out[2] ;
 wire \vgademo.audio_beat_out[3] ;
 wire \vgademo.audio_beat_out[4] ;
 wire \vgademo.audio_kick_frames[0] ;
 wire \vgademo.audio_kick_frames[1] ;
 wire \vgademo.audio_kick_frames[2] ;
 wire \vgademo.audio_snare_frames[0] ;
 wire \vgademo.audio_snare_frames[1] ;
 wire \vgademo.audio_snare_frames[2] ;
 wire \vgademo.audio_snare_frames[3] ;
 wire \vgademo.audio_songpos[0] ;
 wire \vgademo.audio_songpos[1] ;
 wire \vgademo.audio_songpos[2] ;
 wire \vgademo.audio_songpos[3] ;
 wire \vgademo.audio_songpos[4] ;
 wire \vgademo.audio_songpos[5] ;
 wire \vgademo.audio_songpos[6] ;
 wire \vgademo.audio_songpos[7] ;
 wire \vgademo.b_cos[0] ;
 wire \vgademo.b_cos[10] ;
 wire \vgademo.b_cos[11] ;
 wire \vgademo.b_cos[1] ;
 wire \vgademo.b_cos[2] ;
 wire \vgademo.b_cos[3] ;
 wire \vgademo.b_cos[4] ;
 wire \vgademo.b_cos[5] ;
 wire \vgademo.b_cos[6] ;
 wire \vgademo.b_cos[7] ;
 wire \vgademo.b_cos[8] ;
 wire \vgademo.b_cos[9] ;
 wire \vgademo.b_sin[0] ;
 wire \vgademo.b_sin[10] ;
 wire \vgademo.b_sin[11] ;
 wire \vgademo.b_sin[1] ;
 wire \vgademo.b_sin[2] ;
 wire \vgademo.b_sin[3] ;
 wire \vgademo.b_sin[4] ;
 wire \vgademo.b_sin[5] ;
 wire \vgademo.b_sin[6] ;
 wire \vgademo.b_sin[7] ;
 wire \vgademo.b_sin[8] ;
 wire \vgademo.b_sin[9] ;
 wire \vgademo.bayer_j[0] ;
 wire \vgademo.bayer_j[1] ;
 wire \vgademo.h_count[0] ;
 wire \vgademo.h_count[10] ;
 wire \vgademo.h_count[1] ;
 wire \vgademo.h_count[2] ;
 wire \vgademo.h_count[3] ;
 wire \vgademo.h_count[4] ;
 wire \vgademo.h_count[5] ;
 wire \vgademo.h_count[6] ;
 wire \vgademo.h_count[7] ;
 wire \vgademo.h_count[8] ;
 wire \vgademo.h_count[9] ;
 wire \vgademo.linelfsr[0] ;
 wire \vgademo.linelfsr[10] ;
 wire \vgademo.linelfsr[11] ;
 wire \vgademo.linelfsr[12] ;
 wire \vgademo.linelfsr[1] ;
 wire \vgademo.linelfsr[2] ;
 wire \vgademo.linelfsr[3] ;
 wire \vgademo.linelfsr[4] ;
 wire \vgademo.linelfsr[5] ;
 wire \vgademo.linelfsr[6] ;
 wire \vgademo.linelfsr[7] ;
 wire \vgademo.linelfsr[8] ;
 wire \vgademo.linelfsr[9] ;
 wire \vgademo.plane_du[0] ;
 wire \vgademo.plane_du[10] ;
 wire \vgademo.plane_du[1] ;
 wire \vgademo.plane_du[2] ;
 wire \vgademo.plane_du[3] ;
 wire \vgademo.plane_du[4] ;
 wire \vgademo.plane_du[5] ;
 wire \vgademo.plane_du[6] ;
 wire \vgademo.plane_du[7] ;
 wire \vgademo.plane_du[8] ;
 wire \vgademo.plane_du[9] ;
 wire \vgademo.plane_dx[0] ;
 wire \vgademo.plane_dx[1] ;
 wire \vgademo.plane_dx[2] ;
 wire \vgademo.plane_dx_div.d[16] ;
 wire \vgademo.plane_dx_div.d[17] ;
 wire \vgademo.plane_dx_div.d[18] ;
 wire \vgademo.plane_dx_div.d[19] ;
 wire \vgademo.plane_dx_div.d[20] ;
 wire \vgademo.plane_dx_div.d[21] ;
 wire \vgademo.plane_dx_div.d[22] ;
 wire \vgademo.plane_dx_div.d[23] ;
 wire \vgademo.plane_dx_div.d[24] ;
 wire \vgademo.plane_dx_div.i[0] ;
 wire \vgademo.plane_dx_div.i[1] ;
 wire \vgademo.plane_dx_div.i[2] ;
 wire \vgademo.plane_dx_div.i[3] ;
 wire \vgademo.plane_dx_div.q[2] ;
 wire \vgademo.plane_dx_div.q[3] ;
 wire \vgademo.plane_dx_div.q[4] ;
 wire \vgademo.plane_dx_div.q[5] ;
 wire \vgademo.plane_dx_div.q[6] ;
 wire \vgademo.plane_dx_div.q[7] ;
 wire \vgademo.plane_dx_div.q[8] ;
 wire \vgademo.plane_dx_div.q[9] ;
 wire \vgademo.plane_dx_div.r[16] ;
 wire \vgademo.plane_dx_div.r[17] ;
 wire \vgademo.plane_dx_div.r[18] ;
 wire \vgademo.plane_dx_div.r[19] ;
 wire \vgademo.plane_dx_div.r[20] ;
 wire \vgademo.plane_dx_div.r[21] ;
 wire \vgademo.plane_dx_div.r[22] ;
 wire \vgademo.plane_dx_div.r[23] ;
 wire \vgademo.plane_dx_div.r[24] ;
 wire \vgademo.plane_dx_div.r[25] ;
 wire \vgademo.plane_u[0] ;
 wire \vgademo.plane_u[10] ;
 wire \vgademo.plane_u[11] ;
 wire \vgademo.plane_u[12] ;
 wire \vgademo.plane_u[13] ;
 wire \vgademo.plane_u[14] ;
 wire \vgademo.plane_u[15] ;
 wire \vgademo.plane_u[16] ;
 wire \vgademo.plane_u[17] ;
 wire \vgademo.plane_u[18] ;
 wire \vgademo.plane_u[19] ;
 wire \vgademo.plane_u[1] ;
 wire \vgademo.plane_u[20] ;
 wire \vgademo.plane_u[21] ;
 wire \vgademo.plane_u[2] ;
 wire \vgademo.plane_u[3] ;
 wire \vgademo.plane_u[4] ;
 wire \vgademo.plane_u[5] ;
 wire \vgademo.plane_u[6] ;
 wire \vgademo.plane_u[7] ;
 wire \vgademo.plane_u[8] ;
 wire \vgademo.plane_u[9] ;
 wire \vgademo.scanline_audio_sample[0] ;
 wire \vgademo.scanline_audio_sample[1] ;
 wire \vgademo.scanline_audio_sample[2] ;
 wire \vgademo.scanline_audio_sample[3] ;
 wire \vgademo.scanline_audio_sample[4] ;
 wire \vgademo.scanline_audio_sample[5] ;
 wire \vgademo.scanline_audio_sample[6] ;
 wire \vgademo.soundtrack.noise_lfsr[0] ;
 wire \vgademo.soundtrack.noise_lfsr[10] ;
 wire \vgademo.soundtrack.noise_lfsr[11] ;
 wire \vgademo.soundtrack.noise_lfsr[12] ;
 wire \vgademo.soundtrack.noise_lfsr[13] ;
 wire \vgademo.soundtrack.noise_lfsr[14] ;
 wire \vgademo.soundtrack.noise_lfsr[1] ;
 wire \vgademo.soundtrack.noise_lfsr[2] ;
 wire \vgademo.soundtrack.noise_lfsr[3] ;
 wire \vgademo.soundtrack.noise_lfsr[4] ;
 wire \vgademo.soundtrack.noise_lfsr[5] ;
 wire \vgademo.soundtrack.noise_lfsr[6] ;
 wire \vgademo.soundtrack.noise_lfsr[7] ;
 wire \vgademo.soundtrack.noise_lfsr[8] ;
 wire \vgademo.soundtrack.noise_lfsr[9] ;
 wire \vgademo.soundtrack.pulse_osc_p[0] ;
 wire \vgademo.soundtrack.pulse_osc_p[10] ;
 wire \vgademo.soundtrack.pulse_osc_p[11] ;
 wire \vgademo.soundtrack.pulse_osc_p[12] ;
 wire \vgademo.soundtrack.pulse_osc_p[13] ;
 wire \vgademo.soundtrack.pulse_osc_p[1] ;
 wire \vgademo.soundtrack.pulse_osc_p[2] ;
 wire \vgademo.soundtrack.pulse_osc_p[3] ;
 wire \vgademo.soundtrack.pulse_osc_p[4] ;
 wire \vgademo.soundtrack.pulse_osc_p[5] ;
 wire \vgademo.soundtrack.pulse_osc_p[6] ;
 wire \vgademo.soundtrack.pulse_osc_p[7] ;
 wire \vgademo.soundtrack.pulse_osc_p[8] ;
 wire \vgademo.soundtrack.pulse_osc_p[9] ;
 wire \vgademo.soundtrack.pulse_vol[0] ;
 wire \vgademo.soundtrack.pulse_vol[1] ;
 wire \vgademo.soundtrack.pulse_vol[2] ;
 wire \vgademo.soundtrack.pulse_vol[3] ;
 wire \vgademo.soundtrack.sample_div[0] ;
 wire \vgademo.soundtrack.sample_div[1] ;
 wire \vgademo.soundtrack.sample_div[2] ;
 wire \vgademo.soundtrack.sample_div[3] ;
 wire \vgademo.soundtrack.sample_div[4] ;
 wire \vgademo.soundtrack.sample_div[5] ;
 wire \vgademo.soundtrack.sample_div[6] ;
 wire \vgademo.soundtrack.sample_div[7] ;
 wire \vgademo.soundtrack.sample_div[8] ;
 wire \vgademo.soundtrack.sample_div[9] ;
 wire \vgademo.soundtrack.sample_div_[0] ;
 wire \vgademo.soundtrack.sample_div_[1] ;
 wire \vgademo.soundtrack.sample_div_[2] ;
 wire \vgademo.soundtrack.sample_div_[3] ;
 wire \vgademo.soundtrack.sample_div_[4] ;
 wire \vgademo.soundtrack.sample_div_[5] ;
 wire \vgademo.soundtrack.sample_div_[6] ;
 wire \vgademo.soundtrack.sample_div_[7] ;
 wire \vgademo.soundtrack.sample_div_[8] ;
 wire \vgademo.soundtrack.sample_div_[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum[9] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[0] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[10] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[11] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[12] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[13] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[14] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[15] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[1] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[2] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[3] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[4] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[5] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[6] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[7] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[8] ;
 wire \vgademo.soundtrack.sigma_delta_accum_[9] ;
 wire \vgademo.soundtrack.tick_div[0] ;
 wire \vgademo.soundtrack.tick_div[1] ;
 wire \vgademo.soundtrack.tick_div[2] ;
 wire \vgademo.soundtrack.tick_div[3] ;
 wire \vgademo.soundtrack.tick_div[4] ;
 wire \vgademo.soundtrack.tick_div[5] ;
 wire \vgademo.soundtrack.tick_div[6] ;
 wire \vgademo.soundtrack.tick_div[7] ;
 wire \vgademo.soundtrack.tick_div_[0] ;
 wire \vgademo.soundtrack.tri_osc_i[0] ;
 wire \vgademo.soundtrack.tri_osc_i[1] ;
 wire \vgademo.soundtrack.tri_osc_i[2] ;
 wire \vgademo.soundtrack.tri_osc_i[3] ;
 wire \vgademo.soundtrack.tri_osc_i[4] ;
 wire \vgademo.soundtrack.tri_osc_i[5] ;
 wire \vgademo.soundtrack.tri_osc_i[6] ;
 wire \vgademo.soundtrack.tri_osc_i[7] ;
 wire \vgademo.soundtrack.tri_osc_i[8] ;
 wire \vgademo.soundtrack.tri_osc_p[0] ;
 wire \vgademo.soundtrack.tri_osc_p[10] ;
 wire \vgademo.soundtrack.tri_osc_p[11] ;
 wire \vgademo.soundtrack.tri_osc_p[12] ;
 wire \vgademo.soundtrack.tri_osc_p[13] ;
 wire \vgademo.soundtrack.tri_osc_p[14] ;
 wire \vgademo.soundtrack.tri_osc_p[15] ;
 wire \vgademo.soundtrack.tri_osc_p[1] ;
 wire \vgademo.soundtrack.tri_osc_p[2] ;
 wire \vgademo.soundtrack.tri_osc_p[3] ;
 wire \vgademo.soundtrack.tri_osc_p[4] ;
 wire \vgademo.soundtrack.tri_osc_p[5] ;
 wire \vgademo.soundtrack.tri_osc_p[6] ;
 wire \vgademo.soundtrack.tri_osc_p[7] ;
 wire \vgademo.soundtrack.tri_osc_p[8] ;
 wire \vgademo.soundtrack.tri_osc_p[9] ;
 wire \vgademo.v_count[2] ;
 wire \vgademo.v_count[3] ;
 wire \vgademo.v_count[4] ;
 wire \vgademo.v_count[5] ;
 wire \vgademo.v_count[6] ;
 wire \vgademo.v_count[7] ;
 wire \vgademo.v_count[8] ;
 wire \vgademo.v_count[9] ;
 wire \vgademo.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_1 _4773_ (.A(\vgademo.h_count[0] ),
    .X(_4275_));
 sg13g2_buf_1 _4774_ (.A(\vgademo.h_count[1] ),
    .X(_4276_));
 sg13g2_buf_1 _4775_ (.A(\vgademo.h_count[3] ),
    .X(_4277_));
 sg13g2_buf_2 _4776_ (.A(\vgademo.h_count[2] ),
    .X(_4278_));
 sg13g2_inv_2 _4777_ (.Y(_4279_),
    .A(_4278_));
 sg13g2_nor4_2 _4778_ (.A(net127),
    .B(net126),
    .C(net125),
    .Y(_4280_),
    .D(_4279_));
 sg13g2_buf_2 _4779_ (.A(\vgademo.h_count[7] ),
    .X(_4281_));
 sg13g2_inv_1 _4780_ (.Y(_4282_),
    .A(_4281_));
 sg13g2_buf_1 _4781_ (.A(\vgademo.h_count[6] ),
    .X(_4283_));
 sg13g2_buf_1 _4782_ (.A(\vgademo.h_count[4] ),
    .X(_4284_));
 sg13g2_buf_2 _4783_ (.A(\vgademo.h_count[5] ),
    .X(_4285_));
 sg13g2_nand2_1 _4784_ (.Y(_4286_),
    .A(net123),
    .B(_4285_));
 sg13g2_nor3_1 _4785_ (.A(_4282_),
    .B(_4283_),
    .C(_4286_),
    .Y(_4287_));
 sg13g2_buf_2 _4786_ (.A(_0078_),
    .X(_4288_));
 sg13g2_buf_2 _4787_ (.A(\vgademo.h_count[9] ),
    .X(_4289_));
 sg13g2_nor2_1 _4788_ (.A(_4289_),
    .B(\vgademo.h_count[8] ),
    .Y(_4290_));
 sg13g2_inv_1 _4789_ (.Y(_4291_),
    .A(_4290_));
 sg13g2_nor2_1 _4790_ (.A(_4288_),
    .B(_4291_),
    .Y(_4292_));
 sg13g2_nand3_1 _4791_ (.B(_4287_),
    .C(_4292_),
    .A(_4280_),
    .Y(_4293_));
 sg13g2_buf_1 _4792_ (.A(_4293_),
    .X(_4294_));
 sg13g2_nand2_1 _4793_ (.Y(_4295_),
    .A(_4280_),
    .B(_4292_));
 sg13g2_inv_1 _4794_ (.Y(_4296_),
    .A(_4295_));
 sg13g2_nand2_1 _4795_ (.Y(_4297_),
    .A(_4296_),
    .B(_4287_));
 sg13g2_buf_1 _4796_ (.A(_4297_),
    .X(_4298_));
 sg13g2_buf_8 _4797_ (.A(\vgademo.a_scrolly[8] ),
    .X(_4299_));
 sg13g2_buf_8 _4798_ (.A(\vgademo.a_scrolly[9] ),
    .X(_4300_));
 sg13g2_inv_4 _4799_ (.A(_4300_),
    .Y(_4301_));
 sg13g2_nor2_1 _4800_ (.A(_4299_),
    .B(_4301_),
    .Y(_4302_));
 sg13g2_buf_8 _4801_ (.A(\vgademo.a_scrolly[4] ),
    .X(_4303_));
 sg13g2_buf_2 _4802_ (.A(\vgademo.a_scrolly[5] ),
    .X(_4304_));
 sg13g2_nor2_1 _4803_ (.A(_4303_),
    .B(_4304_),
    .Y(_4305_));
 sg13g2_buf_2 _4804_ (.A(_4305_),
    .X(_4306_));
 sg13g2_buf_8 _4805_ (.A(\vgademo.a_scrolly[7] ),
    .X(_4307_));
 sg13g2_buf_8 _4806_ (.A(\vgademo.a_scrolly[6] ),
    .X(_4308_));
 sg13g2_nor2_1 _4807_ (.A(_4307_),
    .B(_4308_),
    .Y(_4309_));
 sg13g2_buf_2 _4808_ (.A(_4309_),
    .X(_4310_));
 sg13g2_nand3_1 _4809_ (.B(_4306_),
    .C(_4310_),
    .A(_4302_),
    .Y(_4311_));
 sg13g2_buf_2 _4810_ (.A(\vgademo.a_scrolly[11] ),
    .X(_4312_));
 sg13g2_buf_2 _4811_ (.A(\vgademo.a_scrolly[10] ),
    .X(_4313_));
 sg13g2_nand3_1 _4812_ (.B(_4313_),
    .C(_4300_),
    .A(_4312_),
    .Y(_4314_));
 sg13g2_inv_1 _4813_ (.Y(_4315_),
    .A(_4314_));
 sg13g2_nand2_1 _4814_ (.Y(_4316_),
    .A(_4311_),
    .B(_4315_));
 sg13g2_buf_2 _4815_ (.A(\vgademo.a_scrolly[12] ),
    .X(_4317_));
 sg13g2_buf_2 _4816_ (.A(\vgademo.a_scrolly[13] ),
    .X(_4318_));
 sg13g2_nor2_2 _4817_ (.A(_4317_),
    .B(_4318_),
    .Y(_4319_));
 sg13g2_nand2_1 _4818_ (.Y(_4320_),
    .A(_4316_),
    .B(_4319_));
 sg13g2_nor2_1 _4819_ (.A(_4307_),
    .B(_4299_),
    .Y(_4321_));
 sg13g2_nor2b_1 _4820_ (.A(_4314_),
    .B_N(_4321_),
    .Y(_4322_));
 sg13g2_inv_2 _4821_ (.Y(_4323_),
    .A(_4303_));
 sg13g2_buf_2 _4822_ (.A(\vgademo.a_scrolly[3] ),
    .X(_4324_));
 sg13g2_nand2_1 _4823_ (.Y(_4325_),
    .A(_4323_),
    .B(_4324_));
 sg13g2_nor2_1 _4824_ (.A(_4308_),
    .B(_4304_),
    .Y(_4326_));
 sg13g2_inv_1 _4825_ (.Y(_4327_),
    .A(_4326_));
 sg13g2_nor2_1 _4826_ (.A(_4325_),
    .B(_4327_),
    .Y(_4328_));
 sg13g2_nand2_1 _4827_ (.Y(_4329_),
    .A(_4322_),
    .B(_4328_));
 sg13g2_nor2b_1 _4828_ (.A(_4320_),
    .B_N(_4329_),
    .Y(_4330_));
 sg13g2_buf_2 _4829_ (.A(_4330_),
    .X(_4331_));
 sg13g2_buf_8 _4830_ (.A(_4303_),
    .X(_4332_));
 sg13g2_nand2_2 _4831_ (.Y(_4333_),
    .A(_4332_),
    .B(_4324_));
 sg13g2_nor2b_2 _4832_ (.A(_4333_),
    .B_N(_4304_),
    .Y(_4334_));
 sg13g2_inv_2 _4833_ (.Y(_4335_),
    .A(_4312_));
 sg13g2_nor2b_1 _4834_ (.A(_4334_),
    .B_N(_4335_),
    .Y(_4336_));
 sg13g2_inv_8 _4835_ (.Y(_4337_),
    .A(_4299_));
 sg13g2_nand2_1 _4836_ (.Y(_4338_),
    .A(_4301_),
    .B(net106));
 sg13g2_inv_4 _4837_ (.A(_4310_),
    .Y(_4339_));
 sg13g2_nor2_2 _4838_ (.A(_4338_),
    .B(_4339_),
    .Y(_4340_));
 sg13g2_inv_2 _4839_ (.Y(_4341_),
    .A(_4313_));
 sg13g2_nand2_1 _4840_ (.Y(_4342_),
    .A(_4317_),
    .B(_4318_));
 sg13g2_a21oi_1 _4841_ (.A1(_4335_),
    .A2(_4341_),
    .Y(_4343_),
    .B1(_4342_));
 sg13g2_inv_1 _4842_ (.Y(_4344_),
    .A(_4343_));
 sg13g2_a21oi_1 _4843_ (.A1(_4336_),
    .A2(_4340_),
    .Y(_4345_),
    .B1(_4344_));
 sg13g2_buf_8 _4844_ (.A(_4308_),
    .X(_4346_));
 sg13g2_inv_8 _4845_ (.Y(_4347_),
    .A(net105));
 sg13g2_buf_8 _4846_ (.A(_4307_),
    .X(_4348_));
 sg13g2_nand2_1 _4847_ (.Y(_4349_),
    .A(_4347_),
    .B(net104));
 sg13g2_nor2_1 _4848_ (.A(_4349_),
    .B(_4338_),
    .Y(_4350_));
 sg13g2_nand2_1 _4849_ (.Y(_4351_),
    .A(_4350_),
    .B(_4334_));
 sg13g2_inv_1 _4850_ (.Y(_4352_),
    .A(_4342_));
 sg13g2_nor2_1 _4851_ (.A(_4300_),
    .B(_4299_),
    .Y(_4353_));
 sg13g2_nand2_1 _4852_ (.Y(_4354_),
    .A(_4307_),
    .B(net105));
 sg13g2_nand2_1 _4853_ (.Y(_4355_),
    .A(_4353_),
    .B(_4354_));
 sg13g2_nor2_1 _4854_ (.A(_4352_),
    .B(_4355_),
    .Y(_4356_));
 sg13g2_nand2_1 _4855_ (.Y(_4357_),
    .A(_4351_),
    .B(_4356_));
 sg13g2_nand2_1 _4856_ (.Y(_4358_),
    .A(_4312_),
    .B(_4313_));
 sg13g2_inv_2 _4857_ (.Y(_4359_),
    .A(_4317_));
 sg13g2_inv_1 _4858_ (.Y(_4360_),
    .A(_4318_));
 sg13g2_a21oi_1 _4859_ (.A1(_4358_),
    .A2(_4359_),
    .Y(_4361_),
    .B1(_4360_));
 sg13g2_nand2_1 _4860_ (.Y(_4362_),
    .A(_4357_),
    .B(_4361_));
 sg13g2_nor2_1 _4861_ (.A(_4345_),
    .B(_4362_),
    .Y(_4363_));
 sg13g2_inv_1 _4862_ (.Y(_4364_),
    .A(_0081_));
 sg13g2_inv_4 _4863_ (.A(_4307_),
    .Y(_4365_));
 sg13g2_nor2_1 _4864_ (.A(_4308_),
    .B(_4365_),
    .Y(_4366_));
 sg13g2_nand2_1 _4865_ (.Y(_4367_),
    .A(_4366_),
    .B(_4306_));
 sg13g2_nor2_1 _4866_ (.A(_0014_),
    .B(_4301_),
    .Y(_4368_));
 sg13g2_nand2_1 _4867_ (.Y(_4369_),
    .A(_4367_),
    .B(_4368_));
 sg13g2_nand2_1 _4868_ (.Y(_4370_),
    .A(_4300_),
    .B(_4299_));
 sg13g2_inv_1 _4869_ (.Y(_4371_),
    .A(_4370_));
 sg13g2_nand2_1 _4870_ (.Y(_4372_),
    .A(_4319_),
    .B(_4335_));
 sg13g2_nor2_1 _4871_ (.A(_4371_),
    .B(_4372_),
    .Y(_4373_));
 sg13g2_nand2_1 _4872_ (.Y(_4374_),
    .A(_4369_),
    .B(_4373_));
 sg13g2_nand3_1 _4873_ (.B(_4335_),
    .C(_4341_),
    .A(_4319_),
    .Y(_4375_));
 sg13g2_buf_1 _4874_ (.A(_4375_),
    .X(_4376_));
 sg13g2_nand2_1 _4875_ (.Y(_4377_),
    .A(_4374_),
    .B(_4376_));
 sg13g2_inv_1 _4876_ (.Y(_4378_),
    .A(_0015_));
 sg13g2_nor3_2 _4877_ (.A(_4317_),
    .B(_4312_),
    .C(_4378_),
    .Y(_4379_));
 sg13g2_nand2_1 _4878_ (.Y(_4380_),
    .A(_4313_),
    .B(_4300_));
 sg13g2_inv_1 _4879_ (.Y(_4381_),
    .A(_4380_));
 sg13g2_buf_1 _4880_ (.A(_4299_),
    .X(_4382_));
 sg13g2_nor2_1 _4881_ (.A(net103),
    .B(_4365_),
    .Y(_4383_));
 sg13g2_nand4_1 _4882_ (.B(_4379_),
    .C(_4381_),
    .A(_4328_),
    .Y(_4384_),
    .D(_4383_));
 sg13g2_nand2_2 _4883_ (.Y(_4385_),
    .A(_4377_),
    .B(_4384_));
 sg13g2_inv_4 _4884_ (.A(_4385_),
    .Y(_4386_));
 sg13g2_nor2_1 _4885_ (.A(_4364_),
    .B(_4386_),
    .Y(_4387_));
 sg13g2_o21ai_1 _4886_ (.B1(_4387_),
    .Y(_4388_),
    .A1(_4331_),
    .A2(_4363_));
 sg13g2_buf_1 _4887_ (.A(\vgademo.bayer_j[0] ),
    .X(_4389_));
 sg13g2_inv_1 _4888_ (.Y(_4390_),
    .A(_4389_));
 sg13g2_nand2b_1 _4889_ (.Y(_4391_),
    .B(_4390_),
    .A_N(_4388_));
 sg13g2_nand2_1 _4890_ (.Y(_4392_),
    .A(_4388_),
    .B(_4389_));
 sg13g2_nand2_1 _4891_ (.Y(_4393_),
    .A(_4391_),
    .B(_4392_));
 sg13g2_xnor2_1 _4892_ (.Y(_4394_),
    .A(_0077_),
    .B(_4393_));
 sg13g2_inv_1 _4893_ (.Y(_4395_),
    .A(_4394_));
 sg13g2_nor2_1 _4894_ (.A(_4298_),
    .B(_4395_),
    .Y(_4396_));
 sg13g2_a21o_1 _4895_ (.A2(_4294_),
    .A1(\vgademo.plane_dx_div.d[16] ),
    .B1(_4396_),
    .X(_0013_));
 sg13g2_nand2_1 _4896_ (.Y(_4397_),
    .A(_4281_),
    .B(net124));
 sg13g2_nor2_1 _4897_ (.A(_4286_),
    .B(_4397_),
    .Y(_4398_));
 sg13g2_inv_1 _4898_ (.Y(_4399_),
    .A(\vgademo.h_count[8] ));
 sg13g2_nor3_1 _4899_ (.A(_4289_),
    .B(_4288_),
    .C(_4399_),
    .Y(_4400_));
 sg13g2_nand3_1 _4900_ (.B(_4398_),
    .C(_4400_),
    .A(_4280_),
    .Y(_4401_));
 sg13g2_buf_1 _4901_ (.A(_4401_),
    .X(_4402_));
 sg13g2_inv_1 _4902_ (.Y(_4403_),
    .A(_4402_));
 sg13g2_buf_1 _4903_ (.A(_4403_),
    .X(_4404_));
 sg13g2_nor2_1 _4904_ (.A(net127),
    .B(net73),
    .Y(_0000_));
 sg13g2_xor2_1 _4905_ (.B(net126),
    .A(_4275_),
    .X(_0002_));
 sg13g2_buf_1 _4906_ (.A(_0051_),
    .X(_4405_));
 sg13g2_nand2_1 _4907_ (.Y(_4406_),
    .A(net127),
    .B(net126));
 sg13g2_xnor2_1 _4908_ (.Y(_4407_),
    .A(_4405_),
    .B(_4406_));
 sg13g2_nor2_1 _4909_ (.A(_4407_),
    .B(net73),
    .Y(_0003_));
 sg13g2_inv_1 _4910_ (.Y(_4408_),
    .A(_0052_));
 sg13g2_nor2_1 _4911_ (.A(_4279_),
    .B(_4406_),
    .Y(_4409_));
 sg13g2_xnor2_1 _4912_ (.Y(_4410_),
    .A(_4408_),
    .B(_4409_));
 sg13g2_nor2_1 _4913_ (.A(_4410_),
    .B(net73),
    .Y(_0004_));
 sg13g2_buf_1 _4914_ (.A(_0053_),
    .X(_4411_));
 sg13g2_inv_1 _4915_ (.Y(_4412_),
    .A(_4411_));
 sg13g2_nand2_1 _4916_ (.Y(_4413_),
    .A(_4409_),
    .B(net125));
 sg13g2_inv_1 _4917_ (.Y(_4414_),
    .A(_4413_));
 sg13g2_nor2_1 _4918_ (.A(_4412_),
    .B(_4414_),
    .Y(_4415_));
 sg13g2_nor2_1 _4919_ (.A(_4411_),
    .B(_4413_),
    .Y(_4416_));
 sg13g2_nor3_1 _4920_ (.A(_4415_),
    .B(_4416_),
    .C(net73),
    .Y(_0005_));
 sg13g2_inv_1 _4921_ (.Y(_4417_),
    .A(net123));
 sg13g2_nor3_1 _4922_ (.A(_4417_),
    .B(_0054_),
    .C(_4413_),
    .Y(_4418_));
 sg13g2_inv_1 _4923_ (.Y(_4419_),
    .A(_0054_));
 sg13g2_a21oi_1 _4924_ (.A1(_4414_),
    .A2(net123),
    .Y(_4420_),
    .B1(_4419_));
 sg13g2_nor3_1 _4925_ (.A(_4418_),
    .B(_4420_),
    .C(net73),
    .Y(_0006_));
 sg13g2_buf_1 _4926_ (.A(_0055_),
    .X(_4421_));
 sg13g2_nor2_1 _4927_ (.A(_4286_),
    .B(_4413_),
    .Y(_4422_));
 sg13g2_inv_1 _4928_ (.Y(_4423_),
    .A(_4422_));
 sg13g2_nand3_1 _4929_ (.B(_4398_),
    .C(_4400_),
    .A(_4280_),
    .Y(_4424_));
 sg13g2_buf_1 _4930_ (.A(_4424_),
    .X(_4425_));
 sg13g2_o21ai_1 _4931_ (.B1(_4425_),
    .Y(_4426_),
    .A1(_4421_),
    .A2(_4423_));
 sg13g2_a21oi_1 _4932_ (.A1(_4421_),
    .A2(_4423_),
    .Y(_0007_),
    .B1(_4426_));
 sg13g2_inv_1 _4933_ (.Y(_4427_),
    .A(_0056_));
 sg13g2_inv_2 _4934_ (.Y(_4428_),
    .A(net124));
 sg13g2_nor2_1 _4935_ (.A(_4428_),
    .B(_4423_),
    .Y(_4429_));
 sg13g2_nor2_1 _4936_ (.A(_4289_),
    .B(_4288_),
    .Y(_4430_));
 sg13g2_nand4_1 _4937_ (.B(\vgademo.h_count[8] ),
    .C(_4398_),
    .A(_4280_),
    .Y(_4431_),
    .D(_4430_));
 sg13g2_buf_1 _4938_ (.A(_4431_),
    .X(_4432_));
 sg13g2_o21ai_1 _4939_ (.B1(_4432_),
    .Y(_4433_),
    .A1(_4427_),
    .A2(_4429_));
 sg13g2_a21oi_1 _4940_ (.A1(_4427_),
    .A2(_4429_),
    .Y(_0008_),
    .B1(_4433_));
 sg13g2_inv_2 _4941_ (.Y(_4434_),
    .A(_0079_));
 sg13g2_nor2_1 _4942_ (.A(_4397_),
    .B(_4423_),
    .Y(_4435_));
 sg13g2_o21ai_1 _4943_ (.B1(_4432_),
    .Y(_4436_),
    .A1(_4434_),
    .A2(_4435_));
 sg13g2_a21oi_1 _4944_ (.A1(_4434_),
    .A2(_4435_),
    .Y(_0009_),
    .B1(_4436_));
 sg13g2_inv_1 _4945_ (.Y(_4437_),
    .A(_0057_));
 sg13g2_nand2_1 _4946_ (.Y(_4438_),
    .A(_4281_),
    .B(\vgademo.h_count[8] ));
 sg13g2_inv_1 _4947_ (.Y(_4439_),
    .A(_4429_));
 sg13g2_nor2_1 _4948_ (.A(_4438_),
    .B(_4439_),
    .Y(_4440_));
 sg13g2_o21ai_1 _4949_ (.B1(_4425_),
    .Y(_4441_),
    .A1(_4437_),
    .A2(_4440_));
 sg13g2_a21oi_1 _4950_ (.A1(_4437_),
    .A2(_4440_),
    .Y(_0010_),
    .B1(_4441_));
 sg13g2_inv_1 _4951_ (.Y(_4442_),
    .A(_4288_));
 sg13g2_inv_1 _4952_ (.Y(_4443_),
    .A(_4289_));
 sg13g2_nor3_1 _4953_ (.A(_4443_),
    .B(_4438_),
    .C(_4439_),
    .Y(_4444_));
 sg13g2_o21ai_1 _4954_ (.B1(_4432_),
    .Y(_4445_),
    .A1(_4442_),
    .A2(_4444_));
 sg13g2_a21oi_1 _4955_ (.A1(_4442_),
    .A2(_4444_),
    .Y(_0001_),
    .B1(_4445_));
 sg13g2_buf_1 _4956_ (.A(\vgademo.v_count[4] ),
    .X(_4446_));
 sg13g2_buf_2 _4957_ (.A(\vgademo.v_count[9] ),
    .X(_4447_));
 sg13g2_buf_2 _4958_ (.A(\vgademo.v_count[5] ),
    .X(_4448_));
 sg13g2_inv_1 _4959_ (.Y(_4449_),
    .A(_4448_));
 sg13g2_buf_1 _4960_ (.A(\vgademo.v_count[8] ),
    .X(_4450_));
 sg13g2_inv_1 _4961_ (.Y(_4451_),
    .A(_4450_));
 sg13g2_nor4_1 _4962_ (.A(net122),
    .B(_4447_),
    .C(_4449_),
    .D(_4451_),
    .Y(_4452_));
 sg13g2_buf_1 _4963_ (.A(\vgademo.v_count[7] ),
    .X(_4453_));
 sg13g2_buf_2 _4964_ (.A(\vgademo.v_count[6] ),
    .X(_4454_));
 sg13g2_buf_1 _4965_ (.A(\vgademo.v_count[2] ),
    .X(_4455_));
 sg13g2_buf_1 _4966_ (.A(\vgademo.bayer_j[1] ),
    .X(_4456_));
 sg13g2_inv_1 _4967_ (.Y(_4457_),
    .A(_4456_));
 sg13g2_buf_1 _4968_ (.A(\vgademo.v_count[3] ),
    .X(_4458_));
 sg13g2_inv_1 _4969_ (.Y(_4459_),
    .A(_4458_));
 sg13g2_nor3_1 _4970_ (.A(_4455_),
    .B(_4457_),
    .C(_4459_),
    .Y(_4460_));
 sg13g2_nand4_1 _4971_ (.B(net121),
    .C(_4454_),
    .A(_4452_),
    .Y(_0012_),
    .D(_4460_));
 sg13g2_buf_1 _4972_ (.A(\vgademo.h_count[10] ),
    .X(_4461_));
 sg13g2_inv_1 _4973_ (.Y(_4462_),
    .A(_4461_));
 sg13g2_nand2_1 _4974_ (.Y(_4463_),
    .A(net125),
    .B(net123));
 sg13g2_nor2_1 _4975_ (.A(net126),
    .B(_4278_),
    .Y(_4464_));
 sg13g2_nor2_1 _4976_ (.A(_4285_),
    .B(net124),
    .Y(_4465_));
 sg13g2_o21ai_1 _4977_ (.B1(_4465_),
    .Y(_4466_),
    .A1(_4463_),
    .A2(_4464_));
 sg13g2_inv_1 _4978_ (.Y(_4467_),
    .A(_4438_));
 sg13g2_a21oi_1 _4979_ (.A1(_4466_),
    .A2(_4467_),
    .Y(_4468_),
    .B1(_4289_));
 sg13g2_inv_1 _4980_ (.Y(_4469_),
    .A(_4406_));
 sg13g2_nand2_1 _4981_ (.Y(_4470_),
    .A(_4469_),
    .B(_4279_));
 sg13g2_nor2_1 _4982_ (.A(net125),
    .B(net123),
    .Y(_4471_));
 sg13g2_nand3_1 _4983_ (.B(_4405_),
    .C(_4471_),
    .A(_4470_),
    .Y(_4472_));
 sg13g2_nor3_1 _4984_ (.A(_4282_),
    .B(_4462_),
    .C(_4291_),
    .Y(_4473_));
 sg13g2_nand4_1 _4985_ (.B(_4285_),
    .C(net124),
    .A(_4472_),
    .Y(_4474_),
    .D(_4473_));
 sg13g2_o21ai_1 _4986_ (.B1(_4461_),
    .Y(_4475_),
    .A1(_4289_),
    .A2(_4434_));
 sg13g2_inv_1 _4987_ (.Y(_4476_),
    .A(_4285_));
 sg13g2_nor4_1 _4988_ (.A(_4277_),
    .B(_4278_),
    .C(_4284_),
    .D(_4476_),
    .Y(_4477_));
 sg13g2_nor2_1 _4989_ (.A(_4397_),
    .B(_4406_),
    .Y(_4478_));
 sg13g2_nand3_1 _4990_ (.B(_4292_),
    .C(_4478_),
    .A(_4477_),
    .Y(_4479_));
 sg13g2_nand3_1 _4991_ (.B(_4475_),
    .C(_4479_),
    .A(_4474_),
    .Y(_4480_));
 sg13g2_o21ai_1 _4992_ (.B1(_4480_),
    .Y(_0011_),
    .A1(_4462_),
    .A2(_4468_));
 sg13g2_nand2_1 _4993_ (.Y(_4481_),
    .A(_4451_),
    .B(_4447_));
 sg13g2_nor3_1 _4994_ (.A(net121),
    .B(_4454_),
    .C(_4481_),
    .Y(_4482_));
 sg13g2_nor2_1 _4995_ (.A(_4456_),
    .B(_4389_),
    .Y(_4483_));
 sg13g2_nand2_1 _4996_ (.Y(_4484_),
    .A(_4458_),
    .B(_4455_));
 sg13g2_inv_1 _4997_ (.Y(_4485_),
    .A(_4484_));
 sg13g2_nor2_1 _4998_ (.A(_4448_),
    .B(net122),
    .Y(_4486_));
 sg13g2_nand4_1 _4999_ (.B(_4483_),
    .C(_4485_),
    .A(_4482_),
    .Y(_4487_),
    .D(_4486_));
 sg13g2_nor2_1 _5000_ (.A(_4425_),
    .B(_4487_),
    .Y(_4488_));
 sg13g2_buf_2 _5001_ (.A(_4488_),
    .X(_4489_));
 sg13g2_inv_1 _5002_ (.Y(_4490_),
    .A(_4489_));
 sg13g2_inv_1 _5003_ (.Y(_4491_),
    .A(\vgademo.a_sin[6] ));
 sg13g2_nor2_1 _5004_ (.A(\vgademo.a_cos[0] ),
    .B(_4491_),
    .Y(_4492_));
 sg13g2_inv_1 _5005_ (.Y(_4493_),
    .A(_4492_));
 sg13g2_o21ai_1 _5006_ (.B1(\vgademo.a_cos[0] ),
    .Y(_4494_),
    .A1(_4491_),
    .A2(_4490_));
 sg13g2_o21ai_1 _5007_ (.B1(_4494_),
    .Y(_0112_),
    .A1(_4490_),
    .A2(_4493_));
 sg13g2_buf_1 _5008_ (.A(\vgademo.a_cos[10] ),
    .X(_4495_));
 sg13g2_inv_1 _5009_ (.Y(_4496_),
    .A(_4495_));
 sg13g2_buf_1 _5010_ (.A(\vgademo.a_sin[14] ),
    .X(_4497_));
 sg13g2_inv_2 _5011_ (.Y(_4498_),
    .A(_4497_));
 sg13g2_nor2_1 _5012_ (.A(_4495_),
    .B(_4498_),
    .Y(_4499_));
 sg13g2_buf_1 _5013_ (.A(_4497_),
    .X(_4500_));
 sg13g2_nor2_1 _5014_ (.A(net102),
    .B(_4496_),
    .Y(_4501_));
 sg13g2_nor2_1 _5015_ (.A(_4499_),
    .B(_4501_),
    .Y(_4502_));
 sg13g2_buf_2 _5016_ (.A(\vgademo.a_cos[8] ),
    .X(_4503_));
 sg13g2_inv_1 _5017_ (.Y(_4504_),
    .A(_4503_));
 sg13g2_buf_1 _5018_ (.A(\vgademo.a_sin[13] ),
    .X(_4505_));
 sg13g2_inv_1 _5019_ (.Y(_4506_),
    .A(_4505_));
 sg13g2_buf_2 _5020_ (.A(\vgademo.a_cos[7] ),
    .X(_4507_));
 sg13g2_nand2_1 _5021_ (.Y(_4508_),
    .A(_4506_),
    .B(_4507_));
 sg13g2_inv_1 _5022_ (.Y(_4509_),
    .A(_4508_));
 sg13g2_a21oi_1 _5023_ (.A1(_4503_),
    .A2(_4498_),
    .Y(_4510_),
    .B1(_4509_));
 sg13g2_buf_1 _5024_ (.A(\vgademo.a_sin[12] ),
    .X(_4511_));
 sg13g2_inv_1 _5025_ (.Y(_4512_),
    .A(_4511_));
 sg13g2_nor2_1 _5026_ (.A(\vgademo.a_cos[6] ),
    .B(_4512_),
    .Y(_4513_));
 sg13g2_buf_1 _5027_ (.A(\vgademo.a_sin[9] ),
    .X(_4514_));
 sg13g2_inv_1 _5028_ (.Y(_4515_),
    .A(\vgademo.a_cos[3] ));
 sg13g2_nor2_1 _5029_ (.A(_4514_),
    .B(_4515_),
    .Y(_4516_));
 sg13g2_inv_1 _5030_ (.Y(_4517_),
    .A(_4514_));
 sg13g2_nor2_1 _5031_ (.A(\vgademo.a_cos[3] ),
    .B(_4517_),
    .Y(_4518_));
 sg13g2_buf_1 _5032_ (.A(\vgademo.a_sin[8] ),
    .X(_4519_));
 sg13g2_inv_1 _5033_ (.Y(_4520_),
    .A(_4519_));
 sg13g2_buf_1 _5034_ (.A(\vgademo.a_sin[7] ),
    .X(_4521_));
 sg13g2_inv_1 _5035_ (.Y(_4522_),
    .A(_4521_));
 sg13g2_xnor2_1 _5036_ (.Y(_4523_),
    .A(_4521_),
    .B(\vgademo.a_cos[1] ));
 sg13g2_nand2_1 _5037_ (.Y(_4524_),
    .A(_4523_),
    .B(_4493_));
 sg13g2_inv_1 _5038_ (.Y(_4525_),
    .A(_4524_));
 sg13g2_a21oi_1 _5039_ (.A1(_4522_),
    .A2(\vgademo.a_cos[1] ),
    .Y(_4526_),
    .B1(_4525_));
 sg13g2_xnor2_1 _5040_ (.Y(_4527_),
    .A(_4519_),
    .B(\vgademo.a_cos[2] ));
 sg13g2_nand2b_1 _5041_ (.Y(_4528_),
    .B(_4527_),
    .A_N(_4526_));
 sg13g2_inv_1 _5042_ (.Y(_4529_),
    .A(_4528_));
 sg13g2_a21oi_1 _5043_ (.A1(_4520_),
    .A2(\vgademo.a_cos[2] ),
    .Y(_4530_),
    .B1(_4529_));
 sg13g2_nor2_1 _5044_ (.A(_4518_),
    .B(_4530_),
    .Y(_4531_));
 sg13g2_nor2_1 _5045_ (.A(_4516_),
    .B(_4531_),
    .Y(_4532_));
 sg13g2_buf_1 _5046_ (.A(\vgademo.a_cos[4] ),
    .X(_4533_));
 sg13g2_inv_1 _5047_ (.Y(_4534_),
    .A(_4533_));
 sg13g2_nor2_1 _5048_ (.A(\vgademo.a_sin[10] ),
    .B(_4534_),
    .Y(_4535_));
 sg13g2_inv_1 _5049_ (.Y(_4536_),
    .A(_4535_));
 sg13g2_inv_1 _5050_ (.Y(_4537_),
    .A(\vgademo.a_sin[10] ));
 sg13g2_nor2_1 _5051_ (.A(_4533_),
    .B(_4537_),
    .Y(_4538_));
 sg13g2_a21oi_1 _5052_ (.A1(_4532_),
    .A2(_4536_),
    .Y(_4539_),
    .B1(_4538_));
 sg13g2_buf_1 _5053_ (.A(\vgademo.a_cos[5] ),
    .X(_4540_));
 sg13g2_buf_1 _5054_ (.A(\vgademo.a_sin[11] ),
    .X(_4541_));
 sg13g2_inv_1 _5055_ (.Y(_4542_),
    .A(_4541_));
 sg13g2_nor2_1 _5056_ (.A(_4540_),
    .B(_4542_),
    .Y(_4543_));
 sg13g2_inv_1 _5057_ (.Y(_4544_),
    .A(_4543_));
 sg13g2_inv_1 _5058_ (.Y(_4545_),
    .A(_4540_));
 sg13g2_nor2_1 _5059_ (.A(_4541_),
    .B(_4545_),
    .Y(_4546_));
 sg13g2_a21oi_1 _5060_ (.A1(_4539_),
    .A2(_4544_),
    .Y(_4547_),
    .B1(_4546_));
 sg13g2_inv_1 _5061_ (.Y(_4548_),
    .A(\vgademo.a_cos[6] ));
 sg13g2_nor2_1 _5062_ (.A(_4511_),
    .B(_4548_),
    .Y(_4549_));
 sg13g2_inv_1 _5063_ (.Y(_4550_),
    .A(_4549_));
 sg13g2_o21ai_1 _5064_ (.B1(_4550_),
    .Y(_4551_),
    .A1(_4513_),
    .A2(_4547_));
 sg13g2_nor2_1 _5065_ (.A(_4507_),
    .B(_4506_),
    .Y(_4552_));
 sg13g2_nor2_1 _5066_ (.A(_4552_),
    .B(_4509_),
    .Y(_4553_));
 sg13g2_nand2_1 _5067_ (.Y(_4554_),
    .A(_4551_),
    .B(_4553_));
 sg13g2_a22oi_1 _5068_ (.Y(_4555_),
    .B1(_4510_),
    .B2(_4554_),
    .A2(net102),
    .A1(_4504_));
 sg13g2_buf_1 _5069_ (.A(\vgademo.a_cos[9] ),
    .X(_4556_));
 sg13g2_xnor2_1 _5070_ (.Y(_4557_),
    .A(_4556_),
    .B(_4497_));
 sg13g2_inv_1 _5071_ (.Y(_4558_),
    .A(_4556_));
 sg13g2_nor2_1 _5072_ (.A(net102),
    .B(_4558_),
    .Y(_4559_));
 sg13g2_a21oi_2 _5073_ (.B1(_4559_),
    .Y(_4560_),
    .A2(_4557_),
    .A1(_4555_));
 sg13g2_xnor2_1 _5074_ (.Y(_4561_),
    .A(_4502_),
    .B(_4560_));
 sg13g2_nor2_1 _5075_ (.A(_4490_),
    .B(_4561_),
    .Y(_4562_));
 sg13g2_a21oi_1 _5076_ (.A1(_4496_),
    .A2(_4490_),
    .Y(_0113_),
    .B1(_4562_));
 sg13g2_buf_2 _5077_ (.A(\vgademo.a_cos[11] ),
    .X(_4563_));
 sg13g2_xnor2_1 _5078_ (.Y(_4564_),
    .A(_4563_),
    .B(net102));
 sg13g2_inv_1 _5079_ (.Y(_4565_),
    .A(_4501_));
 sg13g2_o21ai_1 _5080_ (.B1(_4565_),
    .Y(_4566_),
    .A1(_4499_),
    .A2(_4560_));
 sg13g2_xor2_1 _5081_ (.B(_4566_),
    .A(_4564_),
    .X(_4567_));
 sg13g2_inv_1 _5082_ (.Y(_4568_),
    .A(_4567_));
 sg13g2_inv_1 _5083_ (.Y(_4569_),
    .A(net122));
 sg13g2_inv_1 _5084_ (.Y(_4570_),
    .A(_4483_));
 sg13g2_nor2_1 _5085_ (.A(_4448_),
    .B(_4570_),
    .Y(_4571_));
 sg13g2_nand4_1 _5086_ (.B(_4569_),
    .C(_4485_),
    .A(_4482_),
    .Y(_4572_),
    .D(_4571_));
 sg13g2_nor2_1 _5087_ (.A(_4572_),
    .B(_4432_),
    .Y(_4573_));
 sg13g2_buf_1 _5088_ (.A(_4573_),
    .X(_4574_));
 sg13g2_buf_1 _5089_ (.A(_4574_),
    .X(_4575_));
 sg13g2_buf_1 _5090_ (.A(_4489_),
    .X(_4576_));
 sg13g2_nor2_1 _5091_ (.A(_4563_),
    .B(net71),
    .Y(_4577_));
 sg13g2_a21oi_1 _5092_ (.A1(_4568_),
    .A2(net72),
    .Y(_0114_),
    .B1(_4577_));
 sg13g2_buf_2 _5093_ (.A(\vgademo.a_cos[12] ),
    .X(_4578_));
 sg13g2_xnor2_1 _5094_ (.Y(_0365_),
    .A(_4578_),
    .B(net102));
 sg13g2_xor2_1 _5095_ (.B(_4497_),
    .A(_4503_),
    .X(_0366_));
 sg13g2_nand2_1 _5096_ (.Y(_0367_),
    .A(_4502_),
    .B(_4564_));
 sg13g2_inv_1 _5097_ (.Y(_0368_),
    .A(_0367_));
 sg13g2_nand3b_1 _5098_ (.B(_0368_),
    .C(_4557_),
    .Y(_0369_),
    .A_N(_0366_));
 sg13g2_nor2_1 _5099_ (.A(_4549_),
    .B(_4513_),
    .Y(_0370_));
 sg13g2_nor2b_1 _5100_ (.A(_4547_),
    .B_N(_0370_),
    .Y(_0371_));
 sg13g2_a21oi_1 _5101_ (.A1(_4550_),
    .A2(_4508_),
    .Y(_0372_),
    .B1(_4552_));
 sg13g2_a21oi_1 _5102_ (.A1(_0371_),
    .A2(_4553_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_a21oi_1 _5103_ (.A1(_4504_),
    .A2(_4558_),
    .Y(_0374_),
    .B1(net102));
 sg13g2_inv_1 _5104_ (.Y(_0375_),
    .A(_4563_));
 sg13g2_nor2_1 _5105_ (.A(_4500_),
    .B(_0375_),
    .Y(_0376_));
 sg13g2_a221oi_1 _5106_ (.B2(_0374_),
    .C1(_0376_),
    .B1(_0368_),
    .A1(_4495_),
    .Y(_0377_),
    .A2(_4498_));
 sg13g2_o21ai_1 _5107_ (.B1(_0377_),
    .Y(_0378_),
    .A1(_0369_),
    .A2(_0373_));
 sg13g2_xnor2_1 _5108_ (.Y(_0379_),
    .A(_0365_),
    .B(_0378_));
 sg13g2_nor2_1 _5109_ (.A(_4578_),
    .B(net71),
    .Y(_0380_));
 sg13g2_a21oi_1 _5110_ (.A1(_0379_),
    .A2(net72),
    .Y(_0115_),
    .B1(_0380_));
 sg13g2_buf_1 _5111_ (.A(\vgademo.a_cos[13] ),
    .X(_0381_));
 sg13g2_xnor2_1 _5112_ (.Y(_0382_),
    .A(_0381_),
    .B(net102));
 sg13g2_nand3_1 _5113_ (.B(_4564_),
    .C(_0365_),
    .A(_4566_),
    .Y(_0383_));
 sg13g2_o21ai_1 _5114_ (.B1(_4498_),
    .Y(_0384_),
    .A1(_4563_),
    .A2(_4578_));
 sg13g2_nand2_1 _5115_ (.Y(_0385_),
    .A(_0383_),
    .B(_0384_));
 sg13g2_xnor2_1 _5116_ (.Y(_0386_),
    .A(_0382_),
    .B(_0385_));
 sg13g2_inv_1 _5117_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_nor2_1 _5118_ (.A(_0086_),
    .B(net71),
    .Y(_0388_));
 sg13g2_a21oi_1 _5119_ (.A1(_0387_),
    .A2(net72),
    .Y(_0116_),
    .B1(_0388_));
 sg13g2_nand2_1 _5120_ (.Y(_0389_),
    .A(_0365_),
    .B(_0382_));
 sg13g2_nand2b_1 _5121_ (.Y(_0390_),
    .B(_0368_),
    .A_N(_0389_));
 sg13g2_inv_1 _5122_ (.Y(_0391_),
    .A(_4578_));
 sg13g2_inv_1 _5123_ (.Y(_0392_),
    .A(_0381_));
 sg13g2_a21oi_1 _5124_ (.A1(_0391_),
    .A2(_0392_),
    .Y(_0393_),
    .B1(_4500_));
 sg13g2_nor2_1 _5125_ (.A(_4501_),
    .B(_0376_),
    .Y(_0394_));
 sg13g2_nor2_1 _5126_ (.A(_0394_),
    .B(_0389_),
    .Y(_0395_));
 sg13g2_nor2_1 _5127_ (.A(_0393_),
    .B(_0395_),
    .Y(_0396_));
 sg13g2_o21ai_1 _5128_ (.B1(_0396_),
    .Y(_0397_),
    .A1(_0390_),
    .A2(_4560_));
 sg13g2_buf_1 _5129_ (.A(\vgademo.a_cos[14] ),
    .X(_0398_));
 sg13g2_xor2_1 _5130_ (.B(net102),
    .A(_0398_),
    .X(_0399_));
 sg13g2_nand2b_1 _5131_ (.Y(_0400_),
    .B(_0399_),
    .A_N(_0397_));
 sg13g2_nand2b_1 _5132_ (.Y(_0401_),
    .B(_0397_),
    .A_N(_0399_));
 sg13g2_nand2_1 _5133_ (.Y(_0402_),
    .A(_0400_),
    .B(_0401_));
 sg13g2_buf_1 _5134_ (.A(_0402_),
    .X(_0403_));
 sg13g2_nor2_1 _5135_ (.A(_0398_),
    .B(net71),
    .Y(_0404_));
 sg13g2_a21oi_1 _5136_ (.A1(_0403_),
    .A2(net72),
    .Y(_0117_),
    .B1(_0404_));
 sg13g2_inv_1 _5137_ (.Y(_0405_),
    .A(net121));
 sg13g2_inv_2 _5138_ (.Y(_0406_),
    .A(_4454_));
 sg13g2_nand3_1 _5139_ (.B(_0405_),
    .C(_0406_),
    .A(_4486_),
    .Y(_0407_));
 sg13g2_nor4_1 _5140_ (.A(_4481_),
    .B(_4570_),
    .C(_4484_),
    .D(_0407_),
    .Y(_0408_));
 sg13g2_nand2_1 _5141_ (.Y(_0409_),
    .A(_4403_),
    .B(_0408_));
 sg13g2_buf_2 _5142_ (.A(_0409_),
    .X(_0410_));
 sg13g2_buf_1 _5143_ (.A(_0410_),
    .X(_0411_));
 sg13g2_xnor2_1 _5144_ (.Y(_0412_),
    .A(_4493_),
    .B(_4523_));
 sg13g2_nand2_1 _5145_ (.Y(_0413_),
    .A(net64),
    .B(\vgademo.a_cos[1] ));
 sg13g2_o21ai_1 _5146_ (.B1(_0413_),
    .Y(_0118_),
    .A1(net64),
    .A2(_0412_));
 sg13g2_xor2_1 _5147_ (.B(_4526_),
    .A(_4527_),
    .X(_0414_));
 sg13g2_nor2_1 _5148_ (.A(\vgademo.a_cos[2] ),
    .B(net71),
    .Y(_0415_));
 sg13g2_a21oi_1 _5149_ (.A1(_0414_),
    .A2(net71),
    .Y(_0119_),
    .B1(_0415_));
 sg13g2_nor2_1 _5150_ (.A(_4516_),
    .B(_4518_),
    .Y(_0416_));
 sg13g2_xor2_1 _5151_ (.B(_4530_),
    .A(_0416_),
    .X(_0417_));
 sg13g2_nor2_1 _5152_ (.A(\vgademo.a_cos[3] ),
    .B(net71),
    .Y(_0418_));
 sg13g2_a21oi_1 _5153_ (.A1(_0417_),
    .A2(net72),
    .Y(_0120_),
    .B1(_0418_));
 sg13g2_nor2_1 _5154_ (.A(_4538_),
    .B(_4535_),
    .Y(_0419_));
 sg13g2_xor2_1 _5155_ (.B(_4532_),
    .A(_0419_),
    .X(_0420_));
 sg13g2_buf_1 _5156_ (.A(_4574_),
    .X(_0421_));
 sg13g2_nor2_1 _5157_ (.A(_4533_),
    .B(net70),
    .Y(_0422_));
 sg13g2_a21oi_1 _5158_ (.A1(_0420_),
    .A2(net72),
    .Y(_0121_),
    .B1(_0422_));
 sg13g2_nor2_1 _5159_ (.A(_4546_),
    .B(_4543_),
    .Y(_0423_));
 sg13g2_xnor2_1 _5160_ (.Y(_0424_),
    .A(_0423_),
    .B(_4539_));
 sg13g2_nor2_1 _5161_ (.A(_4540_),
    .B(net71),
    .Y(_0425_));
 sg13g2_a21oi_1 _5162_ (.A1(_0424_),
    .A2(net72),
    .Y(_0122_),
    .B1(_0425_));
 sg13g2_inv_1 _5163_ (.Y(_0426_),
    .A(_0410_));
 sg13g2_xnor2_1 _5164_ (.Y(_0427_),
    .A(_0370_),
    .B(_4547_));
 sg13g2_nand2_1 _5165_ (.Y(_0428_),
    .A(_0427_),
    .B(_0426_));
 sg13g2_o21ai_1 _5166_ (.B1(_0428_),
    .Y(_0123_),
    .A1(_4548_),
    .A2(_0426_));
 sg13g2_xor2_1 _5167_ (.B(_4551_),
    .A(_4553_),
    .X(_0429_));
 sg13g2_inv_1 _5168_ (.Y(_0430_),
    .A(_0429_));
 sg13g2_nor2_1 _5169_ (.A(_4507_),
    .B(_4576_),
    .Y(_0431_));
 sg13g2_a21oi_1 _5170_ (.A1(_0430_),
    .A2(_4575_),
    .Y(_0124_),
    .B1(_0431_));
 sg13g2_xor2_1 _5171_ (.B(_0373_),
    .A(_0366_),
    .X(_0432_));
 sg13g2_inv_1 _5172_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_nor2_1 _5173_ (.A(_4503_),
    .B(_4576_),
    .Y(_0434_));
 sg13g2_a21oi_1 _5174_ (.A1(_0433_),
    .A2(net72),
    .Y(_0125_),
    .B1(_0434_));
 sg13g2_xor2_1 _5175_ (.B(_4555_),
    .A(_4557_),
    .X(_0435_));
 sg13g2_inv_1 _5176_ (.Y(_0436_),
    .A(_0435_));
 sg13g2_buf_1 _5177_ (.A(_4489_),
    .X(_0437_));
 sg13g2_nor2_1 _5178_ (.A(_4556_),
    .B(net69),
    .Y(_0438_));
 sg13g2_a21oi_1 _5179_ (.A1(_0436_),
    .A2(_4575_),
    .Y(_0126_),
    .B1(_0438_));
 sg13g2_xnor2_1 _5180_ (.Y(_0127_),
    .A(\vgademo.a_sin[0] ),
    .B(_0428_));
 sg13g2_nor2_1 _5181_ (.A(_4537_),
    .B(net25),
    .Y(_0439_));
 sg13g2_inv_1 _5182_ (.Y(_0440_),
    .A(net25));
 sg13g2_nor2_1 _5183_ (.A(\vgademo.a_sin[10] ),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_nor2_1 _5184_ (.A(_0439_),
    .B(_0441_),
    .Y(_0442_));
 sg13g2_xnor2_1 _5185_ (.Y(_0443_),
    .A(_4514_),
    .B(net25));
 sg13g2_inv_1 _5186_ (.Y(_0444_),
    .A(_0443_));
 sg13g2_nor2_1 _5187_ (.A(_4520_),
    .B(net25),
    .Y(_0445_));
 sg13g2_nor2_1 _5188_ (.A(_4519_),
    .B(_0440_),
    .Y(_0446_));
 sg13g2_inv_1 _5189_ (.Y(_0447_),
    .A(\vgademo.a_sin[2] ));
 sg13g2_inv_1 _5190_ (.Y(_0448_),
    .A(\vgademo.a_sin[1] ));
 sg13g2_nor2_1 _5191_ (.A(_0448_),
    .B(_0430_),
    .Y(_0449_));
 sg13g2_nand2_1 _5192_ (.Y(_0450_),
    .A(_0427_),
    .B(\vgademo.a_sin[0] ));
 sg13g2_xnor2_1 _5193_ (.Y(_0451_),
    .A(_0448_),
    .B(_0429_));
 sg13g2_inv_1 _5194_ (.Y(_0452_),
    .A(_0451_));
 sg13g2_nor2_1 _5195_ (.A(_0450_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_xnor2_1 _5196_ (.Y(_0454_),
    .A(_0447_),
    .B(_0432_));
 sg13g2_o21ai_1 _5197_ (.B1(_0454_),
    .Y(_0455_),
    .A1(_0449_),
    .A2(_0453_));
 sg13g2_o21ai_1 _5198_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0447_),
    .A2(_0433_));
 sg13g2_inv_1 _5199_ (.Y(_0457_),
    .A(\vgademo.a_sin[3] ));
 sg13g2_nand2_1 _5200_ (.Y(_0458_),
    .A(_0436_),
    .B(_0457_));
 sg13g2_nor2_1 _5201_ (.A(_0457_),
    .B(_0436_),
    .Y(_0459_));
 sg13g2_a21oi_1 _5202_ (.A1(_0456_),
    .A2(_0458_),
    .Y(_0460_),
    .B1(_0459_));
 sg13g2_buf_1 _5203_ (.A(\vgademo.a_sin[4] ),
    .X(_0461_));
 sg13g2_nand2_1 _5204_ (.Y(_0462_),
    .A(_4561_),
    .B(_0461_));
 sg13g2_nor2_1 _5205_ (.A(_0461_),
    .B(_4561_),
    .Y(_0463_));
 sg13g2_a21oi_1 _5206_ (.A1(_0460_),
    .A2(_0462_),
    .Y(_0464_),
    .B1(_0463_));
 sg13g2_inv_1 _5207_ (.Y(_0465_),
    .A(\vgademo.a_sin[5] ));
 sg13g2_nand2_1 _5208_ (.Y(_0466_),
    .A(_4568_),
    .B(_0465_));
 sg13g2_nor2_1 _5209_ (.A(_0465_),
    .B(_4568_),
    .Y(_0467_));
 sg13g2_a21oi_1 _5210_ (.A1(_0464_),
    .A2(_0466_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_inv_1 _5211_ (.Y(_0469_),
    .A(_0468_));
 sg13g2_nand2_1 _5212_ (.Y(_0470_),
    .A(_0379_),
    .B(_4491_));
 sg13g2_nor2_1 _5213_ (.A(_4491_),
    .B(_0379_),
    .Y(_0471_));
 sg13g2_a21oi_1 _5214_ (.A1(_0469_),
    .A2(_0470_),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_inv_1 _5215_ (.Y(_0473_),
    .A(_0472_));
 sg13g2_nor2_1 _5216_ (.A(_4521_),
    .B(_0387_),
    .Y(_0474_));
 sg13g2_inv_1 _5217_ (.Y(_0475_),
    .A(_0474_));
 sg13g2_nor2_1 _5218_ (.A(_4522_),
    .B(_0386_),
    .Y(_0476_));
 sg13g2_a21oi_1 _5219_ (.A1(_0473_),
    .A2(_0475_),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_nor2_1 _5220_ (.A(_0446_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_nor2_1 _5221_ (.A(_0445_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_nor2_1 _5222_ (.A(_0444_),
    .B(_0479_),
    .Y(_0480_));
 sg13g2_a21oi_1 _5223_ (.A1(_4514_),
    .A2(_0440_),
    .Y(_0481_),
    .B1(_0480_));
 sg13g2_xor2_1 _5224_ (.B(_0481_),
    .A(_0442_),
    .X(_0482_));
 sg13g2_nor2_1 _5225_ (.A(\vgademo.a_sin[10] ),
    .B(net69),
    .Y(_0483_));
 sg13g2_a21oi_1 _5226_ (.A1(_0482_),
    .A2(net70),
    .Y(_0128_),
    .B1(_0483_));
 sg13g2_xnor2_1 _5227_ (.Y(_0484_),
    .A(_4541_),
    .B(net25));
 sg13g2_inv_1 _5228_ (.Y(_0485_),
    .A(_0439_));
 sg13g2_o21ai_1 _5229_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0441_),
    .A2(_0481_));
 sg13g2_xnor2_1 _5230_ (.Y(_0487_),
    .A(_0484_),
    .B(_0486_));
 sg13g2_nor2_1 _5231_ (.A(_4541_),
    .B(net69),
    .Y(_0488_));
 sg13g2_a21oi_1 _5232_ (.A1(_0487_),
    .A2(net70),
    .Y(_0129_),
    .B1(_0488_));
 sg13g2_xnor2_1 _5233_ (.Y(_0489_),
    .A(_4511_),
    .B(net25));
 sg13g2_nand2_1 _5234_ (.Y(_0490_),
    .A(_0440_),
    .B(_4541_));
 sg13g2_nand2_1 _5235_ (.Y(_0491_),
    .A(_0485_),
    .B(_0490_));
 sg13g2_nand3b_1 _5236_ (.B(_0442_),
    .C(_0484_),
    .Y(_0492_),
    .A_N(_0481_));
 sg13g2_nand2b_1 _5237_ (.Y(_0493_),
    .B(_0492_),
    .A_N(_0491_));
 sg13g2_xnor2_1 _5238_ (.Y(_0494_),
    .A(_0489_),
    .B(_0493_));
 sg13g2_nor2_1 _5239_ (.A(_4511_),
    .B(net69),
    .Y(_0495_));
 sg13g2_a21oi_1 _5240_ (.A1(_0494_),
    .A2(net70),
    .Y(_0130_),
    .B1(_0495_));
 sg13g2_xnor2_1 _5241_ (.Y(_0496_),
    .A(_4505_),
    .B(net25));
 sg13g2_nor2_1 _5242_ (.A(_4512_),
    .B(_0403_),
    .Y(_0497_));
 sg13g2_nand3_1 _5243_ (.B(_0484_),
    .C(_0489_),
    .A(_0486_),
    .Y(_0498_));
 sg13g2_nand3b_1 _5244_ (.B(_0498_),
    .C(_0490_),
    .Y(_0499_),
    .A_N(_0497_));
 sg13g2_xnor2_1 _5245_ (.Y(_0500_),
    .A(_0496_),
    .B(_0499_));
 sg13g2_nor2_1 _5246_ (.A(_4505_),
    .B(net69),
    .Y(_0501_));
 sg13g2_a21oi_1 _5247_ (.A1(_0500_),
    .A2(net70),
    .Y(_0131_),
    .B1(_0501_));
 sg13g2_nand2_1 _5248_ (.Y(_0502_),
    .A(_0489_),
    .B(_0496_));
 sg13g2_inv_1 _5249_ (.Y(_0503_),
    .A(_0502_));
 sg13g2_a21oi_1 _5250_ (.A1(_0503_),
    .A2(_0491_),
    .Y(_0504_),
    .B1(_0497_));
 sg13g2_o21ai_1 _5251_ (.B1(_0504_),
    .Y(_0505_),
    .A1(_0502_),
    .A2(_0492_));
 sg13g2_nor2_1 _5252_ (.A(_4505_),
    .B(net25),
    .Y(_0506_));
 sg13g2_o21ai_1 _5253_ (.B1(_4489_),
    .Y(_0507_),
    .A1(_0506_),
    .A2(_0505_));
 sg13g2_a21oi_1 _5254_ (.A1(_0440_),
    .A2(_0505_),
    .Y(_0508_),
    .B1(_0507_));
 sg13g2_xnor2_1 _5255_ (.Y(_0132_),
    .A(_4498_),
    .B(_0508_));
 sg13g2_nand2_1 _5256_ (.Y(_0509_),
    .A(_0452_),
    .B(_0450_));
 sg13g2_nand3b_1 _5257_ (.B(_4489_),
    .C(_0509_),
    .Y(_0510_),
    .A_N(_0453_));
 sg13g2_o21ai_1 _5258_ (.B1(_0510_),
    .Y(_0133_),
    .A1(_0448_),
    .A2(_0426_));
 sg13g2_or3_1 _5259_ (.A(_0454_),
    .B(_0449_),
    .C(_0453_),
    .X(_0511_));
 sg13g2_nand3_1 _5260_ (.B(_4574_),
    .C(_0455_),
    .A(_0511_),
    .Y(_0512_));
 sg13g2_o21ai_1 _5261_ (.B1(_0512_),
    .Y(_0134_),
    .A1(_0447_),
    .A2(_0426_));
 sg13g2_nor2b_1 _5262_ (.A(_0459_),
    .B_N(_0458_),
    .Y(_0513_));
 sg13g2_xnor2_1 _5263_ (.Y(_0514_),
    .A(_0513_),
    .B(_0456_));
 sg13g2_nor2_1 _5264_ (.A(\vgademo.a_sin[3] ),
    .B(net69),
    .Y(_0515_));
 sg13g2_a21oi_1 _5265_ (.A1(_0514_),
    .A2(net70),
    .Y(_0135_),
    .B1(_0515_));
 sg13g2_nand2b_1 _5266_ (.Y(_0516_),
    .B(_0462_),
    .A_N(_0463_));
 sg13g2_xnor2_1 _5267_ (.Y(_0517_),
    .A(_0516_),
    .B(_0460_));
 sg13g2_nor2_1 _5268_ (.A(_0461_),
    .B(net69),
    .Y(_0518_));
 sg13g2_a21oi_1 _5269_ (.A1(_0517_),
    .A2(net70),
    .Y(_0136_),
    .B1(_0518_));
 sg13g2_nor2b_1 _5270_ (.A(_0467_),
    .B_N(_0466_),
    .Y(_0519_));
 sg13g2_o21ai_1 _5271_ (.B1(_4489_),
    .Y(_0520_),
    .A1(_0519_),
    .A2(_0464_));
 sg13g2_a21oi_1 _5272_ (.A1(_0464_),
    .A2(_0519_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_a21o_1 _5273_ (.A2(net64),
    .A1(\vgademo.a_sin[5] ),
    .B1(_0521_),
    .X(_0137_));
 sg13g2_nand2b_1 _5274_ (.Y(_0522_),
    .B(_0470_),
    .A_N(_0471_));
 sg13g2_xnor2_1 _5275_ (.Y(_0523_),
    .A(_0522_),
    .B(_0468_));
 sg13g2_nor2_1 _5276_ (.A(\vgademo.a_sin[6] ),
    .B(_0437_),
    .Y(_0524_));
 sg13g2_a21oi_1 _5277_ (.A1(_0523_),
    .A2(_0421_),
    .Y(_0138_),
    .B1(_0524_));
 sg13g2_nor2_1 _5278_ (.A(_0476_),
    .B(_0474_),
    .Y(_0525_));
 sg13g2_xor2_1 _5279_ (.B(_0472_),
    .A(_0525_),
    .X(_0526_));
 sg13g2_nor2_1 _5280_ (.A(_4521_),
    .B(_0437_),
    .Y(_0527_));
 sg13g2_a21oi_1 _5281_ (.A1(_0526_),
    .A2(_0421_),
    .Y(_0139_),
    .B1(_0527_));
 sg13g2_nor2_1 _5282_ (.A(_0445_),
    .B(_0446_),
    .Y(_0528_));
 sg13g2_xor2_1 _5283_ (.B(_0477_),
    .A(_0528_),
    .X(_0529_));
 sg13g2_nor2_1 _5284_ (.A(_4519_),
    .B(net69),
    .Y(_0530_));
 sg13g2_a21oi_1 _5285_ (.A1(_0529_),
    .A2(net70),
    .Y(_0140_),
    .B1(_0530_));
 sg13g2_nand2_1 _5286_ (.Y(_0531_),
    .A(_0479_),
    .B(_0444_));
 sg13g2_nand3b_1 _5287_ (.B(_4489_),
    .C(_0531_),
    .Y(_0532_),
    .A_N(_0480_));
 sg13g2_o21ai_1 _5288_ (.B1(_0532_),
    .Y(_0141_),
    .A1(_4517_),
    .A2(_0426_));
 sg13g2_inv_2 _5289_ (.Y(_0533_),
    .A(net137));
 sg13g2_nor2_1 _5290_ (.A(_0533_),
    .B(_4403_),
    .Y(_0534_));
 sg13g2_buf_1 _5291_ (.A(_0534_),
    .X(_0535_));
 sg13g2_inv_2 _5292_ (.Y(_0536_),
    .A(_0535_));
 sg13g2_buf_1 _5293_ (.A(_0536_),
    .X(_0537_));
 sg13g2_nor3_1 _5294_ (.A(net123),
    .B(_4285_),
    .C(_4397_),
    .Y(_0538_));
 sg13g2_nand2_1 _5295_ (.Y(_0539_),
    .A(_4296_),
    .B(_0538_));
 sg13g2_buf_1 _5296_ (.A(_0539_),
    .X(_0540_));
 sg13g2_buf_1 _5297_ (.A(_0540_),
    .X(_0541_));
 sg13g2_buf_1 _5298_ (.A(net63),
    .X(_0542_));
 sg13g2_inv_1 _5299_ (.Y(_0543_),
    .A(\vgademo.b_sin[7] ));
 sg13g2_nor2_1 _5300_ (.A(\vgademo.b_cos[0] ),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_buf_1 _5301_ (.A(_0540_),
    .X(_0545_));
 sg13g2_nor2_1 _5302_ (.A(_4515_),
    .B(net62),
    .Y(_0546_));
 sg13g2_a21oi_1 _5303_ (.A1(net56),
    .A2(_0544_),
    .Y(_0547_),
    .B1(_0546_));
 sg13g2_nand2_1 _5304_ (.Y(_0548_),
    .A(_0535_),
    .B(\vgademo.b_sin[7] ));
 sg13g2_nor2_1 _5305_ (.A(_0533_),
    .B(_0540_),
    .Y(_0549_));
 sg13g2_buf_1 _5306_ (.A(_0549_),
    .X(_0550_));
 sg13g2_inv_1 _5307_ (.Y(_0551_),
    .A(net55));
 sg13g2_nand3_1 _5308_ (.B(\vgademo.b_cos[0] ),
    .C(_0551_),
    .A(_0548_),
    .Y(_0552_));
 sg13g2_o21ai_1 _5309_ (.B1(_0552_),
    .Y(_0142_),
    .A1(net57),
    .A2(_0547_));
 sg13g2_buf_2 _5310_ (.A(\vgademo.b_cos[10] ),
    .X(_0553_));
 sg13g2_inv_2 _5311_ (.Y(_0554_),
    .A(_0553_));
 sg13g2_buf_1 _5312_ (.A(_0535_),
    .X(_0555_));
 sg13g2_buf_1 _5313_ (.A(net61),
    .X(_0556_));
 sg13g2_inv_1 _5314_ (.Y(_0557_),
    .A(_0540_));
 sg13g2_buf_1 _5315_ (.A(_0557_),
    .X(_0558_));
 sg13g2_buf_1 _5316_ (.A(_0558_),
    .X(_0559_));
 sg13g2_buf_1 _5317_ (.A(\vgademo.b_sin[11] ),
    .X(_0560_));
 sg13g2_xor2_1 _5318_ (.B(_0553_),
    .A(net120),
    .X(_0561_));
 sg13g2_inv_1 _5319_ (.Y(_0562_),
    .A(\vgademo.b_cos[2] ));
 sg13g2_buf_1 _5320_ (.A(\vgademo.b_sin[8] ),
    .X(_0563_));
 sg13g2_inv_1 _5321_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_xnor2_1 _5322_ (.Y(_0565_),
    .A(\vgademo.b_cos[1] ),
    .B(_0563_));
 sg13g2_inv_1 _5323_ (.Y(_0566_),
    .A(_0544_));
 sg13g2_nand2_1 _5324_ (.Y(_0567_),
    .A(_0565_),
    .B(_0566_));
 sg13g2_inv_1 _5325_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_a21oi_1 _5326_ (.A1(\vgademo.b_cos[1] ),
    .A2(_0564_),
    .Y(_0569_),
    .B1(_0568_));
 sg13g2_xnor2_1 _5327_ (.Y(_0570_),
    .A(\vgademo.b_cos[2] ),
    .B(\vgademo.b_sin[9] ));
 sg13g2_nand2b_1 _5328_ (.Y(_0571_),
    .B(_0570_),
    .A_N(_0569_));
 sg13g2_o21ai_1 _5329_ (.B1(_0571_),
    .Y(_0572_),
    .A1(_0562_),
    .A2(\vgademo.b_sin[9] ));
 sg13g2_inv_1 _5330_ (.Y(_0573_),
    .A(\vgademo.b_sin[10] ));
 sg13g2_nor2_1 _5331_ (.A(\vgademo.b_cos[3] ),
    .B(_0573_),
    .Y(_0574_));
 sg13g2_inv_1 _5332_ (.Y(_0575_),
    .A(_0574_));
 sg13g2_inv_1 _5333_ (.Y(_0576_),
    .A(\vgademo.b_cos[3] ));
 sg13g2_nor2_1 _5334_ (.A(\vgademo.b_sin[10] ),
    .B(_0576_),
    .Y(_0577_));
 sg13g2_a21oi_1 _5335_ (.A1(_0572_),
    .A2(_0575_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_inv_1 _5336_ (.Y(_0579_),
    .A(net120));
 sg13g2_nand2_1 _5337_ (.Y(_0580_),
    .A(net101),
    .B(\vgademo.b_cos[4] ));
 sg13g2_nor2_1 _5338_ (.A(\vgademo.b_cos[4] ),
    .B(net101),
    .Y(_0581_));
 sg13g2_a21oi_1 _5339_ (.A1(_0578_),
    .A2(_0580_),
    .Y(_0582_),
    .B1(_0581_));
 sg13g2_inv_1 _5340_ (.Y(_0583_),
    .A(\vgademo.b_cos[5] ));
 sg13g2_nand2_1 _5341_ (.Y(_0584_),
    .A(_0583_),
    .B(net120));
 sg13g2_nand2_1 _5342_ (.Y(_0585_),
    .A(_0582_),
    .B(_0584_));
 sg13g2_nand2_1 _5343_ (.Y(_0586_),
    .A(_0579_),
    .B(\vgademo.b_cos[5] ));
 sg13g2_nand2_1 _5344_ (.Y(_0587_),
    .A(_0585_),
    .B(_0586_));
 sg13g2_buf_2 _5345_ (.A(\vgademo.b_cos[7] ),
    .X(_0588_));
 sg13g2_xnor2_1 _5346_ (.Y(_0589_),
    .A(net120),
    .B(_0588_));
 sg13g2_buf_1 _5347_ (.A(\vgademo.b_cos[6] ),
    .X(_0590_));
 sg13g2_inv_1 _5348_ (.Y(_0591_),
    .A(_0590_));
 sg13g2_nor2_1 _5349_ (.A(net120),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_nor2_1 _5350_ (.A(_0590_),
    .B(net101),
    .Y(_0593_));
 sg13g2_nor2_1 _5351_ (.A(_0592_),
    .B(_0593_),
    .Y(_0594_));
 sg13g2_nand3_1 _5352_ (.B(_0589_),
    .C(_0594_),
    .A(_0587_),
    .Y(_0595_));
 sg13g2_o21ai_1 _5353_ (.B1(net101),
    .Y(_0596_),
    .A1(_0590_),
    .A2(_0588_));
 sg13g2_nand2_1 _5354_ (.Y(_0597_),
    .A(_0595_),
    .B(_0596_));
 sg13g2_buf_1 _5355_ (.A(\vgademo.b_cos[9] ),
    .X(_0598_));
 sg13g2_buf_1 _5356_ (.A(_0598_),
    .X(_0599_));
 sg13g2_xnor2_1 _5357_ (.Y(_0600_),
    .A(net120),
    .B(net100));
 sg13g2_buf_1 _5358_ (.A(\vgademo.b_cos[8] ),
    .X(_0601_));
 sg13g2_xnor2_1 _5359_ (.Y(_0602_),
    .A(_0560_),
    .B(net119));
 sg13g2_nand3_1 _5360_ (.B(_0600_),
    .C(_0602_),
    .A(_0597_),
    .Y(_0603_));
 sg13g2_o21ai_1 _5361_ (.B1(net101),
    .Y(_0604_),
    .A1(net119),
    .A2(net100));
 sg13g2_nand2_1 _5362_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_xor2_1 _5363_ (.B(_0605_),
    .A(_0561_),
    .X(_0606_));
 sg13g2_inv_1 _5364_ (.Y(_0607_),
    .A(_0606_));
 sg13g2_buf_1 _5365_ (.A(_0558_),
    .X(_0608_));
 sg13g2_a21oi_1 _5366_ (.A1(_0392_),
    .A2(net44),
    .Y(_0609_),
    .B1(net57));
 sg13g2_o21ai_1 _5367_ (.B1(_0609_),
    .Y(_0610_),
    .A1(_0559_),
    .A2(_0607_));
 sg13g2_o21ai_1 _5368_ (.B1(_0610_),
    .Y(_0143_),
    .A1(_0554_),
    .A2(net54));
 sg13g2_buf_2 _5369_ (.A(\vgademo.b_cos[11] ),
    .X(_0611_));
 sg13g2_xor2_1 _5370_ (.B(_0611_),
    .A(net120),
    .X(_0612_));
 sg13g2_a21oi_1 _5371_ (.A1(_0582_),
    .A2(_0584_),
    .Y(_0613_),
    .B1(_0592_));
 sg13g2_o21ai_1 _5372_ (.B1(_0586_),
    .Y(_0614_),
    .A1(_0593_),
    .A2(_0613_));
 sg13g2_nand3_1 _5373_ (.B(_0602_),
    .C(_0589_),
    .A(_0614_),
    .Y(_0615_));
 sg13g2_o21ai_1 _5374_ (.B1(net101),
    .Y(_0616_),
    .A1(_0588_),
    .A2(net119));
 sg13g2_nand2_1 _5375_ (.Y(_0617_),
    .A(_0615_),
    .B(_0616_));
 sg13g2_nand2_1 _5376_ (.Y(_0618_),
    .A(_0617_),
    .B(_0600_));
 sg13g2_inv_1 _5377_ (.Y(_0619_),
    .A(_0598_));
 sg13g2_nand2_1 _5378_ (.Y(_0620_),
    .A(_0619_),
    .B(_0554_));
 sg13g2_nand2_1 _5379_ (.Y(_0621_),
    .A(_0620_),
    .B(net101));
 sg13g2_o21ai_1 _5380_ (.B1(_0621_),
    .Y(_0622_),
    .A1(_0561_),
    .A2(_0618_));
 sg13g2_or2_1 _5381_ (.X(_0623_),
    .B(_0622_),
    .A(_0612_));
 sg13g2_nand2_1 _5382_ (.Y(_0624_),
    .A(_0622_),
    .B(_0612_));
 sg13g2_nand2_1 _5383_ (.Y(_0625_),
    .A(_0623_),
    .B(_0624_));
 sg13g2_inv_1 _5384_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_o21ai_1 _5385_ (.B1(_0535_),
    .Y(_0627_),
    .A1(_0398_),
    .A2(net63));
 sg13g2_a21oi_1 _5386_ (.A1(_0626_),
    .A2(net56),
    .Y(_0628_),
    .B1(_0627_));
 sg13g2_a21o_1 _5387_ (.A2(net57),
    .A1(_0611_),
    .B1(_0628_),
    .X(_0144_));
 sg13g2_nor2_1 _5388_ (.A(_0566_),
    .B(_0565_),
    .Y(_0629_));
 sg13g2_o21ai_1 _5389_ (.B1(net62),
    .Y(_0630_),
    .A1(_0568_),
    .A2(_0629_));
 sg13g2_o21ai_1 _5390_ (.B1(_0630_),
    .Y(_0631_),
    .A1(_4533_),
    .A2(net56));
 sg13g2_nor2_1 _5391_ (.A(\vgademo.b_cos[1] ),
    .B(net61),
    .Y(_0632_));
 sg13g2_a21oi_1 _5392_ (.A1(_0631_),
    .A2(net54),
    .Y(_0145_),
    .B1(_0632_));
 sg13g2_xnor2_1 _5393_ (.Y(_0633_),
    .A(_0570_),
    .B(_0569_));
 sg13g2_buf_1 _5394_ (.A(net63),
    .X(_0634_));
 sg13g2_nand2_1 _5395_ (.Y(_0635_),
    .A(_0633_),
    .B(net53));
 sg13g2_a21oi_1 _5396_ (.A1(_4540_),
    .A2(net45),
    .Y(_0636_),
    .B1(net57));
 sg13g2_a22oi_1 _5397_ (.Y(_0146_),
    .B1(_0635_),
    .B2(_0636_),
    .A2(net57),
    .A1(_0562_));
 sg13g2_buf_1 _5398_ (.A(_0558_),
    .X(_0637_));
 sg13g2_nor2_1 _5399_ (.A(_0577_),
    .B(_0574_),
    .Y(_0638_));
 sg13g2_xor2_1 _5400_ (.B(_0572_),
    .A(_0638_),
    .X(_0639_));
 sg13g2_buf_1 _5401_ (.A(_0536_),
    .X(_0640_));
 sg13g2_a21oi_1 _5402_ (.A1(_4548_),
    .A2(net44),
    .Y(_0641_),
    .B1(net52));
 sg13g2_o21ai_1 _5403_ (.B1(_0641_),
    .Y(_0642_),
    .A1(net43),
    .A2(_0639_));
 sg13g2_o21ai_1 _5404_ (.B1(_0642_),
    .Y(_0147_),
    .A1(_0576_),
    .A2(net54));
 sg13g2_buf_1 _5405_ (.A(_0558_),
    .X(_0643_));
 sg13g2_nand2b_1 _5406_ (.Y(_0644_),
    .B(_0580_),
    .A_N(_0581_));
 sg13g2_o21ai_1 _5407_ (.B1(_0540_),
    .Y(_0645_),
    .A1(_0644_),
    .A2(_0578_));
 sg13g2_a21oi_1 _5408_ (.A1(_0578_),
    .A2(_0644_),
    .Y(_0646_),
    .B1(_0645_));
 sg13g2_a21oi_1 _5409_ (.A1(_4507_),
    .A2(net42),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nand2_1 _5410_ (.Y(_0648_),
    .A(net57),
    .B(\vgademo.b_cos[4] ));
 sg13g2_o21ai_1 _5411_ (.B1(_0648_),
    .Y(_0148_),
    .A1(net57),
    .A2(_0647_));
 sg13g2_a21oi_1 _5412_ (.A1(_4503_),
    .A2(_0643_),
    .Y(_0649_),
    .B1(net57));
 sg13g2_nand2_1 _5413_ (.Y(_0650_),
    .A(_0586_),
    .B(_0584_));
 sg13g2_xnor2_1 _5414_ (.Y(_0651_),
    .A(_0650_),
    .B(_0582_));
 sg13g2_nand2_1 _5415_ (.Y(_0652_),
    .A(_0651_),
    .B(net53));
 sg13g2_a22oi_1 _5416_ (.Y(_0149_),
    .B1(_0649_),
    .B2(_0652_),
    .A2(_0537_),
    .A1(_0583_));
 sg13g2_xor2_1 _5417_ (.B(_0587_),
    .A(_0594_),
    .X(_0653_));
 sg13g2_a21oi_1 _5418_ (.A1(_4558_),
    .A2(net44),
    .Y(_0654_),
    .B1(net52));
 sg13g2_o21ai_1 _5419_ (.B1(_0654_),
    .Y(_0655_),
    .A1(net43),
    .A2(_0653_));
 sg13g2_o21ai_1 _5420_ (.B1(_0655_),
    .Y(_0150_),
    .A1(_0591_),
    .A2(net54));
 sg13g2_inv_1 _5421_ (.Y(_0656_),
    .A(_0588_));
 sg13g2_xor2_1 _5422_ (.B(_0614_),
    .A(_0589_),
    .X(_0657_));
 sg13g2_a21oi_1 _5423_ (.A1(_4496_),
    .A2(net44),
    .Y(_0658_),
    .B1(net52));
 sg13g2_o21ai_1 _5424_ (.B1(_0658_),
    .Y(_0659_),
    .A1(net43),
    .A2(_0657_));
 sg13g2_o21ai_1 _5425_ (.B1(_0659_),
    .Y(_0151_),
    .A1(_0656_),
    .A2(net54));
 sg13g2_inv_1 _5426_ (.Y(_0660_),
    .A(net119));
 sg13g2_xor2_1 _5427_ (.B(_0597_),
    .A(_0602_),
    .X(_0661_));
 sg13g2_a21oi_1 _5428_ (.A1(_0375_),
    .A2(net44),
    .Y(_0662_),
    .B1(net52));
 sg13g2_o21ai_1 _5429_ (.B1(_0662_),
    .Y(_0663_),
    .A1(net43),
    .A2(_0661_));
 sg13g2_o21ai_1 _5430_ (.B1(_0663_),
    .Y(_0152_),
    .A1(_0660_),
    .A2(net54));
 sg13g2_xor2_1 _5431_ (.B(_0617_),
    .A(_0600_),
    .X(_0664_));
 sg13g2_a21oi_1 _5432_ (.A1(_0391_),
    .A2(net44),
    .Y(_0665_),
    .B1(net52));
 sg13g2_o21ai_1 _5433_ (.B1(_0665_),
    .Y(_0666_),
    .A1(net43),
    .A2(_0664_));
 sg13g2_o21ai_1 _5434_ (.B1(_0666_),
    .Y(_0153_),
    .A1(_0619_),
    .A2(_0556_));
 sg13g2_inv_1 _5435_ (.Y(_0667_),
    .A(\vgademo.b_sin[0] ));
 sg13g2_xnor2_1 _5436_ (.Y(_0668_),
    .A(_0667_),
    .B(_0657_));
 sg13g2_a21oi_1 _5437_ (.A1(_0457_),
    .A2(_0608_),
    .Y(_0669_),
    .B1(_0640_));
 sg13g2_o21ai_1 _5438_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0637_),
    .A2(_0668_));
 sg13g2_o21ai_1 _5439_ (.B1(_0670_),
    .Y(_0156_),
    .A1(_0667_),
    .A2(_0556_));
 sg13g2_buf_1 _5440_ (.A(_0625_),
    .X(_0671_));
 sg13g2_nor2_1 _5441_ (.A(\vgademo.b_sin[10] ),
    .B(_0671_),
    .Y(_0672_));
 sg13g2_nand2_1 _5442_ (.Y(_0673_),
    .A(net28),
    .B(\vgademo.b_sin[10] ));
 sg13g2_nor2b_1 _5443_ (.A(_0672_),
    .B_N(_0673_),
    .Y(_0674_));
 sg13g2_xnor2_1 _5444_ (.Y(_0675_),
    .A(_0543_),
    .B(net28));
 sg13g2_xnor2_1 _5445_ (.Y(_0676_),
    .A(_0563_),
    .B(net28));
 sg13g2_inv_1 _5446_ (.Y(_0677_),
    .A(\vgademo.b_sin[4] ));
 sg13g2_nor2_1 _5447_ (.A(_0677_),
    .B(_0626_),
    .Y(_0678_));
 sg13g2_nor2_1 _5448_ (.A(\vgademo.b_sin[3] ),
    .B(_0607_),
    .Y(_0679_));
 sg13g2_inv_1 _5449_ (.Y(_0680_),
    .A(\vgademo.b_sin[3] ));
 sg13g2_nor2_1 _5450_ (.A(_0680_),
    .B(_0606_),
    .Y(_0681_));
 sg13g2_xnor2_1 _5451_ (.Y(_0682_),
    .A(\vgademo.b_sin[1] ),
    .B(_0661_));
 sg13g2_nor2b_1 _5452_ (.A(_0667_),
    .B_N(_0657_),
    .Y(_0683_));
 sg13g2_nor2b_1 _5453_ (.A(_0682_),
    .B_N(_0683_),
    .Y(_0684_));
 sg13g2_a21oi_1 _5454_ (.A1(\vgademo.b_sin[1] ),
    .A2(_0661_),
    .Y(_0685_),
    .B1(_0684_));
 sg13g2_nand2_1 _5455_ (.Y(_0686_),
    .A(_0664_),
    .B(\vgademo.b_sin[2] ));
 sg13g2_nor2_1 _5456_ (.A(\vgademo.b_sin[2] ),
    .B(_0664_),
    .Y(_0687_));
 sg13g2_a21oi_1 _5457_ (.A1(_0685_),
    .A2(_0686_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_nor2_1 _5458_ (.A(_0681_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nor2_1 _5459_ (.A(_0679_),
    .B(_0689_),
    .Y(_0690_));
 sg13g2_nor2_1 _5460_ (.A(\vgademo.b_sin[4] ),
    .B(_0625_),
    .Y(_0691_));
 sg13g2_inv_1 _5461_ (.Y(_0692_),
    .A(_0691_));
 sg13g2_o21ai_1 _5462_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0678_),
    .A2(_0690_));
 sg13g2_inv_1 _5463_ (.Y(_0694_),
    .A(_0693_));
 sg13g2_nor2_1 _5464_ (.A(\vgademo.b_sin[5] ),
    .B(net28),
    .Y(_0695_));
 sg13g2_inv_1 _5465_ (.Y(_0696_),
    .A(_0695_));
 sg13g2_inv_1 _5466_ (.Y(_0697_),
    .A(\vgademo.b_sin[5] ));
 sg13g2_nor2_1 _5467_ (.A(_0697_),
    .B(_0626_),
    .Y(_0698_));
 sg13g2_a21oi_1 _5468_ (.A1(_0694_),
    .A2(_0696_),
    .Y(_0699_),
    .B1(_0698_));
 sg13g2_inv_1 _5469_ (.Y(_0700_),
    .A(\vgademo.b_sin[6] ));
 sg13g2_nor2_1 _5470_ (.A(_0700_),
    .B(_0626_),
    .Y(_0701_));
 sg13g2_inv_1 _5471_ (.Y(_0702_),
    .A(_0701_));
 sg13g2_nor2_1 _5472_ (.A(\vgademo.b_sin[6] ),
    .B(net28),
    .Y(_0703_));
 sg13g2_a21oi_1 _5473_ (.A1(_0699_),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_nor2b_1 _5474_ (.A(_0676_),
    .B_N(_0704_),
    .Y(_0705_));
 sg13g2_a22oi_1 _5475_ (.Y(_0706_),
    .B1(_0675_),
    .B2(_0705_),
    .A2(net28),
    .A1(_0563_));
 sg13g2_o21ai_1 _5476_ (.B1(_0706_),
    .Y(_0707_),
    .A1(_0543_),
    .A2(_0626_));
 sg13g2_inv_1 _5477_ (.Y(_0708_),
    .A(\vgademo.b_sin[9] ));
 sg13g2_xnor2_1 _5478_ (.Y(_0709_),
    .A(_0708_),
    .B(_0671_));
 sg13g2_nor2_1 _5479_ (.A(_0708_),
    .B(_0626_),
    .Y(_0710_));
 sg13g2_a21oi_1 _5480_ (.A1(_0707_),
    .A2(_0709_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_xnor2_1 _5481_ (.Y(_0712_),
    .A(_0674_),
    .B(_0711_));
 sg13g2_a21oi_1 _5482_ (.A1(_4506_),
    .A2(net44),
    .Y(_0713_),
    .B1(net52));
 sg13g2_o21ai_1 _5483_ (.B1(_0713_),
    .Y(_0714_),
    .A1(net43),
    .A2(_0712_));
 sg13g2_o21ai_1 _5484_ (.B1(_0714_),
    .Y(_0157_),
    .A1(_0573_),
    .A2(net54));
 sg13g2_xnor2_1 _5485_ (.Y(_0715_),
    .A(net120),
    .B(net28));
 sg13g2_o21ai_1 _5486_ (.B1(_0673_),
    .Y(_0716_),
    .A1(_0672_),
    .A2(_0711_));
 sg13g2_xnor2_1 _5487_ (.Y(_0717_),
    .A(_0715_),
    .B(_0716_));
 sg13g2_a21oi_1 _5488_ (.A1(_4498_),
    .A2(net44),
    .Y(_0718_),
    .B1(net52));
 sg13g2_o21ai_1 _5489_ (.B1(_0718_),
    .Y(_0719_),
    .A1(net43),
    .A2(_0717_));
 sg13g2_o21ai_1 _5490_ (.B1(_0719_),
    .Y(_0158_),
    .A1(net101),
    .A2(net54));
 sg13g2_xor2_1 _5491_ (.B(_0682_),
    .A(_0683_),
    .X(_0720_));
 sg13g2_o21ai_1 _5492_ (.B1(_0535_),
    .Y(_0721_),
    .A1(_0461_),
    .A2(net63));
 sg13g2_a21oi_1 _5493_ (.A1(_0720_),
    .A2(_0542_),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_a21o_1 _5494_ (.A2(_0537_),
    .A1(\vgademo.b_sin[1] ),
    .B1(_0722_),
    .X(_0159_));
 sg13g2_inv_1 _5495_ (.Y(_0723_),
    .A(\vgademo.b_sin[2] ));
 sg13g2_nor2b_1 _5496_ (.A(_0687_),
    .B_N(_0686_),
    .Y(_0724_));
 sg13g2_xnor2_1 _5497_ (.Y(_0725_),
    .A(_0685_),
    .B(_0724_));
 sg13g2_a21oi_1 _5498_ (.A1(_0465_),
    .A2(_0608_),
    .Y(_0726_),
    .B1(_0640_));
 sg13g2_o21ai_1 _5499_ (.B1(_0726_),
    .Y(_0727_),
    .A1(_0637_),
    .A2(_0725_));
 sg13g2_o21ai_1 _5500_ (.B1(_0727_),
    .Y(_0160_),
    .A1(_0723_),
    .A2(net61));
 sg13g2_nor2_1 _5501_ (.A(_0681_),
    .B(_0679_),
    .Y(_0728_));
 sg13g2_xor2_1 _5502_ (.B(_0688_),
    .A(_0728_),
    .X(_0729_));
 sg13g2_buf_1 _5503_ (.A(_0558_),
    .X(_0730_));
 sg13g2_a21oi_1 _5504_ (.A1(_4491_),
    .A2(_0730_),
    .Y(_0731_),
    .B1(net52));
 sg13g2_o21ai_1 _5505_ (.B1(_0731_),
    .Y(_0732_),
    .A1(net43),
    .A2(_0729_));
 sg13g2_o21ai_1 _5506_ (.B1(_0732_),
    .Y(_0161_),
    .A1(_0680_),
    .A2(_0555_));
 sg13g2_nor2_1 _5507_ (.A(_0691_),
    .B(_0678_),
    .Y(_0733_));
 sg13g2_xor2_1 _5508_ (.B(_0690_),
    .A(_0733_),
    .X(_0734_));
 sg13g2_a21oi_1 _5509_ (.A1(_4522_),
    .A2(net41),
    .Y(_0735_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5510_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0643_),
    .A2(_0734_));
 sg13g2_o21ai_1 _5511_ (.B1(_0736_),
    .Y(_0162_),
    .A1(_0677_),
    .A2(_0555_));
 sg13g2_nor2_1 _5512_ (.A(_0695_),
    .B(_0698_),
    .Y(_0737_));
 sg13g2_xnor2_1 _5513_ (.Y(_0738_),
    .A(_0737_),
    .B(_0693_));
 sg13g2_a21oi_1 _5514_ (.A1(_4520_),
    .A2(net41),
    .Y(_0739_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5515_ (.B1(_0739_),
    .Y(_0740_),
    .A1(net42),
    .A2(_0738_));
 sg13g2_o21ai_1 _5516_ (.B1(_0740_),
    .Y(_0163_),
    .A1(_0697_),
    .A2(net61));
 sg13g2_nor2_1 _5517_ (.A(_0703_),
    .B(_0701_),
    .Y(_0741_));
 sg13g2_xnor2_1 _5518_ (.Y(_0742_),
    .A(_0741_),
    .B(_0699_));
 sg13g2_a21oi_1 _5519_ (.A1(_4517_),
    .A2(net41),
    .Y(_0743_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5520_ (.B1(_0743_),
    .Y(_0744_),
    .A1(net42),
    .A2(_0742_));
 sg13g2_o21ai_1 _5521_ (.B1(_0744_),
    .Y(_0164_),
    .A1(_0700_),
    .A2(net61));
 sg13g2_xor2_1 _5522_ (.B(_0704_),
    .A(_0675_),
    .X(_0745_));
 sg13g2_a21oi_1 _5523_ (.A1(_4537_),
    .A2(net41),
    .Y(_0746_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5524_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net42),
    .A2(_0745_));
 sg13g2_o21ai_1 _5525_ (.B1(_0747_),
    .Y(_0165_),
    .A1(_0543_),
    .A2(net61));
 sg13g2_nor2b_1 _5526_ (.A(_0699_),
    .B_N(_0675_),
    .Y(_0748_));
 sg13g2_a21oi_1 _5527_ (.A1(\vgademo.b_sin[7] ),
    .A2(net28),
    .Y(_0749_),
    .B1(_0748_));
 sg13g2_o21ai_1 _5528_ (.B1(_0702_),
    .Y(_0750_),
    .A1(_0703_),
    .A2(_0749_));
 sg13g2_xnor2_1 _5529_ (.Y(_0751_),
    .A(_0676_),
    .B(_0750_));
 sg13g2_a21oi_1 _5530_ (.A1(_4542_),
    .A2(net41),
    .Y(_0752_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5531_ (.B1(_0752_),
    .Y(_0753_),
    .A1(net42),
    .A2(_0751_));
 sg13g2_o21ai_1 _5532_ (.B1(_0753_),
    .Y(_0166_),
    .A1(_0564_),
    .A2(net61));
 sg13g2_xor2_1 _5533_ (.B(_0707_),
    .A(_0709_),
    .X(_0754_));
 sg13g2_a21oi_1 _5534_ (.A1(_4512_),
    .A2(net41),
    .Y(_0755_),
    .B1(_0536_));
 sg13g2_o21ai_1 _5535_ (.B1(_0755_),
    .Y(_0756_),
    .A1(net42),
    .A2(_0754_));
 sg13g2_o21ai_1 _5536_ (.B1(_0756_),
    .Y(_0167_),
    .A1(_0708_),
    .A2(net61));
 sg13g2_buf_1 _5537_ (.A(_4324_),
    .X(_0757_));
 sg13g2_inv_1 _5538_ (.Y(_0758_),
    .A(_4376_));
 sg13g2_nor2_1 _5539_ (.A(_4348_),
    .B(_4347_),
    .Y(_0759_));
 sg13g2_inv_2 _5540_ (.Y(_0760_),
    .A(_4306_));
 sg13g2_nor2_1 _5541_ (.A(_4364_),
    .B(_0760_),
    .Y(_0761_));
 sg13g2_nand4_1 _5542_ (.B(_4353_),
    .C(_0759_),
    .A(_0758_),
    .Y(_0762_),
    .D(_0761_));
 sg13g2_buf_1 _5543_ (.A(\vgademo.audio_songpos[4] ),
    .X(_0763_));
 sg13g2_buf_1 _5544_ (.A(_0763_),
    .X(_0764_));
 sg13g2_buf_1 _5545_ (.A(\vgademo.audio_songpos[6] ),
    .X(_0765_));
 sg13g2_buf_1 _5546_ (.A(\vgademo.audio_songpos[1] ),
    .X(_0766_));
 sg13g2_inv_2 _5547_ (.Y(_0767_),
    .A(net117));
 sg13g2_buf_1 _5548_ (.A(\vgademo.audio_songpos[0] ),
    .X(_0768_));
 sg13g2_inv_2 _5549_ (.Y(_0769_),
    .A(net116));
 sg13g2_nand2_2 _5550_ (.Y(_0770_),
    .A(_0767_),
    .B(_0769_));
 sg13g2_buf_1 _5551_ (.A(\vgademo.audio_songpos[3] ),
    .X(_0771_));
 sg13g2_buf_1 _5552_ (.A(_0771_),
    .X(_0772_));
 sg13g2_buf_2 _5553_ (.A(\vgademo.audio_songpos[2] ),
    .X(_0773_));
 sg13g2_nor2_2 _5554_ (.A(net97),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_buf_1 _5555_ (.A(\vgademo.audio_songpos[5] ),
    .X(_0775_));
 sg13g2_inv_1 _5556_ (.Y(_0776_),
    .A(_0775_));
 sg13g2_buf_1 _5557_ (.A(_0776_),
    .X(_0777_));
 sg13g2_buf_1 _5558_ (.A(\vgademo.audio_songpos[7] ),
    .X(_0778_));
 sg13g2_inv_1 _5559_ (.Y(_0779_),
    .A(_0778_));
 sg13g2_nand3_1 _5560_ (.B(net84),
    .C(_0779_),
    .A(_0774_),
    .Y(_0780_));
 sg13g2_nor4_1 _5561_ (.A(net98),
    .B(net118),
    .C(_0770_),
    .D(_0780_),
    .Y(_0781_));
 sg13g2_nand2_1 _5562_ (.Y(_0782_),
    .A(_0758_),
    .B(_4340_));
 sg13g2_nand3_1 _5563_ (.B(_0781_),
    .C(_0782_),
    .A(_0762_),
    .Y(_0783_));
 sg13g2_nand2_1 _5564_ (.Y(_0784_),
    .A(_0783_),
    .B(_4489_));
 sg13g2_buf_1 _5565_ (.A(_0784_),
    .X(_0785_));
 sg13g2_nand2_1 _5566_ (.Y(_0786_),
    .A(net64),
    .B(net99));
 sg13g2_o21ai_1 _5567_ (.B1(_0786_),
    .Y(_0168_),
    .A1(net99),
    .A2(net60));
 sg13g2_buf_1 _5568_ (.A(_4304_),
    .X(_0787_));
 sg13g2_nand2_1 _5569_ (.Y(_0788_),
    .A(net105),
    .B(_0787_));
 sg13g2_nor2_1 _5570_ (.A(_4333_),
    .B(_0788_),
    .Y(_0789_));
 sg13g2_nand2_1 _5571_ (.Y(_0790_),
    .A(_0789_),
    .B(net104));
 sg13g2_nor2_1 _5572_ (.A(net106),
    .B(_0790_),
    .Y(_0791_));
 sg13g2_nand2_1 _5573_ (.Y(_0792_),
    .A(_0791_),
    .B(_4315_));
 sg13g2_nor2_1 _5574_ (.A(_4359_),
    .B(_0792_),
    .Y(_0793_));
 sg13g2_xnor2_1 _5575_ (.Y(_0794_),
    .A(_4378_),
    .B(_0793_));
 sg13g2_nand2_1 _5576_ (.Y(_0795_),
    .A(net64),
    .B(_4318_));
 sg13g2_o21ai_1 _5577_ (.B1(_0795_),
    .Y(_0169_),
    .A1(_0794_),
    .A2(net60));
 sg13g2_nor2_1 _5578_ (.A(net107),
    .B(_4324_),
    .Y(_0796_));
 sg13g2_inv_1 _5579_ (.Y(_0797_),
    .A(_0796_));
 sg13g2_nand2_1 _5580_ (.Y(_0798_),
    .A(_0797_),
    .B(_4333_));
 sg13g2_nand2_1 _5581_ (.Y(_0799_),
    .A(net64),
    .B(_4332_));
 sg13g2_o21ai_1 _5582_ (.B1(_0799_),
    .Y(_0170_),
    .A1(_0798_),
    .A2(net60));
 sg13g2_xnor2_1 _5583_ (.Y(_0800_),
    .A(_0058_),
    .B(_4333_));
 sg13g2_nand2_1 _5584_ (.Y(_0801_),
    .A(net64),
    .B(net96));
 sg13g2_o21ai_1 _5585_ (.B1(_0801_),
    .Y(_0171_),
    .A1(_0800_),
    .A2(_0785_));
 sg13g2_buf_2 _5586_ (.A(_0024_),
    .X(_0802_));
 sg13g2_inv_1 _5587_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_xnor2_1 _5588_ (.Y(_0804_),
    .A(_0803_),
    .B(_4334_));
 sg13g2_nand2_1 _5589_ (.Y(_0805_),
    .A(net64),
    .B(_4346_));
 sg13g2_o21ai_1 _5590_ (.B1(_0805_),
    .Y(_0172_),
    .A1(_0804_),
    .A2(net60));
 sg13g2_inv_2 _5591_ (.Y(_0806_),
    .A(_0014_));
 sg13g2_xnor2_1 _5592_ (.Y(_0807_),
    .A(_0806_),
    .B(_0789_));
 sg13g2_nand2_1 _5593_ (.Y(_0808_),
    .A(_0411_),
    .B(net104));
 sg13g2_o21ai_1 _5594_ (.B1(_0808_),
    .Y(_0173_),
    .A1(_0807_),
    .A2(_0785_));
 sg13g2_xnor2_1 _5595_ (.Y(_0809_),
    .A(_0029_),
    .B(_0790_));
 sg13g2_nand2_1 _5596_ (.Y(_0810_),
    .A(_0411_),
    .B(net103));
 sg13g2_o21ai_1 _5597_ (.B1(_0810_),
    .Y(_0174_),
    .A1(_0809_),
    .A2(net60));
 sg13g2_inv_1 _5598_ (.Y(_0811_),
    .A(_0059_));
 sg13g2_xnor2_1 _5599_ (.Y(_0812_),
    .A(_0811_),
    .B(_0791_));
 sg13g2_buf_1 _5600_ (.A(_4300_),
    .X(_0813_));
 sg13g2_nand2_1 _5601_ (.Y(_0814_),
    .A(_0410_),
    .B(net95));
 sg13g2_o21ai_1 _5602_ (.B1(_0814_),
    .Y(_0175_),
    .A1(_0812_),
    .A2(net60));
 sg13g2_inv_1 _5603_ (.Y(_0815_),
    .A(_0034_));
 sg13g2_nor2_1 _5604_ (.A(_4370_),
    .B(_0790_),
    .Y(_0816_));
 sg13g2_xnor2_1 _5605_ (.Y(_0817_),
    .A(_0815_),
    .B(_0816_));
 sg13g2_buf_1 _5606_ (.A(_4313_),
    .X(_0818_));
 sg13g2_nand2_1 _5607_ (.Y(_0819_),
    .A(_0410_),
    .B(net94));
 sg13g2_o21ai_1 _5608_ (.B1(_0819_),
    .Y(_0176_),
    .A1(_0817_),
    .A2(net60));
 sg13g2_nand2_1 _5609_ (.Y(_0820_),
    .A(_0816_),
    .B(net94));
 sg13g2_xnor2_1 _5610_ (.Y(_0821_),
    .A(_0037_),
    .B(_0820_));
 sg13g2_nand2_1 _5611_ (.Y(_0822_),
    .A(_0410_),
    .B(_4312_));
 sg13g2_o21ai_1 _5612_ (.B1(_0822_),
    .Y(_0177_),
    .A1(_0821_),
    .A2(net60));
 sg13g2_xnor2_1 _5613_ (.Y(_0823_),
    .A(_0060_),
    .B(_0792_));
 sg13g2_nand2_1 _5614_ (.Y(_0824_),
    .A(_0410_),
    .B(_4317_));
 sg13g2_o21ai_1 _5615_ (.B1(_0824_),
    .Y(_0178_),
    .A1(_0823_),
    .A2(_0784_));
 sg13g2_nor2_1 _5616_ (.A(_0533_),
    .B(_4490_),
    .Y(_0825_));
 sg13g2_buf_1 _5617_ (.A(\vgademo.linelfsr[1] ),
    .X(_0826_));
 sg13g2_inv_1 _5618_ (.Y(_0827_),
    .A(net115));
 sg13g2_buf_1 _5619_ (.A(\vgademo.linelfsr[0] ),
    .X(_0828_));
 sg13g2_buf_1 _5620_ (.A(_0828_),
    .X(_0829_));
 sg13g2_inv_1 _5621_ (.Y(_0830_),
    .A(net93));
 sg13g2_nor2_1 _5622_ (.A(_0549_),
    .B(_0825_),
    .Y(_0831_));
 sg13g2_buf_1 _5623_ (.A(_0831_),
    .X(_0832_));
 sg13g2_nor3_1 _5624_ (.A(_0827_),
    .B(_0830_),
    .C(_0832_),
    .Y(_0833_));
 sg13g2_inv_1 _5625_ (.Y(_0834_),
    .A(_0832_));
 sg13g2_a21oi_1 _5626_ (.A1(_0834_),
    .A2(net115),
    .Y(_0835_),
    .B1(_0829_));
 sg13g2_nor3_1 _5627_ (.A(_0825_),
    .B(_0833_),
    .C(_0835_),
    .Y(_0181_));
 sg13g2_inv_1 _5628_ (.Y(_0836_),
    .A(\vgademo.linelfsr[11] ));
 sg13g2_buf_1 _5629_ (.A(_0832_),
    .X(_0837_));
 sg13g2_nand2_1 _5630_ (.Y(_0838_),
    .A(net39),
    .B(\vgademo.linelfsr[10] ));
 sg13g2_o21ai_1 _5631_ (.B1(_0838_),
    .Y(_0182_),
    .A1(_0836_),
    .A2(_0551_));
 sg13g2_inv_1 _5632_ (.Y(_0839_),
    .A(\vgademo.linelfsr[12] ));
 sg13g2_a22oi_1 _5633_ (.Y(_0183_),
    .B1(_0836_),
    .B2(_0837_),
    .A2(net55),
    .A1(_0839_));
 sg13g2_a22oi_1 _5634_ (.Y(_0184_),
    .B1(_0839_),
    .B2(_0837_),
    .A2(net55),
    .A1(_0830_));
 sg13g2_inv_1 _5635_ (.Y(_0840_),
    .A(\vgademo.linelfsr[2] ));
 sg13g2_a22oi_1 _5636_ (.Y(_0185_),
    .B1(_0827_),
    .B2(net39),
    .A2(net55),
    .A1(_0840_));
 sg13g2_inv_1 _5637_ (.Y(_0841_),
    .A(\vgademo.linelfsr[3] ));
 sg13g2_nand2_1 _5638_ (.Y(_0842_),
    .A(_0832_),
    .B(\vgademo.linelfsr[2] ));
 sg13g2_o21ai_1 _5639_ (.B1(_0842_),
    .Y(_0186_),
    .A1(_0841_),
    .A2(_0551_));
 sg13g2_xnor2_1 _5640_ (.Y(_0843_),
    .A(net93),
    .B(\vgademo.linelfsr[4] ));
 sg13g2_a22oi_1 _5641_ (.Y(_0187_),
    .B1(_0841_),
    .B2(net39),
    .A2(_0843_),
    .A1(net55));
 sg13g2_xnor2_1 _5642_ (.Y(_0844_),
    .A(net93),
    .B(\vgademo.linelfsr[5] ));
 sg13g2_inv_1 _5643_ (.Y(_0845_),
    .A(\vgademo.linelfsr[4] ));
 sg13g2_a22oi_1 _5644_ (.Y(_0188_),
    .B1(_0845_),
    .B2(net39),
    .A2(_0844_),
    .A1(net55));
 sg13g2_inv_1 _5645_ (.Y(_0846_),
    .A(\vgademo.linelfsr[6] ));
 sg13g2_inv_1 _5646_ (.Y(_0847_),
    .A(\vgademo.linelfsr[5] ));
 sg13g2_a22oi_1 _5647_ (.Y(_0189_),
    .B1(_0847_),
    .B2(net39),
    .A2(net55),
    .A1(_0846_));
 sg13g2_xnor2_1 _5648_ (.Y(_0848_),
    .A(net93),
    .B(\vgademo.linelfsr[7] ));
 sg13g2_a22oi_1 _5649_ (.Y(_0190_),
    .B1(_0846_),
    .B2(net39),
    .A2(_0848_),
    .A1(_0550_));
 sg13g2_inv_1 _5650_ (.Y(_0849_),
    .A(\vgademo.linelfsr[8] ));
 sg13g2_inv_1 _5651_ (.Y(_0850_),
    .A(\vgademo.linelfsr[7] ));
 sg13g2_a22oi_1 _5652_ (.Y(_0191_),
    .B1(_0850_),
    .B2(net39),
    .A2(_0550_),
    .A1(_0849_));
 sg13g2_xnor2_1 _5653_ (.Y(_0851_),
    .A(net93),
    .B(\vgademo.linelfsr[9] ));
 sg13g2_nand2_1 _5654_ (.Y(_0852_),
    .A(_0832_),
    .B(\vgademo.linelfsr[8] ));
 sg13g2_o21ai_1 _5655_ (.B1(_0852_),
    .Y(_0192_),
    .A1(_0551_),
    .A2(_0851_));
 sg13g2_inv_1 _5656_ (.Y(_0853_),
    .A(\vgademo.linelfsr[10] ));
 sg13g2_inv_1 _5657_ (.Y(_0854_),
    .A(\vgademo.linelfsr[9] ));
 sg13g2_a22oi_1 _5658_ (.Y(_0193_),
    .B1(_0854_),
    .B2(net39),
    .A2(net55),
    .A1(_0853_));
 sg13g2_buf_1 _5659_ (.A(\vgademo.plane_dx[0] ),
    .X(_0855_));
 sg13g2_inv_1 _5660_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_nor2_1 _5661_ (.A(_4285_),
    .B(_4428_),
    .Y(_0857_));
 sg13g2_nand4_1 _5662_ (.B(_4278_),
    .C(_4471_),
    .A(_4473_),
    .Y(_0858_),
    .D(_0857_));
 sg13g2_nor4_1 _5663_ (.A(net127),
    .B(net126),
    .C(_0533_),
    .D(_0858_),
    .Y(_0859_));
 sg13g2_buf_2 _5664_ (.A(_0859_),
    .X(_0860_));
 sg13g2_buf_1 _5665_ (.A(_0860_),
    .X(_0861_));
 sg13g2_buf_1 _5666_ (.A(_0860_),
    .X(_0862_));
 sg13g2_nor2_1 _5667_ (.A(\vgademo.plane_du[0] ),
    .B(net67),
    .Y(_0863_));
 sg13g2_a21oi_1 _5668_ (.A1(_0856_),
    .A2(net68),
    .Y(_0194_),
    .B1(_0863_));
 sg13g2_buf_1 _5669_ (.A(\vgademo.plane_dx_div.q[9] ),
    .X(_0864_));
 sg13g2_inv_1 _5670_ (.Y(_0865_),
    .A(net114));
 sg13g2_buf_1 _5671_ (.A(\vgademo.plane_du[10] ),
    .X(_0866_));
 sg13g2_nor2_1 _5672_ (.A(_0866_),
    .B(_0862_),
    .Y(_0867_));
 sg13g2_a21oi_1 _5673_ (.A1(_0865_),
    .A2(net68),
    .Y(_0195_),
    .B1(_0867_));
 sg13g2_buf_1 _5674_ (.A(\vgademo.plane_dx[1] ),
    .X(_0868_));
 sg13g2_inv_1 _5675_ (.Y(_0869_),
    .A(_0868_));
 sg13g2_buf_1 _5676_ (.A(_0860_),
    .X(_0870_));
 sg13g2_nor2_1 _5677_ (.A(\vgademo.plane_du[1] ),
    .B(net66),
    .Y(_0871_));
 sg13g2_a21oi_1 _5678_ (.A1(_0869_),
    .A2(net68),
    .Y(_0196_),
    .B1(_0871_));
 sg13g2_buf_1 _5679_ (.A(\vgademo.plane_dx[2] ),
    .X(_0872_));
 sg13g2_inv_1 _5680_ (.Y(_0873_),
    .A(_0872_));
 sg13g2_nor2_1 _5681_ (.A(\vgademo.plane_du[2] ),
    .B(_0870_),
    .Y(_0874_));
 sg13g2_a21oi_1 _5682_ (.A1(_0873_),
    .A2(net68),
    .Y(_0197_),
    .B1(_0874_));
 sg13g2_buf_1 _5683_ (.A(\vgademo.plane_dx_div.q[2] ),
    .X(_0875_));
 sg13g2_inv_1 _5684_ (.Y(_0876_),
    .A(net112));
 sg13g2_buf_1 _5685_ (.A(\vgademo.plane_du[3] ),
    .X(_0877_));
 sg13g2_nor2_1 _5686_ (.A(_0877_),
    .B(_0870_),
    .Y(_0878_));
 sg13g2_a21oi_1 _5687_ (.A1(_0876_),
    .A2(_0861_),
    .Y(_0198_),
    .B1(_0878_));
 sg13g2_buf_2 _5688_ (.A(\vgademo.plane_dx_div.q[3] ),
    .X(_0879_));
 sg13g2_inv_1 _5689_ (.Y(_0880_),
    .A(_0879_));
 sg13g2_buf_2 _5690_ (.A(\vgademo.plane_du[4] ),
    .X(_0881_));
 sg13g2_nor2_1 _5691_ (.A(_0881_),
    .B(net66),
    .Y(_0882_));
 sg13g2_a21oi_1 _5692_ (.A1(_0880_),
    .A2(_0861_),
    .Y(_0199_),
    .B1(_0882_));
 sg13g2_buf_2 _5693_ (.A(\vgademo.plane_dx_div.q[4] ),
    .X(_0883_));
 sg13g2_inv_1 _5694_ (.Y(_0884_),
    .A(_0883_));
 sg13g2_buf_2 _5695_ (.A(\vgademo.plane_du[5] ),
    .X(_0885_));
 sg13g2_nor2_1 _5696_ (.A(_0885_),
    .B(net66),
    .Y(_0886_));
 sg13g2_a21oi_1 _5697_ (.A1(_0884_),
    .A2(net68),
    .Y(_0200_),
    .B1(_0886_));
 sg13g2_buf_2 _5698_ (.A(\vgademo.plane_dx_div.q[5] ),
    .X(_0887_));
 sg13g2_inv_1 _5699_ (.Y(_0888_),
    .A(_0887_));
 sg13g2_buf_2 _5700_ (.A(\vgademo.plane_du[6] ),
    .X(_0889_));
 sg13g2_nor2_1 _5701_ (.A(_0889_),
    .B(net66),
    .Y(_0890_));
 sg13g2_a21oi_1 _5702_ (.A1(_0888_),
    .A2(net68),
    .Y(_0201_),
    .B1(_0890_));
 sg13g2_buf_2 _5703_ (.A(\vgademo.plane_dx_div.q[6] ),
    .X(_0891_));
 sg13g2_inv_1 _5704_ (.Y(_0892_),
    .A(_0891_));
 sg13g2_buf_2 _5705_ (.A(\vgademo.plane_du[7] ),
    .X(_0893_));
 sg13g2_nor2_1 _5706_ (.A(_0893_),
    .B(net66),
    .Y(_0894_));
 sg13g2_a21oi_1 _5707_ (.A1(_0892_),
    .A2(net68),
    .Y(_0202_),
    .B1(_0894_));
 sg13g2_buf_2 _5708_ (.A(\vgademo.plane_dx_div.q[7] ),
    .X(_0895_));
 sg13g2_inv_1 _5709_ (.Y(_0896_),
    .A(_0895_));
 sg13g2_buf_1 _5710_ (.A(\vgademo.plane_du[8] ),
    .X(_0897_));
 sg13g2_nor2_1 _5711_ (.A(_0897_),
    .B(net66),
    .Y(_0898_));
 sg13g2_a21oi_1 _5712_ (.A1(_0896_),
    .A2(net68),
    .Y(_0203_),
    .B1(_0898_));
 sg13g2_buf_1 _5713_ (.A(\vgademo.plane_dx_div.q[8] ),
    .X(_0899_));
 sg13g2_inv_1 _5714_ (.Y(_0900_),
    .A(net110));
 sg13g2_buf_2 _5715_ (.A(\vgademo.plane_du[9] ),
    .X(_0901_));
 sg13g2_nor2_1 _5716_ (.A(_0901_),
    .B(net66),
    .Y(_0902_));
 sg13g2_a21oi_1 _5717_ (.A1(_0900_),
    .A2(_0862_),
    .Y(_0204_),
    .B1(_0902_));
 sg13g2_inv_1 _5718_ (.Y(_0903_),
    .A(\vgademo.plane_dx_div.d[17] ));
 sg13g2_inv_2 _5719_ (.Y(_0904_),
    .A(_4298_));
 sg13g2_buf_1 _5720_ (.A(_0904_),
    .X(_0905_));
 sg13g2_nand2_1 _5721_ (.Y(_0906_),
    .A(_4363_),
    .B(_4323_));
 sg13g2_nand3_1 _5722_ (.B(_4329_),
    .C(_4319_),
    .A(_4316_),
    .Y(_0907_));
 sg13g2_buf_8 _5723_ (.A(_0907_),
    .X(_0908_));
 sg13g2_nand2_1 _5724_ (.Y(_0909_),
    .A(_0906_),
    .B(_0908_));
 sg13g2_a21oi_1 _5725_ (.A1(_4331_),
    .A2(_0017_),
    .Y(_0910_),
    .B1(_4386_));
 sg13g2_nand2_1 _5726_ (.Y(_0911_),
    .A(_0909_),
    .B(_0910_));
 sg13g2_inv_2 _5727_ (.Y(_0912_),
    .A(_0911_));
 sg13g2_nand2_1 _5728_ (.Y(_0913_),
    .A(_0912_),
    .B(_4457_));
 sg13g2_nand2_1 _5729_ (.Y(_0914_),
    .A(_0911_),
    .B(_4456_));
 sg13g2_a21oi_1 _5730_ (.A1(_0913_),
    .A2(_0914_),
    .Y(_0915_),
    .B1(_0016_));
 sg13g2_nand3_1 _5731_ (.B(_0016_),
    .C(_0914_),
    .A(_0913_),
    .Y(_0916_));
 sg13g2_nand2b_1 _5732_ (.Y(_0917_),
    .B(_0916_),
    .A_N(_0915_));
 sg13g2_inv_1 _5733_ (.Y(_0918_),
    .A(_0018_));
 sg13g2_inv_1 _5734_ (.Y(_0919_),
    .A(_0077_));
 sg13g2_nor2_1 _5735_ (.A(_0919_),
    .B(_4393_),
    .Y(_0920_));
 sg13g2_a21oi_1 _5736_ (.A1(_0918_),
    .A2(_4388_),
    .Y(_0921_),
    .B1(_0920_));
 sg13g2_nor2_1 _5737_ (.A(_0917_),
    .B(_0921_),
    .Y(_0922_));
 sg13g2_inv_1 _5738_ (.Y(_0923_),
    .A(_0922_));
 sg13g2_nand2_1 _5739_ (.Y(_0924_),
    .A(_0921_),
    .B(_0917_));
 sg13g2_nand2_1 _5740_ (.Y(_0925_),
    .A(_0923_),
    .B(_0924_));
 sg13g2_inv_1 _5741_ (.Y(_0926_),
    .A(_0925_));
 sg13g2_nand2_1 _5742_ (.Y(_0927_),
    .A(_0926_),
    .B(_0904_));
 sg13g2_o21ai_1 _5743_ (.B1(_0927_),
    .Y(_0205_),
    .A1(_0903_),
    .A2(net51));
 sg13g2_buf_2 _5744_ (.A(\vgademo.audio_kick_frames[2] ),
    .X(_0928_));
 sg13g2_inv_1 _5745_ (.Y(_0929_),
    .A(_0020_));
 sg13g2_nand2_1 _5746_ (.Y(_0930_),
    .A(net107),
    .B(_4304_));
 sg13g2_nand2_1 _5747_ (.Y(_0931_),
    .A(_0760_),
    .B(_0930_));
 sg13g2_nand2b_1 _5748_ (.Y(_0932_),
    .B(_4331_),
    .A_N(_0931_));
 sg13g2_nand2_1 _5749_ (.Y(_0933_),
    .A(_4359_),
    .B(_4318_));
 sg13g2_nor2_1 _5750_ (.A(_4358_),
    .B(_0933_),
    .Y(_0934_));
 sg13g2_nand3_1 _5751_ (.B(_0934_),
    .C(_4334_),
    .A(_4350_),
    .Y(_0935_));
 sg13g2_nand3_1 _5752_ (.B(_4342_),
    .C(_4354_),
    .A(_4353_),
    .Y(_0936_));
 sg13g2_nand2_1 _5753_ (.Y(_0937_),
    .A(_0936_),
    .B(_4361_));
 sg13g2_nand2_1 _5754_ (.Y(_0938_),
    .A(_0935_),
    .B(_0937_));
 sg13g2_buf_8 _5755_ (.A(_0938_),
    .X(_0939_));
 sg13g2_nand2_1 _5756_ (.Y(_0940_),
    .A(_4336_),
    .B(_4340_));
 sg13g2_nand2_1 _5757_ (.Y(_0941_),
    .A(_0940_),
    .B(_4343_));
 sg13g2_inv_2 _5758_ (.Y(_0942_),
    .A(_4304_));
 sg13g2_nand3_1 _5759_ (.B(_0941_),
    .C(_0942_),
    .A(net65),
    .Y(_0943_));
 sg13g2_nand2_1 _5760_ (.Y(_0944_),
    .A(_0932_),
    .B(_0943_));
 sg13g2_nand2_1 _5761_ (.Y(_0945_),
    .A(_0944_),
    .B(_4385_));
 sg13g2_xnor2_1 _5762_ (.Y(_0946_),
    .A(_0929_),
    .B(_0945_));
 sg13g2_buf_1 _5763_ (.A(_0021_),
    .X(_0947_));
 sg13g2_o21ai_1 _5764_ (.B1(_0916_),
    .Y(_0948_),
    .A1(_0947_),
    .A2(_0912_));
 sg13g2_xor2_1 _5765_ (.B(_0948_),
    .A(_0946_),
    .X(_0949_));
 sg13g2_xnor2_1 _5766_ (.Y(_0950_),
    .A(_0928_),
    .B(_0949_));
 sg13g2_xnor2_1 _5767_ (.Y(_0951_),
    .A(_0923_),
    .B(_0950_));
 sg13g2_mux2_1 _5768_ (.A0(\vgademo.plane_dx_div.d[18] ),
    .A1(_0951_),
    .S(net51),
    .X(_0206_));
 sg13g2_inv_1 _5769_ (.Y(_0952_),
    .A(\vgademo.plane_dx_div.d[19] ));
 sg13g2_buf_1 _5770_ (.A(_4298_),
    .X(_0953_));
 sg13g2_nor2b_1 _5771_ (.A(_0923_),
    .B_N(_0950_),
    .Y(_0954_));
 sg13g2_xnor2_1 _5772_ (.Y(_0955_),
    .A(_0802_),
    .B(_4306_));
 sg13g2_a21oi_1 _5773_ (.A1(_4331_),
    .A2(_0955_),
    .Y(_0956_),
    .B1(_4386_));
 sg13g2_nand3_1 _5774_ (.B(_0941_),
    .C(_0803_),
    .A(net65),
    .Y(_0957_));
 sg13g2_nand2_1 _5775_ (.Y(_0958_),
    .A(_0957_),
    .B(_0908_));
 sg13g2_nand2_1 _5776_ (.Y(_0959_),
    .A(_0956_),
    .B(_0958_));
 sg13g2_inv_1 _5777_ (.Y(_0960_),
    .A(_0023_));
 sg13g2_nand2_1 _5778_ (.Y(_0961_),
    .A(_0959_),
    .B(_0960_));
 sg13g2_nand3_1 _5779_ (.B(_0958_),
    .C(_0023_),
    .A(_0956_),
    .Y(_0962_));
 sg13g2_buf_2 _5780_ (.A(_0962_),
    .X(_0963_));
 sg13g2_inv_1 _5781_ (.Y(_0964_),
    .A(_4455_));
 sg13g2_nand3_1 _5782_ (.B(_0964_),
    .C(_4385_),
    .A(_0944_),
    .Y(_0965_));
 sg13g2_inv_2 _5783_ (.Y(_0966_),
    .A(_0965_));
 sg13g2_a21oi_1 _5784_ (.A1(_0961_),
    .A2(_0963_),
    .Y(_0967_),
    .B1(_0966_));
 sg13g2_nand3_1 _5785_ (.B(_0961_),
    .C(_0963_),
    .A(_0966_),
    .Y(_0968_));
 sg13g2_nor2b_1 _5786_ (.A(_0967_),
    .B_N(_0968_),
    .Y(_0969_));
 sg13g2_nor2b_1 _5787_ (.A(_0928_),
    .B_N(_0949_),
    .Y(_0970_));
 sg13g2_a21oi_1 _5788_ (.A1(_0948_),
    .A2(_0946_),
    .Y(_0971_),
    .B1(_0970_));
 sg13g2_xnor2_1 _5789_ (.Y(_0972_),
    .A(_0969_),
    .B(_0971_));
 sg13g2_xor2_1 _5790_ (.B(_0972_),
    .A(_0954_),
    .X(_0973_));
 sg13g2_nor2_1 _5791_ (.A(net59),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_a21oi_1 _5792_ (.A1(_0952_),
    .A2(net59),
    .Y(_0207_),
    .B1(_0974_));
 sg13g2_buf_1 _5793_ (.A(\vgademo.plane_dx_div.d[20] ),
    .X(_0975_));
 sg13g2_nand2_1 _5794_ (.Y(_0976_),
    .A(_4326_),
    .B(_0017_));
 sg13g2_xnor2_1 _5795_ (.Y(_0977_),
    .A(_0806_),
    .B(_0976_));
 sg13g2_nor2_1 _5796_ (.A(_0977_),
    .B(_0908_),
    .Y(_0978_));
 sg13g2_nor2_1 _5797_ (.A(_4386_),
    .B(_0978_),
    .Y(_0979_));
 sg13g2_nand2_1 _5798_ (.Y(_0980_),
    .A(_4339_),
    .B(_4354_));
 sg13g2_o21ai_1 _5799_ (.B1(net65),
    .Y(_0981_),
    .A1(_0980_),
    .A2(_4345_));
 sg13g2_nand2_1 _5800_ (.Y(_0982_),
    .A(_0979_),
    .B(_0981_));
 sg13g2_inv_1 _5801_ (.Y(_0983_),
    .A(_0027_));
 sg13g2_nand2_1 _5802_ (.Y(_0984_),
    .A(_0982_),
    .B(_0983_));
 sg13g2_nand3_1 _5803_ (.B(_0027_),
    .C(_0981_),
    .A(_0979_),
    .Y(_0985_));
 sg13g2_nand2_1 _5804_ (.Y(_0986_),
    .A(_0984_),
    .B(_0985_));
 sg13g2_xnor2_1 _5805_ (.Y(_0987_),
    .A(_0963_),
    .B(_0986_));
 sg13g2_xnor2_1 _5806_ (.Y(_0988_),
    .A(_0967_),
    .B(_0987_));
 sg13g2_nor2b_1 _5807_ (.A(_0971_),
    .B_N(_0969_),
    .Y(_0989_));
 sg13g2_a21o_1 _5808_ (.A2(_0954_),
    .A1(_0972_),
    .B1(_0989_),
    .X(_0990_));
 sg13g2_xor2_1 _5809_ (.B(_0990_),
    .A(_0988_),
    .X(_0991_));
 sg13g2_mux2_1 _5810_ (.A0(_0975_),
    .A1(_0991_),
    .S(_0904_),
    .X(_0208_));
 sg13g2_buf_1 _5811_ (.A(\vgademo.plane_dx_div.d[21] ),
    .X(_0992_));
 sg13g2_inv_1 _5812_ (.Y(_0993_),
    .A(_0992_));
 sg13g2_nand2_1 _5813_ (.Y(_0994_),
    .A(_0986_),
    .B(_0963_));
 sg13g2_inv_1 _5814_ (.Y(_0995_),
    .A(_0985_));
 sg13g2_inv_1 _5815_ (.Y(_0996_),
    .A(_0029_));
 sg13g2_nand2_1 _5816_ (.Y(_0997_),
    .A(_4306_),
    .B(_4347_));
 sg13g2_nand2_1 _5817_ (.Y(_0998_),
    .A(_0997_),
    .B(_4348_));
 sg13g2_xnor2_1 _5818_ (.Y(_0999_),
    .A(_0996_),
    .B(_0998_));
 sg13g2_nor2_1 _5819_ (.A(_0999_),
    .B(_0908_),
    .Y(_1000_));
 sg13g2_nor2_1 _5820_ (.A(_4386_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nor2_1 _5821_ (.A(net106),
    .B(_4310_),
    .Y(_1002_));
 sg13g2_a21oi_1 _5822_ (.A1(_4347_),
    .A2(_4321_),
    .Y(_1003_),
    .B1(_1002_));
 sg13g2_nand2_1 _5823_ (.Y(_1004_),
    .A(_0941_),
    .B(_1003_));
 sg13g2_nand2_1 _5824_ (.Y(_1005_),
    .A(_1004_),
    .B(net65));
 sg13g2_nand2_1 _5825_ (.Y(_1006_),
    .A(_1005_),
    .B(_0908_));
 sg13g2_nand2_1 _5826_ (.Y(_1007_),
    .A(_1001_),
    .B(_1006_));
 sg13g2_xnor2_1 _5827_ (.Y(_1008_),
    .A(_4448_),
    .B(_1007_));
 sg13g2_xnor2_1 _5828_ (.Y(_1009_),
    .A(_0995_),
    .B(_1008_));
 sg13g2_xnor2_1 _5829_ (.Y(_1010_),
    .A(_0994_),
    .B(_1009_));
 sg13g2_nor2b_1 _5830_ (.A(_0987_),
    .B_N(_0967_),
    .Y(_1011_));
 sg13g2_a21o_1 _5831_ (.A2(_0988_),
    .A1(_0990_),
    .B1(_1011_),
    .X(_1012_));
 sg13g2_xor2_1 _5832_ (.B(_1012_),
    .A(_1010_),
    .X(_1013_));
 sg13g2_nor2_1 _5833_ (.A(net59),
    .B(_1013_),
    .Y(_1014_));
 sg13g2_a21oi_1 _5834_ (.A1(_0993_),
    .A2(net59),
    .Y(_0209_),
    .B1(_1014_));
 sg13g2_nand2_1 _5835_ (.Y(_1015_),
    .A(_1008_),
    .B(_0995_));
 sg13g2_buf_1 _5836_ (.A(_0032_),
    .X(_1016_));
 sg13g2_nand2_1 _5837_ (.Y(_1017_),
    .A(_1007_),
    .B(_1016_));
 sg13g2_buf_1 _5838_ (.A(_4301_),
    .X(_1018_));
 sg13g2_nand2_1 _5839_ (.Y(_1019_),
    .A(net104),
    .B(net103));
 sg13g2_nand2b_1 _5840_ (.Y(_1020_),
    .B(_0976_),
    .A_N(_1019_));
 sg13g2_xnor2_1 _5841_ (.Y(_1021_),
    .A(net83),
    .B(_1020_));
 sg13g2_nor2_1 _5842_ (.A(_1021_),
    .B(_0908_),
    .Y(_1022_));
 sg13g2_nor2_1 _5843_ (.A(_4386_),
    .B(_1022_),
    .Y(_1023_));
 sg13g2_a21oi_1 _5844_ (.A1(_4321_),
    .A2(_0802_),
    .Y(_1024_),
    .B1(net83));
 sg13g2_nand3_1 _5845_ (.B(_4301_),
    .C(_0802_),
    .A(_4321_),
    .Y(_1025_));
 sg13g2_nor2b_1 _5846_ (.A(_1024_),
    .B_N(_1025_),
    .Y(_1026_));
 sg13g2_nand2_1 _5847_ (.Y(_1027_),
    .A(_0941_),
    .B(_1026_));
 sg13g2_nand2_1 _5848_ (.Y(_1028_),
    .A(_1027_),
    .B(_0938_));
 sg13g2_nand2_1 _5849_ (.Y(_1029_),
    .A(_1028_),
    .B(_0908_));
 sg13g2_nand2_1 _5850_ (.Y(_1030_),
    .A(_1023_),
    .B(_1029_));
 sg13g2_buf_2 _5851_ (.A(_0031_),
    .X(_1031_));
 sg13g2_nand2_1 _5852_ (.Y(_1032_),
    .A(_1030_),
    .B(_1031_));
 sg13g2_inv_1 _5853_ (.Y(_1033_),
    .A(_1031_));
 sg13g2_nand3_1 _5854_ (.B(_1029_),
    .C(_1033_),
    .A(_1023_),
    .Y(_1034_));
 sg13g2_nand2_1 _5855_ (.Y(_1035_),
    .A(_1032_),
    .B(_1034_));
 sg13g2_xnor2_1 _5856_ (.Y(_1036_),
    .A(_1017_),
    .B(_1035_));
 sg13g2_nor2b_1 _5857_ (.A(_1015_),
    .B_N(_1036_),
    .Y(_1037_));
 sg13g2_nand2b_1 _5858_ (.Y(_1038_),
    .B(_1015_),
    .A_N(_1036_));
 sg13g2_nand2b_1 _5859_ (.Y(_1039_),
    .B(_1038_),
    .A_N(_1037_));
 sg13g2_nor2b_1 _5860_ (.A(_0994_),
    .B_N(_1009_),
    .Y(_1040_));
 sg13g2_a21oi_1 _5861_ (.A1(_1012_),
    .A2(_1010_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_xnor2_1 _5862_ (.Y(_1042_),
    .A(_1039_),
    .B(_1041_));
 sg13g2_buf_1 _5863_ (.A(\vgademo.plane_dx_div.d[22] ),
    .X(_1043_));
 sg13g2_nor2_1 _5864_ (.A(_1043_),
    .B(_0904_),
    .Y(_1044_));
 sg13g2_a21oi_1 _5865_ (.A1(_1042_),
    .A2(net51),
    .Y(_0210_),
    .B1(_1044_));
 sg13g2_inv_1 _5866_ (.Y(_1045_),
    .A(\vgademo.plane_dx_div.d[23] ));
 sg13g2_nand2_1 _5867_ (.Y(_1046_),
    .A(_1035_),
    .B(_1017_));
 sg13g2_nor2_1 _5868_ (.A(_0014_),
    .B(net106),
    .Y(_1047_));
 sg13g2_a21oi_1 _5869_ (.A1(_4367_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(net95));
 sg13g2_xnor2_1 _5870_ (.Y(_1049_),
    .A(_0034_),
    .B(_1048_));
 sg13g2_a21oi_1 _5871_ (.A1(_1049_),
    .A2(_4331_),
    .Y(_1050_),
    .B1(_4386_));
 sg13g2_xnor2_1 _5872_ (.Y(_1051_),
    .A(_0815_),
    .B(_4340_));
 sg13g2_o21ai_1 _5873_ (.B1(net65),
    .Y(_1052_),
    .A1(_1051_),
    .A2(_4345_));
 sg13g2_nand2_1 _5874_ (.Y(_1053_),
    .A(_1052_),
    .B(_0908_));
 sg13g2_nand2_1 _5875_ (.Y(_1054_),
    .A(_1050_),
    .B(_1053_));
 sg13g2_xnor2_1 _5876_ (.Y(_1055_),
    .A(net121),
    .B(_1054_));
 sg13g2_xor2_1 _5877_ (.B(_1055_),
    .A(_1032_),
    .X(_1056_));
 sg13g2_nor2_1 _5878_ (.A(_1046_),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nand2_1 _5879_ (.Y(_1058_),
    .A(_1056_),
    .B(_1046_));
 sg13g2_nor2b_1 _5880_ (.A(_1057_),
    .B_N(_1058_),
    .Y(_1059_));
 sg13g2_a21oi_1 _5881_ (.A1(_1041_),
    .A2(_1038_),
    .Y(_1060_),
    .B1(_1037_));
 sg13g2_xor2_1 _5882_ (.B(_1060_),
    .A(_1059_),
    .X(_1061_));
 sg13g2_nor2_1 _5883_ (.A(net59),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_a21oi_1 _5884_ (.A1(_1045_),
    .A2(net59),
    .Y(_0211_),
    .B1(_1062_));
 sg13g2_nor2b_1 _5885_ (.A(_1055_),
    .B_N(_1032_),
    .Y(_1063_));
 sg13g2_nand2_1 _5886_ (.Y(_1064_),
    .A(_1025_),
    .B(_4313_));
 sg13g2_xor2_1 _5887_ (.B(_1064_),
    .A(_0037_),
    .X(_1065_));
 sg13g2_nand2_1 _5888_ (.Y(_1066_),
    .A(_4363_),
    .B(_1065_));
 sg13g2_nand2_1 _5889_ (.Y(_1067_),
    .A(_1020_),
    .B(net83));
 sg13g2_nand3_1 _5890_ (.B(_4312_),
    .C(net94),
    .A(_1067_),
    .Y(_1068_));
 sg13g2_nand2_1 _5891_ (.Y(_1069_),
    .A(_4331_),
    .B(_1068_));
 sg13g2_nand2_1 _5892_ (.Y(_1070_),
    .A(_1066_),
    .B(_1069_));
 sg13g2_buf_1 _5893_ (.A(_0036_),
    .X(_1071_));
 sg13g2_nand2_1 _5894_ (.Y(_1072_),
    .A(_1070_),
    .B(_1071_));
 sg13g2_inv_1 _5895_ (.Y(_1073_),
    .A(_1071_));
 sg13g2_nand3_1 _5896_ (.B(_1069_),
    .C(_1073_),
    .A(_1066_),
    .Y(_1074_));
 sg13g2_nand2_1 _5897_ (.Y(_1075_),
    .A(_1072_),
    .B(_1074_));
 sg13g2_buf_2 _5898_ (.A(_0038_),
    .X(_1076_));
 sg13g2_nand2_1 _5899_ (.Y(_1077_),
    .A(_1054_),
    .B(_1076_));
 sg13g2_xor2_1 _5900_ (.B(_1077_),
    .A(_1075_),
    .X(_1078_));
 sg13g2_xnor2_1 _5901_ (.Y(_1079_),
    .A(_1063_),
    .B(_1078_));
 sg13g2_o21ai_1 _5902_ (.B1(_1058_),
    .Y(_1080_),
    .A1(_1057_),
    .A2(_1060_));
 sg13g2_xnor2_1 _5903_ (.Y(_1081_),
    .A(_1079_),
    .B(_1080_));
 sg13g2_nor2_1 _5904_ (.A(\vgademo.plane_dx_div.d[24] ),
    .B(_0904_),
    .Y(_1082_));
 sg13g2_a21oi_1 _5905_ (.A1(_1081_),
    .A2(net51),
    .Y(_0212_),
    .B1(_1082_));
 sg13g2_inv_1 _5906_ (.Y(_1083_),
    .A(\vgademo.plane_dx_div.r[16] ));
 sg13g2_nor2_1 _5907_ (.A(\vgademo.plane_dx_div.i[1] ),
    .B(\vgademo.plane_dx_div.i[0] ),
    .Y(_1084_));
 sg13g2_inv_1 _5908_ (.Y(_1085_),
    .A(\vgademo.plane_dx_div.i[3] ));
 sg13g2_nand3b_1 _5909_ (.B(_1084_),
    .C(_1085_),
    .Y(_1086_),
    .A_N(\vgademo.plane_dx_div.i[2] ));
 sg13g2_nor2_1 _5910_ (.A(_1086_),
    .B(_0904_),
    .Y(_1087_));
 sg13g2_buf_1 _5911_ (.A(_1087_),
    .X(_1088_));
 sg13g2_buf_1 _5912_ (.A(net40),
    .X(_1089_));
 sg13g2_nor2_1 _5913_ (.A(net40),
    .B(_0013_),
    .Y(_1090_));
 sg13g2_a21oi_1 _5914_ (.A1(_1083_),
    .A2(_1089_),
    .Y(_0227_),
    .B1(_1090_));
 sg13g2_inv_1 _5915_ (.Y(_1091_),
    .A(\vgademo.plane_dx_div.r[17] ));
 sg13g2_buf_2 _5916_ (.A(\vgademo.plane_dx_div.r[25] ),
    .X(_1092_));
 sg13g2_nor2_1 _5917_ (.A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ),
    .Y(_1093_));
 sg13g2_inv_1 _5918_ (.Y(_1094_),
    .A(_1093_));
 sg13g2_nand2_1 _5919_ (.Y(_1095_),
    .A(\vgademo.plane_dx_div.d[16] ),
    .B(\vgademo.plane_dx_div.d[17] ));
 sg13g2_a21oi_1 _5920_ (.A1(_1094_),
    .A2(_1095_),
    .Y(_1096_),
    .B1(_1092_));
 sg13g2_a21o_1 _5921_ (.A2(_1092_),
    .A1(_0019_),
    .B1(_1096_),
    .X(_1097_));
 sg13g2_xnor2_1 _5922_ (.Y(_1098_),
    .A(_1083_),
    .B(_1097_));
 sg13g2_nand2_1 _5923_ (.Y(_1099_),
    .A(_4298_),
    .B(_1086_));
 sg13g2_buf_1 _5924_ (.A(_1099_),
    .X(_1100_));
 sg13g2_inv_2 _5925_ (.Y(_1101_),
    .A(net50));
 sg13g2_a21oi_1 _5926_ (.A1(_1098_),
    .A2(_1101_),
    .Y(_1102_),
    .B1(_4396_));
 sg13g2_a22oi_1 _5927_ (.Y(_1103_),
    .B1(_1102_),
    .B2(_0927_),
    .A2(_0926_),
    .A1(_4396_));
 sg13g2_a21oi_1 _5928_ (.A1(_1091_),
    .A2(net38),
    .Y(_0228_),
    .B1(_1103_));
 sg13g2_nor2_1 _5929_ (.A(_1083_),
    .B(_1097_),
    .Y(_1104_));
 sg13g2_inv_1 _5930_ (.Y(_1105_),
    .A(_1092_));
 sg13g2_a21oi_1 _5931_ (.A1(_1094_),
    .A2(\vgademo.plane_dx_div.d[18] ),
    .Y(_1106_),
    .B1(_1092_));
 sg13g2_nor2_1 _5932_ (.A(\vgademo.plane_dx_div.d[18] ),
    .B(_1094_),
    .Y(_1107_));
 sg13g2_inv_1 _5933_ (.Y(_1108_),
    .A(_1107_));
 sg13g2_nand2_1 _5934_ (.Y(_1109_),
    .A(_1106_),
    .B(_1108_));
 sg13g2_o21ai_1 _5935_ (.B1(_1109_),
    .Y(_1110_),
    .A1(_1105_),
    .A2(_0022_));
 sg13g2_xnor2_1 _5936_ (.Y(_1111_),
    .A(\vgademo.plane_dx_div.r[17] ),
    .B(_1110_));
 sg13g2_xor2_1 _5937_ (.B(_1111_),
    .A(_1104_),
    .X(_1112_));
 sg13g2_nor2_1 _5938_ (.A(_4395_),
    .B(_0925_),
    .Y(_1113_));
 sg13g2_xnor2_1 _5939_ (.Y(_1114_),
    .A(_1113_),
    .B(_0951_));
 sg13g2_inv_2 _5940_ (.Y(_1115_),
    .A(net40));
 sg13g2_nor2_1 _5941_ (.A(\vgademo.plane_dx_div.r[18] ),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_a221oi_1 _5942_ (.B2(net51),
    .C1(_1116_),
    .B1(_1114_),
    .A1(_1101_),
    .Y(_0229_),
    .A2(_1112_));
 sg13g2_inv_1 _5943_ (.Y(_1117_),
    .A(\vgademo.plane_dx_div.r[19] ));
 sg13g2_nand3b_1 _5944_ (.B(_0903_),
    .C(_0026_),
    .Y(_1118_),
    .A_N(\vgademo.plane_dx_div.d[18] ));
 sg13g2_a21oi_1 _5945_ (.A1(_1118_),
    .A2(\vgademo.plane_dx_div.d[19] ),
    .Y(_1119_),
    .B1(_1092_));
 sg13g2_nand2b_1 _5946_ (.Y(_1120_),
    .B(_0952_),
    .A_N(_1118_));
 sg13g2_nand2_1 _5947_ (.Y(_1121_),
    .A(_1119_),
    .B(_1120_));
 sg13g2_o21ai_1 _5948_ (.B1(_1121_),
    .Y(_1122_),
    .A1(_1105_),
    .A2(_0025_));
 sg13g2_xnor2_1 _5949_ (.Y(_1123_),
    .A(\vgademo.plane_dx_div.r[18] ),
    .B(_1122_));
 sg13g2_nor2b_1 _5950_ (.A(_1111_),
    .B_N(_1104_),
    .Y(_1124_));
 sg13g2_a21oi_1 _5951_ (.A1(\vgademo.plane_dx_div.r[17] ),
    .A2(_1110_),
    .Y(_1125_),
    .B1(_1124_));
 sg13g2_xnor2_1 _5952_ (.Y(_1126_),
    .A(_1123_),
    .B(_1125_));
 sg13g2_nor2_1 _5953_ (.A(_1113_),
    .B(_0951_),
    .Y(_1127_));
 sg13g2_inv_1 _5954_ (.Y(_1128_),
    .A(_1127_));
 sg13g2_nor2_1 _5955_ (.A(_1128_),
    .B(_0973_),
    .Y(_1129_));
 sg13g2_inv_1 _5956_ (.Y(_1130_),
    .A(_1129_));
 sg13g2_nand2_1 _5957_ (.Y(_1131_),
    .A(_0973_),
    .B(_1128_));
 sg13g2_a21oi_1 _5958_ (.A1(_1130_),
    .A2(_1131_),
    .Y(_1132_),
    .B1(net59));
 sg13g2_a221oi_1 _5959_ (.B2(_1126_),
    .C1(_1132_),
    .B1(_1101_),
    .A1(_1117_),
    .Y(_0230_),
    .A2(net38));
 sg13g2_buf_1 _5960_ (.A(_1105_),
    .X(_1133_));
 sg13g2_nor2_1 _5961_ (.A(\vgademo.plane_dx_div.d[19] ),
    .B(_1108_),
    .Y(_1134_));
 sg13g2_inv_1 _5962_ (.Y(_1135_),
    .A(_1134_));
 sg13g2_a21oi_1 _5963_ (.A1(_1135_),
    .A2(_0975_),
    .Y(_1136_),
    .B1(_1092_));
 sg13g2_nor2_1 _5964_ (.A(_0975_),
    .B(_1135_),
    .Y(_1137_));
 sg13g2_inv_1 _5965_ (.Y(_1138_),
    .A(_1137_));
 sg13g2_nand2_1 _5966_ (.Y(_1139_),
    .A(_1136_),
    .B(_1138_));
 sg13g2_o21ai_1 _5967_ (.B1(_1139_),
    .Y(_1140_),
    .A1(net82),
    .A2(_0028_));
 sg13g2_xnor2_1 _5968_ (.Y(_1141_),
    .A(_1117_),
    .B(_1140_));
 sg13g2_nand2_1 _5969_ (.Y(_1142_),
    .A(_1122_),
    .B(\vgademo.plane_dx_div.r[18] ));
 sg13g2_o21ai_1 _5970_ (.B1(_1142_),
    .Y(_1143_),
    .A1(_1123_),
    .A2(_1125_));
 sg13g2_xnor2_1 _5971_ (.Y(_1144_),
    .A(_1141_),
    .B(_1143_));
 sg13g2_xnor2_1 _5972_ (.Y(_1145_),
    .A(_1130_),
    .B(_0991_));
 sg13g2_nor2_1 _5973_ (.A(\vgademo.plane_dx_div.r[20] ),
    .B(_1115_),
    .Y(_1146_));
 sg13g2_a221oi_1 _5974_ (.B2(_0905_),
    .C1(_1146_),
    .B1(_1145_),
    .A1(_1101_),
    .Y(_0231_),
    .A2(_1144_));
 sg13g2_inv_1 _5975_ (.Y(_1147_),
    .A(\vgademo.plane_dx_div.r[21] ));
 sg13g2_o21ai_1 _5976_ (.B1(_0992_),
    .Y(_1148_),
    .A1(_0975_),
    .A2(_1120_));
 sg13g2_nor2_1 _5977_ (.A(_0975_),
    .B(_1120_),
    .Y(_1149_));
 sg13g2_nand2_1 _5978_ (.Y(_1150_),
    .A(_1149_),
    .B(_0993_));
 sg13g2_nand3_1 _5979_ (.B(net82),
    .C(_1150_),
    .A(_1148_),
    .Y(_1151_));
 sg13g2_o21ai_1 _5980_ (.B1(_1151_),
    .Y(_1152_),
    .A1(net82),
    .A2(_0030_));
 sg13g2_xor2_1 _5981_ (.B(_1152_),
    .A(\vgademo.plane_dx_div.r[20] ),
    .X(_1153_));
 sg13g2_nand2_1 _5982_ (.Y(_1154_),
    .A(_1143_),
    .B(_1141_));
 sg13g2_nand2_1 _5983_ (.Y(_1155_),
    .A(_1140_),
    .B(\vgademo.plane_dx_div.r[19] ));
 sg13g2_nand2_1 _5984_ (.Y(_1156_),
    .A(_1154_),
    .B(_1155_));
 sg13g2_xnor2_1 _5985_ (.Y(_1157_),
    .A(_1153_),
    .B(_1156_));
 sg13g2_nor2_1 _5986_ (.A(_1130_),
    .B(_0991_),
    .Y(_1158_));
 sg13g2_inv_1 _5987_ (.Y(_1159_),
    .A(_1158_));
 sg13g2_nor2_1 _5988_ (.A(_1159_),
    .B(_1013_),
    .Y(_1160_));
 sg13g2_inv_1 _5989_ (.Y(_1161_),
    .A(_1160_));
 sg13g2_nand2_1 _5990_ (.Y(_1162_),
    .A(_1013_),
    .B(_1159_));
 sg13g2_a21oi_1 _5991_ (.A1(_1161_),
    .A2(_1162_),
    .Y(_1163_),
    .B1(_0953_));
 sg13g2_a221oi_1 _5992_ (.B2(_1157_),
    .C1(_1163_),
    .B1(_1101_),
    .A1(_1147_),
    .Y(_0232_),
    .A2(_1089_));
 sg13g2_o21ai_1 _5993_ (.B1(_1043_),
    .Y(_1164_),
    .A1(_0992_),
    .A2(_1138_));
 sg13g2_nor3_1 _5994_ (.A(_0992_),
    .B(_1043_),
    .C(_1138_),
    .Y(_1165_));
 sg13g2_inv_1 _5995_ (.Y(_1166_),
    .A(_1165_));
 sg13g2_nand3_1 _5996_ (.B(_1166_),
    .C(net82),
    .A(_1164_),
    .Y(_1167_));
 sg13g2_o21ai_1 _5997_ (.B1(_1167_),
    .Y(_1168_),
    .A1(net82),
    .A2(_0033_));
 sg13g2_xnor2_1 _5998_ (.Y(_1169_),
    .A(_1147_),
    .B(_1168_));
 sg13g2_nand2_1 _5999_ (.Y(_1170_),
    .A(_1156_),
    .B(_1153_));
 sg13g2_nand2_1 _6000_ (.Y(_1171_),
    .A(_1152_),
    .B(\vgademo.plane_dx_div.r[20] ));
 sg13g2_nand2_1 _6001_ (.Y(_1172_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_xnor2_1 _6002_ (.Y(_1173_),
    .A(_1169_),
    .B(_1172_));
 sg13g2_xnor2_1 _6003_ (.Y(_1174_),
    .A(_1160_),
    .B(_1042_));
 sg13g2_nor2_1 _6004_ (.A(\vgademo.plane_dx_div.r[22] ),
    .B(_1115_),
    .Y(_1175_));
 sg13g2_a221oi_1 _6005_ (.B2(_0905_),
    .C1(_1175_),
    .B1(_1174_),
    .A1(_1101_),
    .Y(_0233_),
    .A2(_1173_));
 sg13g2_o21ai_1 _6006_ (.B1(\vgademo.plane_dx_div.d[23] ),
    .Y(_1176_),
    .A1(_1043_),
    .A2(_1150_));
 sg13g2_nor2_1 _6007_ (.A(_1043_),
    .B(_1150_),
    .Y(_1177_));
 sg13g2_nand2_1 _6008_ (.Y(_1178_),
    .A(_1177_),
    .B(_1045_));
 sg13g2_nand3_1 _6009_ (.B(net82),
    .C(_1178_),
    .A(_1176_),
    .Y(_1179_));
 sg13g2_o21ai_1 _6010_ (.B1(_1179_),
    .Y(_1180_),
    .A1(net82),
    .A2(_0035_));
 sg13g2_xor2_1 _6011_ (.B(_1180_),
    .A(\vgademo.plane_dx_div.r[22] ),
    .X(_1181_));
 sg13g2_nand2_1 _6012_ (.Y(_1182_),
    .A(_1172_),
    .B(_1169_));
 sg13g2_nand2_1 _6013_ (.Y(_1183_),
    .A(_1168_),
    .B(\vgademo.plane_dx_div.r[21] ));
 sg13g2_nand2_1 _6014_ (.Y(_1184_),
    .A(_1182_),
    .B(_1183_));
 sg13g2_xor2_1 _6015_ (.B(_1184_),
    .A(_1181_),
    .X(_1185_));
 sg13g2_nor2b_1 _6016_ (.A(_1161_),
    .B_N(_1042_),
    .Y(_1186_));
 sg13g2_inv_1 _6017_ (.Y(_1187_),
    .A(_1186_));
 sg13g2_nand2_1 _6018_ (.Y(_1188_),
    .A(_1187_),
    .B(_1061_));
 sg13g2_nor2_1 _6019_ (.A(_1061_),
    .B(_1187_),
    .Y(_1189_));
 sg13g2_nor2_1 _6020_ (.A(_0953_),
    .B(_1189_),
    .Y(_1190_));
 sg13g2_a22oi_1 _6021_ (.Y(_1191_),
    .B1(_1188_),
    .B2(_1190_),
    .A2(_1185_),
    .A1(_4294_));
 sg13g2_nor2_1 _6022_ (.A(\vgademo.plane_dx_div.r[23] ),
    .B(_1115_),
    .Y(_1192_));
 sg13g2_a21oi_1 _6023_ (.A1(_1191_),
    .A2(_1115_),
    .Y(_0234_),
    .B1(_1192_));
 sg13g2_inv_1 _6024_ (.Y(_1193_),
    .A(\vgademo.plane_dx_div.r[24] ));
 sg13g2_o21ai_1 _6025_ (.B1(\vgademo.plane_dx_div.d[24] ),
    .Y(_1194_),
    .A1(\vgademo.plane_dx_div.d[23] ),
    .A2(_1166_));
 sg13g2_nand3b_1 _6026_ (.B(_1165_),
    .C(_1045_),
    .Y(_1195_),
    .A_N(\vgademo.plane_dx_div.d[24] ));
 sg13g2_nand3_1 _6027_ (.B(_1195_),
    .C(_1133_),
    .A(_1194_),
    .Y(_1196_));
 sg13g2_o21ai_1 _6028_ (.B1(_1196_),
    .Y(_1197_),
    .A1(_1133_),
    .A2(_0039_));
 sg13g2_xor2_1 _6029_ (.B(_1197_),
    .A(\vgademo.plane_dx_div.r[23] ),
    .X(_1198_));
 sg13g2_nand2_1 _6030_ (.Y(_1199_),
    .A(_1184_),
    .B(_1181_));
 sg13g2_nand2_1 _6031_ (.Y(_1200_),
    .A(_1180_),
    .B(\vgademo.plane_dx_div.r[22] ));
 sg13g2_nand2_1 _6032_ (.Y(_1201_),
    .A(_1199_),
    .B(_1200_));
 sg13g2_xor2_1 _6033_ (.B(_1201_),
    .A(_1198_),
    .X(_1202_));
 sg13g2_a21oi_1 _6034_ (.A1(_1202_),
    .A2(_4294_),
    .Y(_1203_),
    .B1(_1088_));
 sg13g2_a21oi_1 _6035_ (.A1(_1081_),
    .A2(_1189_),
    .Y(_1204_),
    .B1(_4298_));
 sg13g2_o21ai_1 _6036_ (.B1(_1204_),
    .Y(_1205_),
    .A1(_1081_),
    .A2(_1189_));
 sg13g2_a22oi_1 _6037_ (.Y(_0235_),
    .B1(_1203_),
    .B2(_1205_),
    .A2(net38),
    .A1(_1193_));
 sg13g2_o21ai_1 _6038_ (.B1(net82),
    .Y(_1206_),
    .A1(\vgademo.plane_dx_div.d[24] ),
    .A2(_1178_));
 sg13g2_xnor2_1 _6039_ (.Y(_1207_),
    .A(_1193_),
    .B(_1206_));
 sg13g2_nand2_1 _6040_ (.Y(_1208_),
    .A(_1201_),
    .B(_1198_));
 sg13g2_nand2_1 _6041_ (.Y(_1209_),
    .A(_1197_),
    .B(\vgademo.plane_dx_div.r[23] ));
 sg13g2_nand2_1 _6042_ (.Y(_1210_),
    .A(_1208_),
    .B(_1209_));
 sg13g2_xnor2_1 _6043_ (.Y(_1211_),
    .A(_1207_),
    .B(_1210_));
 sg13g2_a21oi_1 _6044_ (.A1(_4294_),
    .A2(_1211_),
    .Y(_1212_),
    .B1(_1204_));
 sg13g2_nor2_1 _6045_ (.A(_1092_),
    .B(_1115_),
    .Y(_1213_));
 sg13g2_a21oi_1 _6046_ (.A1(_1212_),
    .A2(_1115_),
    .Y(_0236_),
    .B1(_1213_));
 sg13g2_nand2_1 _6047_ (.Y(_1214_),
    .A(\vgademo.plane_u[0] ),
    .B(\vgademo.plane_du[0] ));
 sg13g2_a21oi_1 _6048_ (.A1(_4471_),
    .A2(_4476_),
    .Y(_1215_),
    .B1(_4428_));
 sg13g2_nand2_1 _6049_ (.Y(_1216_),
    .A(_0858_),
    .B(_4475_));
 sg13g2_a21oi_1 _6050_ (.A1(_4473_),
    .A2(_1215_),
    .Y(_1217_),
    .B1(_1216_));
 sg13g2_a21oi_1 _6051_ (.A1(_1217_),
    .A2(net143),
    .Y(_1218_),
    .B1(_0549_));
 sg13g2_buf_1 _6052_ (.A(_1218_),
    .X(_1219_));
 sg13g2_buf_1 _6053_ (.A(_1219_),
    .X(_1220_));
 sg13g2_a21oi_1 _6054_ (.A1(net53),
    .A2(_1214_),
    .Y(_1221_),
    .B1(net37));
 sg13g2_inv_1 _6055_ (.Y(_1222_),
    .A(_1219_));
 sg13g2_a21oi_1 _6056_ (.A1(_1222_),
    .A2(\vgademo.plane_du[0] ),
    .Y(_1223_),
    .B1(\vgademo.plane_u[0] ));
 sg13g2_nor2_1 _6057_ (.A(_1221_),
    .B(_1223_),
    .Y(_0237_));
 sg13g2_buf_1 _6058_ (.A(\vgademo.plane_u[10] ),
    .X(_1224_));
 sg13g2_inv_1 _6059_ (.Y(_1225_),
    .A(_1224_));
 sg13g2_buf_1 _6060_ (.A(_1219_),
    .X(_1226_));
 sg13g2_buf_1 _6061_ (.A(net36),
    .X(_1227_));
 sg13g2_nor2_1 _6062_ (.A(net113),
    .B(net112),
    .Y(_1228_));
 sg13g2_nand2_1 _6063_ (.Y(_1229_),
    .A(net113),
    .B(_0875_));
 sg13g2_nor2b_1 _6064_ (.A(_1228_),
    .B_N(_1229_),
    .Y(_1230_));
 sg13g2_xnor2_1 _6065_ (.Y(_1231_),
    .A(_0891_),
    .B(_1230_));
 sg13g2_nor2_1 _6066_ (.A(_0868_),
    .B(net113),
    .Y(_1232_));
 sg13g2_nand2_1 _6067_ (.Y(_1233_),
    .A(_0868_),
    .B(net113));
 sg13g2_o21ai_1 _6068_ (.B1(_1233_),
    .Y(_1234_),
    .A1(_0888_),
    .A2(_1232_));
 sg13g2_nor2b_1 _6069_ (.A(_1231_),
    .B_N(_1234_),
    .Y(_1235_));
 sg13g2_nand2b_1 _6070_ (.Y(_1236_),
    .B(_1231_),
    .A_N(_1234_));
 sg13g2_nand2b_1 _6071_ (.Y(_1237_),
    .B(_1236_),
    .A_N(_1235_));
 sg13g2_inv_1 _6072_ (.Y(_1238_),
    .A(_1237_));
 sg13g2_nor2_1 _6073_ (.A(_0868_),
    .B(_1105_),
    .Y(_1239_));
 sg13g2_inv_1 _6074_ (.Y(_1240_),
    .A(_1239_));
 sg13g2_nor2_1 _6075_ (.A(_1092_),
    .B(_0869_),
    .Y(_1241_));
 sg13g2_a21oi_1 _6076_ (.A1(_1240_),
    .A2(_0883_),
    .Y(_1242_),
    .B1(_1241_));
 sg13g2_nor2b_1 _6077_ (.A(_1232_),
    .B_N(_1233_),
    .Y(_1243_));
 sg13g2_xnor2_1 _6078_ (.Y(_1244_),
    .A(_0887_),
    .B(_1243_));
 sg13g2_xor2_1 _6079_ (.B(_1244_),
    .A(_1242_),
    .X(_1245_));
 sg13g2_nand2_1 _6080_ (.Y(_1246_),
    .A(_0855_),
    .B(_0879_));
 sg13g2_nor2_1 _6081_ (.A(_1241_),
    .B(_1239_),
    .Y(_1247_));
 sg13g2_xnor2_1 _6082_ (.Y(_1248_),
    .A(_0883_),
    .B(_1247_));
 sg13g2_nor2_1 _6083_ (.A(_1246_),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_nor2_1 _6084_ (.A(_1242_),
    .B(_1244_),
    .Y(_1250_));
 sg13g2_a21oi_1 _6085_ (.A1(_1245_),
    .A2(_1249_),
    .Y(_1251_),
    .B1(_1250_));
 sg13g2_xnor2_1 _6086_ (.Y(_1252_),
    .A(_1238_),
    .B(_1251_));
 sg13g2_inv_1 _6087_ (.Y(_1253_),
    .A(_1252_));
 sg13g2_xor2_1 _6088_ (.B(_1245_),
    .A(_1249_),
    .X(_1254_));
 sg13g2_nand2_1 _6089_ (.Y(_1255_),
    .A(_1253_),
    .B(_1254_));
 sg13g2_inv_1 _6090_ (.Y(_1256_),
    .A(_1254_));
 sg13g2_nand2_1 _6091_ (.Y(_1257_),
    .A(_1252_),
    .B(_1256_));
 sg13g2_nand2_1 _6092_ (.Y(_1258_),
    .A(_1255_),
    .B(_1257_));
 sg13g2_inv_1 _6093_ (.Y(_1259_),
    .A(_1258_));
 sg13g2_inv_1 _6094_ (.Y(_1260_),
    .A(_1246_));
 sg13g2_xnor2_1 _6095_ (.Y(_1261_),
    .A(_1260_),
    .B(_1248_));
 sg13g2_nor2_1 _6096_ (.A(_0855_),
    .B(_0879_),
    .Y(_1262_));
 sg13g2_nor2_1 _6097_ (.A(_1262_),
    .B(_1260_),
    .Y(_1263_));
 sg13g2_nor2_1 _6098_ (.A(net113),
    .B(_1240_),
    .Y(_1264_));
 sg13g2_inv_1 _6099_ (.Y(_1265_),
    .A(_1264_));
 sg13g2_nor3_1 _6100_ (.A(net112),
    .B(_1263_),
    .C(_1265_),
    .Y(_1266_));
 sg13g2_nor2_1 _6101_ (.A(_1266_),
    .B(_1261_),
    .Y(_1267_));
 sg13g2_o21ai_1 _6102_ (.B1(_1256_),
    .Y(_1268_),
    .A1(_1261_),
    .A2(_1267_));
 sg13g2_nand2_1 _6103_ (.Y(_1269_),
    .A(_1259_),
    .B(_1268_));
 sg13g2_xor2_1 _6104_ (.B(_0879_),
    .A(net112),
    .X(_1270_));
 sg13g2_xnor2_1 _6105_ (.Y(_1271_),
    .A(_0895_),
    .B(_1270_));
 sg13g2_o21ai_1 _6106_ (.B1(_1229_),
    .Y(_1272_),
    .A1(_0892_),
    .A2(_1228_));
 sg13g2_nor2b_1 _6107_ (.A(_1271_),
    .B_N(_1272_),
    .Y(_1273_));
 sg13g2_inv_1 _6108_ (.Y(_1274_),
    .A(_1273_));
 sg13g2_nand2b_1 _6109_ (.Y(_1275_),
    .B(_1271_),
    .A_N(_1272_));
 sg13g2_nand2_1 _6110_ (.Y(_1276_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_inv_1 _6111_ (.Y(_1277_),
    .A(_1251_));
 sg13g2_a21o_1 _6112_ (.A2(_1236_),
    .A1(_1277_),
    .B1(_1235_),
    .X(_1278_));
 sg13g2_buf_1 _6113_ (.A(_1278_),
    .X(_1279_));
 sg13g2_xnor2_1 _6114_ (.Y(_1280_),
    .A(_1276_),
    .B(_1279_));
 sg13g2_xnor2_1 _6115_ (.Y(_1281_),
    .A(_0856_),
    .B(_1280_));
 sg13g2_xnor2_1 _6116_ (.Y(_1282_),
    .A(_1253_),
    .B(_1281_));
 sg13g2_o21ai_1 _6117_ (.B1(_1281_),
    .Y(_1283_),
    .A1(_1253_),
    .A2(_1256_));
 sg13g2_o21ai_1 _6118_ (.B1(_1283_),
    .Y(_1284_),
    .A1(_1269_),
    .A2(_1282_));
 sg13g2_nor2_1 _6119_ (.A(_0855_),
    .B(_1280_),
    .Y(_1285_));
 sg13g2_inv_1 _6120_ (.Y(_1286_),
    .A(_1285_));
 sg13g2_xor2_1 _6121_ (.B(_0883_),
    .A(_0879_),
    .X(_1287_));
 sg13g2_xnor2_1 _6122_ (.Y(_1288_),
    .A(\vgademo.plane_dx_div.q[8] ),
    .B(_1287_));
 sg13g2_nand2_1 _6123_ (.Y(_1289_),
    .A(_1270_),
    .B(_0895_));
 sg13g2_o21ai_1 _6124_ (.B1(_1289_),
    .Y(_1290_),
    .A1(_0876_),
    .A2(_0880_));
 sg13g2_nor2b_1 _6125_ (.A(_1288_),
    .B_N(_1290_),
    .Y(_1291_));
 sg13g2_inv_1 _6126_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nand2b_1 _6127_ (.Y(_1293_),
    .B(_1288_),
    .A_N(_1290_));
 sg13g2_nand2_1 _6128_ (.Y(_1294_),
    .A(_1292_),
    .B(_1293_));
 sg13g2_a21oi_1 _6129_ (.A1(_1279_),
    .A2(_1275_),
    .Y(_1295_),
    .B1(_1273_));
 sg13g2_xor2_1 _6130_ (.B(_1295_),
    .A(_1294_),
    .X(_1296_));
 sg13g2_xnor2_1 _6131_ (.Y(_1297_),
    .A(_0868_),
    .B(_1296_));
 sg13g2_nor2_1 _6132_ (.A(_1286_),
    .B(_1297_),
    .Y(_1298_));
 sg13g2_inv_1 _6133_ (.Y(_1299_),
    .A(_1298_));
 sg13g2_nand2_1 _6134_ (.Y(_1300_),
    .A(_1297_),
    .B(_1286_));
 sg13g2_nand2_1 _6135_ (.Y(_1301_),
    .A(_1299_),
    .B(_1300_));
 sg13g2_nand2b_1 _6136_ (.Y(_1302_),
    .B(_1301_),
    .A_N(_1284_));
 sg13g2_inv_1 _6137_ (.Y(_1303_),
    .A(_1301_));
 sg13g2_nand2_1 _6138_ (.Y(_1304_),
    .A(_1303_),
    .B(_1284_));
 sg13g2_nand3_1 _6139_ (.B(net45),
    .C(_1304_),
    .A(_1302_),
    .Y(_1305_));
 sg13g2_nor2_1 _6140_ (.A(_1224_),
    .B(_0866_),
    .Y(_1306_));
 sg13g2_nand2_1 _6141_ (.Y(_1307_),
    .A(_1224_),
    .B(_0866_));
 sg13g2_nor2b_1 _6142_ (.A(_1306_),
    .B_N(_1307_),
    .Y(_1308_));
 sg13g2_nor2_1 _6143_ (.A(\vgademo.plane_u[9] ),
    .B(_0901_),
    .Y(_1309_));
 sg13g2_nor2_1 _6144_ (.A(\vgademo.plane_u[5] ),
    .B(_0885_),
    .Y(_1310_));
 sg13g2_nor2_1 _6145_ (.A(\vgademo.plane_u[4] ),
    .B(_0881_),
    .Y(_1311_));
 sg13g2_xor2_1 _6146_ (.B(\vgademo.plane_du[1] ),
    .A(\vgademo.plane_u[1] ),
    .X(_1312_));
 sg13g2_inv_1 _6147_ (.Y(_1313_),
    .A(_1312_));
 sg13g2_nand2_1 _6148_ (.Y(_1314_),
    .A(\vgademo.plane_u[1] ),
    .B(\vgademo.plane_du[1] ));
 sg13g2_o21ai_1 _6149_ (.B1(_1314_),
    .Y(_1315_),
    .A1(_1214_),
    .A2(_1313_));
 sg13g2_nor2_1 _6150_ (.A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ),
    .Y(_1316_));
 sg13g2_inv_1 _6151_ (.Y(_1317_),
    .A(_1316_));
 sg13g2_nand2_1 _6152_ (.Y(_1318_),
    .A(\vgademo.plane_u[2] ),
    .B(\vgademo.plane_du[2] ));
 sg13g2_inv_1 _6153_ (.Y(_1319_),
    .A(_1318_));
 sg13g2_a21oi_1 _6154_ (.A1(_1315_),
    .A2(_1317_),
    .Y(_1320_),
    .B1(_1319_));
 sg13g2_nand2_1 _6155_ (.Y(_1321_),
    .A(\vgademo.plane_u[3] ),
    .B(_0877_));
 sg13g2_nor2_1 _6156_ (.A(\vgademo.plane_u[3] ),
    .B(_0877_),
    .Y(_1322_));
 sg13g2_a21oi_1 _6157_ (.A1(_1320_),
    .A2(_1321_),
    .Y(_1323_),
    .B1(_1322_));
 sg13g2_inv_1 _6158_ (.Y(_1324_),
    .A(_1323_));
 sg13g2_nand2_1 _6159_ (.Y(_1325_),
    .A(\vgademo.plane_u[4] ),
    .B(_0881_));
 sg13g2_o21ai_1 _6160_ (.B1(_1325_),
    .Y(_1326_),
    .A1(_1311_),
    .A2(_1324_));
 sg13g2_inv_1 _6161_ (.Y(_1327_),
    .A(_1326_));
 sg13g2_nand2_1 _6162_ (.Y(_1328_),
    .A(\vgademo.plane_u[5] ),
    .B(_0885_));
 sg13g2_o21ai_1 _6163_ (.B1(_1328_),
    .Y(_1329_),
    .A1(_1310_),
    .A2(_1327_));
 sg13g2_buf_1 _6164_ (.A(_1329_),
    .X(_1330_));
 sg13g2_nor2_1 _6165_ (.A(\vgademo.plane_u[7] ),
    .B(_0893_),
    .Y(_1331_));
 sg13g2_nand2_1 _6166_ (.Y(_1332_),
    .A(\vgademo.plane_u[7] ),
    .B(_0893_));
 sg13g2_inv_1 _6167_ (.Y(_1333_),
    .A(_1332_));
 sg13g2_nor2_1 _6168_ (.A(_1331_),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_inv_1 _6169_ (.Y(_1335_),
    .A(_1334_));
 sg13g2_nor2_1 _6170_ (.A(\vgademo.plane_u[6] ),
    .B(_0889_),
    .Y(_1336_));
 sg13g2_nand2_1 _6171_ (.Y(_1337_),
    .A(\vgademo.plane_u[6] ),
    .B(_0889_));
 sg13g2_inv_1 _6172_ (.Y(_1338_),
    .A(_1337_));
 sg13g2_nor2_1 _6173_ (.A(_1336_),
    .B(_1338_),
    .Y(_1339_));
 sg13g2_nor2b_1 _6174_ (.A(_1335_),
    .B_N(_1339_),
    .Y(_1340_));
 sg13g2_a21oi_1 _6175_ (.A1(_1337_),
    .A2(_1332_),
    .Y(_1341_),
    .B1(_1331_));
 sg13g2_a21oi_1 _6176_ (.A1(_1330_),
    .A2(_1340_),
    .Y(_1342_),
    .B1(_1341_));
 sg13g2_inv_1 _6177_ (.Y(_1343_),
    .A(_1342_));
 sg13g2_nor2_1 _6178_ (.A(\vgademo.plane_u[8] ),
    .B(net111),
    .Y(_1344_));
 sg13g2_nand2_1 _6179_ (.Y(_1345_),
    .A(\vgademo.plane_u[8] ),
    .B(net111));
 sg13g2_inv_1 _6180_ (.Y(_1346_),
    .A(_1345_));
 sg13g2_nor2_1 _6181_ (.A(_1344_),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_nand2_1 _6182_ (.Y(_1348_),
    .A(_1343_),
    .B(_1347_));
 sg13g2_nand2_1 _6183_ (.Y(_1349_),
    .A(\vgademo.plane_u[9] ),
    .B(_0901_));
 sg13g2_nand3_1 _6184_ (.B(_1345_),
    .C(_1349_),
    .A(_1348_),
    .Y(_1350_));
 sg13g2_nand2b_1 _6185_ (.Y(_1351_),
    .B(_1350_),
    .A_N(_1309_));
 sg13g2_xnor2_1 _6186_ (.Y(_1352_),
    .A(_1308_),
    .B(_1351_));
 sg13g2_a21oi_1 _6187_ (.A1(_1352_),
    .A2(_0634_),
    .Y(_1353_),
    .B1(_1220_));
 sg13g2_a22oi_1 _6188_ (.Y(_0238_),
    .B1(_1305_),
    .B2(_1353_),
    .A2(net32),
    .A1(_1225_));
 sg13g2_buf_1 _6189_ (.A(net36),
    .X(_1354_));
 sg13g2_o21ai_1 _6190_ (.B1(_1307_),
    .Y(_1355_),
    .A1(_1306_),
    .A2(_1351_));
 sg13g2_inv_1 _6191_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_nor2_1 _6192_ (.A(_0041_),
    .B(_1356_),
    .Y(_1357_));
 sg13g2_nor2_1 _6193_ (.A(_0558_),
    .B(_1357_),
    .Y(_1358_));
 sg13g2_nand2_1 _6194_ (.Y(_1359_),
    .A(_1356_),
    .B(_0041_));
 sg13g2_nand2_1 _6195_ (.Y(_1360_),
    .A(_1245_),
    .B(_1261_));
 sg13g2_xnor2_1 _6196_ (.Y(_1361_),
    .A(_1261_),
    .B(_1254_));
 sg13g2_inv_1 _6197_ (.Y(_1362_),
    .A(_1267_));
 sg13g2_nand2_1 _6198_ (.Y(_1363_),
    .A(_1361_),
    .B(_1362_));
 sg13g2_inv_1 _6199_ (.Y(_1364_),
    .A(_1363_));
 sg13g2_a22oi_1 _6200_ (.Y(_1365_),
    .B1(_1364_),
    .B2(_1259_),
    .A2(_1360_),
    .A1(_1252_));
 sg13g2_nor2_1 _6201_ (.A(_1365_),
    .B(_1282_),
    .Y(_1366_));
 sg13g2_inv_1 _6202_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_inv_1 _6203_ (.Y(_1368_),
    .A(_1281_));
 sg13g2_nor2_1 _6204_ (.A(_1252_),
    .B(_1368_),
    .Y(_1369_));
 sg13g2_inv_1 _6205_ (.Y(_1370_),
    .A(_1369_));
 sg13g2_nand3_1 _6206_ (.B(_1299_),
    .C(_1370_),
    .A(_1367_),
    .Y(_1371_));
 sg13g2_nand2_1 _6207_ (.Y(_1372_),
    .A(_1371_),
    .B(_1300_));
 sg13g2_nor2_1 _6208_ (.A(_0868_),
    .B(_1296_),
    .Y(_1373_));
 sg13g2_inv_1 _6209_ (.Y(_1374_),
    .A(_1373_));
 sg13g2_nand2_1 _6210_ (.Y(_1375_),
    .A(_0884_),
    .B(_0888_));
 sg13g2_nand2_1 _6211_ (.Y(_1376_),
    .A(_0883_),
    .B(_0887_));
 sg13g2_a21oi_1 _6212_ (.A1(_1375_),
    .A2(_1376_),
    .Y(_1377_),
    .B1(net114));
 sg13g2_nand3_1 _6213_ (.B(net114),
    .C(_1376_),
    .A(_1375_),
    .Y(_1378_));
 sg13g2_nand2b_1 _6214_ (.Y(_1379_),
    .B(_1378_),
    .A_N(_1377_));
 sg13g2_nand2_1 _6215_ (.Y(_1380_),
    .A(_1287_),
    .B(net110));
 sg13g2_o21ai_1 _6216_ (.B1(_1380_),
    .Y(_1381_),
    .A1(_0880_),
    .A2(_0884_));
 sg13g2_nor2b_1 _6217_ (.A(_1379_),
    .B_N(_1381_),
    .Y(_1382_));
 sg13g2_nor2b_1 _6218_ (.A(_1381_),
    .B_N(_1379_),
    .Y(_1383_));
 sg13g2_nor2_1 _6219_ (.A(_1382_),
    .B(_1383_),
    .Y(_1384_));
 sg13g2_nor2b_1 _6220_ (.A(_1276_),
    .B_N(_1279_),
    .Y(_1385_));
 sg13g2_nor3_1 _6221_ (.A(_1273_),
    .B(_1291_),
    .C(_1385_),
    .Y(_1386_));
 sg13g2_nor2b_1 _6222_ (.A(_1386_),
    .B_N(_1293_),
    .Y(_1387_));
 sg13g2_xor2_1 _6223_ (.B(_1387_),
    .A(_1384_),
    .X(_1388_));
 sg13g2_xnor2_1 _6224_ (.Y(_1389_),
    .A(net113),
    .B(_1388_));
 sg13g2_xnor2_1 _6225_ (.Y(_1390_),
    .A(_1374_),
    .B(_1389_));
 sg13g2_nor2_1 _6226_ (.A(_1372_),
    .B(_1390_),
    .Y(_1391_));
 sg13g2_inv_1 _6227_ (.Y(_1392_),
    .A(_1391_));
 sg13g2_a21oi_1 _6228_ (.A1(_1390_),
    .A2(_1372_),
    .Y(_1393_),
    .B1(net63));
 sg13g2_a22oi_1 _6229_ (.Y(_1394_),
    .B1(_1392_),
    .B2(_1393_),
    .A2(_1359_),
    .A1(_1358_));
 sg13g2_nand2_1 _6230_ (.Y(_1395_),
    .A(_1354_),
    .B(\vgademo.plane_u[11] ));
 sg13g2_o21ai_1 _6231_ (.B1(_1395_),
    .Y(_0239_),
    .A1(_1354_),
    .A2(_1394_));
 sg13g2_buf_1 _6232_ (.A(\vgademo.plane_u[12] ),
    .X(_1396_));
 sg13g2_inv_1 _6233_ (.Y(_1397_),
    .A(_1396_));
 sg13g2_nor2_1 _6234_ (.A(net113),
    .B(_1388_),
    .Y(_1398_));
 sg13g2_inv_1 _6235_ (.Y(_1399_),
    .A(_1398_));
 sg13g2_xor2_1 _6236_ (.B(_0891_),
    .A(_0887_),
    .X(_1400_));
 sg13g2_nand2_1 _6237_ (.Y(_1401_),
    .A(_1378_),
    .B(_1376_));
 sg13g2_xnor2_1 _6238_ (.Y(_1402_),
    .A(_1400_),
    .B(_1401_));
 sg13g2_nor2_1 _6239_ (.A(_1294_),
    .B(_1295_),
    .Y(_1403_));
 sg13g2_nor3_1 _6240_ (.A(_1291_),
    .B(_1382_),
    .C(_1403_),
    .Y(_1404_));
 sg13g2_nor2_1 _6241_ (.A(_1383_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_xnor2_1 _6242_ (.Y(_1406_),
    .A(_1402_),
    .B(_1405_));
 sg13g2_xnor2_1 _6243_ (.Y(_1407_),
    .A(net112),
    .B(_1406_));
 sg13g2_nor2_1 _6244_ (.A(_1399_),
    .B(_1407_),
    .Y(_1408_));
 sg13g2_inv_1 _6245_ (.Y(_1409_),
    .A(_1408_));
 sg13g2_nand2_1 _6246_ (.Y(_1410_),
    .A(_1407_),
    .B(_1399_));
 sg13g2_nand2_1 _6247_ (.Y(_1411_),
    .A(_1409_),
    .B(_1410_));
 sg13g2_nor2_1 _6248_ (.A(_1374_),
    .B(_1389_),
    .Y(_1412_));
 sg13g2_nor2_1 _6249_ (.A(_1298_),
    .B(_1412_),
    .Y(_1413_));
 sg13g2_a22oi_1 _6250_ (.Y(_1414_),
    .B1(_1304_),
    .B2(_1413_),
    .A2(_1389_),
    .A1(_1374_));
 sg13g2_xnor2_1 _6251_ (.Y(_1415_),
    .A(_1411_),
    .B(_1414_));
 sg13g2_xor2_1 _6252_ (.B(_1357_),
    .A(_0042_),
    .X(_1416_));
 sg13g2_o21ai_1 _6253_ (.B1(_1222_),
    .Y(_1417_),
    .A1(net41),
    .A2(_1416_));
 sg13g2_a21oi_1 _6254_ (.A1(net45),
    .A2(_1415_),
    .Y(_1418_),
    .B1(_1417_));
 sg13g2_a21oi_1 _6255_ (.A1(_1397_),
    .A2(net32),
    .Y(_0240_),
    .B1(_1418_));
 sg13g2_inv_1 _6256_ (.Y(_1419_),
    .A(\vgademo.plane_u[13] ));
 sg13g2_inv_1 _6257_ (.Y(_1420_),
    .A(\vgademo.plane_u[11] ));
 sg13g2_nor3_1 _6258_ (.A(_1420_),
    .B(_1397_),
    .C(_1356_),
    .Y(_1421_));
 sg13g2_inv_1 _6259_ (.Y(_1422_),
    .A(_1421_));
 sg13g2_o21ai_1 _6260_ (.B1(_0540_),
    .Y(_1423_),
    .A1(_0043_),
    .A2(_1422_));
 sg13g2_a21oi_1 _6261_ (.A1(_0043_),
    .A2(_1422_),
    .Y(_1424_),
    .B1(_1423_));
 sg13g2_inv_1 _6262_ (.Y(_1425_),
    .A(_1412_));
 sg13g2_nand2_1 _6263_ (.Y(_1426_),
    .A(_1409_),
    .B(_1425_));
 sg13g2_o21ai_1 _6264_ (.B1(_1410_),
    .Y(_1427_),
    .A1(_1426_),
    .A2(_1391_));
 sg13g2_inv_1 _6265_ (.Y(_1428_),
    .A(_1427_));
 sg13g2_nor2_1 _6266_ (.A(net112),
    .B(_1406_),
    .Y(_1429_));
 sg13g2_nand2_1 _6267_ (.Y(_1430_),
    .A(_0892_),
    .B(_0896_));
 sg13g2_nand2_1 _6268_ (.Y(_1431_),
    .A(_0891_),
    .B(_0895_));
 sg13g2_nand2_1 _6269_ (.Y(_1432_),
    .A(_0887_),
    .B(_0891_));
 sg13g2_inv_1 _6270_ (.Y(_1433_),
    .A(_1432_));
 sg13g2_a21oi_1 _6271_ (.A1(_1430_),
    .A2(_1431_),
    .Y(_1434_),
    .B1(_1433_));
 sg13g2_nor2_1 _6272_ (.A(_0895_),
    .B(_1432_),
    .Y(_1435_));
 sg13g2_inv_1 _6273_ (.Y(_1436_),
    .A(_1435_));
 sg13g2_nand2b_1 _6274_ (.Y(_1437_),
    .B(_1436_),
    .A_N(_1434_));
 sg13g2_nor3_1 _6275_ (.A(_1383_),
    .B(_1402_),
    .C(_1404_),
    .Y(_1438_));
 sg13g2_a21o_1 _6276_ (.A2(_1400_),
    .A1(_1401_),
    .B1(_1438_),
    .X(_1439_));
 sg13g2_xnor2_1 _6277_ (.Y(_1440_),
    .A(_1437_),
    .B(_1439_));
 sg13g2_xnor2_1 _6278_ (.Y(_1441_),
    .A(_0879_),
    .B(_1440_));
 sg13g2_xnor2_1 _6279_ (.Y(_1442_),
    .A(_1429_),
    .B(_1441_));
 sg13g2_nor2_1 _6280_ (.A(_1428_),
    .B(_1442_),
    .Y(_1443_));
 sg13g2_nand2_1 _6281_ (.Y(_1444_),
    .A(_1442_),
    .B(_1428_));
 sg13g2_inv_1 _6282_ (.Y(_1445_),
    .A(_1444_));
 sg13g2_nor3_1 _6283_ (.A(net63),
    .B(_1443_),
    .C(_1445_),
    .Y(_1446_));
 sg13g2_nor3_1 _6284_ (.A(net36),
    .B(_1424_),
    .C(_1446_),
    .Y(_1447_));
 sg13g2_a21oi_1 _6285_ (.A1(_1419_),
    .A2(net32),
    .Y(_0241_),
    .B1(_1447_));
 sg13g2_buf_1 _6286_ (.A(\vgademo.plane_u[14] ),
    .X(_1448_));
 sg13g2_inv_1 _6287_ (.Y(_1449_),
    .A(_1448_));
 sg13g2_nand2_1 _6288_ (.Y(_1450_),
    .A(_1396_),
    .B(\vgademo.plane_u[13] ));
 sg13g2_nor3_1 _6289_ (.A(_0041_),
    .B(_1450_),
    .C(_1356_),
    .Y(_1451_));
 sg13g2_xnor2_1 _6290_ (.Y(_1452_),
    .A(_0044_),
    .B(_1451_));
 sg13g2_nor2_1 _6291_ (.A(_0879_),
    .B(_1440_),
    .Y(_1453_));
 sg13g2_inv_1 _6292_ (.Y(_1454_),
    .A(_1453_));
 sg13g2_nor2_1 _6293_ (.A(net110),
    .B(_1431_),
    .Y(_1455_));
 sg13g2_inv_1 _6294_ (.Y(_1456_),
    .A(_1431_));
 sg13g2_xor2_1 _6295_ (.B(net110),
    .A(_0895_),
    .X(_1457_));
 sg13g2_nor2_1 _6296_ (.A(_1456_),
    .B(_1457_),
    .Y(_1458_));
 sg13g2_nor2_1 _6297_ (.A(_1455_),
    .B(_1458_),
    .Y(_1459_));
 sg13g2_inv_1 _6298_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_nand2b_1 _6299_ (.Y(_1461_),
    .B(_1439_),
    .A_N(_1437_));
 sg13g2_nand2_1 _6300_ (.Y(_1462_),
    .A(_1461_),
    .B(_1436_));
 sg13g2_xnor2_1 _6301_ (.Y(_1463_),
    .A(_1460_),
    .B(_1462_));
 sg13g2_xnor2_1 _6302_ (.Y(_1464_),
    .A(_0883_),
    .B(_1463_));
 sg13g2_nor2_1 _6303_ (.A(_1454_),
    .B(_1464_),
    .Y(_1465_));
 sg13g2_inv_1 _6304_ (.Y(_1466_),
    .A(_1465_));
 sg13g2_nand2_1 _6305_ (.Y(_1467_),
    .A(_1464_),
    .B(_1454_));
 sg13g2_nand2_1 _6306_ (.Y(_1468_),
    .A(_1466_),
    .B(_1467_));
 sg13g2_nor2b_1 _6307_ (.A(_1441_),
    .B_N(_1429_),
    .Y(_1469_));
 sg13g2_nor2_1 _6308_ (.A(_1469_),
    .B(_1445_),
    .Y(_1470_));
 sg13g2_nor2_1 _6309_ (.A(_1468_),
    .B(_1470_),
    .Y(_1471_));
 sg13g2_nor2_1 _6310_ (.A(_0541_),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_nand2_1 _6311_ (.Y(_1473_),
    .A(_1470_),
    .B(_1468_));
 sg13g2_a221oi_1 _6312_ (.B2(_1473_),
    .C1(net36),
    .B1(_1472_),
    .A1(_0542_),
    .Y(_1474_),
    .A2(_1452_));
 sg13g2_a21oi_1 _6313_ (.A1(_1449_),
    .A2(net32),
    .Y(_0242_),
    .B1(_1474_));
 sg13g2_buf_1 _6314_ (.A(\vgademo.plane_u[15] ),
    .X(_1475_));
 sg13g2_inv_1 _6315_ (.Y(_1476_),
    .A(_1475_));
 sg13g2_nor3_1 _6316_ (.A(_1419_),
    .B(_1449_),
    .C(_1422_),
    .Y(_1477_));
 sg13g2_xnor2_1 _6317_ (.Y(_1478_),
    .A(_0045_),
    .B(_1477_));
 sg13g2_inv_1 _6318_ (.Y(_1479_),
    .A(_1467_));
 sg13g2_a21oi_1 _6319_ (.A1(_1470_),
    .A2(_1466_),
    .Y(_1480_),
    .B1(_1479_));
 sg13g2_inv_1 _6320_ (.Y(_1481_),
    .A(_1480_));
 sg13g2_nor2_1 _6321_ (.A(_0883_),
    .B(_1463_),
    .Y(_1482_));
 sg13g2_inv_1 _6322_ (.Y(_1483_),
    .A(_1482_));
 sg13g2_nor3_1 _6323_ (.A(net114),
    .B(_0896_),
    .C(_0900_),
    .Y(_1484_));
 sg13g2_nor2_1 _6324_ (.A(net110),
    .B(net114),
    .Y(_1485_));
 sg13g2_inv_1 _6325_ (.Y(_1486_),
    .A(_1485_));
 sg13g2_nand2_1 _6326_ (.Y(_1487_),
    .A(_0899_),
    .B(net114));
 sg13g2_nand2_1 _6327_ (.Y(_1488_),
    .A(_1486_),
    .B(_1487_));
 sg13g2_o21ai_1 _6328_ (.B1(_1488_),
    .Y(_1489_),
    .A1(_0896_),
    .A2(_0900_));
 sg13g2_nor2b_1 _6329_ (.A(_1484_),
    .B_N(_1489_),
    .Y(_1490_));
 sg13g2_o21ai_1 _6330_ (.B1(_1457_),
    .Y(_1491_),
    .A1(_1433_),
    .A2(_1456_));
 sg13g2_o21ai_1 _6331_ (.B1(_1491_),
    .Y(_1492_),
    .A1(_1460_),
    .A2(_1461_));
 sg13g2_xor2_1 _6332_ (.B(_1492_),
    .A(_1490_),
    .X(_1493_));
 sg13g2_xnor2_1 _6333_ (.Y(_1494_),
    .A(_0887_),
    .B(_1493_));
 sg13g2_nor2_1 _6334_ (.A(_1483_),
    .B(_1494_),
    .Y(_1495_));
 sg13g2_inv_1 _6335_ (.Y(_1496_),
    .A(_1495_));
 sg13g2_nand2_1 _6336_ (.Y(_1497_),
    .A(_1494_),
    .B(_1483_));
 sg13g2_nand2_1 _6337_ (.Y(_1498_),
    .A(_1496_),
    .B(_1497_));
 sg13g2_a21oi_1 _6338_ (.A1(_1481_),
    .A2(_1498_),
    .Y(_1499_),
    .B1(_0541_));
 sg13g2_nor2b_1 _6339_ (.A(_1498_),
    .B_N(_1480_),
    .Y(_1500_));
 sg13g2_inv_1 _6340_ (.Y(_1501_),
    .A(_1500_));
 sg13g2_a221oi_1 _6341_ (.B2(_1501_),
    .C1(net36),
    .B1(_1499_),
    .A1(net62),
    .Y(_1502_),
    .A2(_1478_));
 sg13g2_a21oi_1 _6342_ (.A1(_1476_),
    .A2(net32),
    .Y(_0243_),
    .B1(_1502_));
 sg13g2_inv_1 _6343_ (.Y(_1503_),
    .A(\vgademo.plane_u[16] ));
 sg13g2_nor2_1 _6344_ (.A(_0887_),
    .B(_1493_),
    .Y(_1504_));
 sg13g2_inv_1 _6345_ (.Y(_1505_),
    .A(_1504_));
 sg13g2_nor2_1 _6346_ (.A(net110),
    .B(_0865_),
    .Y(_1506_));
 sg13g2_nand2_1 _6347_ (.Y(_1507_),
    .A(_1490_),
    .B(_1459_));
 sg13g2_inv_1 _6348_ (.Y(_1508_),
    .A(_1462_));
 sg13g2_a21oi_1 _6349_ (.A1(_1455_),
    .A2(net114),
    .Y(_1509_),
    .B1(_1484_));
 sg13g2_o21ai_1 _6350_ (.B1(_1509_),
    .Y(_1510_),
    .A1(_1507_),
    .A2(_1508_));
 sg13g2_xor2_1 _6351_ (.B(_1510_),
    .A(_1506_),
    .X(_1511_));
 sg13g2_xnor2_1 _6352_ (.Y(_1512_),
    .A(_0891_),
    .B(_1511_));
 sg13g2_nor2_1 _6353_ (.A(_1505_),
    .B(_1512_),
    .Y(_1513_));
 sg13g2_nand2_1 _6354_ (.Y(_1514_),
    .A(_1512_),
    .B(_1505_));
 sg13g2_inv_1 _6355_ (.Y(_1515_),
    .A(_1514_));
 sg13g2_nor2_1 _6356_ (.A(_1513_),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_nand2_1 _6357_ (.Y(_1517_),
    .A(_1496_),
    .B(_1466_));
 sg13g2_o21ai_1 _6358_ (.B1(_1497_),
    .Y(_1518_),
    .A1(_1471_),
    .A2(_1517_));
 sg13g2_xnor2_1 _6359_ (.Y(_1519_),
    .A(_1516_),
    .B(_1518_));
 sg13g2_nand3_1 _6360_ (.B(_1448_),
    .C(_1475_),
    .A(_1451_),
    .Y(_1520_));
 sg13g2_xnor2_1 _6361_ (.Y(_1521_),
    .A(_0046_),
    .B(_1520_));
 sg13g2_o21ai_1 _6362_ (.B1(_1222_),
    .Y(_1522_),
    .A1(_0730_),
    .A2(_1521_));
 sg13g2_a21oi_1 _6363_ (.A1(_1519_),
    .A2(net45),
    .Y(_1523_),
    .B1(_1522_));
 sg13g2_a21oi_1 _6364_ (.A1(_1503_),
    .A2(net32),
    .Y(_0244_),
    .B1(_1523_));
 sg13g2_inv_1 _6365_ (.Y(_1524_),
    .A(\vgademo.plane_u[17] ));
 sg13g2_inv_1 _6366_ (.Y(_1525_),
    .A(_0047_));
 sg13g2_nand3_1 _6367_ (.B(_1475_),
    .C(\vgademo.plane_u[16] ),
    .A(_1477_),
    .Y(_1526_));
 sg13g2_xnor2_1 _6368_ (.Y(_1527_),
    .A(_1525_),
    .B(_1526_));
 sg13g2_a21oi_1 _6369_ (.A1(_1527_),
    .A2(net53),
    .Y(_1528_),
    .B1(_1220_));
 sg13g2_nor2_1 _6370_ (.A(_1495_),
    .B(_1513_),
    .Y(_1529_));
 sg13g2_a21oi_1 _6371_ (.A1(_1501_),
    .A2(_1529_),
    .Y(_1530_),
    .B1(_1515_));
 sg13g2_inv_1 _6372_ (.Y(_1531_),
    .A(_1530_));
 sg13g2_o21ai_1 _6373_ (.B1(net114),
    .Y(_1532_),
    .A1(_0899_),
    .A2(_1492_));
 sg13g2_xnor2_1 _6374_ (.Y(_1533_),
    .A(_0895_),
    .B(_1532_));
 sg13g2_inv_1 _6375_ (.Y(_1534_),
    .A(_1533_));
 sg13g2_nand2b_1 _6376_ (.Y(_1535_),
    .B(_0892_),
    .A_N(_1511_));
 sg13g2_xnor2_1 _6377_ (.Y(_1536_),
    .A(_1534_),
    .B(_1535_));
 sg13g2_a21oi_1 _6378_ (.A1(_1531_),
    .A2(_1536_),
    .Y(_1537_),
    .B1(net62));
 sg13g2_nor2_1 _6379_ (.A(_1536_),
    .B(_1531_),
    .Y(_1538_));
 sg13g2_inv_1 _6380_ (.Y(_1539_),
    .A(_1538_));
 sg13g2_nand2_1 _6381_ (.Y(_1540_),
    .A(_1537_),
    .B(_1539_));
 sg13g2_a22oi_1 _6382_ (.Y(_0245_),
    .B1(_1528_),
    .B2(_1540_),
    .A2(net32),
    .A1(_1524_));
 sg13g2_inv_1 _6383_ (.Y(_1541_),
    .A(\vgademo.plane_u[18] ));
 sg13g2_nor3_1 _6384_ (.A(_1503_),
    .B(_1524_),
    .C(_1520_),
    .Y(_1542_));
 sg13g2_xnor2_1 _6385_ (.Y(_1543_),
    .A(_0048_),
    .B(_1542_));
 sg13g2_a21oi_1 _6386_ (.A1(_1543_),
    .A2(net53),
    .Y(_1544_),
    .B1(net36));
 sg13g2_inv_1 _6387_ (.Y(_1545_),
    .A(_1457_));
 sg13g2_a22oi_1 _6388_ (.Y(_1546_),
    .B1(_1545_),
    .B2(_1532_),
    .A2(_0864_),
    .A1(net110));
 sg13g2_nor2_1 _6389_ (.A(_1534_),
    .B(_1535_),
    .Y(_1547_));
 sg13g2_inv_1 _6390_ (.Y(_1548_),
    .A(_1547_));
 sg13g2_nand2_1 _6391_ (.Y(_1549_),
    .A(_1539_),
    .B(_1548_));
 sg13g2_inv_1 _6392_ (.Y(_1550_),
    .A(_1549_));
 sg13g2_nor2_1 _6393_ (.A(_1546_),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_inv_1 _6394_ (.Y(_1552_),
    .A(_1551_));
 sg13g2_nand2_1 _6395_ (.Y(_1553_),
    .A(_1550_),
    .B(_1546_));
 sg13g2_nand3_1 _6396_ (.B(_0559_),
    .C(_1553_),
    .A(_1552_),
    .Y(_1554_));
 sg13g2_a22oi_1 _6397_ (.Y(_0246_),
    .B1(_1544_),
    .B2(_1554_),
    .A2(net32),
    .A1(_1541_));
 sg13g2_inv_1 _6398_ (.Y(_1555_),
    .A(\vgademo.plane_u[19] ));
 sg13g2_nand2_1 _6399_ (.Y(_1556_),
    .A(\vgademo.plane_u[17] ),
    .B(\vgademo.plane_u[18] ));
 sg13g2_nor2_1 _6400_ (.A(_1556_),
    .B(_1526_),
    .Y(_1557_));
 sg13g2_xnor2_1 _6401_ (.Y(_1558_),
    .A(_0049_),
    .B(_1557_));
 sg13g2_a21oi_1 _6402_ (.A1(_1558_),
    .A2(net53),
    .Y(_1559_),
    .B1(net36));
 sg13g2_o21ai_1 _6403_ (.B1(_1552_),
    .Y(_1560_),
    .A1(_1506_),
    .A2(_1484_));
 sg13g2_a21oi_1 _6404_ (.A1(_1551_),
    .A2(_1488_),
    .Y(_1561_),
    .B1(_0545_));
 sg13g2_nand2_1 _6405_ (.Y(_1562_),
    .A(_1560_),
    .B(_1561_));
 sg13g2_a22oi_1 _6406_ (.Y(_0247_),
    .B1(_1559_),
    .B2(_1562_),
    .A2(_1227_),
    .A1(_1555_));
 sg13g2_xnor2_1 _6407_ (.Y(_1563_),
    .A(_1214_),
    .B(_1312_));
 sg13g2_nor2_1 _6408_ (.A(_0856_),
    .B(net62),
    .Y(_1564_));
 sg13g2_a21oi_1 _6409_ (.A1(net56),
    .A2(_1563_),
    .Y(_1565_),
    .B1(_1564_));
 sg13g2_nand2_1 _6410_ (.Y(_1566_),
    .A(net37),
    .B(\vgademo.plane_u[1] ));
 sg13g2_o21ai_1 _6411_ (.B1(_1566_),
    .Y(_0248_),
    .A1(net31),
    .A2(_1565_));
 sg13g2_inv_1 _6412_ (.Y(_1567_),
    .A(\vgademo.plane_u[20] ));
 sg13g2_nor2_1 _6413_ (.A(_1487_),
    .B(_1549_),
    .Y(_1568_));
 sg13g2_a21oi_1 _6414_ (.A1(_1551_),
    .A2(_1485_),
    .Y(_1569_),
    .B1(_1568_));
 sg13g2_inv_1 _6415_ (.Y(_1570_),
    .A(_0050_));
 sg13g2_nor4_1 _6416_ (.A(_1503_),
    .B(_1555_),
    .C(_1556_),
    .D(_1520_),
    .Y(_1571_));
 sg13g2_xnor2_1 _6417_ (.Y(_1572_),
    .A(_1570_),
    .B(_1571_));
 sg13g2_a21oi_1 _6418_ (.A1(_1572_),
    .A2(_0545_),
    .Y(_1573_),
    .B1(_1226_));
 sg13g2_o21ai_1 _6419_ (.B1(_1573_),
    .Y(_1574_),
    .A1(_0634_),
    .A2(_1569_));
 sg13g2_o21ai_1 _6420_ (.B1(_1574_),
    .Y(_0249_),
    .A1(_1567_),
    .A2(_1222_));
 sg13g2_inv_1 _6421_ (.Y(_1575_),
    .A(\vgademo.plane_u[21] ));
 sg13g2_nor4_1 _6422_ (.A(_1555_),
    .B(_1567_),
    .C(_1556_),
    .D(_1526_),
    .Y(_1576_));
 sg13g2_xnor2_1 _6423_ (.Y(_1577_),
    .A(_1575_),
    .B(_1576_));
 sg13g2_a21oi_1 _6424_ (.A1(_1577_),
    .A2(net56),
    .Y(_1578_),
    .B1(_1226_));
 sg13g2_o21ai_1 _6425_ (.B1(net45),
    .Y(_1579_),
    .A1(_1486_),
    .A2(_1552_));
 sg13g2_a22oi_1 _6426_ (.Y(_0250_),
    .B1(_1578_),
    .B2(_1579_),
    .A2(_1227_),
    .A1(_1575_));
 sg13g2_nor2_1 _6427_ (.A(_1316_),
    .B(_1319_),
    .Y(_1580_));
 sg13g2_xnor2_1 _6428_ (.Y(_1581_),
    .A(_1580_),
    .B(_1315_));
 sg13g2_nor2_1 _6429_ (.A(_1247_),
    .B(net62),
    .Y(_1582_));
 sg13g2_a21oi_1 _6430_ (.A1(_1581_),
    .A2(net56),
    .Y(_1583_),
    .B1(_1582_));
 sg13g2_mux2_1 _6431_ (.A0(_1583_),
    .A1(\vgademo.plane_u[2] ),
    .S(net31),
    .X(_0251_));
 sg13g2_nor2b_1 _6432_ (.A(_1322_),
    .B_N(_1321_),
    .Y(_1584_));
 sg13g2_xnor2_1 _6433_ (.Y(_1585_),
    .A(_1584_),
    .B(_1320_));
 sg13g2_nor2_1 _6434_ (.A(_0873_),
    .B(_1239_),
    .Y(_1586_));
 sg13g2_nor3_1 _6435_ (.A(_1264_),
    .B(_1586_),
    .C(net63),
    .Y(_1587_));
 sg13g2_a21oi_1 _6436_ (.A1(_1585_),
    .A2(net56),
    .Y(_1588_),
    .B1(_1587_));
 sg13g2_nand2_1 _6437_ (.Y(_1589_),
    .A(net37),
    .B(\vgademo.plane_u[3] ));
 sg13g2_o21ai_1 _6438_ (.B1(_1589_),
    .Y(_0252_),
    .A1(net31),
    .A2(_1588_));
 sg13g2_nor2_1 _6439_ (.A(net112),
    .B(_1265_),
    .Y(_1590_));
 sg13g2_nor2_1 _6440_ (.A(_0876_),
    .B(_1264_),
    .Y(_1591_));
 sg13g2_o21ai_1 _6441_ (.B1(net41),
    .Y(_1592_),
    .A1(_1590_),
    .A2(_1591_));
 sg13g2_nand2_1 _6442_ (.Y(_1593_),
    .A(_1222_),
    .B(_1592_));
 sg13g2_nor2b_1 _6443_ (.A(_1311_),
    .B_N(_1325_),
    .Y(_1594_));
 sg13g2_o21ai_1 _6444_ (.B1(net62),
    .Y(_1595_),
    .A1(_1594_),
    .A2(_1324_));
 sg13g2_a21oi_1 _6445_ (.A1(_1324_),
    .A2(_1594_),
    .Y(_1596_),
    .B1(_1595_));
 sg13g2_nand2_1 _6446_ (.Y(_1597_),
    .A(net37),
    .B(\vgademo.plane_u[4] ));
 sg13g2_o21ai_1 _6447_ (.B1(_1597_),
    .Y(_0253_),
    .A1(_1593_),
    .A2(_1596_));
 sg13g2_inv_1 _6448_ (.Y(_1598_),
    .A(\vgademo.plane_u[5] ));
 sg13g2_nor2b_1 _6449_ (.A(_1590_),
    .B_N(_1263_),
    .Y(_1599_));
 sg13g2_nor3_1 _6450_ (.A(_1266_),
    .B(_1599_),
    .C(net62),
    .Y(_1600_));
 sg13g2_nor2_1 _6451_ (.A(_1600_),
    .B(net37),
    .Y(_1601_));
 sg13g2_nor2b_1 _6452_ (.A(_1310_),
    .B_N(_1328_),
    .Y(_1602_));
 sg13g2_a21oi_1 _6453_ (.A1(_1326_),
    .A2(_1602_),
    .Y(_1603_),
    .B1(net42));
 sg13g2_o21ai_1 _6454_ (.B1(_1603_),
    .Y(_1604_),
    .A1(_1326_),
    .A2(_1602_));
 sg13g2_a22oi_1 _6455_ (.Y(_0254_),
    .B1(_1601_),
    .B2(_1604_),
    .A2(net31),
    .A1(_1598_));
 sg13g2_inv_1 _6456_ (.Y(_1605_),
    .A(\vgademo.plane_u[6] ));
 sg13g2_nor2_1 _6457_ (.A(_1263_),
    .B(_1590_),
    .Y(_1606_));
 sg13g2_xnor2_1 _6458_ (.Y(_1607_),
    .A(_1262_),
    .B(_1248_));
 sg13g2_xnor2_1 _6459_ (.Y(_1608_),
    .A(_1606_),
    .B(_1607_));
 sg13g2_a21oi_1 _6460_ (.A1(net45),
    .A2(_1608_),
    .Y(_1609_),
    .B1(net36));
 sg13g2_a21oi_1 _6461_ (.A1(_1330_),
    .A2(_1339_),
    .Y(_1610_),
    .B1(net42));
 sg13g2_o21ai_1 _6462_ (.B1(_1610_),
    .Y(_1611_),
    .A1(_1339_),
    .A2(_1330_));
 sg13g2_a22oi_1 _6463_ (.Y(_0255_),
    .B1(_1609_),
    .B2(_1611_),
    .A2(net31),
    .A1(_1605_));
 sg13g2_inv_1 _6464_ (.Y(_1612_),
    .A(\vgademo.plane_u[7] ));
 sg13g2_nand2b_1 _6465_ (.Y(_1613_),
    .B(_1267_),
    .A_N(_1361_));
 sg13g2_nand3_1 _6466_ (.B(net45),
    .C(_1363_),
    .A(_1613_),
    .Y(_1614_));
 sg13g2_inv_1 _6467_ (.Y(_1615_),
    .A(_1330_));
 sg13g2_o21ai_1 _6468_ (.B1(_1337_),
    .Y(_1616_),
    .A1(_1336_),
    .A2(_1615_));
 sg13g2_xnor2_1 _6469_ (.Y(_1617_),
    .A(_1335_),
    .B(_1616_));
 sg13g2_a21oi_1 _6470_ (.A1(_1617_),
    .A2(net53),
    .Y(_1618_),
    .B1(net37));
 sg13g2_a22oi_1 _6471_ (.Y(_0256_),
    .B1(_1614_),
    .B2(_1618_),
    .A2(net31),
    .A1(_1612_));
 sg13g2_inv_1 _6472_ (.Y(_1619_),
    .A(\vgademo.plane_u[8] ));
 sg13g2_nand2b_1 _6473_ (.Y(_1620_),
    .B(_1258_),
    .A_N(_1268_));
 sg13g2_nand3_1 _6474_ (.B(net45),
    .C(_1620_),
    .A(_1269_),
    .Y(_1621_));
 sg13g2_xnor2_1 _6475_ (.Y(_1622_),
    .A(_1347_),
    .B(_1342_));
 sg13g2_a21oi_1 _6476_ (.A1(_1622_),
    .A2(net53),
    .Y(_1623_),
    .B1(net37));
 sg13g2_a22oi_1 _6477_ (.Y(_0257_),
    .B1(_1621_),
    .B2(_1623_),
    .A2(net31),
    .A1(_1619_));
 sg13g2_a21oi_1 _6478_ (.A1(_1282_),
    .A2(_1365_),
    .Y(_1624_),
    .B1(net63));
 sg13g2_nor2b_1 _6479_ (.A(_1309_),
    .B_N(_1349_),
    .Y(_1625_));
 sg13g2_a221oi_1 _6480_ (.B2(_1334_),
    .C1(_1333_),
    .B1(_1616_),
    .A1(\vgademo.plane_u[8] ),
    .Y(_1626_),
    .A2(net111));
 sg13g2_nor2_1 _6481_ (.A(_1344_),
    .B(_1626_),
    .Y(_1627_));
 sg13g2_xor2_1 _6482_ (.B(_1627_),
    .A(_1625_),
    .X(_1628_));
 sg13g2_a22oi_1 _6483_ (.Y(_1629_),
    .B1(net56),
    .B2(_1628_),
    .A2(_1624_),
    .A1(_1367_));
 sg13g2_nand2_1 _6484_ (.Y(_1630_),
    .A(net37),
    .B(\vgademo.plane_u[9] ));
 sg13g2_o21ai_1 _6485_ (.B1(_1630_),
    .Y(_0258_),
    .A1(net31),
    .A2(_1629_));
 sg13g2_inv_1 _6486_ (.Y(_1631_),
    .A(\vgademo.scanline_audio_sample[0] ));
 sg13g2_buf_2 _6487_ (.A(\vgademo.soundtrack.tri_osc_p[15] ),
    .X(_1632_));
 sg13g2_buf_1 _6488_ (.A(_1632_),
    .X(_1633_));
 sg13g2_buf_1 _6489_ (.A(\vgademo.soundtrack.tri_osc_p[10] ),
    .X(_1634_));
 sg13g2_xor2_1 _6490_ (.B(_1634_),
    .A(net92),
    .X(_1635_));
 sg13g2_buf_2 _6491_ (.A(\vgademo.audio_snare_frames[3] ),
    .X(_1636_));
 sg13g2_buf_1 _6492_ (.A(_1636_),
    .X(_1637_));
 sg13g2_buf_1 _6493_ (.A(\vgademo.audio_snare_frames[2] ),
    .X(_1638_));
 sg13g2_buf_1 _6494_ (.A(_1638_),
    .X(_1639_));
 sg13g2_buf_1 _6495_ (.A(\vgademo.soundtrack.noise_lfsr[12] ),
    .X(_1640_));
 sg13g2_buf_1 _6496_ (.A(\vgademo.audio_snare_frames[0] ),
    .X(_1641_));
 sg13g2_mux2_1 _6497_ (.A0(\vgademo.soundtrack.noise_lfsr[11] ),
    .A1(_1640_),
    .S(_1641_),
    .X(_1642_));
 sg13g2_buf_1 _6498_ (.A(\vgademo.audio_snare_frames[1] ),
    .X(_1643_));
 sg13g2_inv_1 _6499_ (.Y(_1644_),
    .A(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_nor2_1 _6500_ (.A(_1641_),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_a21oi_1 _6501_ (.A1(_1641_),
    .A2(\vgademo.soundtrack.noise_lfsr[10] ),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_nor2_1 _6502_ (.A(_1643_),
    .B(_1646_),
    .Y(_1647_));
 sg13g2_a21oi_1 _6503_ (.A1(_1642_),
    .A2(net109),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_nor2_1 _6504_ (.A(_1639_),
    .B(_1648_),
    .Y(_1649_));
 sg13g2_inv_1 _6505_ (.Y(_1650_),
    .A(_1649_));
 sg13g2_nor2_1 _6506_ (.A(net91),
    .B(_1650_),
    .Y(_1651_));
 sg13g2_buf_1 _6507_ (.A(\vgademo.soundtrack.pulse_vol[1] ),
    .X(_1652_));
 sg13g2_nor2_1 _6508_ (.A(_1652_),
    .B(\vgademo.soundtrack.pulse_vol[2] ),
    .Y(_1653_));
 sg13g2_nand2_1 _6509_ (.Y(_1654_),
    .A(_1652_),
    .B(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_inv_1 _6510_ (.Y(_1655_),
    .A(_1654_));
 sg13g2_nor2_1 _6511_ (.A(_1653_),
    .B(_1655_),
    .Y(_1656_));
 sg13g2_inv_1 _6512_ (.Y(_1657_),
    .A(_1656_));
 sg13g2_buf_1 _6513_ (.A(\vgademo.soundtrack.pulse_vol[0] ),
    .X(_1658_));
 sg13g2_inv_1 _6514_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_nand2b_1 _6515_ (.Y(_1660_),
    .B(_1659_),
    .A_N(_1652_));
 sg13g2_inv_2 _6516_ (.Y(_1661_),
    .A(_0773_));
 sg13g2_nor2_1 _6517_ (.A(net116),
    .B(_0767_),
    .Y(_1662_));
 sg13g2_inv_1 _6518_ (.Y(_1663_),
    .A(_1662_));
 sg13g2_nand2_1 _6519_ (.Y(_1664_),
    .A(net117),
    .B(_0773_));
 sg13g2_nand2_1 _6520_ (.Y(_1665_),
    .A(_0769_),
    .B(_0771_));
 sg13g2_nor2_1 _6521_ (.A(_1664_),
    .B(_1665_),
    .Y(_1666_));
 sg13g2_a21oi_1 _6522_ (.A1(_1661_),
    .A2(_1663_),
    .Y(_1667_),
    .B1(_1666_));
 sg13g2_nand2_1 _6523_ (.Y(_1668_),
    .A(net117),
    .B(net116));
 sg13g2_buf_2 _6524_ (.A(_1668_),
    .X(_1669_));
 sg13g2_nand2_1 _6525_ (.Y(_1670_),
    .A(_0770_),
    .B(_1669_));
 sg13g2_nor2_1 _6526_ (.A(net97),
    .B(_1661_),
    .Y(_1671_));
 sg13g2_nand2_1 _6527_ (.Y(_1672_),
    .A(_1670_),
    .B(_1671_));
 sg13g2_a21o_1 _6528_ (.A2(_1672_),
    .A1(_1667_),
    .B1(_0763_),
    .X(_1673_));
 sg13g2_inv_1 _6529_ (.Y(_1674_),
    .A(_0763_));
 sg13g2_nor2_1 _6530_ (.A(net97),
    .B(_1674_),
    .Y(_1675_));
 sg13g2_buf_2 _6531_ (.A(_1675_),
    .X(_1676_));
 sg13g2_nand2_1 _6532_ (.Y(_1677_),
    .A(_1670_),
    .B(_1661_));
 sg13g2_nand2_1 _6533_ (.Y(_1678_),
    .A(_0763_),
    .B(_0772_));
 sg13g2_inv_1 _6534_ (.Y(_1679_),
    .A(_1678_));
 sg13g2_nand2_2 _6535_ (.Y(_1680_),
    .A(_1662_),
    .B(_0773_));
 sg13g2_nand2_1 _6536_ (.Y(_1681_),
    .A(_1677_),
    .B(_1680_));
 sg13g2_a22oi_1 _6537_ (.Y(_1682_),
    .B1(_1679_),
    .B2(_1681_),
    .A2(_1677_),
    .A1(_1676_));
 sg13g2_buf_1 _6538_ (.A(_0775_),
    .X(_1683_));
 sg13g2_nand3_1 _6539_ (.B(_1682_),
    .C(net89),
    .A(_1673_),
    .Y(_1684_));
 sg13g2_nand2_1 _6540_ (.Y(_1685_),
    .A(_1684_),
    .B(_0778_));
 sg13g2_nor2_2 _6541_ (.A(_0773_),
    .B(_0767_),
    .Y(_1686_));
 sg13g2_nand2_1 _6542_ (.Y(_1687_),
    .A(_1686_),
    .B(net116));
 sg13g2_nand2_1 _6543_ (.Y(_1688_),
    .A(_1680_),
    .B(_1687_));
 sg13g2_a22oi_1 _6544_ (.Y(_1689_),
    .B1(_1679_),
    .B2(_1688_),
    .A2(_1676_),
    .A1(_1662_));
 sg13g2_buf_1 _6545_ (.A(_0773_),
    .X(_1690_));
 sg13g2_nor2_1 _6546_ (.A(net116),
    .B(net88),
    .Y(_1691_));
 sg13g2_nand2_1 _6547_ (.Y(_1692_),
    .A(net117),
    .B(net97));
 sg13g2_inv_1 _6548_ (.Y(_1693_),
    .A(_1692_));
 sg13g2_inv_1 _6549_ (.Y(_1694_),
    .A(_0770_));
 sg13g2_nor2_1 _6550_ (.A(_1693_),
    .B(_1694_),
    .Y(_1695_));
 sg13g2_nor2_1 _6551_ (.A(_0763_),
    .B(_0774_),
    .Y(_1696_));
 sg13g2_o21ai_1 _6552_ (.B1(_1696_),
    .Y(_1697_),
    .A1(_1691_),
    .A2(_1695_));
 sg13g2_a21oi_1 _6553_ (.A1(_1689_),
    .A2(_1697_),
    .Y(_1698_),
    .B1(net89));
 sg13g2_nand2_1 _6554_ (.Y(_1699_),
    .A(_0767_),
    .B(net116));
 sg13g2_nor2_1 _6555_ (.A(net88),
    .B(_1699_),
    .Y(_1700_));
 sg13g2_buf_1 _6556_ (.A(_1674_),
    .X(_1701_));
 sg13g2_inv_1 _6557_ (.Y(_1702_),
    .A(_0771_));
 sg13g2_nor2_1 _6558_ (.A(net117),
    .B(_0773_),
    .Y(_1703_));
 sg13g2_nor2_1 _6559_ (.A(_1702_),
    .B(_1703_),
    .Y(_1704_));
 sg13g2_inv_1 _6560_ (.Y(_1705_),
    .A(_1704_));
 sg13g2_a22oi_1 _6561_ (.Y(_1706_),
    .B1(net81),
    .B2(_1705_),
    .A2(_1679_),
    .A1(_1700_));
 sg13g2_nand2_1 _6562_ (.Y(_1707_),
    .A(_1706_),
    .B(_0776_));
 sg13g2_o21ai_1 _6563_ (.B1(_0775_),
    .Y(_1708_),
    .A1(_1694_),
    .A2(_1696_));
 sg13g2_nand3_1 _6564_ (.B(_0765_),
    .C(_1708_),
    .A(_1707_),
    .Y(_1709_));
 sg13g2_nand2_1 _6565_ (.Y(_1710_),
    .A(net118),
    .B(_0778_));
 sg13g2_buf_2 _6566_ (.A(_1710_),
    .X(_1711_));
 sg13g2_nand2_1 _6567_ (.Y(_1712_),
    .A(_1709_),
    .B(_1711_));
 sg13g2_o21ai_1 _6568_ (.B1(_1712_),
    .Y(_1713_),
    .A1(_1685_),
    .A2(_1698_));
 sg13g2_mux2_1 _6569_ (.A0(_0062_),
    .A1(_0061_),
    .S(_1713_),
    .X(_1714_));
 sg13g2_buf_1 _6570_ (.A(_1714_),
    .X(_1715_));
 sg13g2_nand2_1 _6571_ (.Y(_1716_),
    .A(net108),
    .B(_1652_));
 sg13g2_o21ai_1 _6572_ (.B1(_1716_),
    .Y(_1717_),
    .A1(_1660_),
    .A2(_1715_));
 sg13g2_nor2b_1 _6573_ (.A(_1657_),
    .B_N(_1717_),
    .Y(_1718_));
 sg13g2_buf_2 _6574_ (.A(\vgademo.soundtrack.pulse_vol[3] ),
    .X(_1719_));
 sg13g2_inv_2 _6575_ (.Y(_1720_),
    .A(_1719_));
 sg13g2_nand2_1 _6576_ (.Y(_1721_),
    .A(_1718_),
    .B(_1720_));
 sg13g2_xor2_1 _6577_ (.B(_1721_),
    .A(_1651_),
    .X(_1722_));
 sg13g2_xor2_1 _6578_ (.B(_1722_),
    .A(_1635_),
    .X(_1723_));
 sg13g2_xnor2_1 _6579_ (.Y(_1724_),
    .A(net92),
    .B(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_nand2_1 _6580_ (.Y(_1725_),
    .A(_1715_),
    .B(net108));
 sg13g2_buf_2 _6581_ (.A(_1725_),
    .X(_1726_));
 sg13g2_inv_1 _6582_ (.Y(_1727_),
    .A(\vgademo.soundtrack.pulse_vol[2] ));
 sg13g2_nor3_1 _6583_ (.A(_1652_),
    .B(_1719_),
    .C(_1727_),
    .Y(_1728_));
 sg13g2_buf_1 _6584_ (.A(net109),
    .X(_1729_));
 sg13g2_buf_1 _6585_ (.A(_1641_),
    .X(_1730_));
 sg13g2_inv_1 _6586_ (.Y(_1731_),
    .A(\vgademo.soundtrack.noise_lfsr[10] ));
 sg13g2_nand2_1 _6587_ (.Y(_1732_),
    .A(net86),
    .B(\vgademo.soundtrack.noise_lfsr[11] ));
 sg13g2_o21ai_1 _6588_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net86),
    .A2(_1731_));
 sg13g2_buf_1 _6589_ (.A(_1641_),
    .X(_1734_));
 sg13g2_nand2_1 _6590_ (.Y(_1735_),
    .A(_1644_),
    .B(net85));
 sg13g2_o21ai_1 _6591_ (.B1(_1735_),
    .Y(_1736_),
    .A1(net85),
    .A2(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_nor2_1 _6592_ (.A(net109),
    .B(_1736_),
    .Y(_1737_));
 sg13g2_a21oi_1 _6593_ (.A1(_1729_),
    .A2(_1733_),
    .Y(_1738_),
    .B1(_1737_));
 sg13g2_inv_1 _6594_ (.Y(_1739_),
    .A(_1638_));
 sg13g2_buf_1 _6595_ (.A(_1739_),
    .X(_1740_));
 sg13g2_nor2_1 _6596_ (.A(net109),
    .B(_1730_),
    .Y(_1741_));
 sg13g2_a21oi_1 _6597_ (.A1(_1741_),
    .A2(_1640_),
    .Y(_1742_),
    .B1(_1739_));
 sg13g2_a21o_1 _6598_ (.A2(net80),
    .A1(_1738_),
    .B1(_1742_),
    .X(_1743_));
 sg13g2_nor2_1 _6599_ (.A(net91),
    .B(_1743_),
    .Y(_1744_));
 sg13g2_a21oi_1 _6600_ (.A1(_1726_),
    .A2(_1728_),
    .Y(_1745_),
    .B1(_1744_));
 sg13g2_nand3_1 _6601_ (.B(_1728_),
    .C(_1744_),
    .A(_1726_),
    .Y(_1746_));
 sg13g2_o21ai_1 _6602_ (.B1(_1746_),
    .Y(_1747_),
    .A1(_1724_),
    .A2(_1745_));
 sg13g2_nor2b_1 _6603_ (.A(_1723_),
    .B_N(_1747_),
    .Y(_1748_));
 sg13g2_nand2b_1 _6604_ (.Y(_1749_),
    .B(_1723_),
    .A_N(_1747_));
 sg13g2_nor2b_1 _6605_ (.A(_1748_),
    .B_N(_1749_),
    .Y(_1750_));
 sg13g2_nor2b_1 _6606_ (.A(_1745_),
    .B_N(_1746_),
    .Y(_1751_));
 sg13g2_xor2_1 _6607_ (.B(_1751_),
    .A(_1724_),
    .X(_1752_));
 sg13g2_inv_1 _6608_ (.Y(_1753_),
    .A(\vgademo.soundtrack.noise_lfsr[7] ));
 sg13g2_nand2_1 _6609_ (.Y(_1754_),
    .A(net85),
    .B(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_o21ai_1 _6610_ (.B1(_1754_),
    .Y(_1755_),
    .A1(net85),
    .A2(_1753_));
 sg13g2_nor2_1 _6611_ (.A(net87),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_a21oi_1 _6612_ (.A1(net87),
    .A2(_1646_),
    .Y(_1757_),
    .B1(_1756_));
 sg13g2_inv_2 _6613_ (.Y(_1758_),
    .A(_1643_));
 sg13g2_nand2_1 _6614_ (.Y(_1759_),
    .A(_1642_),
    .B(_1758_));
 sg13g2_a21oi_1 _6615_ (.A1(_1759_),
    .A2(net90),
    .Y(_1760_),
    .B1(_1637_));
 sg13g2_o21ai_1 _6616_ (.B1(_1760_),
    .Y(_1761_),
    .A1(net90),
    .A2(_1757_));
 sg13g2_nor4_1 _6617_ (.A(net108),
    .B(_1719_),
    .C(_1654_),
    .D(_1715_),
    .Y(_1762_));
 sg13g2_a21o_1 _6618_ (.A2(_1728_),
    .A1(net108),
    .B1(_1762_),
    .X(_1763_));
 sg13g2_nor2b_1 _6619_ (.A(_1761_),
    .B_N(_1763_),
    .Y(_1764_));
 sg13g2_xor2_1 _6620_ (.B(_1763_),
    .A(_1761_),
    .X(_1765_));
 sg13g2_buf_1 _6621_ (.A(\vgademo.soundtrack.tri_osc_p[8] ),
    .X(_1766_));
 sg13g2_xor2_1 _6622_ (.B(_1766_),
    .A(net92),
    .X(_1767_));
 sg13g2_nor2b_1 _6623_ (.A(_1765_),
    .B_N(_1767_),
    .Y(_1768_));
 sg13g2_nor2_1 _6624_ (.A(_1764_),
    .B(_1768_),
    .Y(_1769_));
 sg13g2_nor2_1 _6625_ (.A(_1752_),
    .B(_1769_),
    .Y(_1770_));
 sg13g2_xor2_1 _6626_ (.B(_1765_),
    .A(_1767_),
    .X(_1771_));
 sg13g2_inv_1 _6627_ (.Y(_1772_),
    .A(net85));
 sg13g2_nand2_1 _6628_ (.Y(_1773_),
    .A(net109),
    .B(_1640_));
 sg13g2_inv_1 _6629_ (.Y(_1774_),
    .A(_1773_));
 sg13g2_a22oi_1 _6630_ (.Y(_1775_),
    .B1(_1758_),
    .B2(_1733_),
    .A2(_1774_),
    .A1(_1772_));
 sg13g2_nand2_1 _6631_ (.Y(_1776_),
    .A(_1753_),
    .B(net85));
 sg13g2_o21ai_1 _6632_ (.B1(_1776_),
    .Y(_1777_),
    .A1(_1734_),
    .A2(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_mux2_1 _6633_ (.A0(_1777_),
    .A1(_1736_),
    .S(net109),
    .X(_1778_));
 sg13g2_a21o_1 _6634_ (.A2(net80),
    .A1(_1778_),
    .B1(_1637_),
    .X(_1779_));
 sg13g2_a21oi_1 _6635_ (.A1(net90),
    .A2(_1775_),
    .Y(_1780_),
    .B1(_1779_));
 sg13g2_nand3_1 _6636_ (.B(_1720_),
    .C(_1655_),
    .A(_1726_),
    .Y(_1781_));
 sg13g2_xor2_1 _6637_ (.B(_1781_),
    .A(_1780_),
    .X(_1782_));
 sg13g2_buf_1 _6638_ (.A(\vgademo.soundtrack.tri_osc_p[7] ),
    .X(_1783_));
 sg13g2_xor2_1 _6639_ (.B(_1783_),
    .A(net92),
    .X(_1784_));
 sg13g2_nand2b_1 _6640_ (.Y(_1785_),
    .B(_1784_),
    .A_N(_1782_));
 sg13g2_nand2b_1 _6641_ (.Y(_1786_),
    .B(_1780_),
    .A_N(_1781_));
 sg13g2_nand2_1 _6642_ (.Y(_1787_),
    .A(_1785_),
    .B(_1786_));
 sg13g2_nor2b_1 _6643_ (.A(_1771_),
    .B_N(_1787_),
    .Y(_1788_));
 sg13g2_nand2_1 _6644_ (.Y(_1789_),
    .A(_1717_),
    .B(_1657_));
 sg13g2_inv_1 _6645_ (.Y(_1790_),
    .A(_1789_));
 sg13g2_nor2_1 _6646_ (.A(_1720_),
    .B(_1654_),
    .Y(_1791_));
 sg13g2_nor2_1 _6647_ (.A(_1719_),
    .B(_1655_),
    .Y(_1792_));
 sg13g2_nor2_1 _6648_ (.A(_1791_),
    .B(_1792_),
    .Y(_1793_));
 sg13g2_nand2_1 _6649_ (.Y(_1794_),
    .A(_1790_),
    .B(_1793_));
 sg13g2_nand2_1 _6650_ (.Y(_1795_),
    .A(_1648_),
    .B(net90));
 sg13g2_inv_1 _6651_ (.Y(_1796_),
    .A(\vgademo.soundtrack.noise_lfsr[5] ));
 sg13g2_nor2_1 _6652_ (.A(_1641_),
    .B(_1796_),
    .Y(_1797_));
 sg13g2_a21oi_1 _6653_ (.A1(_1734_),
    .A2(\vgademo.soundtrack.noise_lfsr[6] ),
    .Y(_1798_),
    .B1(_1797_));
 sg13g2_nor2_1 _6654_ (.A(net109),
    .B(_1798_),
    .Y(_1799_));
 sg13g2_a21oi_1 _6655_ (.A1(net109),
    .A2(_1755_),
    .Y(_1800_),
    .B1(_1799_));
 sg13g2_nand2_1 _6656_ (.Y(_1801_),
    .A(_1800_),
    .B(net80));
 sg13g2_inv_2 _6657_ (.Y(_1802_),
    .A(_1636_));
 sg13g2_nand3_1 _6658_ (.B(_1801_),
    .C(_1802_),
    .A(_1795_),
    .Y(_1803_));
 sg13g2_nand2_1 _6659_ (.Y(_1804_),
    .A(_1794_),
    .B(_1803_));
 sg13g2_buf_1 _6660_ (.A(\vgademo.soundtrack.tri_osc_p[6] ),
    .X(_1805_));
 sg13g2_xor2_1 _6661_ (.B(_1805_),
    .A(net92),
    .X(_1806_));
 sg13g2_nor2_1 _6662_ (.A(_1803_),
    .B(_1794_),
    .Y(_1807_));
 sg13g2_a21oi_1 _6663_ (.A1(_1804_),
    .A2(_1806_),
    .Y(_1808_),
    .B1(_1807_));
 sg13g2_xor2_1 _6664_ (.B(_1782_),
    .A(_1784_),
    .X(_1809_));
 sg13g2_nand2_1 _6665_ (.Y(_1810_),
    .A(_1726_),
    .B(_1653_));
 sg13g2_inv_1 _6666_ (.Y(_1811_),
    .A(_1810_));
 sg13g2_nand2_1 _6667_ (.Y(_1812_),
    .A(_1811_),
    .B(_1719_));
 sg13g2_nand3_1 _6668_ (.B(net80),
    .C(_1640_),
    .A(_1741_),
    .Y(_1813_));
 sg13g2_nand2_1 _6669_ (.Y(_1814_),
    .A(_1738_),
    .B(net90));
 sg13g2_nand2_1 _6670_ (.Y(_1815_),
    .A(net85),
    .B(\vgademo.soundtrack.noise_lfsr[5] ));
 sg13g2_o21ai_1 _6671_ (.B1(_1815_),
    .Y(_1816_),
    .A1(net86),
    .A2(_0063_));
 sg13g2_nor2_1 _6672_ (.A(_1758_),
    .B(_1777_),
    .Y(_1817_));
 sg13g2_a21oi_1 _6673_ (.A1(_1758_),
    .A2(_1816_),
    .Y(_1818_),
    .B1(_1817_));
 sg13g2_nand2_1 _6674_ (.Y(_1819_),
    .A(_1818_),
    .B(net80));
 sg13g2_a21oi_1 _6675_ (.A1(_1814_),
    .A2(_1819_),
    .Y(_1820_),
    .B1(_1636_));
 sg13g2_a21oi_1 _6676_ (.A1(net91),
    .A2(_1813_),
    .Y(_1821_),
    .B1(_1820_));
 sg13g2_nor2b_1 _6677_ (.A(_1812_),
    .B_N(_1821_),
    .Y(_1822_));
 sg13g2_xor2_1 _6678_ (.B(_1812_),
    .A(_1821_),
    .X(_1823_));
 sg13g2_buf_1 _6679_ (.A(\vgademo.soundtrack.tri_osc_p[5] ),
    .X(_1824_));
 sg13g2_xor2_1 _6680_ (.B(_1824_),
    .A(_1632_),
    .X(_1825_));
 sg13g2_nor2b_1 _6681_ (.A(_1823_),
    .B_N(_1825_),
    .Y(_1826_));
 sg13g2_nor2_1 _6682_ (.A(_1822_),
    .B(_1826_),
    .Y(_1827_));
 sg13g2_nor2b_1 _6683_ (.A(_1807_),
    .B_N(_1804_),
    .Y(_1828_));
 sg13g2_xnor2_1 _6684_ (.Y(_1829_),
    .A(_1806_),
    .B(_1828_));
 sg13g2_nor2_1 _6685_ (.A(_1827_),
    .B(_1829_),
    .Y(_1830_));
 sg13g2_nand3_1 _6686_ (.B(_1727_),
    .C(_1716_),
    .A(_1660_),
    .Y(_1831_));
 sg13g2_a21oi_1 _6687_ (.A1(_1715_),
    .A2(_1659_),
    .Y(_1832_),
    .B1(_1831_));
 sg13g2_nand2_1 _6688_ (.Y(_1833_),
    .A(_1832_),
    .B(_1719_));
 sg13g2_nand3_1 _6689_ (.B(_1758_),
    .C(net80),
    .A(_1642_),
    .Y(_1834_));
 sg13g2_nand2_1 _6690_ (.Y(_1835_),
    .A(_1757_),
    .B(_1639_));
 sg13g2_nor2_1 _6691_ (.A(net85),
    .B(\vgademo.soundtrack.noise_lfsr[3] ),
    .Y(_1836_));
 sg13g2_a21oi_1 _6692_ (.A1(net86),
    .A2(_0063_),
    .Y(_1837_),
    .B1(_1836_));
 sg13g2_nor2_1 _6693_ (.A(net87),
    .B(_1837_),
    .Y(_1838_));
 sg13g2_a21oi_1 _6694_ (.A1(net87),
    .A2(_1798_),
    .Y(_1839_),
    .B1(_1838_));
 sg13g2_a21oi_1 _6695_ (.A1(_1839_),
    .A2(_1740_),
    .Y(_1840_),
    .B1(_1636_));
 sg13g2_a22oi_1 _6696_ (.Y(_1841_),
    .B1(_1835_),
    .B2(_1840_),
    .A2(_1834_),
    .A1(_1636_));
 sg13g2_nor2b_1 _6697_ (.A(_1833_),
    .B_N(_1841_),
    .Y(_1842_));
 sg13g2_xor2_1 _6698_ (.B(_1833_),
    .A(_1841_),
    .X(_1843_));
 sg13g2_buf_1 _6699_ (.A(\vgademo.soundtrack.tri_osc_p[4] ),
    .X(_1844_));
 sg13g2_xor2_1 _6700_ (.B(_1844_),
    .A(_1632_),
    .X(_1845_));
 sg13g2_nor2b_1 _6701_ (.A(_1843_),
    .B_N(_1845_),
    .Y(_1846_));
 sg13g2_nor2_1 _6702_ (.A(_1842_),
    .B(_1846_),
    .Y(_1847_));
 sg13g2_xor2_1 _6703_ (.B(_1823_),
    .A(_1825_),
    .X(_1848_));
 sg13g2_nand3_1 _6704_ (.B(_1652_),
    .C(_1727_),
    .A(_1726_),
    .Y(_1849_));
 sg13g2_inv_1 _6705_ (.Y(_1850_),
    .A(_1849_));
 sg13g2_nand2_1 _6706_ (.Y(_1851_),
    .A(_1850_),
    .B(_1719_));
 sg13g2_nand2b_1 _6707_ (.Y(_1852_),
    .B(_1740_),
    .A_N(_1775_));
 sg13g2_nor2_1 _6708_ (.A(_1758_),
    .B(_1816_),
    .Y(_1853_));
 sg13g2_mux2_1 _6709_ (.A0(\vgademo.soundtrack.noise_lfsr[2] ),
    .A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .S(net86),
    .X(_1854_));
 sg13g2_nor2_1 _6710_ (.A(net87),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_o21ai_1 _6711_ (.B1(_1739_),
    .Y(_1856_),
    .A1(_1853_),
    .A2(_1855_));
 sg13g2_nand2_1 _6712_ (.Y(_1857_),
    .A(_1778_),
    .B(net90));
 sg13g2_nand3_1 _6713_ (.B(_1857_),
    .C(_1802_),
    .A(_1856_),
    .Y(_1858_));
 sg13g2_o21ai_1 _6714_ (.B1(_1858_),
    .Y(_1859_),
    .A1(_1802_),
    .A2(_1852_));
 sg13g2_nor2b_1 _6715_ (.A(_1851_),
    .B_N(_1859_),
    .Y(_1860_));
 sg13g2_xor2_1 _6716_ (.B(_1851_),
    .A(_1859_),
    .X(_1861_));
 sg13g2_buf_1 _6717_ (.A(\vgademo.soundtrack.tri_osc_p[3] ),
    .X(_1862_));
 sg13g2_xor2_1 _6718_ (.B(_1862_),
    .A(_1632_),
    .X(_1863_));
 sg13g2_nor2b_1 _6719_ (.A(_1861_),
    .B_N(_1863_),
    .Y(_1864_));
 sg13g2_nor2_1 _6720_ (.A(_1860_),
    .B(_1864_),
    .Y(_1865_));
 sg13g2_xor2_1 _6721_ (.B(_1843_),
    .A(_1845_),
    .X(_1866_));
 sg13g2_nand2_1 _6722_ (.Y(_1867_),
    .A(_1718_),
    .B(_1793_));
 sg13g2_nand2_1 _6723_ (.Y(_1868_),
    .A(_1800_),
    .B(net90));
 sg13g2_mux2_1 _6724_ (.A0(\vgademo.soundtrack.noise_lfsr[1] ),
    .A1(\vgademo.soundtrack.noise_lfsr[2] ),
    .S(net86),
    .X(_1869_));
 sg13g2_nand2_1 _6725_ (.Y(_1870_),
    .A(_1869_),
    .B(_1758_));
 sg13g2_nand2_1 _6726_ (.Y(_1871_),
    .A(_1837_),
    .B(net87));
 sg13g2_nand3_1 _6727_ (.B(_1739_),
    .C(_1871_),
    .A(_1870_),
    .Y(_1872_));
 sg13g2_nand3_1 _6728_ (.B(_1872_),
    .C(_1802_),
    .A(_1868_),
    .Y(_1873_));
 sg13g2_o21ai_1 _6729_ (.B1(_1873_),
    .Y(_1874_),
    .A1(_1802_),
    .A2(_1650_));
 sg13g2_nor2b_1 _6730_ (.A(_1867_),
    .B_N(_1874_),
    .Y(_1875_));
 sg13g2_xor2_1 _6731_ (.B(_1867_),
    .A(_1874_),
    .X(_1876_));
 sg13g2_buf_1 _6732_ (.A(\vgademo.soundtrack.tri_osc_p[2] ),
    .X(_1877_));
 sg13g2_xor2_1 _6733_ (.B(_1877_),
    .A(_1632_),
    .X(_1878_));
 sg13g2_nor2b_1 _6734_ (.A(_1876_),
    .B_N(_1878_),
    .Y(_1879_));
 sg13g2_nor2_1 _6735_ (.A(_1875_),
    .B(_1879_),
    .Y(_1880_));
 sg13g2_xor2_1 _6736_ (.B(_1861_),
    .A(_1863_),
    .X(_1881_));
 sg13g2_xor2_1 _6737_ (.B(_1880_),
    .A(_1881_),
    .X(_1882_));
 sg13g2_xor2_1 _6738_ (.B(_1876_),
    .A(_1878_),
    .X(_1883_));
 sg13g2_buf_1 _6739_ (.A(\vgademo.soundtrack.tri_osc_p[1] ),
    .X(_1884_));
 sg13g2_xor2_1 _6740_ (.B(_1884_),
    .A(_1632_),
    .X(_1885_));
 sg13g2_inv_1 _6741_ (.Y(_1886_),
    .A(_1885_));
 sg13g2_nand2_1 _6742_ (.Y(_1887_),
    .A(_1818_),
    .B(net90));
 sg13g2_nand2_1 _6743_ (.Y(_1888_),
    .A(_1772_),
    .B(\vgademo.soundtrack.noise_lfsr[0] ));
 sg13g2_nand2_1 _6744_ (.Y(_1889_),
    .A(net86),
    .B(\vgademo.soundtrack.noise_lfsr[1] ));
 sg13g2_a21oi_1 _6745_ (.A1(_1888_),
    .A2(_1889_),
    .Y(_1890_),
    .B1(net87));
 sg13g2_a21oi_1 _6746_ (.A1(_1854_),
    .A2(net87),
    .Y(_1891_),
    .B1(_1890_));
 sg13g2_nand2_1 _6747_ (.Y(_1892_),
    .A(_1891_),
    .B(_1739_));
 sg13g2_a21oi_1 _6748_ (.A1(_1887_),
    .A2(_1892_),
    .Y(_1893_),
    .B1(_1636_));
 sg13g2_a21oi_1 _6749_ (.A1(_1743_),
    .A2(_1636_),
    .Y(_1894_),
    .B1(_1893_));
 sg13g2_nor3_1 _6750_ (.A(_1652_),
    .B(_1720_),
    .C(_1727_),
    .Y(_1895_));
 sg13g2_nand2_1 _6751_ (.Y(_1896_),
    .A(_1726_),
    .B(_1895_));
 sg13g2_xor2_1 _6752_ (.B(_1896_),
    .A(_1894_),
    .X(_1897_));
 sg13g2_nand3_1 _6753_ (.B(_1895_),
    .C(_1894_),
    .A(_1726_),
    .Y(_1898_));
 sg13g2_o21ai_1 _6754_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_1886_),
    .A2(_1897_));
 sg13g2_nor2b_1 _6755_ (.A(_1883_),
    .B_N(_1899_),
    .Y(_1900_));
 sg13g2_nand2_1 _6756_ (.Y(_1901_),
    .A(_1882_),
    .B(_1900_));
 sg13g2_o21ai_1 _6757_ (.B1(_1901_),
    .Y(_1902_),
    .A1(_1880_),
    .A2(_1881_));
 sg13g2_xor2_1 _6758_ (.B(_1865_),
    .A(_1866_),
    .X(_1903_));
 sg13g2_nand2_1 _6759_ (.Y(_1904_),
    .A(_1902_),
    .B(_1903_));
 sg13g2_o21ai_1 _6760_ (.B1(_1904_),
    .Y(_1905_),
    .A1(_1865_),
    .A2(_1866_));
 sg13g2_xor2_1 _6761_ (.B(_1848_),
    .A(_1847_),
    .X(_1906_));
 sg13g2_nand2_1 _6762_ (.Y(_1907_),
    .A(_1905_),
    .B(_1906_));
 sg13g2_o21ai_1 _6763_ (.B1(_1907_),
    .Y(_1908_),
    .A1(_1847_),
    .A2(_1848_));
 sg13g2_xnor2_1 _6764_ (.Y(_1909_),
    .A(_1827_),
    .B(_1829_));
 sg13g2_inv_1 _6765_ (.Y(_1910_),
    .A(_1909_));
 sg13g2_nand2_1 _6766_ (.Y(_1911_),
    .A(_1908_),
    .B(_1910_));
 sg13g2_nand2b_1 _6767_ (.Y(_1912_),
    .B(_1911_),
    .A_N(_1830_));
 sg13g2_xor2_1 _6768_ (.B(_1808_),
    .A(_1809_),
    .X(_1913_));
 sg13g2_nand2_1 _6769_ (.Y(_1914_),
    .A(_1912_),
    .B(_1913_));
 sg13g2_o21ai_1 _6770_ (.B1(_1914_),
    .Y(_1915_),
    .A1(_1808_),
    .A2(_1809_));
 sg13g2_xnor2_1 _6771_ (.Y(_1916_),
    .A(_1787_),
    .B(_1771_));
 sg13g2_nand2_1 _6772_ (.Y(_1917_),
    .A(_1915_),
    .B(_1916_));
 sg13g2_nand2b_1 _6773_ (.Y(_1918_),
    .B(_1917_),
    .A_N(_1788_));
 sg13g2_nor2_1 _6774_ (.A(_1770_),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_nand2_1 _6775_ (.Y(_1920_),
    .A(_1769_),
    .B(_1752_));
 sg13g2_nor2b_1 _6776_ (.A(_1919_),
    .B_N(_1920_),
    .Y(_1921_));
 sg13g2_xor2_1 _6777_ (.B(_1921_),
    .A(_1750_),
    .X(_1922_));
 sg13g2_nand2_1 _6778_ (.Y(_1923_),
    .A(_1922_),
    .B(_0860_));
 sg13g2_o21ai_1 _6779_ (.B1(_1923_),
    .Y(_0261_),
    .A1(_1631_),
    .A2(net67));
 sg13g2_buf_1 _6780_ (.A(\vgademo.soundtrack.tri_osc_p[11] ),
    .X(_1924_));
 sg13g2_xor2_1 _6781_ (.B(_1924_),
    .A(net92),
    .X(_1925_));
 sg13g2_nor2_1 _6782_ (.A(net91),
    .B(_1852_),
    .Y(_1926_));
 sg13g2_nand2_1 _6783_ (.Y(_1927_),
    .A(_1850_),
    .B(_1720_));
 sg13g2_xor2_1 _6784_ (.B(_1927_),
    .A(_1926_),
    .X(_1928_));
 sg13g2_xor2_1 _6785_ (.B(_1928_),
    .A(_1925_),
    .X(_1929_));
 sg13g2_nor2b_1 _6786_ (.A(_1721_),
    .B_N(_1651_),
    .Y(_1930_));
 sg13g2_nor2b_1 _6787_ (.A(_1722_),
    .B_N(_1635_),
    .Y(_1931_));
 sg13g2_nor2_1 _6788_ (.A(_1930_),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_nor2_1 _6789_ (.A(_1929_),
    .B(_1932_),
    .Y(_1933_));
 sg13g2_inv_1 _6790_ (.Y(_1934_),
    .A(_1933_));
 sg13g2_nand2_1 _6791_ (.Y(_1935_),
    .A(_1932_),
    .B(_1929_));
 sg13g2_nand2_1 _6792_ (.Y(_1936_),
    .A(_1934_),
    .B(_1935_));
 sg13g2_nor2b_1 _6793_ (.A(_1770_),
    .B_N(_1920_),
    .Y(_1937_));
 sg13g2_nand2_1 _6794_ (.Y(_1938_),
    .A(_1937_),
    .B(_1750_));
 sg13g2_inv_1 _6795_ (.Y(_1939_),
    .A(_1918_));
 sg13g2_a21oi_1 _6796_ (.A1(_1770_),
    .A2(_1749_),
    .Y(_1940_),
    .B1(_1748_));
 sg13g2_o21ai_1 _6797_ (.B1(_1940_),
    .Y(_1941_),
    .A1(_1938_),
    .A2(_1939_));
 sg13g2_xnor2_1 _6798_ (.Y(_1942_),
    .A(_1936_),
    .B(_1941_));
 sg13g2_inv_1 _6799_ (.Y(_1943_),
    .A(_1942_));
 sg13g2_nor2_1 _6800_ (.A(\vgademo.scanline_audio_sample[1] ),
    .B(net66),
    .Y(_1944_));
 sg13g2_a21oi_1 _6801_ (.A1(_1943_),
    .A2(net67),
    .Y(_0262_),
    .B1(_1944_));
 sg13g2_inv_1 _6802_ (.Y(_1945_),
    .A(\vgademo.scanline_audio_sample[2] ));
 sg13g2_xor2_1 _6803_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .A(net92),
    .X(_1946_));
 sg13g2_nor2_1 _6804_ (.A(net91),
    .B(_1834_),
    .Y(_1947_));
 sg13g2_nand2_1 _6805_ (.Y(_1948_),
    .A(_1832_),
    .B(_1720_));
 sg13g2_xor2_1 _6806_ (.B(_1948_),
    .A(_1947_),
    .X(_1949_));
 sg13g2_xor2_1 _6807_ (.B(_1949_),
    .A(_1946_),
    .X(_1950_));
 sg13g2_nor2b_1 _6808_ (.A(_1927_),
    .B_N(_1926_),
    .Y(_1951_));
 sg13g2_nor2b_1 _6809_ (.A(_1928_),
    .B_N(_1925_),
    .Y(_1952_));
 sg13g2_nor2_1 _6810_ (.A(_1951_),
    .B(_1952_),
    .Y(_1953_));
 sg13g2_xnor2_1 _6811_ (.Y(_1954_),
    .A(_1950_),
    .B(_1953_));
 sg13g2_nand2_1 _6812_ (.Y(_1955_),
    .A(_1921_),
    .B(_1750_));
 sg13g2_o21ai_1 _6813_ (.B1(_1935_),
    .Y(_1956_),
    .A1(_1933_),
    .A2(_1748_));
 sg13g2_o21ai_1 _6814_ (.B1(_1956_),
    .Y(_1957_),
    .A1(_1936_),
    .A2(_1955_));
 sg13g2_xnor2_1 _6815_ (.Y(_1958_),
    .A(_1954_),
    .B(_1957_));
 sg13g2_nand2_1 _6816_ (.Y(_1959_),
    .A(_1958_),
    .B(_0860_));
 sg13g2_o21ai_1 _6817_ (.B1(_1959_),
    .Y(_0263_),
    .A1(_1945_),
    .A2(net67));
 sg13g2_nor2b_1 _6818_ (.A(_1948_),
    .B_N(_1947_),
    .Y(_1960_));
 sg13g2_nor2b_1 _6819_ (.A(_1949_),
    .B_N(_1946_),
    .Y(_1961_));
 sg13g2_nor2_1 _6820_ (.A(_1960_),
    .B(_1961_),
    .Y(_1962_));
 sg13g2_xor2_1 _6821_ (.B(\vgademo.soundtrack.tri_osc_p[13] ),
    .A(net92),
    .X(_1963_));
 sg13g2_nor2_1 _6822_ (.A(net91),
    .B(_1813_),
    .Y(_1964_));
 sg13g2_nand2_1 _6823_ (.Y(_1965_),
    .A(_1811_),
    .B(_1720_));
 sg13g2_xor2_1 _6824_ (.B(_1965_),
    .A(_1964_),
    .X(_1966_));
 sg13g2_xor2_1 _6825_ (.B(_1966_),
    .A(_1963_),
    .X(_1967_));
 sg13g2_nor2_1 _6826_ (.A(_1962_),
    .B(_1967_),
    .Y(_1968_));
 sg13g2_inv_1 _6827_ (.Y(_1969_),
    .A(_1968_));
 sg13g2_nand2_1 _6828_ (.Y(_1970_),
    .A(_1967_),
    .B(_1962_));
 sg13g2_nand2_1 _6829_ (.Y(_1971_),
    .A(_1969_),
    .B(_1970_));
 sg13g2_inv_1 _6830_ (.Y(_1972_),
    .A(_1971_));
 sg13g2_inv_1 _6831_ (.Y(_1973_),
    .A(_1954_));
 sg13g2_nor2_1 _6832_ (.A(_1954_),
    .B(_1936_),
    .Y(_1974_));
 sg13g2_nor2_1 _6833_ (.A(_1950_),
    .B(_1953_),
    .Y(_1975_));
 sg13g2_a221oi_1 _6834_ (.B2(_1974_),
    .C1(_1975_),
    .B1(_1941_),
    .A1(_1933_),
    .Y(_1976_),
    .A2(_1973_));
 sg13g2_xnor2_1 _6835_ (.Y(_1977_),
    .A(_1972_),
    .B(_1976_));
 sg13g2_inv_1 _6836_ (.Y(_1978_),
    .A(_1977_));
 sg13g2_buf_2 _6837_ (.A(\vgademo.scanline_audio_sample[3] ),
    .X(_1979_));
 sg13g2_nor2_1 _6838_ (.A(_1979_),
    .B(_0860_),
    .Y(_1980_));
 sg13g2_a21oi_1 _6839_ (.A1(_1978_),
    .A2(net67),
    .Y(_0264_),
    .B1(_1980_));
 sg13g2_buf_1 _6840_ (.A(\vgademo.scanline_audio_sample[4] ),
    .X(_1981_));
 sg13g2_xnor2_1 _6841_ (.Y(_1982_),
    .A(\vgademo.soundtrack.tri_osc_p[14] ),
    .B(_1633_));
 sg13g2_nand2_1 _6842_ (.Y(_1983_),
    .A(_1790_),
    .B(_1792_));
 sg13g2_xor2_1 _6843_ (.B(_1983_),
    .A(_1982_),
    .X(_1984_));
 sg13g2_nor2b_1 _6844_ (.A(_1965_),
    .B_N(_1964_),
    .Y(_1985_));
 sg13g2_nand2b_1 _6845_ (.Y(_1986_),
    .B(_1963_),
    .A_N(_1966_));
 sg13g2_nor2b_1 _6846_ (.A(_1985_),
    .B_N(_1986_),
    .Y(_1987_));
 sg13g2_nor2_1 _6847_ (.A(_1984_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_and2_1 _6848_ (.A(_1987_),
    .B(_1984_),
    .X(_1989_));
 sg13g2_nor2_1 _6849_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_));
 sg13g2_nor2_1 _6850_ (.A(_1971_),
    .B(_1954_),
    .Y(_1991_));
 sg13g2_a21oi_1 _6851_ (.A1(_1975_),
    .A2(_1970_),
    .Y(_1992_),
    .B1(_1968_));
 sg13g2_inv_1 _6852_ (.Y(_1993_),
    .A(_1992_));
 sg13g2_a21oi_1 _6853_ (.A1(_1957_),
    .A2(_1991_),
    .Y(_1994_),
    .B1(_1993_));
 sg13g2_xnor2_1 _6854_ (.Y(_1995_),
    .A(_1990_),
    .B(_1994_));
 sg13g2_mux2_1 _6855_ (.A0(_1981_),
    .A1(_1995_),
    .S(net67),
    .X(_0265_));
 sg13g2_nand2_1 _6856_ (.Y(_1996_),
    .A(_1983_),
    .B(_1982_));
 sg13g2_nand2_1 _6857_ (.Y(_1997_),
    .A(_1990_),
    .B(_1972_));
 sg13g2_a21oi_1 _6858_ (.A1(_1990_),
    .A2(_1968_),
    .Y(_1998_),
    .B1(_1988_));
 sg13g2_o21ai_1 _6859_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_1997_),
    .A2(_1976_));
 sg13g2_nor2_1 _6860_ (.A(_1996_),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_inv_1 _6861_ (.Y(_2001_),
    .A(_2000_));
 sg13g2_nand2_1 _6862_ (.Y(_2002_),
    .A(_1999_),
    .B(_1996_));
 sg13g2_nand2_1 _6863_ (.Y(_2003_),
    .A(_2001_),
    .B(_2002_));
 sg13g2_inv_1 _6864_ (.Y(_2004_),
    .A(_2003_));
 sg13g2_buf_1 _6865_ (.A(\vgademo.scanline_audio_sample[5] ),
    .X(_2005_));
 sg13g2_nor2_1 _6866_ (.A(_2005_),
    .B(_0860_),
    .Y(_2006_));
 sg13g2_a21oi_1 _6867_ (.A1(_2004_),
    .A2(net67),
    .Y(_0266_),
    .B1(_2006_));
 sg13g2_nor2_1 _6868_ (.A(\vgademo.scanline_audio_sample[6] ),
    .B(_0860_),
    .Y(_2007_));
 sg13g2_a21oi_1 _6869_ (.A1(_2000_),
    .A2(net67),
    .Y(_0267_),
    .B1(_2007_));
 sg13g2_buf_1 _6870_ (.A(\vgademo.audio_beat_out[0] ),
    .X(_2008_));
 sg13g2_inv_1 _6871_ (.Y(_2009_),
    .A(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_inv_1 _6872_ (.Y(_2010_),
    .A(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_inv_1 _6873_ (.Y(_2011_),
    .A(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_inv_1 _6874_ (.Y(_2012_),
    .A(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_inv_1 _6875_ (.Y(_2013_),
    .A(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_inv_1 _6876_ (.Y(_2014_),
    .A(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_inv_1 _6877_ (.Y(_2015_),
    .A(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_inv_1 _6878_ (.Y(_2016_),
    .A(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_inv_1 _6879_ (.Y(_2017_),
    .A(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_nand2_1 _6880_ (.Y(_2018_),
    .A(\vgademo.soundtrack.sample_div[1] ),
    .B(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_nor3_2 _6881_ (.A(_2016_),
    .B(_2017_),
    .C(_2018_),
    .Y(_2019_));
 sg13g2_nand2_1 _6882_ (.Y(_2020_),
    .A(_2019_),
    .B(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_nor2b_1 _6883_ (.A(_2020_),
    .B_N(\vgademo.soundtrack.sample_div[5] ),
    .Y(_2021_));
 sg13g2_nand2_1 _6884_ (.Y(_2022_),
    .A(_2021_),
    .B(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_nor2b_1 _6885_ (.A(_2022_),
    .B_N(\vgademo.soundtrack.sample_div[7] ),
    .Y(_2023_));
 sg13g2_nand2_1 _6886_ (.Y(_2024_),
    .A(_2023_),
    .B(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_nor2b_1 _6887_ (.A(_2024_),
    .B_N(\vgademo.soundtrack.sample_div[9] ),
    .Y(_2025_));
 sg13g2_inv_1 _6888_ (.Y(_2026_),
    .A(_2025_));
 sg13g2_nor2_1 _6889_ (.A(_2015_),
    .B(_2026_),
    .Y(_2027_));
 sg13g2_nand2_1 _6890_ (.Y(_2028_),
    .A(_2027_),
    .B(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_nor2_1 _6891_ (.A(_2014_),
    .B(_2028_),
    .Y(_2029_));
 sg13g2_inv_1 _6892_ (.Y(_2030_),
    .A(_2029_));
 sg13g2_nor2_1 _6893_ (.A(_2013_),
    .B(_2030_),
    .Y(_2031_));
 sg13g2_inv_1 _6894_ (.Y(_2032_),
    .A(_2031_));
 sg13g2_nor2_1 _6895_ (.A(_2012_),
    .B(_2032_),
    .Y(_2033_));
 sg13g2_inv_1 _6896_ (.Y(_2034_),
    .A(_2033_));
 sg13g2_nor2_1 _6897_ (.A(_2011_),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_inv_1 _6898_ (.Y(_2036_),
    .A(_2035_));
 sg13g2_nor2_1 _6899_ (.A(_2010_),
    .B(_2036_),
    .Y(_2037_));
 sg13g2_inv_1 _6900_ (.Y(_2038_),
    .A(_2037_));
 sg13g2_nor2_1 _6901_ (.A(_2009_),
    .B(_2038_),
    .Y(_2039_));
 sg13g2_buf_1 _6902_ (.A(\vgademo.audio_beat_out[3] ),
    .X(_2040_));
 sg13g2_buf_1 _6903_ (.A(\vgademo.audio_beat_out[2] ),
    .X(_2041_));
 sg13g2_nor2_1 _6904_ (.A(\vgademo.audio_beat_out[1] ),
    .B(_2008_),
    .Y(_2042_));
 sg13g2_inv_1 _6905_ (.Y(_2043_),
    .A(_2042_));
 sg13g2_nor4_2 _6906_ (.A(_2040_),
    .B(_2041_),
    .C(\vgademo.audio_beat_out[4] ),
    .Y(_2044_),
    .D(_2043_));
 sg13g2_buf_1 _6907_ (.A(_2044_),
    .X(_2045_));
 sg13g2_inv_1 _6908_ (.Y(_2046_),
    .A(_2039_));
 sg13g2_nor2_2 _6909_ (.A(_2045_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_nor2_1 _6910_ (.A(_2008_),
    .B(_2047_),
    .Y(_2048_));
 sg13g2_a21oi_1 _6911_ (.A1(_2008_),
    .A2(_2039_),
    .Y(_0268_),
    .B1(_2048_));
 sg13g2_buf_1 _6912_ (.A(_2025_),
    .X(_2049_));
 sg13g2_nand2_1 _6913_ (.Y(_2050_),
    .A(\vgademo.soundtrack.tick_div[5] ),
    .B(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_nand4_1 _6914_ (.B(\vgademo.soundtrack.tick_div[2] ),
    .C(\vgademo.soundtrack.tick_div[1] ),
    .A(\vgademo.soundtrack.tick_div[3] ),
    .Y(_2051_),
    .D(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_nor4_1 _6915_ (.A(_2009_),
    .B(_2010_),
    .C(_2050_),
    .D(_2051_),
    .Y(_2052_));
 sg13g2_nand2_2 _6916_ (.Y(_2053_),
    .A(net58),
    .B(_2052_));
 sg13g2_nand2_1 _6917_ (.Y(_2054_),
    .A(\vgademo.audio_beat_out[1] ),
    .B(_2008_));
 sg13g2_a22oi_1 _6918_ (.Y(_2055_),
    .B1(_0769_),
    .B2(net76),
    .A2(_2054_),
    .A1(_2043_));
 sg13g2_nand2_1 _6919_ (.Y(_2056_),
    .A(_2053_),
    .B(\vgademo.audio_beat_out[1] ));
 sg13g2_o21ai_1 _6920_ (.B1(_2056_),
    .Y(_0269_),
    .A1(_2053_),
    .A2(_2055_));
 sg13g2_xnor2_1 _6921_ (.Y(_2057_),
    .A(_0080_),
    .B(_2054_));
 sg13g2_inv_1 _6922_ (.Y(_2058_),
    .A(_2047_));
 sg13g2_nand2_1 _6923_ (.Y(_2059_),
    .A(_2053_),
    .B(_2041_));
 sg13g2_o21ai_1 _6924_ (.B1(_2059_),
    .Y(_0270_),
    .A1(_2057_),
    .A2(_2058_));
 sg13g2_inv_1 _6925_ (.Y(_2060_),
    .A(_2044_));
 sg13g2_inv_1 _6926_ (.Y(_2061_),
    .A(_2028_));
 sg13g2_nor3_1 _6927_ (.A(_2013_),
    .B(_2014_),
    .C(_2050_),
    .Y(_2062_));
 sg13g2_nand4_1 _6928_ (.B(\vgademo.soundtrack.tick_div[7] ),
    .C(\vgademo.soundtrack.tick_div[6] ),
    .A(_2061_),
    .Y(_2063_),
    .D(_2062_));
 sg13g2_nor2_1 _6929_ (.A(net75),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_buf_1 _6930_ (.A(_2064_),
    .X(_2065_));
 sg13g2_inv_1 _6931_ (.Y(_2066_),
    .A(_2065_));
 sg13g2_inv_1 _6932_ (.Y(_2067_),
    .A(_2063_));
 sg13g2_inv_1 _6933_ (.Y(_2068_),
    .A(_2041_));
 sg13g2_nor2_1 _6934_ (.A(_2068_),
    .B(_2054_),
    .Y(_2069_));
 sg13g2_nand2_1 _6935_ (.Y(_2070_),
    .A(_2067_),
    .B(_2069_));
 sg13g2_nand2_1 _6936_ (.Y(_2071_),
    .A(_2066_),
    .B(_2070_));
 sg13g2_nor2_1 _6937_ (.A(_2040_),
    .B(_2071_),
    .Y(_2072_));
 sg13g2_inv_1 _6938_ (.Y(_2073_),
    .A(_2070_));
 sg13g2_nor3_1 _6939_ (.A(net116),
    .B(net75),
    .C(_2046_),
    .Y(_2074_));
 sg13g2_a21oi_1 _6940_ (.A1(_2040_),
    .A2(_2073_),
    .Y(_2075_),
    .B1(_2074_));
 sg13g2_nor2b_1 _6941_ (.A(_2072_),
    .B_N(_2075_),
    .Y(_0271_));
 sg13g2_inv_1 _6942_ (.Y(_2076_),
    .A(_2040_));
 sg13g2_o21ai_1 _6943_ (.B1(\vgademo.audio_beat_out[4] ),
    .Y(_2077_),
    .A1(_2076_),
    .A2(_2070_));
 sg13g2_o21ai_1 _6944_ (.B1(_2077_),
    .Y(_0272_),
    .A1(\vgademo.audio_beat_out[4] ),
    .A2(_2075_));
 sg13g2_inv_1 _6945_ (.Y(_2078_),
    .A(\vgademo.audio_kick_frames[0] ));
 sg13g2_nor3_1 _6946_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(_0928_),
    .C(_0919_),
    .Y(_2079_));
 sg13g2_buf_2 _6947_ (.A(_2079_),
    .X(_2080_));
 sg13g2_inv_1 _6948_ (.Y(_2081_),
    .A(_2080_));
 sg13g2_nor2_1 _6949_ (.A(_2081_),
    .B(_2044_),
    .Y(_2082_));
 sg13g2_nand2_1 _6950_ (.Y(_2083_),
    .A(_1669_),
    .B(_1664_));
 sg13g2_inv_1 _6951_ (.Y(_2084_),
    .A(_1669_));
 sg13g2_nand2_1 _6952_ (.Y(_2085_),
    .A(_2084_),
    .B(_1690_));
 sg13g2_buf_2 _6953_ (.A(_2085_),
    .X(_2086_));
 sg13g2_buf_1 _6954_ (.A(_1702_),
    .X(_2087_));
 sg13g2_nand2_1 _6955_ (.Y(_2088_),
    .A(_2086_),
    .B(_2087_));
 sg13g2_nand2_1 _6956_ (.Y(_2089_),
    .A(_0768_),
    .B(net88));
 sg13g2_nor2_1 _6957_ (.A(_1692_),
    .B(_2089_),
    .Y(_2090_));
 sg13g2_inv_1 _6958_ (.Y(_2091_),
    .A(_2090_));
 sg13g2_nand2_1 _6959_ (.Y(_2092_),
    .A(_2088_),
    .B(_2091_));
 sg13g2_inv_1 _6960_ (.Y(_2093_),
    .A(_2092_));
 sg13g2_nand2_1 _6961_ (.Y(_2094_),
    .A(_2093_),
    .B(_1677_));
 sg13g2_o21ai_1 _6962_ (.B1(_2094_),
    .Y(_2095_),
    .A1(_2083_),
    .A2(_2093_));
 sg13g2_nor2_1 _6963_ (.A(_0763_),
    .B(_2090_),
    .Y(_2096_));
 sg13g2_nor2_1 _6964_ (.A(_1678_),
    .B(_2086_),
    .Y(_2097_));
 sg13g2_nor2_2 _6965_ (.A(_2096_),
    .B(_2097_),
    .Y(_2098_));
 sg13g2_inv_1 _6966_ (.Y(_2099_),
    .A(_2098_));
 sg13g2_nor2_1 _6967_ (.A(net84),
    .B(_1678_),
    .Y(_2100_));
 sg13g2_inv_1 _6968_ (.Y(_2101_),
    .A(_2100_));
 sg13g2_nor2_1 _6969_ (.A(_2086_),
    .B(_2101_),
    .Y(_2102_));
 sg13g2_buf_1 _6970_ (.A(net89),
    .X(_2103_));
 sg13g2_nor2_1 _6971_ (.A(_2103_),
    .B(_2097_),
    .Y(_2104_));
 sg13g2_nor2_1 _6972_ (.A(_2102_),
    .B(_2104_),
    .Y(_2105_));
 sg13g2_nor2_1 _6973_ (.A(_2099_),
    .B(_2105_),
    .Y(_2106_));
 sg13g2_inv_1 _6974_ (.Y(_2107_),
    .A(_2105_));
 sg13g2_nor2_1 _6975_ (.A(_2099_),
    .B(_2107_),
    .Y(_2108_));
 sg13g2_nand2_1 _6976_ (.Y(_2109_),
    .A(_1671_),
    .B(_0766_));
 sg13g2_inv_1 _6977_ (.Y(_2110_),
    .A(net118));
 sg13g2_xnor2_1 _6978_ (.Y(_2111_),
    .A(_2110_),
    .B(_2102_));
 sg13g2_buf_1 _6979_ (.A(_2111_),
    .X(_2112_));
 sg13g2_a21o_1 _6980_ (.A2(_2109_),
    .A1(_1669_),
    .B1(_2112_),
    .X(_2113_));
 sg13g2_a22oi_1 _6981_ (.Y(_2114_),
    .B1(_2108_),
    .B2(_2113_),
    .A2(_2106_),
    .A1(_2095_));
 sg13g2_nand2_1 _6982_ (.Y(_2115_),
    .A(_1669_),
    .B(net81));
 sg13g2_a21o_1 _6983_ (.A2(_2115_),
    .A1(_2114_),
    .B1(net75),
    .X(_2116_));
 sg13g2_inv_1 _6984_ (.Y(_2117_),
    .A(_2053_));
 sg13g2_nand2_1 _6985_ (.Y(_2118_),
    .A(_2116_),
    .B(_2117_));
 sg13g2_buf_2 _6986_ (.A(_2118_),
    .X(_2119_));
 sg13g2_nor2_1 _6987_ (.A(_2082_),
    .B(_2119_),
    .Y(_2120_));
 sg13g2_o21ai_1 _6988_ (.B1(_2120_),
    .Y(_2121_),
    .A1(_2078_),
    .A2(net76));
 sg13g2_o21ai_1 _6989_ (.B1(_2121_),
    .Y(_0273_),
    .A1(_2078_),
    .A2(_2120_));
 sg13g2_inv_1 _6990_ (.Y(_2122_),
    .A(_2120_));
 sg13g2_nor2_1 _6991_ (.A(net76),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_inv_1 _6992_ (.Y(_2124_),
    .A(\vgademo.audio_kick_frames[1] ));
 sg13g2_nor2_1 _6993_ (.A(\vgademo.audio_kick_frames[0] ),
    .B(_2124_),
    .Y(_2125_));
 sg13g2_a22oi_1 _6994_ (.Y(_0274_),
    .B1(_2124_),
    .B2(_2121_),
    .A2(_2125_),
    .A1(_2123_));
 sg13g2_inv_1 _6995_ (.Y(_2126_),
    .A(_0928_));
 sg13g2_nor2_1 _6996_ (.A(\vgademo.audio_kick_frames[1] ),
    .B(\vgademo.audio_kick_frames[0] ),
    .Y(_2127_));
 sg13g2_xnor2_1 _6997_ (.Y(_2128_),
    .A(_0928_),
    .B(_2127_));
 sg13g2_a22oi_1 _6998_ (.Y(_0275_),
    .B1(_2128_),
    .B2(_2123_),
    .A2(_2122_),
    .A1(_2126_));
 sg13g2_buf_1 _6999_ (.A(net58),
    .X(_2129_));
 sg13g2_buf_1 _7000_ (.A(net58),
    .X(_2130_));
 sg13g2_nor2_1 _7001_ (.A(_0087_),
    .B(net48),
    .Y(_2131_));
 sg13g2_a21oi_1 _7002_ (.A1(\vgademo.soundtrack.noise_lfsr[1] ),
    .A2(net49),
    .Y(_0276_),
    .B1(_2131_));
 sg13g2_nor2_1 _7003_ (.A(_0088_),
    .B(net48),
    .Y(_2132_));
 sg13g2_a21oi_1 _7004_ (.A1(\vgademo.soundtrack.noise_lfsr[11] ),
    .A2(net49),
    .Y(_0277_),
    .B1(_2132_));
 sg13g2_nor2_1 _7005_ (.A(_0089_),
    .B(net48),
    .Y(_2133_));
 sg13g2_a21oi_1 _7006_ (.A1(_1640_),
    .A2(net49),
    .Y(_0278_),
    .B1(_2133_));
 sg13g2_mux2_1 _7007_ (.A0(_0090_),
    .A1(_0085_),
    .S(net48),
    .X(_0279_));
 sg13g2_xnor2_1 _7008_ (.Y(_2134_),
    .A(\vgademo.soundtrack.noise_lfsr[0] ),
    .B(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_nor2_1 _7009_ (.A(\vgademo.soundtrack.noise_lfsr[13] ),
    .B(net58),
    .Y(_2135_));
 sg13g2_a21oi_1 _7010_ (.A1(net49),
    .A2(_2134_),
    .Y(_0280_),
    .B1(_2135_));
 sg13g2_mux2_1 _7011_ (.A0(\vgademo.soundtrack.noise_lfsr[14] ),
    .A1(\vgademo.soundtrack.noise_lfsr[0] ),
    .S(net48),
    .X(_0281_));
 sg13g2_nor2_1 _7012_ (.A(_0091_),
    .B(_2049_),
    .Y(_2136_));
 sg13g2_a21oi_1 _7013_ (.A1(\vgademo.soundtrack.noise_lfsr[2] ),
    .A2(net49),
    .Y(_0282_),
    .B1(_2136_));
 sg13g2_nor2_1 _7014_ (.A(_0092_),
    .B(_2049_),
    .Y(_2137_));
 sg13g2_a21oi_1 _7015_ (.A1(\vgademo.soundtrack.noise_lfsr[3] ),
    .A2(net49),
    .Y(_0283_),
    .B1(_2137_));
 sg13g2_mux2_1 _7016_ (.A0(_0093_),
    .A1(_0063_),
    .S(net48),
    .X(_0284_));
 sg13g2_nor2_1 _7017_ (.A(\vgademo.soundtrack.noise_lfsr[4] ),
    .B(net58),
    .Y(_2138_));
 sg13g2_a21oi_1 _7018_ (.A1(_1796_),
    .A2(_2129_),
    .Y(_0285_),
    .B1(_2138_));
 sg13g2_mux2_1 _7019_ (.A0(_0094_),
    .A1(_0084_),
    .S(_2130_),
    .X(_0286_));
 sg13g2_nor2_1 _7020_ (.A(\vgademo.soundtrack.noise_lfsr[6] ),
    .B(net58),
    .Y(_2139_));
 sg13g2_a21oi_1 _7021_ (.A1(_1753_),
    .A2(_2129_),
    .Y(_0287_),
    .B1(_2139_));
 sg13g2_mux2_1 _7022_ (.A0(_0095_),
    .A1(_0083_),
    .S(_2130_),
    .X(_0288_));
 sg13g2_nor2_1 _7023_ (.A(\vgademo.soundtrack.noise_lfsr[8] ),
    .B(net58),
    .Y(_2140_));
 sg13g2_a21oi_1 _7024_ (.A1(_1644_),
    .A2(net49),
    .Y(_0289_),
    .B1(_2140_));
 sg13g2_nor2_1 _7025_ (.A(\vgademo.soundtrack.noise_lfsr[9] ),
    .B(net58),
    .Y(_2141_));
 sg13g2_a21oi_1 _7026_ (.A1(_1731_),
    .A2(net49),
    .Y(_0290_),
    .B1(_2141_));
 sg13g2_buf_1 _7027_ (.A(net81),
    .X(_2142_));
 sg13g2_nor2_2 _7028_ (.A(net117),
    .B(_1661_),
    .Y(_2143_));
 sg13g2_inv_1 _7029_ (.Y(_2144_),
    .A(_1699_));
 sg13g2_nor2_1 _7030_ (.A(_2143_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_o21ai_1 _7031_ (.B1(_2145_),
    .Y(_2146_),
    .A1(net77),
    .A2(_2092_));
 sg13g2_nor2_1 _7032_ (.A(_2144_),
    .B(_2092_),
    .Y(_2147_));
 sg13g2_nand2_1 _7033_ (.Y(_2148_),
    .A(_2147_),
    .B(_1680_));
 sg13g2_nand3_1 _7034_ (.B(_2112_),
    .C(_2148_),
    .A(_2146_),
    .Y(_2149_));
 sg13g2_a21oi_1 _7035_ (.A1(_1699_),
    .A2(_1665_),
    .Y(_2150_),
    .B1(_1691_));
 sg13g2_nand3b_1 _7036_ (.B(_2098_),
    .C(_2150_),
    .Y(_2151_),
    .A_N(_2112_));
 sg13g2_a21oi_1 _7037_ (.A1(_2149_),
    .A2(_2151_),
    .Y(_2152_),
    .B1(_2107_));
 sg13g2_inv_1 _7038_ (.Y(_2153_),
    .A(_2145_));
 sg13g2_inv_1 _7039_ (.Y(_2154_),
    .A(_1703_));
 sg13g2_nor2_1 _7040_ (.A(net79),
    .B(_2154_),
    .Y(_2155_));
 sg13g2_inv_1 _7041_ (.Y(_2156_),
    .A(_2155_));
 sg13g2_nand2_1 _7042_ (.Y(_2157_),
    .A(_2156_),
    .B(_1699_));
 sg13g2_a22oi_1 _7043_ (.Y(_2158_),
    .B1(_2157_),
    .B2(_2106_),
    .A2(_2153_),
    .A1(_2099_));
 sg13g2_nand2_1 _7044_ (.Y(_2159_),
    .A(_2158_),
    .B(_2045_));
 sg13g2_a21oi_1 _7045_ (.A1(net75),
    .A2(_2054_),
    .Y(_2160_),
    .B1(_2063_));
 sg13g2_o21ai_1 _7046_ (.B1(_2160_),
    .Y(_2161_),
    .A1(_2152_),
    .A2(_2159_));
 sg13g2_buf_2 _7047_ (.A(_2161_),
    .X(_2162_));
 sg13g2_nand2_1 _7048_ (.Y(_2163_),
    .A(_1729_),
    .B(net86));
 sg13g2_nor2_1 _7049_ (.A(net80),
    .B(_2163_),
    .Y(_2164_));
 sg13g2_nand2_1 _7050_ (.Y(_2165_),
    .A(_2164_),
    .B(net91));
 sg13g2_a21oi_1 _7051_ (.A1(_1730_),
    .A2(_2165_),
    .Y(_2166_),
    .B1(net76));
 sg13g2_nand2_1 _7052_ (.Y(_2167_),
    .A(_2162_),
    .B(_0096_));
 sg13g2_o21ai_1 _7053_ (.B1(_2167_),
    .Y(_0291_),
    .A1(_2162_),
    .A2(_2166_));
 sg13g2_nand2b_1 _7054_ (.Y(_2168_),
    .B(_2163_),
    .A_N(_1741_));
 sg13g2_a21oi_1 _7055_ (.A1(_2165_),
    .A2(_2168_),
    .Y(_2169_),
    .B1(net76));
 sg13g2_nand2_1 _7056_ (.Y(_2170_),
    .A(_2162_),
    .B(_0097_));
 sg13g2_o21ai_1 _7057_ (.B1(_2170_),
    .Y(_0292_),
    .A1(_2162_),
    .A2(_2169_));
 sg13g2_nand2_1 _7058_ (.Y(_2171_),
    .A(_2164_),
    .B(_1802_));
 sg13g2_nand2_1 _7059_ (.Y(_2172_),
    .A(_2163_),
    .B(net80));
 sg13g2_nand3_1 _7060_ (.B(_2171_),
    .C(_2172_),
    .A(net75),
    .Y(_2173_));
 sg13g2_mux2_1 _7061_ (.A0(_2173_),
    .A1(_0098_),
    .S(_2162_),
    .X(_0293_));
 sg13g2_o21ai_1 _7062_ (.B1(net75),
    .Y(_2174_),
    .A1(net91),
    .A2(_2164_));
 sg13g2_mux2_1 _7063_ (.A0(_2174_),
    .A1(_0099_),
    .S(_2162_),
    .X(_0294_));
 sg13g2_inv_1 _7064_ (.Y(_2175_),
    .A(audio));
 sg13g2_inv_1 _7065_ (.Y(_2176_),
    .A(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_nor2_1 _7066_ (.A(_2176_),
    .B(_2000_),
    .Y(_2177_));
 sg13g2_nor2_1 _7067_ (.A(_0533_),
    .B(_2177_),
    .Y(_2178_));
 sg13g2_inv_1 _7068_ (.Y(_2179_),
    .A(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_nor2_1 _7069_ (.A(_2179_),
    .B(_2004_),
    .Y(_2180_));
 sg13g2_inv_1 _7070_ (.Y(_2181_),
    .A(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_nor2_1 _7071_ (.A(_2181_),
    .B(_1978_),
    .Y(_2182_));
 sg13g2_inv_1 _7072_ (.Y(_2183_),
    .A(_2182_));
 sg13g2_nand2_1 _7073_ (.Y(_2184_),
    .A(_1995_),
    .B(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_nor2_1 _7074_ (.A(\vgademo.soundtrack.sigma_delta_accum[13] ),
    .B(_1995_),
    .Y(_2185_));
 sg13g2_a21oi_1 _7075_ (.A1(_2183_),
    .A2(_2184_),
    .Y(_2186_),
    .B1(_2185_));
 sg13g2_nand2b_1 _7076_ (.Y(_2187_),
    .B(_2184_),
    .A_N(_2185_));
 sg13g2_inv_1 _7077_ (.Y(_2188_),
    .A(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_xnor2_1 _7078_ (.Y(_2189_),
    .A(_1937_),
    .B(_1918_));
 sg13g2_xnor2_1 _7079_ (.Y(_2190_),
    .A(_2188_),
    .B(_2189_));
 sg13g2_inv_1 _7080_ (.Y(_2191_),
    .A(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_xnor2_1 _7081_ (.Y(_2192_),
    .A(_1913_),
    .B(_1912_));
 sg13g2_nor2_1 _7082_ (.A(_2191_),
    .B(_2192_),
    .Y(_2193_));
 sg13g2_inv_1 _7083_ (.Y(_2194_),
    .A(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_xnor2_1 _7084_ (.Y(_2195_),
    .A(_1910_),
    .B(_1908_));
 sg13g2_nor2_1 _7085_ (.A(_2194_),
    .B(_2195_),
    .Y(_2196_));
 sg13g2_xnor2_1 _7086_ (.Y(_2197_),
    .A(_2194_),
    .B(_2195_));
 sg13g2_inv_1 _7087_ (.Y(_2198_),
    .A(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_xnor2_1 _7088_ (.Y(_2199_),
    .A(_1903_),
    .B(_1902_));
 sg13g2_xnor2_1 _7089_ (.Y(_2200_),
    .A(\vgademo.soundtrack.sigma_delta_accum[3] ),
    .B(_2199_));
 sg13g2_xor2_1 _7090_ (.B(_1883_),
    .A(_1899_),
    .X(_2201_));
 sg13g2_inv_1 _7091_ (.Y(_2202_),
    .A(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_nand2_1 _7092_ (.Y(_2203_),
    .A(_2201_),
    .B(_2202_));
 sg13g2_xnor2_1 _7093_ (.Y(_2204_),
    .A(_1886_),
    .B(_1897_));
 sg13g2_nor2b_1 _7094_ (.A(_2204_),
    .B_N(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .Y(_2205_));
 sg13g2_nor2_1 _7095_ (.A(_2202_),
    .B(_2201_),
    .Y(_2206_));
 sg13g2_a21oi_1 _7096_ (.A1(_2203_),
    .A2(_2205_),
    .Y(_2207_),
    .B1(_2206_));
 sg13g2_xnor2_1 _7097_ (.Y(_2208_),
    .A(_1900_),
    .B(_1882_));
 sg13g2_xor2_1 _7098_ (.B(_2208_),
    .A(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .X(_2209_));
 sg13g2_nand2b_1 _7099_ (.Y(_2210_),
    .B(\vgademo.soundtrack.sigma_delta_accum[2] ),
    .A_N(_2208_));
 sg13g2_o21ai_1 _7100_ (.B1(_2210_),
    .Y(_2211_),
    .A1(_2207_),
    .A2(_2209_));
 sg13g2_nand2_1 _7101_ (.Y(_2212_),
    .A(_2200_),
    .B(_2211_));
 sg13g2_o21ai_1 _7102_ (.B1(_2212_),
    .Y(_2213_),
    .A1(_2198_),
    .A2(_2199_));
 sg13g2_xnor2_1 _7103_ (.Y(_2214_),
    .A(_1906_),
    .B(_1905_));
 sg13g2_inv_1 _7104_ (.Y(_2215_),
    .A(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_nand2_1 _7105_ (.Y(_2216_),
    .A(_2214_),
    .B(_2215_));
 sg13g2_nor2_1 _7106_ (.A(_2215_),
    .B(_2214_),
    .Y(_2217_));
 sg13g2_a21o_1 _7107_ (.A2(_2216_),
    .A1(_2213_),
    .B1(_2217_),
    .X(_2218_));
 sg13g2_nand2b_1 _7108_ (.Y(_2219_),
    .B(_2218_),
    .A_N(_2197_));
 sg13g2_nand2b_1 _7109_ (.Y(_2220_),
    .B(_2219_),
    .A_N(_2196_));
 sg13g2_nor2_1 _7110_ (.A(_2193_),
    .B(_2220_),
    .Y(_2221_));
 sg13g2_nand2_1 _7111_ (.Y(_2222_),
    .A(_2192_),
    .B(_2191_));
 sg13g2_nor2b_1 _7112_ (.A(_2221_),
    .B_N(_2222_),
    .Y(_2223_));
 sg13g2_xnor2_1 _7113_ (.Y(_2224_),
    .A(_1916_),
    .B(_1915_));
 sg13g2_inv_1 _7114_ (.Y(_2225_),
    .A(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_nand2_1 _7115_ (.Y(_2226_),
    .A(_2224_),
    .B(_2225_));
 sg13g2_nor2_1 _7116_ (.A(_2225_),
    .B(_2224_),
    .Y(_2227_));
 sg13g2_a21oi_1 _7117_ (.A1(_2223_),
    .A2(_2226_),
    .Y(_2228_),
    .B1(_2227_));
 sg13g2_nor2_1 _7118_ (.A(_2188_),
    .B(_2189_),
    .Y(_2229_));
 sg13g2_inv_1 _7119_ (.Y(_2230_),
    .A(_2229_));
 sg13g2_o21ai_1 _7120_ (.B1(_2230_),
    .Y(_2231_),
    .A1(_2190_),
    .A2(_2228_));
 sg13g2_inv_1 _7121_ (.Y(_2232_),
    .A(_2231_));
 sg13g2_nand2_1 _7122_ (.Y(_2233_),
    .A(_1922_),
    .B(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_nor2_1 _7123_ (.A(\vgademo.soundtrack.sigma_delta_accum[9] ),
    .B(_1922_),
    .Y(_2234_));
 sg13g2_a21oi_1 _7124_ (.A1(_2232_),
    .A2(_2233_),
    .Y(_2235_),
    .B1(_2234_));
 sg13g2_nor2_1 _7125_ (.A(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .B(_1942_),
    .Y(_2236_));
 sg13g2_nor2b_1 _7126_ (.A(_1943_),
    .B_N(\vgademo.soundtrack.sigma_delta_accum[10] ),
    .Y(_2237_));
 sg13g2_nor2_1 _7127_ (.A(_2236_),
    .B(_2237_),
    .Y(_2238_));
 sg13g2_nand2_1 _7128_ (.Y(_2239_),
    .A(_2235_),
    .B(_2238_));
 sg13g2_nand2_1 _7129_ (.Y(_2240_),
    .A(_1958_),
    .B(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_inv_1 _7130_ (.Y(_2241_),
    .A(_2240_));
 sg13g2_nor2_1 _7131_ (.A(_2237_),
    .B(_2241_),
    .Y(_2242_));
 sg13g2_nor2_1 _7132_ (.A(\vgademo.soundtrack.sigma_delta_accum[11] ),
    .B(_1958_),
    .Y(_2243_));
 sg13g2_a21oi_1 _7133_ (.A1(_2239_),
    .A2(_2242_),
    .Y(_2244_),
    .B1(_2243_));
 sg13g2_nor2_1 _7134_ (.A(\vgademo.soundtrack.sigma_delta_accum[12] ),
    .B(_1977_),
    .Y(_2245_));
 sg13g2_nor2_1 _7135_ (.A(_2245_),
    .B(_2182_),
    .Y(_2246_));
 sg13g2_nand2_1 _7136_ (.Y(_2247_),
    .A(_2244_),
    .B(_2246_));
 sg13g2_nor2_1 _7137_ (.A(_2187_),
    .B(_2247_),
    .Y(_2248_));
 sg13g2_nor2_1 _7138_ (.A(_2186_),
    .B(_2248_),
    .Y(_2249_));
 sg13g2_nand2b_1 _7139_ (.Y(_2250_),
    .B(_2249_),
    .A_N(_2180_));
 sg13g2_nand2_1 _7140_ (.Y(_2251_),
    .A(_2000_),
    .B(_2176_));
 sg13g2_nor2_1 _7141_ (.A(\vgademo.soundtrack.sigma_delta_accum[14] ),
    .B(_2003_),
    .Y(_2252_));
 sg13g2_inv_1 _7142_ (.Y(_2253_),
    .A(_2252_));
 sg13g2_nand3_1 _7143_ (.B(_2251_),
    .C(_2253_),
    .A(_2250_),
    .Y(_2254_));
 sg13g2_a22oi_1 _7144_ (.Y(_0295_),
    .B1(_2178_),
    .B2(_2254_),
    .A2(_2175_),
    .A1(_0533_));
 sg13g2_nor2_1 _7145_ (.A(_0774_),
    .B(_1704_),
    .Y(_2255_));
 sg13g2_o21ai_1 _7146_ (.B1(net84),
    .Y(_2256_),
    .A1(net81),
    .A2(_2255_));
 sg13g2_inv_1 _7147_ (.Y(_2257_),
    .A(_2096_));
 sg13g2_nand2_1 _7148_ (.Y(_2258_),
    .A(_2256_),
    .B(_2257_));
 sg13g2_nor2_1 _7149_ (.A(_0778_),
    .B(_2110_),
    .Y(_2259_));
 sg13g2_a221oi_1 _7150_ (.B2(_2259_),
    .C1(_2041_),
    .B1(_2258_),
    .A1(_2142_),
    .Y(_2260_),
    .A2(_2110_));
 sg13g2_inv_1 _7151_ (.Y(_2261_),
    .A(_1676_));
 sg13g2_nor2_1 _7152_ (.A(net79),
    .B(_1686_),
    .Y(_2262_));
 sg13g2_nor2_1 _7153_ (.A(_0769_),
    .B(_2143_),
    .Y(_2263_));
 sg13g2_inv_1 _7154_ (.Y(_2264_),
    .A(_1670_));
 sg13g2_a22oi_1 _7155_ (.Y(_2265_),
    .B1(_0774_),
    .B2(_2264_),
    .A2(_2263_),
    .A1(_2262_));
 sg13g2_a21oi_1 _7156_ (.A1(_2265_),
    .A2(net81),
    .Y(_2266_),
    .B1(net84));
 sg13g2_o21ai_1 _7157_ (.B1(_2266_),
    .Y(_2267_),
    .A1(_1680_),
    .A2(_2261_));
 sg13g2_nand2_1 _7158_ (.Y(_2268_),
    .A(_2089_),
    .B(net79));
 sg13g2_o21ai_1 _7159_ (.B1(_1705_),
    .Y(_2269_),
    .A1(_1686_),
    .A2(_2268_));
 sg13g2_nor2_2 _7160_ (.A(net89),
    .B(net81),
    .Y(_2270_));
 sg13g2_a21oi_1 _7161_ (.A1(_2269_),
    .A2(_2270_),
    .Y(_2271_),
    .B1(_1711_));
 sg13g2_nand2_1 _7162_ (.Y(_2272_),
    .A(_2267_),
    .B(_2271_));
 sg13g2_a21oi_1 _7163_ (.A1(_1680_),
    .A2(_1676_),
    .Y(_2273_),
    .B1(_0777_));
 sg13g2_inv_1 _7164_ (.Y(_2274_),
    .A(_2273_));
 sg13g2_nor2_1 _7165_ (.A(_1690_),
    .B(_1669_),
    .Y(_2275_));
 sg13g2_nor2_1 _7166_ (.A(_1661_),
    .B(_1670_),
    .Y(_2276_));
 sg13g2_inv_1 _7167_ (.Y(_2277_),
    .A(_2276_));
 sg13g2_nor2_1 _7168_ (.A(_1702_),
    .B(_2143_),
    .Y(_2278_));
 sg13g2_a21oi_1 _7169_ (.A1(_2277_),
    .A2(_2087_),
    .Y(_2279_),
    .B1(_2278_));
 sg13g2_nor3_1 _7170_ (.A(net98),
    .B(_2275_),
    .C(_2279_),
    .Y(_2280_));
 sg13g2_inv_1 _7171_ (.Y(_2281_),
    .A(_1711_));
 sg13g2_o21ai_1 _7172_ (.B1(_2281_),
    .Y(_2282_),
    .A1(_2274_),
    .A2(_2280_));
 sg13g2_nand3_1 _7173_ (.B(net118),
    .C(_2270_),
    .A(_2255_),
    .Y(_2283_));
 sg13g2_nand3_1 _7174_ (.B(_1711_),
    .C(_2101_),
    .A(_2283_),
    .Y(_2284_));
 sg13g2_nand2_1 _7175_ (.Y(_2285_),
    .A(_2282_),
    .B(_2284_));
 sg13g2_inv_1 _7176_ (.Y(_2286_),
    .A(_2285_));
 sg13g2_a22oi_1 _7177_ (.Y(_2287_),
    .B1(_2041_),
    .B2(_2286_),
    .A2(_2272_),
    .A1(_2260_));
 sg13g2_o21ai_1 _7178_ (.B1(_0764_),
    .Y(_2288_),
    .A1(_1671_),
    .A2(_1694_));
 sg13g2_nand2_1 _7179_ (.Y(_2289_),
    .A(_2288_),
    .B(_2257_));
 sg13g2_nand2_1 _7180_ (.Y(_2290_),
    .A(_2289_),
    .B(net89));
 sg13g2_inv_1 _7181_ (.Y(_2291_),
    .A(_2259_));
 sg13g2_nor3_1 _7182_ (.A(_1701_),
    .B(_0774_),
    .C(_1666_),
    .Y(_2292_));
 sg13g2_nor2_1 _7183_ (.A(net89),
    .B(_2292_),
    .Y(_2293_));
 sg13g2_nor2_1 _7184_ (.A(_2291_),
    .B(_2293_),
    .Y(_2294_));
 sg13g2_nor2_1 _7185_ (.A(_1671_),
    .B(_1693_),
    .Y(_2295_));
 sg13g2_nand2_1 _7186_ (.Y(_2296_),
    .A(_1669_),
    .B(_1661_));
 sg13g2_a21oi_1 _7187_ (.A1(_2295_),
    .A2(_2296_),
    .Y(_2297_),
    .B1(_1701_));
 sg13g2_nand2b_1 _7188_ (.Y(_2298_),
    .B(_1683_),
    .A_N(_2297_));
 sg13g2_nand2_1 _7189_ (.Y(_2299_),
    .A(_2262_),
    .B(_2086_));
 sg13g2_nand3_1 _7190_ (.B(_1672_),
    .C(_0764_),
    .A(_2299_),
    .Y(_2300_));
 sg13g2_nand3_1 _7191_ (.B(net84),
    .C(_2257_),
    .A(_2300_),
    .Y(_2301_));
 sg13g2_o21ai_1 _7192_ (.B1(_2301_),
    .Y(_2302_),
    .A1(_2298_),
    .A2(_2280_));
 sg13g2_a22oi_1 _7193_ (.Y(_2303_),
    .B1(_2281_),
    .B2(_2302_),
    .A2(_2294_),
    .A1(_2290_));
 sg13g2_nand3_1 _7194_ (.B(_1683_),
    .C(_1678_),
    .A(_2257_),
    .Y(_2304_));
 sg13g2_nor2_1 _7195_ (.A(_2143_),
    .B(_1686_),
    .Y(_2305_));
 sg13g2_nor3_1 _7196_ (.A(net98),
    .B(net79),
    .C(_2305_),
    .Y(_2306_));
 sg13g2_a21oi_1 _7197_ (.A1(_2306_),
    .A2(_0777_),
    .Y(_2307_),
    .B1(_2291_));
 sg13g2_nor2_1 _7198_ (.A(_2115_),
    .B(_1705_),
    .Y(_2308_));
 sg13g2_nor3_1 _7199_ (.A(net117),
    .B(net98),
    .C(_2268_),
    .Y(_2309_));
 sg13g2_o21ai_1 _7200_ (.B1(net84),
    .Y(_2310_),
    .A1(_2308_),
    .A2(_2309_));
 sg13g2_inv_1 _7201_ (.Y(_2311_),
    .A(_2270_));
 sg13g2_a21o_1 _7202_ (.A2(_1705_),
    .A1(_2088_),
    .B1(_2311_),
    .X(_2312_));
 sg13g2_nand3_1 _7203_ (.B(_2312_),
    .C(_2274_),
    .A(_2310_),
    .Y(_2313_));
 sg13g2_nand2_1 _7204_ (.Y(_2314_),
    .A(_2261_),
    .B(net89));
 sg13g2_a21oi_1 _7205_ (.A1(_2314_),
    .A2(_2311_),
    .Y(_2315_),
    .B1(net118));
 sg13g2_a221oi_1 _7206_ (.B2(_2281_),
    .C1(_2315_),
    .B1(_2313_),
    .A1(_2304_),
    .Y(_2316_),
    .A2(_2307_));
 sg13g2_mux2_1 _7207_ (.A0(_2303_),
    .A1(_2316_),
    .S(_2068_),
    .X(_2317_));
 sg13g2_buf_1 _7208_ (.A(_2317_),
    .X(_2318_));
 sg13g2_inv_1 _7209_ (.Y(_2319_),
    .A(_1688_));
 sg13g2_a221oi_1 _7210_ (.B2(_1676_),
    .C1(_2280_),
    .B1(_2319_),
    .A1(net98),
    .Y(_2320_),
    .A2(_2278_));
 sg13g2_nand3_1 _7211_ (.B(_2103_),
    .C(net118),
    .A(_2320_),
    .Y(_2321_));
 sg13g2_nor2_1 _7212_ (.A(net97),
    .B(_0769_),
    .Y(_2322_));
 sg13g2_nand3_1 _7213_ (.B(net81),
    .C(net118),
    .A(_2143_),
    .Y(_2323_));
 sg13g2_o21ai_1 _7214_ (.B1(net84),
    .Y(_2324_),
    .A1(_2322_),
    .A2(_2323_));
 sg13g2_nand3_1 _7215_ (.B(_0778_),
    .C(_2324_),
    .A(_2321_),
    .Y(_2325_));
 sg13g2_nand2_1 _7216_ (.Y(_2326_),
    .A(_2110_),
    .B(net89));
 sg13g2_nand3_1 _7217_ (.B(_2283_),
    .C(_2326_),
    .A(_2290_),
    .Y(_2327_));
 sg13g2_a21oi_1 _7218_ (.A1(_2327_),
    .A2(_0779_),
    .Y(_2328_),
    .B1(_2068_));
 sg13g2_nand2_1 _7219_ (.Y(_2329_),
    .A(_2325_),
    .B(_2328_));
 sg13g2_o21ai_1 _7220_ (.B1(_2310_),
    .Y(_2330_),
    .A1(net81),
    .A2(_2269_));
 sg13g2_a21oi_1 _7221_ (.A1(_2086_),
    .A2(_2100_),
    .Y(_2331_),
    .B1(_1711_));
 sg13g2_o21ai_1 _7222_ (.B1(_2331_),
    .Y(_2332_),
    .A1(_2266_),
    .A2(_2330_));
 sg13g2_nand2b_1 _7223_ (.Y(_2333_),
    .B(_1676_),
    .A_N(_2326_));
 sg13g2_o21ai_1 _7224_ (.B1(_2304_),
    .Y(_2334_),
    .A1(_2306_),
    .A2(_2256_));
 sg13g2_nand2_1 _7225_ (.Y(_2335_),
    .A(_2334_),
    .B(_2259_));
 sg13g2_nand3_1 _7226_ (.B(_2333_),
    .C(_2335_),
    .A(_2332_),
    .Y(_2336_));
 sg13g2_nand2_1 _7227_ (.Y(_2337_),
    .A(_2336_),
    .B(_2068_));
 sg13g2_nand2_1 _7228_ (.Y(_2338_),
    .A(_2329_),
    .B(_2337_));
 sg13g2_buf_2 _7229_ (.A(_2338_),
    .X(_2339_));
 sg13g2_a21o_1 _7230_ (.A2(_2318_),
    .A1(_2287_),
    .B1(_2339_),
    .X(_2340_));
 sg13g2_buf_1 _7231_ (.A(_2340_),
    .X(_2341_));
 sg13g2_inv_1 _7232_ (.Y(_2342_),
    .A(_2287_));
 sg13g2_nand2_1 _7233_ (.Y(_2343_),
    .A(_2318_),
    .B(_2342_));
 sg13g2_nand2_1 _7234_ (.Y(_2344_),
    .A(_2339_),
    .B(_2343_));
 sg13g2_nand2_1 _7235_ (.Y(_2345_),
    .A(_2341_),
    .B(_2344_));
 sg13g2_nor2_1 _7236_ (.A(_0533_),
    .B(_2026_),
    .Y(_2346_));
 sg13g2_buf_2 _7237_ (.A(_2346_),
    .X(_2347_));
 sg13g2_buf_1 _7238_ (.A(_2347_),
    .X(_2348_));
 sg13g2_nand2_1 _7239_ (.Y(_2349_),
    .A(_2345_),
    .B(net35));
 sg13g2_xnor2_1 _7240_ (.Y(_0296_),
    .A(\vgademo.soundtrack.pulse_osc_p[0] ),
    .B(_2349_));
 sg13g2_and2_1 _7241_ (.A(_2345_),
    .B(\vgademo.soundtrack.pulse_osc_p[0] ),
    .X(_2350_));
 sg13g2_inv_1 _7242_ (.Y(_2351_),
    .A(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_xnor2_1 _7243_ (.Y(_2352_),
    .A(_2351_),
    .B(_2341_));
 sg13g2_nand2_1 _7244_ (.Y(_2353_),
    .A(_2350_),
    .B(_2352_));
 sg13g2_nand2_1 _7245_ (.Y(_2354_),
    .A(_2341_),
    .B(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_nand2_1 _7246_ (.Y(_2355_),
    .A(_2353_),
    .B(_2354_));
 sg13g2_nand2b_1 _7247_ (.Y(_2356_),
    .B(_2342_),
    .A_N(_2318_));
 sg13g2_nand2_1 _7248_ (.Y(_2357_),
    .A(_2356_),
    .B(_2339_));
 sg13g2_inv_1 _7249_ (.Y(_2358_),
    .A(_2339_));
 sg13g2_nand2_1 _7250_ (.Y(_2359_),
    .A(_2358_),
    .B(_2343_));
 sg13g2_nand2_1 _7251_ (.Y(_2360_),
    .A(_2357_),
    .B(_2359_));
 sg13g2_inv_1 _7252_ (.Y(_2361_),
    .A(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_nand2_1 _7253_ (.Y(_2362_),
    .A(_2360_),
    .B(_2361_));
 sg13g2_nor2_1 _7254_ (.A(_2361_),
    .B(_2360_),
    .Y(_2363_));
 sg13g2_a21oi_1 _7255_ (.A1(_2355_),
    .A2(_2362_),
    .Y(_2364_),
    .B1(_2363_));
 sg13g2_inv_1 _7256_ (.Y(_2365_),
    .A(_2364_));
 sg13g2_nand2_1 _7257_ (.Y(_2366_),
    .A(_2341_),
    .B(_2356_));
 sg13g2_inv_1 _7258_ (.Y(_2367_),
    .A(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_nand2_1 _7259_ (.Y(_2368_),
    .A(_2366_),
    .B(_2367_));
 sg13g2_nand3_1 _7260_ (.B(\vgademo.soundtrack.pulse_osc_p[4] ),
    .C(_2356_),
    .A(_2341_),
    .Y(_2369_));
 sg13g2_nand2_1 _7261_ (.Y(_2370_),
    .A(_2368_),
    .B(_2369_));
 sg13g2_nor2_1 _7262_ (.A(_2342_),
    .B(_2318_),
    .Y(_2371_));
 sg13g2_nor2_1 _7263_ (.A(_2371_),
    .B(_2344_),
    .Y(_2372_));
 sg13g2_a21oi_1 _7264_ (.A1(_2358_),
    .A2(_2371_),
    .Y(_2373_),
    .B1(_2372_));
 sg13g2_nor2_1 _7265_ (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(_2373_),
    .Y(_2374_));
 sg13g2_nand2_1 _7266_ (.Y(_2375_),
    .A(_2373_),
    .B(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_nand2b_1 _7267_ (.Y(_2376_),
    .B(_2375_),
    .A_N(_2374_));
 sg13g2_nor2_1 _7268_ (.A(_2370_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_o21ai_1 _7269_ (.B1(_2369_),
    .Y(_2378_),
    .A1(_2375_),
    .A2(_2370_));
 sg13g2_a21oi_1 _7270_ (.A1(_2365_),
    .A2(_2377_),
    .Y(_2379_),
    .B1(_2378_));
 sg13g2_inv_1 _7271_ (.Y(_2380_),
    .A(_2379_));
 sg13g2_nand2b_1 _7272_ (.Y(_2381_),
    .B(_2359_),
    .A_N(_2371_));
 sg13g2_inv_1 _7273_ (.Y(_2382_),
    .A(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_nand2_1 _7274_ (.Y(_2383_),
    .A(_2381_),
    .B(_2382_));
 sg13g2_nor2_1 _7275_ (.A(_2382_),
    .B(_2381_),
    .Y(_2384_));
 sg13g2_a21oi_1 _7276_ (.A1(_2380_),
    .A2(_2383_),
    .Y(_2385_),
    .B1(_2384_));
 sg13g2_inv_1 _7277_ (.Y(_2386_),
    .A(_2385_));
 sg13g2_inv_1 _7278_ (.Y(_2387_),
    .A(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_nor2_1 _7279_ (.A(_2387_),
    .B(_2358_),
    .Y(_2388_));
 sg13g2_nor2_1 _7280_ (.A(\vgademo.soundtrack.pulse_osc_p[6] ),
    .B(_2339_),
    .Y(_2389_));
 sg13g2_inv_1 _7281_ (.Y(_2390_),
    .A(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_xnor2_1 _7282_ (.Y(_2391_),
    .A(_2390_),
    .B(_2339_));
 sg13g2_nor3_1 _7283_ (.A(_2388_),
    .B(_2389_),
    .C(_2391_),
    .Y(_2392_));
 sg13g2_a21oi_1 _7284_ (.A1(_2339_),
    .A2(_2387_),
    .Y(_2393_),
    .B1(_2390_));
 sg13g2_a21oi_1 _7285_ (.A1(_2386_),
    .A2(_2392_),
    .Y(_2394_),
    .B1(_2393_));
 sg13g2_inv_1 _7286_ (.Y(_2395_),
    .A(_2394_));
 sg13g2_nand4_1 _7287_ (.B(\vgademo.soundtrack.pulse_osc_p[9] ),
    .C(\vgademo.soundtrack.pulse_osc_p[8] ),
    .A(_2395_),
    .Y(_2396_),
    .D(_2347_));
 sg13g2_xnor2_1 _7288_ (.Y(_0297_),
    .A(\vgademo.soundtrack.pulse_osc_p[10] ),
    .B(_2396_));
 sg13g2_inv_1 _7289_ (.Y(_2397_),
    .A(_2347_));
 sg13g2_nor2_1 _7290_ (.A(_0064_),
    .B(_2394_),
    .Y(_2398_));
 sg13g2_inv_1 _7291_ (.Y(_2399_),
    .A(_2398_));
 sg13g2_nor2_1 _7292_ (.A(_2397_),
    .B(_2399_),
    .Y(_2400_));
 sg13g2_nand2_1 _7293_ (.Y(_2401_),
    .A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .B(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_inv_1 _7294_ (.Y(_2402_),
    .A(_2401_));
 sg13g2_nand2_1 _7295_ (.Y(_2403_),
    .A(_2400_),
    .B(_2402_));
 sg13g2_xnor2_1 _7296_ (.Y(_0298_),
    .A(\vgademo.soundtrack.pulse_osc_p[11] ),
    .B(_2403_));
 sg13g2_nand4_1 _7297_ (.B(\vgademo.soundtrack.pulse_osc_p[8] ),
    .C(\vgademo.soundtrack.pulse_osc_p[11] ),
    .A(_2395_),
    .Y(_2404_),
    .D(_2402_));
 sg13g2_xnor2_1 _7298_ (.Y(_2405_),
    .A(_0062_),
    .B(_2404_));
 sg13g2_buf_1 _7299_ (.A(net35),
    .X(_2406_));
 sg13g2_buf_1 _7300_ (.A(_2347_),
    .X(_2407_));
 sg13g2_nor2_1 _7301_ (.A(\vgademo.soundtrack.pulse_osc_p[12] ),
    .B(net34),
    .Y(_2408_));
 sg13g2_a21oi_1 _7302_ (.A1(_2405_),
    .A2(net30),
    .Y(_0299_),
    .B1(_2408_));
 sg13g2_nand3_1 _7303_ (.B(\vgademo.soundtrack.pulse_osc_p[11] ),
    .C(\vgademo.soundtrack.pulse_osc_p[12] ),
    .A(_2402_),
    .Y(_2409_));
 sg13g2_nor2_1 _7304_ (.A(_2409_),
    .B(_2399_),
    .Y(_2410_));
 sg13g2_xor2_1 _7305_ (.B(_2410_),
    .A(_0061_),
    .X(_2411_));
 sg13g2_buf_1 _7306_ (.A(_2347_),
    .X(_2412_));
 sg13g2_nor2_1 _7307_ (.A(\vgademo.soundtrack.pulse_osc_p[13] ),
    .B(net33),
    .Y(_2413_));
 sg13g2_a21oi_1 _7308_ (.A1(_2411_),
    .A2(net30),
    .Y(_0300_),
    .B1(_2413_));
 sg13g2_nor2_1 _7309_ (.A(_2352_),
    .B(_2350_),
    .Y(_2414_));
 sg13g2_nand3b_1 _7310_ (.B(_2348_),
    .C(_2353_),
    .Y(_2415_),
    .A_N(_2414_));
 sg13g2_o21ai_1 _7311_ (.B1(_2415_),
    .Y(_0301_),
    .A1(_2351_),
    .A2(net34));
 sg13g2_nor2b_1 _7312_ (.A(_2363_),
    .B_N(_2362_),
    .Y(_2416_));
 sg13g2_xnor2_1 _7313_ (.Y(_2417_),
    .A(_2416_),
    .B(_2355_));
 sg13g2_nor2_1 _7314_ (.A(\vgademo.soundtrack.pulse_osc_p[2] ),
    .B(net33),
    .Y(_2418_));
 sg13g2_a21oi_1 _7315_ (.A1(_2417_),
    .A2(net30),
    .Y(_0302_),
    .B1(_2418_));
 sg13g2_xnor2_1 _7316_ (.Y(_2419_),
    .A(_2376_),
    .B(_2364_));
 sg13g2_nor2_1 _7317_ (.A(\vgademo.soundtrack.pulse_osc_p[3] ),
    .B(net33),
    .Y(_2420_));
 sg13g2_a21oi_1 _7318_ (.A1(_2419_),
    .A2(net30),
    .Y(_0303_),
    .B1(_2420_));
 sg13g2_a21oi_1 _7319_ (.A1(_2364_),
    .A2(_2375_),
    .Y(_2421_),
    .B1(_2374_));
 sg13g2_xor2_1 _7320_ (.B(_2421_),
    .A(_2370_),
    .X(_2422_));
 sg13g2_nor2_1 _7321_ (.A(\vgademo.soundtrack.pulse_osc_p[4] ),
    .B(net33),
    .Y(_2423_));
 sg13g2_a21oi_1 _7322_ (.A1(_2422_),
    .A2(net30),
    .Y(_0304_),
    .B1(_2423_));
 sg13g2_nand2b_1 _7323_ (.Y(_2424_),
    .B(_2383_),
    .A_N(_2384_));
 sg13g2_xnor2_1 _7324_ (.Y(_2425_),
    .A(_2424_),
    .B(_2379_));
 sg13g2_nor2_1 _7325_ (.A(\vgademo.soundtrack.pulse_osc_p[5] ),
    .B(_2412_),
    .Y(_2426_));
 sg13g2_a21oi_1 _7326_ (.A1(_2425_),
    .A2(_2406_),
    .Y(_0305_),
    .B1(_2426_));
 sg13g2_nor2_1 _7327_ (.A(_2389_),
    .B(_2388_),
    .Y(_2427_));
 sg13g2_a21oi_1 _7328_ (.A1(_2386_),
    .A2(_2427_),
    .Y(_2428_),
    .B1(_2397_));
 sg13g2_o21ai_1 _7329_ (.B1(_2428_),
    .Y(_2429_),
    .A1(_2427_),
    .A2(_2386_));
 sg13g2_o21ai_1 _7330_ (.B1(_2429_),
    .Y(_0306_),
    .A1(_2387_),
    .A2(_2407_));
 sg13g2_inv_1 _7331_ (.Y(_2430_),
    .A(_2389_));
 sg13g2_a21oi_1 _7332_ (.A1(_2386_),
    .A2(_2430_),
    .Y(_2431_),
    .B1(_2388_));
 sg13g2_xnor2_1 _7333_ (.Y(_2432_),
    .A(_2391_),
    .B(_2431_));
 sg13g2_nor2_1 _7334_ (.A(\vgademo.soundtrack.pulse_osc_p[7] ),
    .B(_2412_),
    .Y(_2433_));
 sg13g2_a21oi_1 _7335_ (.A1(_2432_),
    .A2(_2406_),
    .Y(_0307_),
    .B1(_2433_));
 sg13g2_inv_1 _7336_ (.Y(_2434_),
    .A(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_nand2_1 _7337_ (.Y(_2435_),
    .A(_2394_),
    .B(_0064_));
 sg13g2_nand3_1 _7338_ (.B(_2348_),
    .C(_2435_),
    .A(_2399_),
    .Y(_2436_));
 sg13g2_o21ai_1 _7339_ (.B1(_2436_),
    .Y(_0308_),
    .A1(_2434_),
    .A2(_2407_));
 sg13g2_xor2_1 _7340_ (.B(_2400_),
    .A(\vgademo.soundtrack.pulse_osc_p[9] ),
    .X(_0309_));
 sg13g2_nor2_1 _7341_ (.A(net97),
    .B(_2084_),
    .Y(_2437_));
 sg13g2_o21ai_1 _7342_ (.B1(_2437_),
    .Y(_2438_),
    .A1(net88),
    .A2(_0770_));
 sg13g2_a21oi_1 _7343_ (.A1(_2148_),
    .A2(_2438_),
    .Y(_2439_),
    .B1(_2098_));
 sg13g2_nand3_1 _7344_ (.B(net78),
    .C(net118),
    .A(_2097_),
    .Y(_2440_));
 sg13g2_xnor2_1 _7345_ (.Y(_2441_),
    .A(_0779_),
    .B(_2440_));
 sg13g2_nand3_1 _7346_ (.B(_2264_),
    .C(_2109_),
    .A(_2098_),
    .Y(_2442_));
 sg13g2_nand2_1 _7347_ (.Y(_2443_),
    .A(_2441_),
    .B(_2442_));
 sg13g2_inv_1 _7348_ (.Y(_2444_),
    .A(_2441_));
 sg13g2_a21oi_1 _7349_ (.A1(_0768_),
    .A2(net88),
    .Y(_2445_),
    .B1(net77));
 sg13g2_nand2b_1 _7350_ (.Y(_2446_),
    .B(_1665_),
    .A_N(_2322_));
 sg13g2_nor3_1 _7351_ (.A(net98),
    .B(_1661_),
    .C(_1693_),
    .Y(_2447_));
 sg13g2_a22oi_1 _7352_ (.Y(_2448_),
    .B1(_2446_),
    .B2(_2447_),
    .A2(_2445_),
    .A1(_2153_));
 sg13g2_a21oi_1 _7353_ (.A1(_2444_),
    .A2(_2448_),
    .Y(_2449_),
    .B1(_2107_));
 sg13g2_o21ai_1 _7354_ (.B1(_2449_),
    .Y(_2450_),
    .A1(_2439_),
    .A2(_2443_));
 sg13g2_a21oi_1 _7355_ (.A1(_1663_),
    .A2(_1664_),
    .Y(_2451_),
    .B1(_0772_));
 sg13g2_nand2_1 _7356_ (.Y(_2452_),
    .A(_2086_),
    .B(_0770_));
 sg13g2_nor2_1 _7357_ (.A(_2142_),
    .B(_2092_),
    .Y(_2453_));
 sg13g2_a22oi_1 _7358_ (.Y(_2454_),
    .B1(_2452_),
    .B2(_2453_),
    .A2(_2451_),
    .A1(_2099_));
 sg13g2_a21oi_1 _7359_ (.A1(_2444_),
    .A2(_2454_),
    .Y(_2455_),
    .B1(_2105_));
 sg13g2_a21oi_1 _7360_ (.A1(_2147_),
    .A2(net77),
    .Y(_2456_),
    .B1(_2437_));
 sg13g2_nand3_1 _7361_ (.B(_2154_),
    .C(_2277_),
    .A(_2453_),
    .Y(_2457_));
 sg13g2_nand3_1 _7362_ (.B(_2456_),
    .C(_2457_),
    .A(_2441_),
    .Y(_2458_));
 sg13g2_nand2_1 _7363_ (.Y(_2459_),
    .A(_2455_),
    .B(_2458_));
 sg13g2_nand3_1 _7364_ (.B(_2459_),
    .C(_2112_),
    .A(_2450_),
    .Y(_2460_));
 sg13g2_inv_1 _7365_ (.Y(_2461_),
    .A(_2108_));
 sg13g2_a21oi_1 _7366_ (.A1(_2461_),
    .A2(_2147_),
    .Y(_2462_),
    .B1(_2112_));
 sg13g2_o21ai_1 _7367_ (.B1(_1669_),
    .Y(_2463_),
    .A1(net79),
    .A2(_2108_));
 sg13g2_a21oi_1 _7368_ (.A1(_2462_),
    .A2(_2463_),
    .Y(_2464_),
    .B1(net75));
 sg13g2_nand2_1 _7369_ (.Y(_2465_),
    .A(_2460_),
    .B(_2464_));
 sg13g2_nand2_1 _7370_ (.Y(_2466_),
    .A(_2071_),
    .B(_2465_));
 sg13g2_buf_2 _7371_ (.A(_2466_),
    .X(_2467_));
 sg13g2_inv_1 _7372_ (.Y(_2468_),
    .A(_1791_));
 sg13g2_a21oi_1 _7373_ (.A1(net108),
    .A2(_2468_),
    .Y(_2469_),
    .B1(net76));
 sg13g2_nand2_1 _7374_ (.Y(_2470_),
    .A(_2467_),
    .B(_0100_));
 sg13g2_o21ai_1 _7375_ (.B1(_2470_),
    .Y(_0310_),
    .A1(_2467_),
    .A2(_2469_));
 sg13g2_a22oi_1 _7376_ (.Y(_2471_),
    .B1(net108),
    .B2(_1791_),
    .A2(_1716_),
    .A1(_1660_));
 sg13g2_nor2_1 _7377_ (.A(net76),
    .B(_2471_),
    .Y(_2472_));
 sg13g2_nand2_1 _7378_ (.Y(_2473_),
    .A(_2467_),
    .B(_0101_));
 sg13g2_o21ai_1 _7379_ (.B1(_2473_),
    .Y(_0311_),
    .A1(_2467_),
    .A2(_2472_));
 sg13g2_nand3_1 _7380_ (.B(_2468_),
    .C(net108),
    .A(_1657_),
    .Y(_2474_));
 sg13g2_nand2_1 _7381_ (.Y(_2475_),
    .A(_1659_),
    .B(_1727_));
 sg13g2_nand3_1 _7382_ (.B(_2474_),
    .C(_2475_),
    .A(net75),
    .Y(_2476_));
 sg13g2_mux2_1 _7383_ (.A0(_2476_),
    .A1(_0102_),
    .S(_2467_),
    .X(_0312_));
 sg13g2_a21oi_1 _7384_ (.A1(_1655_),
    .A2(net108),
    .Y(_2477_),
    .B1(_1719_));
 sg13g2_nor2_1 _7385_ (.A(_2477_),
    .B(net76),
    .Y(_2478_));
 sg13g2_nand2_1 _7386_ (.Y(_2479_),
    .A(_2467_),
    .B(_0103_));
 sg13g2_o21ai_1 _7387_ (.B1(_2479_),
    .Y(_0313_),
    .A1(_2467_),
    .A2(_2478_));
 sg13g2_inv_1 _7388_ (.Y(_2480_),
    .A(_0104_));
 sg13g2_a21oi_1 _7389_ (.A1(_2480_),
    .A2(_2066_),
    .Y(_0314_),
    .B1(_2074_));
 sg13g2_buf_1 _7390_ (.A(_2065_),
    .X(_2481_));
 sg13g2_nor2_1 _7391_ (.A(_0105_),
    .B(_2481_),
    .Y(_2482_));
 sg13g2_a21oi_1 _7392_ (.A1(_2264_),
    .A2(net29),
    .Y(_0315_),
    .B1(_2482_));
 sg13g2_nand2_1 _7393_ (.Y(_2483_),
    .A(_2086_),
    .B(_2296_));
 sg13g2_mux2_1 _7394_ (.A0(_0106_),
    .A1(_2483_),
    .S(net29),
    .X(_0316_));
 sg13g2_nor2_1 _7395_ (.A(_0107_),
    .B(net29),
    .Y(_2484_));
 sg13g2_a21oi_1 _7396_ (.A1(_2093_),
    .A2(net29),
    .Y(_0317_),
    .B1(_2484_));
 sg13g2_nor2_1 _7397_ (.A(_0108_),
    .B(net29),
    .Y(_2485_));
 sg13g2_a21oi_1 _7398_ (.A1(net29),
    .A2(_2098_),
    .Y(_0318_),
    .B1(_2485_));
 sg13g2_nor2_1 _7399_ (.A(_0109_),
    .B(_2065_),
    .Y(_2486_));
 sg13g2_a21oi_1 _7400_ (.A1(net29),
    .A2(_2105_),
    .Y(_0319_),
    .B1(_2486_));
 sg13g2_nor2_1 _7401_ (.A(_0110_),
    .B(_2065_),
    .Y(_2487_));
 sg13g2_a21oi_1 _7402_ (.A1(net29),
    .A2(_2112_),
    .Y(_0320_),
    .B1(_2487_));
 sg13g2_nor2_1 _7403_ (.A(_0111_),
    .B(_2065_),
    .Y(_2488_));
 sg13g2_a21oi_1 _7404_ (.A1(_2481_),
    .A2(_2444_),
    .Y(_0321_),
    .B1(_2488_));
 sg13g2_nand2_1 _7405_ (.Y(_2489_),
    .A(net48),
    .B(\vgademo.soundtrack.tick_div_[0] ));
 sg13g2_o21ai_1 _7406_ (.B1(_2489_),
    .Y(_0322_),
    .A1(_2015_),
    .A2(net48));
 sg13g2_xor2_1 _7407_ (.B(_2027_),
    .A(\vgademo.soundtrack.tick_div[1] ),
    .X(_0323_));
 sg13g2_xnor2_1 _7408_ (.Y(_0324_),
    .A(\vgademo.soundtrack.tick_div[2] ),
    .B(_2028_));
 sg13g2_xnor2_1 _7409_ (.Y(_0325_),
    .A(_2013_),
    .B(_2029_));
 sg13g2_xnor2_1 _7410_ (.Y(_0326_),
    .A(_2012_),
    .B(_2031_));
 sg13g2_xnor2_1 _7411_ (.Y(_0327_),
    .A(_2011_),
    .B(_2033_));
 sg13g2_xnor2_1 _7412_ (.Y(_0328_),
    .A(_2010_),
    .B(_2035_));
 sg13g2_xnor2_1 _7413_ (.Y(_0329_),
    .A(_2009_),
    .B(_2037_));
 sg13g2_buf_1 _7414_ (.A(\vgademo.soundtrack.tri_osc_i[0] ),
    .X(_2490_));
 sg13g2_inv_1 _7415_ (.Y(_2491_),
    .A(_2490_));
 sg13g2_inv_1 _7416_ (.Y(_2492_),
    .A(_2119_));
 sg13g2_buf_1 _7417_ (.A(_2081_),
    .X(_2493_));
 sg13g2_buf_2 _7418_ (.A(\vgademo.soundtrack.tri_osc_i[3] ),
    .X(_2494_));
 sg13g2_xnor2_1 _7419_ (.Y(_2495_),
    .A(_2490_),
    .B(_2494_));
 sg13g2_inv_1 _7420_ (.Y(_2496_),
    .A(_1686_));
 sg13g2_nand2_1 _7421_ (.Y(_2497_),
    .A(_1664_),
    .B(net79));
 sg13g2_nand2_1 _7422_ (.Y(_2498_),
    .A(_2497_),
    .B(net77));
 sg13g2_inv_1 _7423_ (.Y(_2499_),
    .A(_2498_));
 sg13g2_nand2b_1 _7424_ (.Y(_2500_),
    .B(_2499_),
    .A_N(_2262_));
 sg13g2_o21ai_1 _7425_ (.B1(_2500_),
    .Y(_2501_),
    .A1(_2496_),
    .A2(_2261_));
 sg13g2_a21oi_1 _7426_ (.A1(_2143_),
    .A2(_1676_),
    .Y(_2502_),
    .B1(net78));
 sg13g2_a21o_1 _7427_ (.A2(net78),
    .A1(_2501_),
    .B1(_2502_),
    .X(_2503_));
 sg13g2_buf_1 _7428_ (.A(_2503_),
    .X(_2504_));
 sg13g2_nand2_1 _7429_ (.Y(_2505_),
    .A(_2496_),
    .B(_1676_));
 sg13g2_a22oi_1 _7430_ (.Y(_2506_),
    .B1(_2270_),
    .B2(_2156_),
    .A2(net78),
    .A1(_2505_));
 sg13g2_buf_1 _7431_ (.A(_2506_),
    .X(_2507_));
 sg13g2_nand2_1 _7432_ (.Y(_2508_),
    .A(_2496_),
    .B(net77));
 sg13g2_a21oi_1 _7433_ (.A1(_2262_),
    .A2(net98),
    .Y(_2509_),
    .B1(net84));
 sg13g2_a22oi_1 _7434_ (.Y(_2510_),
    .B1(_2500_),
    .B2(_2509_),
    .A2(_2508_),
    .A1(_2502_));
 sg13g2_buf_1 _7435_ (.A(_2510_),
    .X(_2511_));
 sg13g2_inv_1 _7436_ (.Y(_2512_),
    .A(_2511_));
 sg13g2_a21o_1 _7437_ (.A2(_2507_),
    .A1(_2504_),
    .B1(_2512_),
    .X(_2513_));
 sg13g2_buf_1 _7438_ (.A(_2513_),
    .X(_2514_));
 sg13g2_inv_1 _7439_ (.Y(_2515_),
    .A(_2507_));
 sg13g2_o21ai_1 _7440_ (.B1(_2512_),
    .Y(_2516_),
    .A1(_2515_),
    .A2(_2504_));
 sg13g2_nand2_1 _7441_ (.Y(_2517_),
    .A(_2514_),
    .B(_2516_));
 sg13g2_mux2_1 _7442_ (.A0(_2295_),
    .A1(_2305_),
    .S(net98),
    .X(_2518_));
 sg13g2_inv_1 _7443_ (.Y(_2519_),
    .A(_2518_));
 sg13g2_a22oi_1 _7444_ (.Y(_2520_),
    .B1(_1692_),
    .B2(_2497_),
    .A2(net77),
    .A1(_2154_));
 sg13g2_nor3_1 _7445_ (.A(net78),
    .B(_2499_),
    .C(_2520_),
    .Y(_2521_));
 sg13g2_a21oi_1 _7446_ (.A1(_2519_),
    .A2(net78),
    .Y(_2522_),
    .B1(_2521_));
 sg13g2_buf_2 _7447_ (.A(_2522_),
    .X(_2523_));
 sg13g2_a21oi_1 _7448_ (.A1(_2517_),
    .A2(_2523_),
    .Y(_2524_),
    .B1(net74));
 sg13g2_a21oi_1 _7449_ (.A1(net74),
    .A2(_2495_),
    .Y(_2525_),
    .B1(_2524_));
 sg13g2_nand3_1 _7450_ (.B(_2060_),
    .C(_2492_),
    .A(_2525_),
    .Y(_2526_));
 sg13g2_o21ai_1 _7451_ (.B1(_2526_),
    .Y(_0330_),
    .A1(_2491_),
    .A2(_2492_));
 sg13g2_buf_1 _7452_ (.A(\vgademo.soundtrack.tri_osc_i[1] ),
    .X(_2527_));
 sg13g2_inv_1 _7453_ (.Y(_2528_),
    .A(_2527_));
 sg13g2_inv_1 _7454_ (.Y(_2529_),
    .A(_2494_));
 sg13g2_nor2_1 _7455_ (.A(_2490_),
    .B(_2529_),
    .Y(_2530_));
 sg13g2_buf_2 _7456_ (.A(\vgademo.soundtrack.tri_osc_i[4] ),
    .X(_2531_));
 sg13g2_xnor2_1 _7457_ (.Y(_2532_),
    .A(_2527_),
    .B(_2531_));
 sg13g2_xor2_1 _7458_ (.B(_2532_),
    .A(_2530_),
    .X(_2533_));
 sg13g2_inv_2 _7459_ (.Y(_2534_),
    .A(_2523_));
 sg13g2_nand2_1 _7460_ (.Y(_2535_),
    .A(_2517_),
    .B(_2534_));
 sg13g2_a21oi_1 _7461_ (.A1(_2514_),
    .A2(_2523_),
    .Y(_2536_),
    .B1(net74));
 sg13g2_a22oi_1 _7462_ (.Y(_2537_),
    .B1(_2535_),
    .B2(_2536_),
    .A2(_2533_),
    .A1(net74));
 sg13g2_nand2_1 _7463_ (.Y(_2538_),
    .A(_2047_),
    .B(_2537_));
 sg13g2_o21ai_1 _7464_ (.B1(_2538_),
    .Y(_0331_),
    .A1(_2528_),
    .A2(_2492_));
 sg13g2_buf_1 _7465_ (.A(\vgademo.soundtrack.tri_osc_i[2] ),
    .X(_2539_));
 sg13g2_buf_2 _7466_ (.A(\vgademo.soundtrack.tri_osc_i[5] ),
    .X(_2540_));
 sg13g2_xnor2_1 _7467_ (.Y(_2541_),
    .A(_2539_),
    .B(_2540_));
 sg13g2_nand2b_1 _7468_ (.Y(_2542_),
    .B(_2532_),
    .A_N(_2530_));
 sg13g2_o21ai_1 _7469_ (.B1(_2542_),
    .Y(_2543_),
    .A1(_2528_),
    .A2(_2531_));
 sg13g2_xor2_1 _7470_ (.B(_2543_),
    .A(_2541_),
    .X(_2544_));
 sg13g2_nor2_1 _7471_ (.A(_2507_),
    .B(_2504_),
    .Y(_2545_));
 sg13g2_nand2_1 _7472_ (.Y(_2546_),
    .A(_2545_),
    .B(_2512_));
 sg13g2_a21oi_1 _7473_ (.A1(_2514_),
    .A2(_2534_),
    .Y(_2547_),
    .B1(_2493_));
 sg13g2_o21ai_1 _7474_ (.B1(_2547_),
    .Y(_2548_),
    .A1(_2534_),
    .A2(_2546_));
 sg13g2_o21ai_1 _7475_ (.B1(_2548_),
    .Y(_2549_),
    .A1(_2080_),
    .A2(_2544_));
 sg13g2_nand2_1 _7476_ (.Y(_2550_),
    .A(_2119_),
    .B(_2539_));
 sg13g2_o21ai_1 _7477_ (.B1(_2550_),
    .Y(_0332_),
    .A1(_2549_),
    .A2(_2058_));
 sg13g2_nor2b_1 _7478_ (.A(_2540_),
    .B_N(_2539_),
    .Y(_2551_));
 sg13g2_a21oi_1 _7479_ (.A1(_2543_),
    .A2(_2541_),
    .Y(_2552_),
    .B1(_2551_));
 sg13g2_inv_1 _7480_ (.Y(_2553_),
    .A(_2552_));
 sg13g2_buf_1 _7481_ (.A(\vgademo.soundtrack.tri_osc_i[6] ),
    .X(_2554_));
 sg13g2_xnor2_1 _7482_ (.Y(_2555_),
    .A(_2494_),
    .B(_2554_));
 sg13g2_nand2_1 _7483_ (.Y(_2556_),
    .A(_2553_),
    .B(_2555_));
 sg13g2_inv_1 _7484_ (.Y(_2557_),
    .A(_2555_));
 sg13g2_a21oi_1 _7485_ (.A1(_2552_),
    .A2(_2557_),
    .Y(_2558_),
    .B1(_2080_));
 sg13g2_a21oi_1 _7486_ (.A1(_2546_),
    .A2(_2534_),
    .Y(_2559_),
    .B1(net74));
 sg13g2_nor2b_1 _7487_ (.A(_2507_),
    .B_N(_2504_),
    .Y(_2560_));
 sg13g2_nand2_1 _7488_ (.Y(_2561_),
    .A(_2560_),
    .B(_2511_));
 sg13g2_o21ai_1 _7489_ (.B1(_2561_),
    .Y(_2562_),
    .A1(_2560_),
    .A2(_2516_));
 sg13g2_nand2_1 _7490_ (.Y(_2563_),
    .A(_2562_),
    .B(_2523_));
 sg13g2_a22oi_1 _7491_ (.Y(_2564_),
    .B1(_2559_),
    .B2(_2563_),
    .A2(_2558_),
    .A1(_2556_));
 sg13g2_nand2_1 _7492_ (.Y(_2565_),
    .A(_2119_),
    .B(_2494_));
 sg13g2_o21ai_1 _7493_ (.B1(_2565_),
    .Y(_0333_),
    .A1(_2564_),
    .A2(_2058_));
 sg13g2_buf_2 _7494_ (.A(\vgademo.soundtrack.tri_osc_i[7] ),
    .X(_2566_));
 sg13g2_xnor2_1 _7495_ (.Y(_2567_),
    .A(_2531_),
    .B(_2566_));
 sg13g2_o21ai_1 _7496_ (.B1(_2556_),
    .Y(_2568_),
    .A1(_2529_),
    .A2(_2554_));
 sg13g2_xor2_1 _7497_ (.B(_2568_),
    .A(_2567_),
    .X(_2569_));
 sg13g2_nand2_1 _7498_ (.Y(_2570_),
    .A(_2514_),
    .B(_2546_));
 sg13g2_inv_1 _7499_ (.Y(_2571_),
    .A(_2570_));
 sg13g2_a21oi_1 _7500_ (.A1(_2571_),
    .A2(_2523_),
    .Y(_2572_),
    .B1(_2081_));
 sg13g2_o21ai_1 _7501_ (.B1(_2572_),
    .Y(_2573_),
    .A1(_2523_),
    .A2(_2562_));
 sg13g2_o21ai_1 _7502_ (.B1(_2573_),
    .Y(_2574_),
    .A1(_2080_),
    .A2(_2569_));
 sg13g2_nand2_1 _7503_ (.Y(_2575_),
    .A(_2119_),
    .B(_2531_));
 sg13g2_o21ai_1 _7504_ (.B1(_2575_),
    .Y(_0334_),
    .A1(_2574_),
    .A2(_2058_));
 sg13g2_buf_2 _7505_ (.A(\vgademo.soundtrack.tri_osc_i[8] ),
    .X(_2576_));
 sg13g2_xnor2_1 _7506_ (.Y(_2577_),
    .A(_2540_),
    .B(_2576_));
 sg13g2_inv_1 _7507_ (.Y(_2578_),
    .A(_2531_));
 sg13g2_nand2_1 _7508_ (.Y(_2579_),
    .A(_2568_),
    .B(_2567_));
 sg13g2_o21ai_1 _7509_ (.B1(_2579_),
    .Y(_2580_),
    .A1(_2578_),
    .A2(_2566_));
 sg13g2_xor2_1 _7510_ (.B(_2580_),
    .A(_2577_),
    .X(_2581_));
 sg13g2_nor3_1 _7511_ (.A(_2511_),
    .B(_2534_),
    .C(_2560_),
    .Y(_2582_));
 sg13g2_nor2_1 _7512_ (.A(_2493_),
    .B(_2582_),
    .Y(_2583_));
 sg13g2_o21ai_1 _7513_ (.B1(_2583_),
    .Y(_2584_),
    .A1(_2523_),
    .A2(_2570_));
 sg13g2_o21ai_1 _7514_ (.B1(_2584_),
    .Y(_2585_),
    .A1(_2080_),
    .A2(_2581_));
 sg13g2_nand2_1 _7515_ (.Y(_2586_),
    .A(_2119_),
    .B(_2540_));
 sg13g2_o21ai_1 _7516_ (.B1(_2586_),
    .Y(_0335_),
    .A1(_2585_),
    .A2(_2058_));
 sg13g2_inv_1 _7517_ (.Y(_2587_),
    .A(_2554_));
 sg13g2_a21oi_1 _7518_ (.A1(_2560_),
    .A2(_2534_),
    .Y(_2588_),
    .B1(_2511_));
 sg13g2_inv_1 _7519_ (.Y(_2589_),
    .A(_2540_));
 sg13g2_nand2_1 _7520_ (.Y(_2590_),
    .A(_2580_),
    .B(_2577_));
 sg13g2_o21ai_1 _7521_ (.B1(_2590_),
    .Y(_2591_),
    .A1(_2589_),
    .A2(_2576_));
 sg13g2_nand2b_1 _7522_ (.Y(_2592_),
    .B(_2587_),
    .A_N(_2591_));
 sg13g2_nand2_1 _7523_ (.Y(_2593_),
    .A(_2591_),
    .B(_2554_));
 sg13g2_a21oi_1 _7524_ (.A1(_2592_),
    .A2(_2593_),
    .Y(_2594_),
    .B1(_2080_));
 sg13g2_a21oi_1 _7525_ (.A1(_2080_),
    .A2(_2588_),
    .Y(_2595_),
    .B1(_2594_));
 sg13g2_a22oi_1 _7526_ (.Y(_0336_),
    .B1(_2595_),
    .B2(_2047_),
    .A2(_2119_),
    .A1(_2587_));
 sg13g2_inv_1 _7527_ (.Y(_2596_),
    .A(_2566_));
 sg13g2_xnor2_1 _7528_ (.Y(_2597_),
    .A(_2596_),
    .B(_2592_));
 sg13g2_nand3_1 _7529_ (.B(_2060_),
    .C(net74),
    .A(_2597_),
    .Y(_2598_));
 sg13g2_nand2_1 _7530_ (.Y(_2599_),
    .A(_2534_),
    .B(_2512_));
 sg13g2_nand2_1 _7531_ (.Y(_2600_),
    .A(_2523_),
    .B(_2511_));
 sg13g2_nand3_1 _7532_ (.B(_2082_),
    .C(_2600_),
    .A(_2599_),
    .Y(_2601_));
 sg13g2_nand3_1 _7533_ (.B(_2492_),
    .C(_2601_),
    .A(_2598_),
    .Y(_2602_));
 sg13g2_o21ai_1 _7534_ (.B1(_2602_),
    .Y(_0337_),
    .A1(_2596_),
    .A2(_2492_));
 sg13g2_inv_1 _7535_ (.Y(_2603_),
    .A(_2576_));
 sg13g2_o21ai_1 _7536_ (.B1(_2576_),
    .Y(_2604_),
    .A1(_2566_),
    .A2(_2592_));
 sg13g2_a21oi_1 _7537_ (.A1(_2534_),
    .A2(_2511_),
    .Y(_2605_),
    .B1(net74));
 sg13g2_a21o_1 _7538_ (.A2(net74),
    .A1(_2604_),
    .B1(_2605_),
    .X(_2606_));
 sg13g2_a22oi_1 _7539_ (.Y(_0338_),
    .B1(_2047_),
    .B2(_2606_),
    .A2(_2119_),
    .A1(_2603_));
 sg13g2_nand2_1 _7540_ (.Y(_2607_),
    .A(net35),
    .B(_2490_));
 sg13g2_xnor2_1 _7541_ (.Y(_0339_),
    .A(\vgademo.soundtrack.tri_osc_p[0] ),
    .B(_2607_));
 sg13g2_inv_1 _7542_ (.Y(_2608_),
    .A(_1783_));
 sg13g2_nor2_1 _7543_ (.A(_2540_),
    .B(_1824_),
    .Y(_2609_));
 sg13g2_nand2_1 _7544_ (.Y(_2610_),
    .A(_2490_),
    .B(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_xor2_1 _7545_ (.B(_1884_),
    .A(_2527_),
    .X(_2611_));
 sg13g2_inv_1 _7546_ (.Y(_2612_),
    .A(_2611_));
 sg13g2_nand2_1 _7547_ (.Y(_2613_),
    .A(_2527_),
    .B(_1884_));
 sg13g2_o21ai_1 _7548_ (.B1(_2613_),
    .Y(_2614_),
    .A1(_2610_),
    .A2(_2612_));
 sg13g2_xor2_1 _7549_ (.B(_1877_),
    .A(_2539_),
    .X(_2615_));
 sg13g2_and2_1 _7550_ (.A(_2614_),
    .B(_2615_),
    .X(_2616_));
 sg13g2_a21oi_1 _7551_ (.A1(_2539_),
    .A2(_1877_),
    .Y(_2617_),
    .B1(_2616_));
 sg13g2_nand2_1 _7552_ (.Y(_2618_),
    .A(_2494_),
    .B(_1862_));
 sg13g2_nor2_1 _7553_ (.A(_2494_),
    .B(_1862_),
    .Y(_2619_));
 sg13g2_a21oi_1 _7554_ (.A1(_2617_),
    .A2(_2618_),
    .Y(_2620_),
    .B1(_2619_));
 sg13g2_nor2_1 _7555_ (.A(_2531_),
    .B(_1844_),
    .Y(_2621_));
 sg13g2_inv_1 _7556_ (.Y(_2622_),
    .A(_2621_));
 sg13g2_nand2_1 _7557_ (.Y(_2623_),
    .A(_2531_),
    .B(_1844_));
 sg13g2_inv_1 _7558_ (.Y(_2624_),
    .A(_2623_));
 sg13g2_a21oi_1 _7559_ (.A1(_2620_),
    .A2(_2622_),
    .Y(_2625_),
    .B1(_2624_));
 sg13g2_nand2_1 _7560_ (.Y(_2626_),
    .A(_2540_),
    .B(_1824_));
 sg13g2_o21ai_1 _7561_ (.B1(_2626_),
    .Y(_2627_),
    .A1(_2609_),
    .A2(_2625_));
 sg13g2_nor2_1 _7562_ (.A(_2554_),
    .B(_1805_),
    .Y(_2628_));
 sg13g2_inv_1 _7563_ (.Y(_2629_),
    .A(_2628_));
 sg13g2_nand2_1 _7564_ (.Y(_2630_),
    .A(_2554_),
    .B(_1805_));
 sg13g2_inv_1 _7565_ (.Y(_2631_),
    .A(_2630_));
 sg13g2_a221oi_1 _7566_ (.B2(_2629_),
    .C1(_2631_),
    .B1(_2627_),
    .A1(_2566_),
    .Y(_2632_),
    .A2(_1783_));
 sg13g2_a21oi_1 _7567_ (.A1(_2596_),
    .A2(_2608_),
    .Y(_2633_),
    .B1(_2632_));
 sg13g2_xor2_1 _7568_ (.B(_1766_),
    .A(_2576_),
    .X(_2634_));
 sg13g2_and2_1 _7569_ (.A(_2633_),
    .B(_2634_),
    .X(_2635_));
 sg13g2_a21oi_1 _7570_ (.A1(_2576_),
    .A2(_1766_),
    .Y(_2636_),
    .B1(_2635_));
 sg13g2_nor2_1 _7571_ (.A(_0065_),
    .B(_2636_),
    .Y(_2637_));
 sg13g2_nand2_1 _7572_ (.Y(_2638_),
    .A(_2637_),
    .B(_2347_));
 sg13g2_xnor2_1 _7573_ (.Y(_0340_),
    .A(_1634_),
    .B(_2638_));
 sg13g2_inv_1 _7574_ (.Y(_2639_),
    .A(_2636_));
 sg13g2_nand4_1 _7575_ (.B(_1634_),
    .C(\vgademo.soundtrack.tri_osc_p[9] ),
    .A(_2639_),
    .Y(_2640_),
    .D(_2347_));
 sg13g2_xnor2_1 _7576_ (.Y(_0341_),
    .A(_1924_),
    .B(_2640_));
 sg13g2_inv_1 _7577_ (.Y(_2641_),
    .A(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_inv_1 _7578_ (.Y(_2642_),
    .A(_1924_));
 sg13g2_inv_1 _7579_ (.Y(_2643_),
    .A(_1634_));
 sg13g2_nor3_1 _7580_ (.A(_2642_),
    .B(_2643_),
    .C(_2638_),
    .Y(_2644_));
 sg13g2_xnor2_1 _7581_ (.Y(_0342_),
    .A(_2641_),
    .B(_2644_));
 sg13g2_nor3_1 _7582_ (.A(_2641_),
    .B(_2642_),
    .C(_2640_),
    .Y(_2645_));
 sg13g2_xor2_1 _7583_ (.B(_2645_),
    .A(\vgademo.soundtrack.tri_osc_p[13] ),
    .X(_0343_));
 sg13g2_inv_1 _7584_ (.Y(_2646_),
    .A(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_nand3_1 _7585_ (.B(\vgademo.soundtrack.tri_osc_p[12] ),
    .C(_1924_),
    .A(\vgademo.soundtrack.tri_osc_p[13] ),
    .Y(_2647_));
 sg13g2_nor3_1 _7586_ (.A(_2643_),
    .B(_2647_),
    .C(_2638_),
    .Y(_2648_));
 sg13g2_xnor2_1 _7587_ (.Y(_0344_),
    .A(_2646_),
    .B(_2648_));
 sg13g2_nor3_1 _7588_ (.A(_2646_),
    .B(_2647_),
    .C(_2640_),
    .Y(_2649_));
 sg13g2_xor2_1 _7589_ (.B(_2649_),
    .A(_1633_),
    .X(_0345_));
 sg13g2_xor2_1 _7590_ (.B(_2611_),
    .A(_2610_),
    .X(_2650_));
 sg13g2_nor2_1 _7591_ (.A(_1884_),
    .B(net33),
    .Y(_2651_));
 sg13g2_a21oi_1 _7592_ (.A1(net30),
    .A2(_2650_),
    .Y(_0346_),
    .B1(_2651_));
 sg13g2_xnor2_1 _7593_ (.Y(_2652_),
    .A(_2615_),
    .B(_2614_));
 sg13g2_nor2_1 _7594_ (.A(_1877_),
    .B(net33),
    .Y(_2653_));
 sg13g2_a21oi_1 _7595_ (.A1(net30),
    .A2(_2652_),
    .Y(_0347_),
    .B1(_2653_));
 sg13g2_nand2b_1 _7596_ (.Y(_2654_),
    .B(_2618_),
    .A_N(_2619_));
 sg13g2_xnor2_1 _7597_ (.Y(_2655_),
    .A(_2654_),
    .B(_2617_));
 sg13g2_nor2_1 _7598_ (.A(_1862_),
    .B(net33),
    .Y(_2656_));
 sg13g2_a21oi_1 _7599_ (.A1(net30),
    .A2(_2655_),
    .Y(_0348_),
    .B1(_2656_));
 sg13g2_nor2_1 _7600_ (.A(_2621_),
    .B(_2624_),
    .Y(_2657_));
 sg13g2_xnor2_1 _7601_ (.Y(_2658_),
    .A(_2657_),
    .B(_2620_));
 sg13g2_nor2_1 _7602_ (.A(_1844_),
    .B(net33),
    .Y(_2659_));
 sg13g2_a21oi_1 _7603_ (.A1(_2658_),
    .A2(net34),
    .Y(_0349_),
    .B1(_2659_));
 sg13g2_nand2b_1 _7604_ (.Y(_2660_),
    .B(_2626_),
    .A_N(_2609_));
 sg13g2_xnor2_1 _7605_ (.Y(_2661_),
    .A(_2660_),
    .B(_2625_));
 sg13g2_nor2_1 _7606_ (.A(_1824_),
    .B(net35),
    .Y(_2662_));
 sg13g2_a21oi_1 _7607_ (.A1(_2661_),
    .A2(net34),
    .Y(_0350_),
    .B1(_2662_));
 sg13g2_nor2_1 _7608_ (.A(_2628_),
    .B(_2631_),
    .Y(_2663_));
 sg13g2_xnor2_1 _7609_ (.Y(_2664_),
    .A(_2663_),
    .B(_2627_));
 sg13g2_nor2_1 _7610_ (.A(_1805_),
    .B(net35),
    .Y(_2665_));
 sg13g2_a21oi_1 _7611_ (.A1(_2664_),
    .A2(net34),
    .Y(_0351_),
    .B1(_2665_));
 sg13g2_xor2_1 _7612_ (.B(_1783_),
    .A(_2566_),
    .X(_2666_));
 sg13g2_a21oi_1 _7613_ (.A1(_2627_),
    .A2(_2629_),
    .Y(_2667_),
    .B1(_2631_));
 sg13g2_xor2_1 _7614_ (.B(_2667_),
    .A(_2666_),
    .X(_2668_));
 sg13g2_nor2_1 _7615_ (.A(_1783_),
    .B(net35),
    .Y(_2669_));
 sg13g2_a21oi_1 _7616_ (.A1(_2668_),
    .A2(net34),
    .Y(_0352_),
    .B1(_2669_));
 sg13g2_xnor2_1 _7617_ (.Y(_2670_),
    .A(_2634_),
    .B(_2633_));
 sg13g2_nor2_1 _7618_ (.A(_1766_),
    .B(net35),
    .Y(_2671_));
 sg13g2_a21oi_1 _7619_ (.A1(_2670_),
    .A2(net34),
    .Y(_0353_),
    .B1(_2671_));
 sg13g2_xnor2_1 _7620_ (.Y(_2672_),
    .A(_0065_),
    .B(_2636_));
 sg13g2_nor2_1 _7621_ (.A(\vgademo.soundtrack.tri_osc_p[9] ),
    .B(net35),
    .Y(_2673_));
 sg13g2_a21oi_1 _7622_ (.A1(_2672_),
    .A2(net34),
    .Y(_0354_),
    .B1(_2673_));
 sg13g2_nor2b_1 _7623_ (.A(_4425_),
    .B_N(_4487_),
    .Y(_2674_));
 sg13g2_inv_2 _7624_ (.Y(_2675_),
    .A(_2674_));
 sg13g2_nor2_1 _7625_ (.A(_4390_),
    .B(_4425_),
    .Y(_2676_));
 sg13g2_a21oi_1 _7626_ (.A1(_2675_),
    .A2(_4390_),
    .Y(_0355_),
    .B1(_2676_));
 sg13g2_nand2_1 _7627_ (.Y(_2677_),
    .A(_4456_),
    .B(_4389_));
 sg13g2_nand3_1 _7628_ (.B(_4570_),
    .C(_2677_),
    .A(net73),
    .Y(_2678_));
 sg13g2_o21ai_1 _7629_ (.B1(_2678_),
    .Y(_0356_),
    .A1(_4457_),
    .A2(net73));
 sg13g2_xnor2_1 _7630_ (.Y(_2679_),
    .A(_0020_),
    .B(_2677_));
 sg13g2_nand2_1 _7631_ (.Y(_2680_),
    .A(_4402_),
    .B(_4455_));
 sg13g2_o21ai_1 _7632_ (.B1(_2680_),
    .Y(_0357_),
    .A1(_2679_),
    .A2(_2675_));
 sg13g2_nor2_1 _7633_ (.A(_0964_),
    .B(_2677_),
    .Y(_2681_));
 sg13g2_xnor2_1 _7634_ (.Y(_2682_),
    .A(_0960_),
    .B(_2681_));
 sg13g2_nand2_1 _7635_ (.Y(_2683_),
    .A(_4402_),
    .B(_4458_));
 sg13g2_o21ai_1 _7636_ (.B1(_2683_),
    .Y(_0358_),
    .A1(_2682_),
    .A2(_2675_));
 sg13g2_nor2_1 _7637_ (.A(_4484_),
    .B(_2677_),
    .Y(_2684_));
 sg13g2_xnor2_1 _7638_ (.Y(_2685_),
    .A(_0983_),
    .B(_2684_));
 sg13g2_nand2_1 _7639_ (.Y(_2686_),
    .A(_4402_),
    .B(net122));
 sg13g2_o21ai_1 _7640_ (.B1(_2686_),
    .Y(_0359_),
    .A1(_2685_),
    .A2(_2675_));
 sg13g2_nand2_1 _7641_ (.Y(_2687_),
    .A(_2684_),
    .B(net122));
 sg13g2_a21oi_1 _7642_ (.A1(_1016_),
    .A2(_2687_),
    .Y(_2688_),
    .B1(_2675_));
 sg13g2_o21ai_1 _7643_ (.B1(_2688_),
    .Y(_2689_),
    .A1(_1016_),
    .A2(_2687_));
 sg13g2_o21ai_1 _7644_ (.B1(_2689_),
    .Y(_0360_),
    .A1(_4449_),
    .A2(net73));
 sg13g2_nor2_1 _7645_ (.A(_4449_),
    .B(_2687_),
    .Y(_2690_));
 sg13g2_inv_1 _7646_ (.Y(_2691_),
    .A(_2690_));
 sg13g2_a21oi_1 _7647_ (.A1(_1031_),
    .A2(_2691_),
    .Y(_2692_),
    .B1(_2675_));
 sg13g2_o21ai_1 _7648_ (.B1(_2692_),
    .Y(_2693_),
    .A1(_1031_),
    .A2(_2691_));
 sg13g2_o21ai_1 _7649_ (.B1(_2693_),
    .Y(_0361_),
    .A1(_0406_),
    .A2(_4404_));
 sg13g2_nor2_1 _7650_ (.A(_0406_),
    .B(_2691_),
    .Y(_2694_));
 sg13g2_xor2_1 _7651_ (.B(_2694_),
    .A(_1076_),
    .X(_2695_));
 sg13g2_nand2_1 _7652_ (.Y(_2696_),
    .A(_4402_),
    .B(net121));
 sg13g2_o21ai_1 _7653_ (.B1(_2696_),
    .Y(_0362_),
    .A1(_2675_),
    .A2(_2695_));
 sg13g2_nand2_1 _7654_ (.Y(_2697_),
    .A(_2694_),
    .B(net121));
 sg13g2_xnor2_1 _7655_ (.Y(_2698_),
    .A(_1071_),
    .B(_2697_));
 sg13g2_nand2_1 _7656_ (.Y(_2699_),
    .A(_4402_),
    .B(_4450_));
 sg13g2_o21ai_1 _7657_ (.B1(_2699_),
    .Y(_0363_),
    .A1(_2675_),
    .A2(_2698_));
 sg13g2_inv_1 _7658_ (.Y(_2700_),
    .A(_4447_));
 sg13g2_nor3_1 _7659_ (.A(_4451_),
    .B(_0040_),
    .C(_2697_),
    .Y(_2701_));
 sg13g2_o21ai_1 _7660_ (.B1(_0040_),
    .Y(_2702_),
    .A1(_4451_),
    .A2(_2697_));
 sg13g2_nand3b_1 _7661_ (.B(_2702_),
    .C(_2674_),
    .Y(_2703_),
    .A_N(_2701_));
 sg13g2_o21ai_1 _7662_ (.B1(_2703_),
    .Y(_0364_),
    .A1(_2700_),
    .A2(_4404_));
 sg13g2_a21o_1 _7663_ (.A2(_1086_),
    .A1(_0082_),
    .B1(net51),
    .X(_0213_));
 sg13g2_nand2_1 _7664_ (.Y(_2704_),
    .A(\vgademo.plane_dx_div.i[1] ),
    .B(\vgademo.plane_dx_div.i[0] ));
 sg13g2_inv_1 _7665_ (.Y(_2705_),
    .A(_2704_));
 sg13g2_nor3_1 _7666_ (.A(_1084_),
    .B(_2705_),
    .C(net51),
    .Y(_0214_));
 sg13g2_o21ai_1 _7667_ (.B1(net59),
    .Y(_2706_),
    .A1(\vgademo.plane_dx_div.i[2] ),
    .A2(_2705_));
 sg13g2_nand2_1 _7668_ (.Y(_2707_),
    .A(_2705_),
    .B(\vgademo.plane_dx_div.i[2] ));
 sg13g2_nor2b_1 _7669_ (.A(_2706_),
    .B_N(_2707_),
    .Y(_0215_));
 sg13g2_xnor2_1 _7670_ (.Y(_2708_),
    .A(_1085_),
    .B(_2707_));
 sg13g2_nor2_1 _7671_ (.A(_2708_),
    .B(net51),
    .Y(_0216_));
 sg13g2_a22oi_1 _7672_ (.Y(_0217_),
    .B1(_0869_),
    .B2(net38),
    .A2(_0856_),
    .A1(_1101_));
 sg13g2_nand2_1 _7673_ (.Y(_2709_),
    .A(net38),
    .B(net113));
 sg13g2_o21ai_1 _7674_ (.B1(_2709_),
    .Y(_0218_),
    .A1(_0869_),
    .A2(net50));
 sg13g2_nand2_1 _7675_ (.Y(_2710_),
    .A(net38),
    .B(net112));
 sg13g2_o21ai_1 _7676_ (.B1(_2710_),
    .Y(_0219_),
    .A1(_0873_),
    .A2(net50));
 sg13g2_nand2_1 _7677_ (.Y(_2711_),
    .A(net38),
    .B(_0879_));
 sg13g2_o21ai_1 _7678_ (.B1(_2711_),
    .Y(_0220_),
    .A1(_0876_),
    .A2(net50));
 sg13g2_nand2_1 _7679_ (.Y(_2712_),
    .A(net38),
    .B(_0883_));
 sg13g2_o21ai_1 _7680_ (.B1(_2712_),
    .Y(_0221_),
    .A1(_0880_),
    .A2(_1100_));
 sg13g2_nand2_1 _7681_ (.Y(_2713_),
    .A(net40),
    .B(_0887_));
 sg13g2_o21ai_1 _7682_ (.B1(_2713_),
    .Y(_0222_),
    .A1(_0884_),
    .A2(net50));
 sg13g2_nand2_1 _7683_ (.Y(_2714_),
    .A(net40),
    .B(_0891_));
 sg13g2_o21ai_1 _7684_ (.B1(_2714_),
    .Y(_0223_),
    .A1(_0888_),
    .A2(_1100_));
 sg13g2_nand2_1 _7685_ (.Y(_2715_),
    .A(net40),
    .B(_0895_));
 sg13g2_o21ai_1 _7686_ (.B1(_2715_),
    .Y(_0224_),
    .A1(_0892_),
    .A2(net50));
 sg13g2_nand2_1 _7687_ (.Y(_2716_),
    .A(net40),
    .B(net110));
 sg13g2_o21ai_1 _7688_ (.B1(_2716_),
    .Y(_0225_),
    .A1(_0896_),
    .A2(net50));
 sg13g2_nand2_1 _7689_ (.Y(_2717_),
    .A(net40),
    .B(_0864_));
 sg13g2_o21ai_1 _7690_ (.B1(_2717_),
    .Y(_0226_),
    .A1(_0900_),
    .A2(net50));
 sg13g2_nand3_1 _7691_ (.B(_1074_),
    .C(_2700_),
    .A(_1072_),
    .Y(_2718_));
 sg13g2_nor2_1 _7692_ (.A(_1035_),
    .B(_2718_),
    .Y(_2719_));
 sg13g2_nand2_1 _7693_ (.Y(_2720_),
    .A(_2719_),
    .B(_1055_));
 sg13g2_nand2_1 _7694_ (.Y(_2721_),
    .A(_0945_),
    .B(_4455_));
 sg13g2_nand2_1 _7695_ (.Y(_2722_),
    .A(_2721_),
    .B(_0965_));
 sg13g2_nand2_1 _7696_ (.Y(_2723_),
    .A(_0961_),
    .B(_0963_));
 sg13g2_nor2_1 _7697_ (.A(_2722_),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_inv_1 _7698_ (.Y(_2725_),
    .A(_1016_));
 sg13g2_nand3_1 _7699_ (.B(_1006_),
    .C(_2725_),
    .A(_1001_),
    .Y(_2726_));
 sg13g2_nand2_1 _7700_ (.Y(_2727_),
    .A(_1017_),
    .B(_2726_));
 sg13g2_nor2_1 _7701_ (.A(_0986_),
    .B(_2727_),
    .Y(_2728_));
 sg13g2_nand2_1 _7702_ (.Y(_2729_),
    .A(_2724_),
    .B(_2728_));
 sg13g2_nor2_1 _7703_ (.A(_2720_),
    .B(_2729_),
    .Y(_2730_));
 sg13g2_nand3_1 _7704_ (.B(_4392_),
    .C(_0914_),
    .A(_0913_),
    .Y(_2731_));
 sg13g2_nand2_1 _7705_ (.Y(_2732_),
    .A(_0912_),
    .B(_0947_));
 sg13g2_nand2_1 _7706_ (.Y(_2733_),
    .A(_2731_),
    .B(_2732_));
 sg13g2_nand2_1 _7707_ (.Y(_2734_),
    .A(_1054_),
    .B(_0405_));
 sg13g2_nand2_1 _7708_ (.Y(_2735_),
    .A(_1030_),
    .B(_0406_));
 sg13g2_a21oi_1 _7709_ (.A1(_2734_),
    .A2(_2735_),
    .Y(_2736_),
    .B1(_2718_));
 sg13g2_nand3_1 _7710_ (.B(net121),
    .C(_1053_),
    .A(_1050_),
    .Y(_2737_));
 sg13g2_nand2_1 _7711_ (.Y(_2738_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_nor2_1 _7712_ (.A(_4450_),
    .B(_4447_),
    .Y(_2739_));
 sg13g2_nand2_1 _7713_ (.Y(_2740_),
    .A(_1070_),
    .B(_2739_));
 sg13g2_nand2_1 _7714_ (.Y(_2741_),
    .A(_2738_),
    .B(_2740_));
 sg13g2_a21oi_1 _7715_ (.A1(_2730_),
    .A2(_2733_),
    .Y(_2742_),
    .B1(_2741_));
 sg13g2_nand3_1 _7716_ (.B(_0958_),
    .C(_4459_),
    .A(_0956_),
    .Y(_2743_));
 sg13g2_nand2_1 _7717_ (.Y(_2744_),
    .A(_0968_),
    .B(_2743_));
 sg13g2_nand2_1 _7718_ (.Y(_2745_),
    .A(_2744_),
    .B(_2728_));
 sg13g2_nor2_1 _7719_ (.A(net122),
    .B(_0982_),
    .Y(_2746_));
 sg13g2_nor2b_1 _7720_ (.A(_2727_),
    .B_N(_2746_),
    .Y(_2747_));
 sg13g2_a21oi_1 _7721_ (.A1(_4449_),
    .A2(_1007_),
    .Y(_2748_),
    .B1(_2747_));
 sg13g2_nand2_1 _7722_ (.Y(_2749_),
    .A(_2745_),
    .B(_2748_));
 sg13g2_nand2b_1 _7723_ (.Y(_2750_),
    .B(_2749_),
    .A_N(_2720_));
 sg13g2_nand2_2 _7724_ (.Y(_2751_),
    .A(_2742_),
    .B(_2750_));
 sg13g2_nand3b_1 _7725_ (.B(_2730_),
    .C(_4391_),
    .Y(_2752_),
    .A_N(_2731_));
 sg13g2_buf_2 _7726_ (.A(_2752_),
    .X(_2753_));
 sg13g2_nand2_2 _7727_ (.Y(_2754_),
    .A(_2751_),
    .B(_2753_));
 sg13g2_buf_8 _7728_ (.A(_2754_),
    .X(_2755_));
 sg13g2_buf_1 _7729_ (.A(net27),
    .X(_2756_));
 sg13g2_nor2_1 _7730_ (.A(_2725_),
    .B(_2756_),
    .Y(_2757_));
 sg13g2_a21oi_1 _7731_ (.A1(_0071_),
    .A2(net24),
    .Y(_2758_),
    .B1(_2757_));
 sg13g2_xnor2_1 _7732_ (.Y(_2759_),
    .A(_0554_),
    .B(_2758_));
 sg13g2_nor2b_1 _7733_ (.A(net27),
    .B_N(_0947_),
    .Y(_2760_));
 sg13g2_a21oi_1 _7734_ (.A1(_0068_),
    .A2(net24),
    .Y(_2761_),
    .B1(_2760_));
 sg13g2_inv_1 _7735_ (.Y(_2762_),
    .A(_2761_));
 sg13g2_inv_4 _7736_ (.A(_2754_),
    .Y(_2763_));
 sg13g2_buf_1 _7737_ (.A(_2763_),
    .X(_2764_));
 sg13g2_nor2_1 _7738_ (.A(_4389_),
    .B(_0583_),
    .Y(_2765_));
 sg13g2_nand2b_1 _7739_ (.Y(_2766_),
    .B(\vgademo.b_cos[5] ),
    .A_N(\vgademo.plane_du[2] ));
 sg13g2_a21oi_1 _7740_ (.A1(net23),
    .A2(_4389_),
    .Y(_2767_),
    .B1(_2766_));
 sg13g2_a21oi_1 _7741_ (.A1(net23),
    .A2(_2765_),
    .Y(_2768_),
    .B1(_2767_));
 sg13g2_o21ai_1 _7742_ (.B1(_2768_),
    .Y(_2769_),
    .A1(_0591_),
    .A2(_2761_));
 sg13g2_o21ai_1 _7743_ (.B1(_2769_),
    .Y(_2770_),
    .A1(_0590_),
    .A2(_2762_));
 sg13g2_nor2_1 _7744_ (.A(_0929_),
    .B(net27),
    .Y(_2771_));
 sg13g2_a21oi_1 _7745_ (.A1(_0067_),
    .A2(net24),
    .Y(_2772_),
    .B1(_2771_));
 sg13g2_nand2b_1 _7746_ (.Y(_2773_),
    .B(_0588_),
    .A_N(_2772_));
 sg13g2_nand2_1 _7747_ (.Y(_2774_),
    .A(_2770_),
    .B(_2773_));
 sg13g2_nand2_1 _7748_ (.Y(_2775_),
    .A(_2772_),
    .B(_0656_));
 sg13g2_nand2_1 _7749_ (.Y(_2776_),
    .A(_2774_),
    .B(_2775_));
 sg13g2_nor2_1 _7750_ (.A(_0960_),
    .B(net24),
    .Y(_2777_));
 sg13g2_a21oi_1 _7751_ (.A1(_0069_),
    .A2(net24),
    .Y(_2778_),
    .B1(_2777_));
 sg13g2_xnor2_1 _7752_ (.Y(_2779_),
    .A(net119),
    .B(_2778_));
 sg13g2_nor2b_1 _7753_ (.A(net119),
    .B_N(_2778_),
    .Y(_2780_));
 sg13g2_a21o_1 _7754_ (.A2(_2779_),
    .A1(_2776_),
    .B1(_2780_),
    .X(_2781_));
 sg13g2_nor2_1 _7755_ (.A(_0983_),
    .B(_2756_),
    .Y(_2782_));
 sg13g2_a21oi_1 _7756_ (.A1(_0070_),
    .A2(net24),
    .Y(_2783_),
    .B1(_2782_));
 sg13g2_xnor2_1 _7757_ (.Y(_2784_),
    .A(_0598_),
    .B(_2783_));
 sg13g2_nor2b_1 _7758_ (.A(_0598_),
    .B_N(_2783_),
    .Y(_2785_));
 sg13g2_a21o_1 _7759_ (.A2(_2784_),
    .A1(_2781_),
    .B1(_2785_),
    .X(_2786_));
 sg13g2_xnor2_1 _7760_ (.Y(_2787_),
    .A(_2759_),
    .B(_2786_));
 sg13g2_nand2_1 _7761_ (.Y(_2788_),
    .A(net27),
    .B(_0042_));
 sg13g2_xor2_1 _7762_ (.B(_4278_),
    .A(_4276_),
    .X(_2789_));
 sg13g2_nand3_1 _7763_ (.B(_2753_),
    .C(_2789_),
    .A(_2751_),
    .Y(_2790_));
 sg13g2_nand2_1 _7764_ (.Y(_2791_),
    .A(_4365_),
    .B(_4382_));
 sg13g2_nor3_1 _7765_ (.A(net94),
    .B(net83),
    .C(_2791_),
    .Y(_2792_));
 sg13g2_nor2_1 _7766_ (.A(_4346_),
    .B(_0942_),
    .Y(_2793_));
 sg13g2_nand4_1 _7767_ (.B(_4379_),
    .C(_0796_),
    .A(_2792_),
    .Y(_2794_),
    .D(_2793_));
 sg13g2_nand2_1 _7768_ (.Y(_2795_),
    .A(_4364_),
    .B(_0787_));
 sg13g2_nand3_1 _7769_ (.B(_4310_),
    .C(_0930_),
    .A(_2795_),
    .Y(_2796_));
 sg13g2_a21oi_1 _7770_ (.A1(_2796_),
    .A2(_4371_),
    .Y(_2797_),
    .B1(_4376_));
 sg13g2_nand2_2 _7771_ (.Y(_2798_),
    .A(_2794_),
    .B(_2797_));
 sg13g2_inv_1 _7772_ (.Y(_2799_),
    .A(_2798_));
 sg13g2_nor2_2 _7773_ (.A(net65),
    .B(_2799_),
    .Y(_2800_));
 sg13g2_nand3_1 _7774_ (.B(_2790_),
    .C(_2800_),
    .A(_2788_),
    .Y(_2801_));
 sg13g2_xnor2_1 _7775_ (.Y(_2802_),
    .A(_0052_),
    .B(_4464_));
 sg13g2_nand3b_1 _7776_ (.B(_2751_),
    .C(_2753_),
    .Y(_2803_),
    .A_N(_2802_));
 sg13g2_nand2_1 _7777_ (.Y(_2804_),
    .A(net27),
    .B(_0043_));
 sg13g2_nand2_1 _7778_ (.Y(_2805_),
    .A(_2803_),
    .B(_2804_));
 sg13g2_xnor2_1 _7779_ (.Y(_2806_),
    .A(_2800_),
    .B(_2805_));
 sg13g2_xnor2_1 _7780_ (.Y(_2807_),
    .A(_2801_),
    .B(_2806_));
 sg13g2_inv_1 _7781_ (.Y(_2808_),
    .A(_0044_));
 sg13g2_nand2_1 _7782_ (.Y(_2809_),
    .A(_2754_),
    .B(_2808_));
 sg13g2_inv_1 _7783_ (.Y(_2810_),
    .A(net125));
 sg13g2_nand2_1 _7784_ (.Y(_2811_),
    .A(_4464_),
    .B(_2810_));
 sg13g2_xnor2_1 _7785_ (.Y(_2812_),
    .A(_4412_),
    .B(_2811_));
 sg13g2_nand3_1 _7786_ (.B(_2753_),
    .C(_2812_),
    .A(_2751_),
    .Y(_2813_));
 sg13g2_nand2_1 _7787_ (.Y(_2814_),
    .A(_2809_),
    .B(_2813_));
 sg13g2_inv_1 _7788_ (.Y(_2815_),
    .A(_2800_));
 sg13g2_nand3_1 _7789_ (.B(_0760_),
    .C(_4366_),
    .A(_4302_),
    .Y(_2816_));
 sg13g2_inv_1 _7790_ (.Y(_2817_),
    .A(_4354_));
 sg13g2_a21oi_1 _7791_ (.A1(_2817_),
    .A2(net95),
    .Y(_2818_),
    .B1(_4371_));
 sg13g2_nand2_1 _7792_ (.Y(_2819_),
    .A(_2816_),
    .B(_2818_));
 sg13g2_nor2_1 _7793_ (.A(_0818_),
    .B(_2819_),
    .Y(_2820_));
 sg13g2_inv_1 _7794_ (.Y(_2821_),
    .A(_2820_));
 sg13g2_nor2_1 _7795_ (.A(_4335_),
    .B(_0933_),
    .Y(_2822_));
 sg13g2_a21oi_1 _7796_ (.A1(_2821_),
    .A2(_2822_),
    .Y(_2823_),
    .B1(_4352_));
 sg13g2_inv_1 _7797_ (.Y(_2824_),
    .A(_2823_));
 sg13g2_inv_1 _7798_ (.Y(_2825_),
    .A(_0759_));
 sg13g2_o21ai_1 _7799_ (.B1(_1002_),
    .Y(_2826_),
    .A1(_0760_),
    .A2(_2825_));
 sg13g2_nand4_1 _7800_ (.B(_4335_),
    .C(_1018_),
    .A(_2826_),
    .Y(_2827_),
    .D(_4319_));
 sg13g2_nand2_1 _7801_ (.Y(_2828_),
    .A(_2827_),
    .B(_4376_));
 sg13g2_nand3_1 _7802_ (.B(_4382_),
    .C(_4324_),
    .A(_0759_),
    .Y(_2829_));
 sg13g2_nor3_1 _7803_ (.A(net95),
    .B(_0760_),
    .C(_2829_),
    .Y(_2830_));
 sg13g2_nand3_1 _7804_ (.B(_0818_),
    .C(_4379_),
    .A(_2830_),
    .Y(_2831_));
 sg13g2_nand2_2 _7805_ (.Y(_2832_),
    .A(_2828_),
    .B(_2831_));
 sg13g2_inv_2 _7806_ (.Y(_2833_),
    .A(_2832_));
 sg13g2_a22oi_1 _7807_ (.Y(_2834_),
    .B1(_0081_),
    .B2(_2833_),
    .A2(net99),
    .A1(_2824_));
 sg13g2_nor2b_1 _7808_ (.A(_2815_),
    .B_N(_2834_),
    .Y(_2835_));
 sg13g2_nand2_2 _7809_ (.Y(_2836_),
    .A(_2814_),
    .B(_2835_));
 sg13g2_inv_1 _7810_ (.Y(_2837_),
    .A(_2835_));
 sg13g2_nand3_1 _7811_ (.B(_2813_),
    .C(_2837_),
    .A(_2809_),
    .Y(_2838_));
 sg13g2_nand2_1 _7812_ (.Y(_2839_),
    .A(_2836_),
    .B(_2838_));
 sg13g2_nand2_1 _7813_ (.Y(_2840_),
    .A(_2788_),
    .B(_2790_));
 sg13g2_a21oi_2 _7814_ (.B1(_2815_),
    .Y(_2841_),
    .A2(_2840_),
    .A1(_2805_));
 sg13g2_xnor2_1 _7815_ (.Y(_2842_),
    .A(_2839_),
    .B(_2841_));
 sg13g2_nand2_1 _7816_ (.Y(_2843_),
    .A(_2807_),
    .B(_2842_));
 sg13g2_xnor2_1 _7817_ (.Y(_2844_),
    .A(_2837_),
    .B(_2814_));
 sg13g2_nand2_1 _7818_ (.Y(_2845_),
    .A(_2841_),
    .B(_2844_));
 sg13g2_nand2_1 _7819_ (.Y(_2846_),
    .A(_2845_),
    .B(_2836_));
 sg13g2_inv_1 _7820_ (.Y(_2847_),
    .A(_0045_));
 sg13g2_nand2_1 _7821_ (.Y(_2848_),
    .A(_2755_),
    .B(_2847_));
 sg13g2_nor2_1 _7822_ (.A(net123),
    .B(_2811_),
    .Y(_2849_));
 sg13g2_xnor2_1 _7823_ (.Y(_2850_),
    .A(_4285_),
    .B(_2849_));
 sg13g2_nand3_1 _7824_ (.B(_2753_),
    .C(_2850_),
    .A(_2751_),
    .Y(_2851_));
 sg13g2_nand2_1 _7825_ (.Y(_2852_),
    .A(_2848_),
    .B(_2851_));
 sg13g2_inv_1 _7826_ (.Y(_2853_),
    .A(_0017_));
 sg13g2_nor2_1 _7827_ (.A(_2853_),
    .B(_2832_),
    .Y(_2854_));
 sg13g2_nor2_1 _7828_ (.A(net65),
    .B(_2823_),
    .Y(_2855_));
 sg13g2_a21oi_1 _7829_ (.A1(_2855_),
    .A2(_0798_),
    .Y(_2856_),
    .B1(_2833_));
 sg13g2_nor3_1 _7830_ (.A(_2799_),
    .B(_2854_),
    .C(_2856_),
    .Y(_2857_));
 sg13g2_nand2_1 _7831_ (.Y(_2858_),
    .A(_2852_),
    .B(_2857_));
 sg13g2_inv_1 _7832_ (.Y(_2859_),
    .A(_2857_));
 sg13g2_nand3_1 _7833_ (.B(_2851_),
    .C(_2859_),
    .A(_2848_),
    .Y(_2860_));
 sg13g2_buf_2 _7834_ (.A(_2860_),
    .X(_2861_));
 sg13g2_nand2_2 _7835_ (.Y(_2862_),
    .A(_2858_),
    .B(_2861_));
 sg13g2_inv_1 _7836_ (.Y(_2863_),
    .A(_2862_));
 sg13g2_nand2_1 _7837_ (.Y(_2864_),
    .A(_2846_),
    .B(_2863_));
 sg13g2_nand3_1 _7838_ (.B(_2862_),
    .C(_2836_),
    .A(_2845_),
    .Y(_2865_));
 sg13g2_nand2_1 _7839_ (.Y(_2866_),
    .A(_2864_),
    .B(_2865_));
 sg13g2_buf_2 _7840_ (.A(_2866_),
    .X(_2867_));
 sg13g2_nor2_1 _7841_ (.A(_2843_),
    .B(_2867_),
    .Y(_2868_));
 sg13g2_inv_1 _7842_ (.Y(_2869_),
    .A(_2868_));
 sg13g2_nand2_1 _7843_ (.Y(_2870_),
    .A(_2867_),
    .B(_2843_));
 sg13g2_nand2_1 _7844_ (.Y(_2871_),
    .A(_2869_),
    .B(_2870_));
 sg13g2_nand2_1 _7845_ (.Y(_2872_),
    .A(_2836_),
    .B(_2858_));
 sg13g2_inv_1 _7846_ (.Y(_2873_),
    .A(_2872_));
 sg13g2_nand2_1 _7847_ (.Y(_2874_),
    .A(_2845_),
    .B(_2873_));
 sg13g2_inv_1 _7848_ (.Y(_2875_),
    .A(net99));
 sg13g2_nor2_1 _7849_ (.A(_0942_),
    .B(_0796_),
    .Y(_2876_));
 sg13g2_a21o_1 _7850_ (.A2(_4306_),
    .A1(_2875_),
    .B1(_2876_),
    .X(_2877_));
 sg13g2_o21ai_1 _7851_ (.B1(_2824_),
    .Y(_2878_),
    .A1(net65),
    .A2(_2877_));
 sg13g2_nand2_1 _7852_ (.Y(_2879_),
    .A(_2833_),
    .B(net96));
 sg13g2_nand3_1 _7853_ (.B(_2879_),
    .C(_2798_),
    .A(_2878_),
    .Y(_2880_));
 sg13g2_nor2_1 _7854_ (.A(_4476_),
    .B(_2849_),
    .Y(_2881_));
 sg13g2_xnor2_1 _7855_ (.Y(_2882_),
    .A(_4428_),
    .B(_2881_));
 sg13g2_nand2_1 _7856_ (.Y(_2883_),
    .A(_2763_),
    .B(_2882_));
 sg13g2_nand2b_1 _7857_ (.Y(_2884_),
    .B(_2754_),
    .A_N(_0046_));
 sg13g2_nand2_1 _7858_ (.Y(_2885_),
    .A(_2883_),
    .B(_2884_));
 sg13g2_xnor2_1 _7859_ (.Y(_2886_),
    .A(_2880_),
    .B(_2885_));
 sg13g2_nand3_1 _7860_ (.B(_2886_),
    .C(_2861_),
    .A(_2874_),
    .Y(_2887_));
 sg13g2_nor2_1 _7861_ (.A(_2862_),
    .B(_2839_),
    .Y(_2888_));
 sg13g2_nand2_1 _7862_ (.Y(_2889_),
    .A(_2888_),
    .B(_2841_));
 sg13g2_inv_4 _7863_ (.A(_2886_),
    .Y(_2890_));
 sg13g2_nand2_1 _7864_ (.Y(_2891_),
    .A(_2872_),
    .B(_2861_));
 sg13g2_nand3_1 _7865_ (.B(_2890_),
    .C(_2891_),
    .A(_2889_),
    .Y(_2892_));
 sg13g2_nand2_1 _7866_ (.Y(_2893_),
    .A(_2887_),
    .B(_2892_));
 sg13g2_buf_1 _7867_ (.A(_2893_),
    .X(_2894_));
 sg13g2_nand2_1 _7868_ (.Y(_2895_),
    .A(_2871_),
    .B(net19));
 sg13g2_inv_2 _7869_ (.Y(_2896_),
    .A(_2842_));
 sg13g2_nand2_1 _7870_ (.Y(_2897_),
    .A(_2867_),
    .B(_2896_));
 sg13g2_nand3_1 _7871_ (.B(_2865_),
    .C(_2842_),
    .A(_2864_),
    .Y(_2898_));
 sg13g2_buf_1 _7872_ (.A(_2898_),
    .X(_2899_));
 sg13g2_nand2_1 _7873_ (.Y(_2900_),
    .A(_2897_),
    .B(_2899_));
 sg13g2_nand3_1 _7874_ (.B(_2890_),
    .C(_2861_),
    .A(_2874_),
    .Y(_2901_));
 sg13g2_nand3_1 _7875_ (.B(_2886_),
    .C(_2891_),
    .A(_2889_),
    .Y(_2902_));
 sg13g2_nand2_1 _7876_ (.Y(_2903_),
    .A(_2901_),
    .B(_2902_));
 sg13g2_buf_2 _7877_ (.A(_2903_),
    .X(_2904_));
 sg13g2_nand2_1 _7878_ (.Y(_2905_),
    .A(_2900_),
    .B(_2904_));
 sg13g2_nand2_1 _7879_ (.Y(_2906_),
    .A(_2881_),
    .B(net124));
 sg13g2_xnor2_1 _7880_ (.Y(_2907_),
    .A(_4427_),
    .B(_2906_));
 sg13g2_nand2b_1 _7881_ (.Y(_2908_),
    .B(net23),
    .A_N(_2907_));
 sg13g2_nand2_1 _7882_ (.Y(_2909_),
    .A(_2755_),
    .B(_1525_));
 sg13g2_xnor2_1 _7883_ (.Y(_2910_),
    .A(_0802_),
    .B(_2876_));
 sg13g2_o21ai_1 _7884_ (.B1(_2824_),
    .Y(_2911_),
    .A1(_0939_),
    .A2(_2910_));
 sg13g2_nand2_1 _7885_ (.Y(_2912_),
    .A(_4327_),
    .B(_0788_));
 sg13g2_nand2_1 _7886_ (.Y(_2913_),
    .A(_2833_),
    .B(_2912_));
 sg13g2_nand3_1 _7887_ (.B(_2913_),
    .C(_2798_),
    .A(_2911_),
    .Y(_2914_));
 sg13g2_a21oi_1 _7888_ (.A1(_2908_),
    .A2(_2909_),
    .Y(_2915_),
    .B1(_2914_));
 sg13g2_nand3_1 _7889_ (.B(_2914_),
    .C(_2909_),
    .A(_2908_),
    .Y(_2916_));
 sg13g2_nor2b_1 _7890_ (.A(_2915_),
    .B_N(_2916_),
    .Y(_2917_));
 sg13g2_inv_2 _7891_ (.Y(_2918_),
    .A(_2917_));
 sg13g2_nor2_1 _7892_ (.A(_2862_),
    .B(_2890_),
    .Y(_2919_));
 sg13g2_nand2_1 _7893_ (.Y(_2920_),
    .A(_2846_),
    .B(_2919_));
 sg13g2_a21oi_1 _7894_ (.A1(_2883_),
    .A2(_2884_),
    .Y(_2921_),
    .B1(_2880_));
 sg13g2_inv_1 _7895_ (.Y(_2922_),
    .A(_2858_));
 sg13g2_nand2_1 _7896_ (.Y(_2923_),
    .A(_2886_),
    .B(_2922_));
 sg13g2_nand2b_1 _7897_ (.Y(_2924_),
    .B(_2923_),
    .A_N(_2921_));
 sg13g2_inv_2 _7898_ (.Y(_2925_),
    .A(_2924_));
 sg13g2_nand2_1 _7899_ (.Y(_2926_),
    .A(_2920_),
    .B(_2925_));
 sg13g2_xnor2_1 _7900_ (.Y(_2927_),
    .A(_2918_),
    .B(_2926_));
 sg13g2_buf_8 _7901_ (.A(_2927_),
    .X(_2928_));
 sg13g2_nand3_1 _7902_ (.B(_2905_),
    .C(net17),
    .A(_2895_),
    .Y(_2929_));
 sg13g2_nand2_1 _7903_ (.Y(_2930_),
    .A(_2846_),
    .B(_2862_));
 sg13g2_nand3_1 _7904_ (.B(_2863_),
    .C(_2836_),
    .A(_2845_),
    .Y(_2931_));
 sg13g2_nand2_1 _7905_ (.Y(_2932_),
    .A(_2930_),
    .B(_2931_));
 sg13g2_nor2_2 _7906_ (.A(_2842_),
    .B(_2807_),
    .Y(_2933_));
 sg13g2_inv_4 _7907_ (.A(_2933_),
    .Y(_2934_));
 sg13g2_nand2_1 _7908_ (.Y(_2935_),
    .A(_2932_),
    .B(_2934_));
 sg13g2_nand2_1 _7909_ (.Y(_2936_),
    .A(_2867_),
    .B(_2933_));
 sg13g2_nand2_1 _7910_ (.Y(_2937_),
    .A(_2935_),
    .B(_2936_));
 sg13g2_nand2_1 _7911_ (.Y(_2938_),
    .A(_2937_),
    .B(_2894_));
 sg13g2_nand2_1 _7912_ (.Y(_2939_),
    .A(_2926_),
    .B(_2917_));
 sg13g2_nand3_1 _7913_ (.B(_2925_),
    .C(_2918_),
    .A(_2920_),
    .Y(_2940_));
 sg13g2_nand2_1 _7914_ (.Y(_2941_),
    .A(_2939_),
    .B(_2940_));
 sg13g2_buf_2 _7915_ (.A(_2941_),
    .X(_2942_));
 sg13g2_buf_1 _7916_ (.A(_2942_),
    .X(_2943_));
 sg13g2_nand2_1 _7917_ (.Y(_2944_),
    .A(_2904_),
    .B(_2932_));
 sg13g2_nand3_1 _7918_ (.B(_2943_),
    .C(_2944_),
    .A(_2938_),
    .Y(_2945_));
 sg13g2_o21ai_1 _7919_ (.B1(_0056_),
    .Y(_2946_),
    .A1(_4281_),
    .A2(_2906_));
 sg13g2_xnor2_1 _7920_ (.Y(_2947_),
    .A(_4434_),
    .B(_2946_));
 sg13g2_nor2_1 _7921_ (.A(_2947_),
    .B(net27),
    .Y(_2948_));
 sg13g2_a21oi_1 _7922_ (.A1(_0048_),
    .A2(net27),
    .Y(_2949_),
    .B1(_2948_));
 sg13g2_nand4_1 _7923_ (.B(_4325_),
    .C(_0802_),
    .A(_0760_),
    .Y(_2950_),
    .D(_0930_));
 sg13g2_xnor2_1 _7924_ (.Y(_2951_),
    .A(_4365_),
    .B(_0997_));
 sg13g2_nor2_1 _7925_ (.A(_2950_),
    .B(_2951_),
    .Y(_2952_));
 sg13g2_nand2_1 _7926_ (.Y(_2953_),
    .A(_2951_),
    .B(_2950_));
 sg13g2_nand3b_1 _7927_ (.B(_2824_),
    .C(_2953_),
    .Y(_2954_),
    .A_N(_2952_));
 sg13g2_xnor2_1 _7928_ (.Y(_2955_),
    .A(_0806_),
    .B(_0788_));
 sg13g2_nand2_1 _7929_ (.Y(_2956_),
    .A(_2833_),
    .B(_2955_));
 sg13g2_nand3_1 _7930_ (.B(_2800_),
    .C(_2956_),
    .A(_2954_),
    .Y(_2957_));
 sg13g2_nand2b_1 _7931_ (.Y(_2958_),
    .B(_2957_),
    .A_N(_2949_));
 sg13g2_nand2b_1 _7932_ (.Y(_2959_),
    .B(_2949_),
    .A_N(_2957_));
 sg13g2_nand2_1 _7933_ (.Y(_2960_),
    .A(_2958_),
    .B(_2959_));
 sg13g2_nor3_1 _7934_ (.A(_2890_),
    .B(_2891_),
    .C(_2918_),
    .Y(_2961_));
 sg13g2_a21oi_1 _7935_ (.A1(_2921_),
    .A2(_2916_),
    .Y(_2962_),
    .B1(_2915_));
 sg13g2_nor2b_1 _7936_ (.A(_2961_),
    .B_N(_2962_),
    .Y(_2963_));
 sg13g2_nand4_1 _7937_ (.B(_2917_),
    .C(_2886_),
    .A(_2888_),
    .Y(_2964_),
    .D(_2841_));
 sg13g2_nand2_1 _7938_ (.Y(_2965_),
    .A(_2963_),
    .B(_2964_));
 sg13g2_xnor2_1 _7939_ (.Y(_2966_),
    .A(_2960_),
    .B(_2965_));
 sg13g2_buf_1 _7940_ (.A(_2966_),
    .X(_2967_));
 sg13g2_xor2_1 _7941_ (.B(_2952_),
    .A(_0999_),
    .X(_2968_));
 sg13g2_a21oi_1 _7942_ (.A1(_2855_),
    .A2(_2968_),
    .Y(_2969_),
    .B1(_2833_));
 sg13g2_nor2_1 _7943_ (.A(_0806_),
    .B(_2912_),
    .Y(_2970_));
 sg13g2_nand2_1 _7944_ (.Y(_2971_),
    .A(_4310_),
    .B(_0058_));
 sg13g2_xnor2_1 _7945_ (.Y(_2972_),
    .A(_4337_),
    .B(_2971_));
 sg13g2_nor2b_1 _7946_ (.A(_2970_),
    .B_N(_2972_),
    .Y(_2973_));
 sg13g2_nor2b_1 _7947_ (.A(_2972_),
    .B_N(_2970_),
    .Y(_2974_));
 sg13g2_o21ai_1 _7948_ (.B1(_2833_),
    .Y(_2975_),
    .A1(_2973_),
    .A2(_2974_));
 sg13g2_nand3b_1 _7949_ (.B(_2798_),
    .C(_2975_),
    .Y(_2976_),
    .A_N(_2969_));
 sg13g2_nand3_1 _7950_ (.B(_4282_),
    .C(_4399_),
    .A(_2906_),
    .Y(_2977_));
 sg13g2_nand2_1 _7951_ (.Y(_2978_),
    .A(_2977_),
    .B(_4289_));
 sg13g2_nand2b_1 _7952_ (.Y(_2979_),
    .B(_4443_),
    .A_N(_2977_));
 sg13g2_a21oi_1 _7953_ (.A1(_2978_),
    .A2(_2979_),
    .Y(_2980_),
    .B1(net27));
 sg13g2_a21oi_1 _7954_ (.A1(_0049_),
    .A2(net24),
    .Y(_2981_),
    .B1(_2980_));
 sg13g2_inv_1 _7955_ (.Y(_2982_),
    .A(_2981_));
 sg13g2_nor2_1 _7956_ (.A(_2976_),
    .B(_2982_),
    .Y(_2983_));
 sg13g2_nand2_1 _7957_ (.Y(_2984_),
    .A(_2982_),
    .B(_2976_));
 sg13g2_inv_1 _7958_ (.Y(_2985_),
    .A(_2984_));
 sg13g2_nor2_2 _7959_ (.A(_2983_),
    .B(_2985_),
    .Y(_2986_));
 sg13g2_nor2_1 _7960_ (.A(_2918_),
    .B(_2960_),
    .Y(_2987_));
 sg13g2_nand2_1 _7961_ (.Y(_2988_),
    .A(_2958_),
    .B(_2915_));
 sg13g2_nand2_1 _7962_ (.Y(_2989_),
    .A(_2988_),
    .B(_2959_));
 sg13g2_a21oi_1 _7963_ (.A1(_2987_),
    .A2(_2924_),
    .Y(_2990_),
    .B1(_2989_));
 sg13g2_nand3_1 _7964_ (.B(_2846_),
    .C(_2919_),
    .A(_2987_),
    .Y(_2991_));
 sg13g2_nand2_1 _7965_ (.Y(_2992_),
    .A(_2990_),
    .B(_2991_));
 sg13g2_xnor2_1 _7966_ (.Y(_2993_),
    .A(_2986_),
    .B(_2992_));
 sg13g2_buf_8 _7967_ (.A(_2993_),
    .X(_2994_));
 sg13g2_nor2_1 _7968_ (.A(net16),
    .B(_2994_),
    .Y(_2995_));
 sg13g2_nand3_1 _7969_ (.B(_2945_),
    .C(_2995_),
    .A(_2929_),
    .Y(_2996_));
 sg13g2_nand2_1 _7970_ (.Y(_2997_),
    .A(_2773_),
    .B(_2775_));
 sg13g2_xnor2_1 _7971_ (.Y(_2998_),
    .A(_2997_),
    .B(_2770_));
 sg13g2_inv_2 _7972_ (.Y(_2999_),
    .A(_2998_));
 sg13g2_buf_1 _7973_ (.A(_2999_),
    .X(_3000_));
 sg13g2_nor2_1 _7974_ (.A(_2933_),
    .B(_2867_),
    .Y(_3001_));
 sg13g2_nor2_1 _7975_ (.A(_2904_),
    .B(_3001_),
    .Y(_3002_));
 sg13g2_nor2_1 _7976_ (.A(_2942_),
    .B(_3002_),
    .Y(_3003_));
 sg13g2_inv_1 _7977_ (.Y(_3004_),
    .A(_3003_));
 sg13g2_nand2_1 _7978_ (.Y(_3005_),
    .A(_2897_),
    .B(_2904_));
 sg13g2_nand2_1 _7979_ (.Y(_3006_),
    .A(_2942_),
    .B(_3005_));
 sg13g2_nand2_1 _7980_ (.Y(_3007_),
    .A(_3004_),
    .B(_3006_));
 sg13g2_nand2_1 _7981_ (.Y(_3008_),
    .A(_3007_),
    .B(_2994_));
 sg13g2_inv_2 _7982_ (.Y(_3009_),
    .A(_3008_));
 sg13g2_nor2_1 _7983_ (.A(net20),
    .B(_3009_),
    .Y(_3010_));
 sg13g2_nand2_1 _7984_ (.Y(_3011_),
    .A(_2893_),
    .B(_2867_));
 sg13g2_nand3_1 _7985_ (.B(_2900_),
    .C(_3011_),
    .A(_2927_),
    .Y(_3012_));
 sg13g2_nand3_1 _7986_ (.B(_2942_),
    .C(_2944_),
    .A(_2937_),
    .Y(_3013_));
 sg13g2_nand2_1 _7987_ (.Y(_3014_),
    .A(_3012_),
    .B(_3013_));
 sg13g2_xor2_1 _7988_ (.B(_2992_),
    .A(_2986_),
    .X(_3015_));
 sg13g2_nand3_1 _7989_ (.B(_3015_),
    .C(net16),
    .A(_3014_),
    .Y(_3016_));
 sg13g2_nand3_1 _7990_ (.B(_3010_),
    .C(_3016_),
    .A(_2996_),
    .Y(_3017_));
 sg13g2_a21oi_1 _7991_ (.A1(_2938_),
    .A2(_2942_),
    .Y(_3018_),
    .B1(net16));
 sg13g2_nand2_1 _7992_ (.Y(_3019_),
    .A(_2868_),
    .B(net19));
 sg13g2_nand3_1 _7993_ (.B(_2927_),
    .C(_3019_),
    .A(_2905_),
    .Y(_3020_));
 sg13g2_nand2_1 _7994_ (.Y(_3021_),
    .A(_3018_),
    .B(_3020_));
 sg13g2_nand2_1 _7995_ (.Y(_3022_),
    .A(_3014_),
    .B(net16));
 sg13g2_nor2_1 _7996_ (.A(_2998_),
    .B(_2994_),
    .Y(_3023_));
 sg13g2_buf_2 _7997_ (.A(_3023_),
    .X(_3024_));
 sg13g2_nand3_1 _7998_ (.B(_3022_),
    .C(_3024_),
    .A(_3021_),
    .Y(_3025_));
 sg13g2_xor2_1 _7999_ (.B(_2776_),
    .A(_2779_),
    .X(_3026_));
 sg13g2_buf_1 _8000_ (.A(_3026_),
    .X(_3027_));
 sg13g2_inv_1 _8001_ (.Y(_3028_),
    .A(net18));
 sg13g2_a21oi_1 _8002_ (.A1(_3017_),
    .A2(_3025_),
    .Y(_3029_),
    .B1(_3028_));
 sg13g2_nand2_1 _8003_ (.Y(_3030_),
    .A(_3021_),
    .B(_3022_));
 sg13g2_nor2_2 _8004_ (.A(_2999_),
    .B(_2994_),
    .Y(_3031_));
 sg13g2_a21oi_1 _8005_ (.A1(_3030_),
    .A2(_3031_),
    .Y(_3032_),
    .B1(net18));
 sg13g2_nor2_1 _8006_ (.A(net19),
    .B(_2942_),
    .Y(_3033_));
 sg13g2_nand3_1 _8007_ (.B(_2868_),
    .C(_3033_),
    .A(_2994_),
    .Y(_3034_));
 sg13g2_inv_1 _8008_ (.Y(_3035_),
    .A(_3034_));
 sg13g2_a21oi_1 _8009_ (.A1(_3014_),
    .A2(_3024_),
    .Y(_3036_),
    .B1(_3035_));
 sg13g2_nand2_1 _8010_ (.Y(_3037_),
    .A(_3032_),
    .B(_3036_));
 sg13g2_xnor2_1 _8011_ (.Y(_3038_),
    .A(_2784_),
    .B(_2781_));
 sg13g2_buf_2 _8012_ (.A(_3038_),
    .X(_3039_));
 sg13g2_nand2_1 _8013_ (.Y(_3040_),
    .A(_3037_),
    .B(_3039_));
 sg13g2_nor2_1 _8014_ (.A(_3029_),
    .B(_3040_),
    .Y(_3041_));
 sg13g2_nor2_1 _8015_ (.A(_2787_),
    .B(_3041_),
    .Y(_3042_));
 sg13g2_nand2_1 _8016_ (.Y(_3043_),
    .A(_2899_),
    .B(_2894_));
 sg13g2_nor2b_1 _8017_ (.A(_3043_),
    .B_N(_2936_),
    .Y(_3044_));
 sg13g2_inv_1 _8018_ (.Y(_3045_),
    .A(_3044_));
 sg13g2_nor2_1 _8019_ (.A(_2842_),
    .B(_2932_),
    .Y(_3046_));
 sg13g2_nor2_1 _8020_ (.A(_2893_),
    .B(_3046_),
    .Y(_3047_));
 sg13g2_nor2_1 _8021_ (.A(_3047_),
    .B(_2927_),
    .Y(_3048_));
 sg13g2_nand2_1 _8022_ (.Y(_3049_),
    .A(_3045_),
    .B(_3048_));
 sg13g2_nor2_1 _8023_ (.A(_2934_),
    .B(_2932_),
    .Y(_3050_));
 sg13g2_nor2_1 _8024_ (.A(net19),
    .B(_3050_),
    .Y(_3051_));
 sg13g2_nand2_1 _8025_ (.Y(_3052_),
    .A(_3051_),
    .B(_2899_));
 sg13g2_nand2_1 _8026_ (.Y(_3053_),
    .A(_3003_),
    .B(_3052_));
 sg13g2_nand2_1 _8027_ (.Y(_3054_),
    .A(_3049_),
    .B(_3053_));
 sg13g2_nand2_1 _8028_ (.Y(_3055_),
    .A(_3054_),
    .B(_2999_));
 sg13g2_nand3_1 _8029_ (.B(net19),
    .C(_2897_),
    .A(_2869_),
    .Y(_3056_));
 sg13g2_nand2_1 _8030_ (.Y(_3057_),
    .A(_3056_),
    .B(net15));
 sg13g2_nand2_1 _8031_ (.Y(_3058_),
    .A(_2935_),
    .B(_2904_));
 sg13g2_nand2_1 _8032_ (.Y(_3059_),
    .A(net17),
    .B(_3058_));
 sg13g2_nand2_1 _8033_ (.Y(_3060_),
    .A(_3057_),
    .B(_3059_));
 sg13g2_nand2_1 _8034_ (.Y(_3061_),
    .A(_3060_),
    .B(_3031_));
 sg13g2_nand2_1 _8035_ (.Y(_3062_),
    .A(_3055_),
    .B(_3061_));
 sg13g2_nand2_1 _8036_ (.Y(_3063_),
    .A(_3062_),
    .B(net16));
 sg13g2_nand2_1 _8037_ (.Y(_3064_),
    .A(_3063_),
    .B(_3008_));
 sg13g2_nand2_1 _8038_ (.Y(_3065_),
    .A(_3064_),
    .B(_3028_));
 sg13g2_nand2_1 _8039_ (.Y(_3066_),
    .A(_3002_),
    .B(_2936_));
 sg13g2_nand2_1 _8040_ (.Y(_3067_),
    .A(_3048_),
    .B(_3066_));
 sg13g2_nand2_1 _8041_ (.Y(_3068_),
    .A(_3047_),
    .B(_2899_));
 sg13g2_nand2_1 _8042_ (.Y(_3069_),
    .A(_3003_),
    .B(_3068_));
 sg13g2_nand2_1 _8043_ (.Y(_3070_),
    .A(_3067_),
    .B(_3069_));
 sg13g2_nand2_1 _8044_ (.Y(_3071_),
    .A(_3070_),
    .B(_3015_));
 sg13g2_nor2_1 _8045_ (.A(_2904_),
    .B(_2937_),
    .Y(_3072_));
 sg13g2_nand2_1 _8046_ (.Y(_3073_),
    .A(_3072_),
    .B(_2928_));
 sg13g2_nor2_1 _8047_ (.A(net19),
    .B(_2900_),
    .Y(_3074_));
 sg13g2_nand2_1 _8048_ (.Y(_3075_),
    .A(_3074_),
    .B(net15));
 sg13g2_nand3_1 _8049_ (.B(_3075_),
    .C(_2994_),
    .A(_3073_),
    .Y(_3076_));
 sg13g2_nand2_1 _8050_ (.Y(_3077_),
    .A(_3071_),
    .B(_3076_));
 sg13g2_nor2_1 _8051_ (.A(net20),
    .B(_2995_),
    .Y(_3078_));
 sg13g2_nand2_1 _8052_ (.Y(_3079_),
    .A(_3077_),
    .B(_3078_));
 sg13g2_nand3_1 _8053_ (.B(_3051_),
    .C(_2899_),
    .A(_2928_),
    .Y(_3080_));
 sg13g2_nand2_1 _8054_ (.Y(_3081_),
    .A(_3044_),
    .B(net15));
 sg13g2_nand3_1 _8055_ (.B(_3081_),
    .C(net16),
    .A(_3080_),
    .Y(_3082_));
 sg13g2_nand2b_1 _8056_ (.Y(_3083_),
    .B(_3024_),
    .A_N(_3082_));
 sg13g2_nand2_1 _8057_ (.Y(_3084_),
    .A(_3079_),
    .B(_3083_));
 sg13g2_nand2_1 _8058_ (.Y(_3085_),
    .A(_3084_),
    .B(_3027_));
 sg13g2_inv_1 _8059_ (.Y(_3086_),
    .A(_2996_));
 sg13g2_a21oi_1 _8060_ (.A1(_3009_),
    .A2(_3000_),
    .Y(_3087_),
    .B1(_3086_));
 sg13g2_nand3_1 _8061_ (.B(_3085_),
    .C(_3087_),
    .A(_3065_),
    .Y(_3088_));
 sg13g2_inv_1 _8062_ (.Y(_3089_),
    .A(_3039_));
 sg13g2_nand2_1 _8063_ (.Y(_3090_),
    .A(_3088_),
    .B(_3089_));
 sg13g2_nand2_1 _8064_ (.Y(_3091_),
    .A(_3042_),
    .B(_3090_));
 sg13g2_nor2_1 _8065_ (.A(_3011_),
    .B(net17),
    .Y(_3092_));
 sg13g2_nor3_1 _8066_ (.A(net19),
    .B(net15),
    .C(_2871_),
    .Y(_3093_));
 sg13g2_nor3_1 _8067_ (.A(_3015_),
    .B(_3092_),
    .C(_3093_),
    .Y(_3094_));
 sg13g2_a21oi_1 _8068_ (.A1(_3094_),
    .A2(_3000_),
    .Y(_3095_),
    .B1(_3028_));
 sg13g2_nand2_1 _8069_ (.Y(_3096_),
    .A(_3071_),
    .B(_3034_));
 sg13g2_nand2_1 _8070_ (.Y(_3097_),
    .A(_3096_),
    .B(_2998_));
 sg13g2_nand2_1 _8071_ (.Y(_3098_),
    .A(_3072_),
    .B(net15));
 sg13g2_nand2_1 _8072_ (.Y(_3099_),
    .A(_3074_),
    .B(net17));
 sg13g2_nand3_1 _8073_ (.B(_3099_),
    .C(_2967_),
    .A(_3098_),
    .Y(_3100_));
 sg13g2_inv_2 _8074_ (.Y(_3101_),
    .A(_2967_));
 sg13g2_nand3_1 _8075_ (.B(_3081_),
    .C(_3101_),
    .A(_3080_),
    .Y(_3102_));
 sg13g2_nand2_1 _8076_ (.Y(_3103_),
    .A(_3100_),
    .B(_3102_));
 sg13g2_nand2_1 _8077_ (.Y(_3104_),
    .A(_3103_),
    .B(_3024_));
 sg13g2_nand3_1 _8078_ (.B(_3097_),
    .C(_3104_),
    .A(_3095_),
    .Y(_3105_));
 sg13g2_nand2b_1 _8079_ (.Y(_3106_),
    .B(_3033_),
    .A_N(_2937_));
 sg13g2_nand3_1 _8080_ (.B(_3081_),
    .C(_3101_),
    .A(_3106_),
    .Y(_3107_));
 sg13g2_nand2_1 _8081_ (.Y(_3108_),
    .A(_3100_),
    .B(_3107_));
 sg13g2_nand2_1 _8082_ (.Y(_3109_),
    .A(_3108_),
    .B(_3031_));
 sg13g2_nand3_1 _8083_ (.B(_3019_),
    .C(_3058_),
    .A(net17),
    .Y(_3110_));
 sg13g2_o21ai_1 _8084_ (.B1(_2943_),
    .Y(_3111_),
    .A1(_2904_),
    .A2(_3050_));
 sg13g2_nand2_1 _8085_ (.Y(_3112_),
    .A(_3110_),
    .B(_3111_));
 sg13g2_nand2_1 _8086_ (.Y(_3113_),
    .A(_3112_),
    .B(_3101_));
 sg13g2_nand2_1 _8087_ (.Y(_3114_),
    .A(_3113_),
    .B(_3082_));
 sg13g2_nand2_1 _8088_ (.Y(_3115_),
    .A(_3114_),
    .B(_3024_));
 sg13g2_nor2_1 _8089_ (.A(net18),
    .B(_3094_),
    .Y(_3116_));
 sg13g2_nand3_1 _8090_ (.B(_3115_),
    .C(_3116_),
    .A(_3109_),
    .Y(_3117_));
 sg13g2_nand3_1 _8091_ (.B(_3117_),
    .C(_3089_),
    .A(_3105_),
    .Y(_3118_));
 sg13g2_nor2_1 _8092_ (.A(net15),
    .B(_3005_),
    .Y(_3119_));
 sg13g2_a21oi_1 _8093_ (.A1(net15),
    .A2(_3002_),
    .Y(_3120_),
    .B1(_3119_));
 sg13g2_nand2_1 _8094_ (.Y(_3121_),
    .A(_3120_),
    .B(net20));
 sg13g2_nand3b_1 _8095_ (.B(net15),
    .C(net19),
    .Y(_3122_),
    .A_N(_2870_));
 sg13g2_nand2b_1 _8096_ (.Y(_3123_),
    .B(net17),
    .A_N(_2944_));
 sg13g2_nand3_1 _8097_ (.B(_2998_),
    .C(_3123_),
    .A(_3122_),
    .Y(_3124_));
 sg13g2_nor2_1 _8098_ (.A(net18),
    .B(_2994_),
    .Y(_3125_));
 sg13g2_nand3_1 _8099_ (.B(_3124_),
    .C(_3125_),
    .A(_3121_),
    .Y(_3126_));
 sg13g2_nand2_1 _8100_ (.Y(_3127_),
    .A(_3101_),
    .B(net20));
 sg13g2_nor2_1 _8101_ (.A(_2934_),
    .B(_3092_),
    .Y(_3128_));
 sg13g2_a21oi_1 _8102_ (.A1(_3127_),
    .A2(_3128_),
    .Y(_3129_),
    .B1(_3028_));
 sg13g2_nand2_1 _8103_ (.Y(_3130_),
    .A(_3092_),
    .B(_2896_));
 sg13g2_a21oi_1 _8104_ (.A1(_3130_),
    .A2(_3123_),
    .Y(_3131_),
    .B1(_2994_));
 sg13g2_nand2_1 _8105_ (.Y(_3132_),
    .A(_3129_),
    .B(_3131_));
 sg13g2_nand3_1 _8106_ (.B(_3132_),
    .C(_3034_),
    .A(_3126_),
    .Y(_3133_));
 sg13g2_inv_1 _8107_ (.Y(_3134_),
    .A(_2787_));
 sg13g2_a21oi_1 _8108_ (.A1(_3133_),
    .A2(_3039_),
    .Y(_3135_),
    .B1(_3134_));
 sg13g2_xnor2_1 _8109_ (.Y(_3136_),
    .A(_0553_),
    .B(_0611_));
 sg13g2_buf_1 _8110_ (.A(_3136_),
    .X(_3137_));
 sg13g2_inv_1 _8111_ (.Y(_3138_),
    .A(_3137_));
 sg13g2_buf_1 _8112_ (.A(net24),
    .X(_3139_));
 sg13g2_nor2_1 _8113_ (.A(_0406_),
    .B(net22),
    .Y(_3140_));
 sg13g2_a21oi_1 _8114_ (.A1(net111),
    .A2(net22),
    .Y(_3141_),
    .B1(_3140_));
 sg13g2_xnor2_1 _8115_ (.Y(_3142_),
    .A(_3138_),
    .B(_3141_));
 sg13g2_nand2_1 _8116_ (.Y(_3143_),
    .A(_2786_),
    .B(_2759_));
 sg13g2_nand2_1 _8117_ (.Y(_3144_),
    .A(_2758_),
    .B(_0553_));
 sg13g2_nand2_1 _8118_ (.Y(_3145_),
    .A(_3143_),
    .B(_3144_));
 sg13g2_xnor2_1 _8119_ (.Y(_3146_),
    .A(_3142_),
    .B(_3145_));
 sg13g2_inv_1 _8120_ (.Y(_3147_),
    .A(_3146_));
 sg13g2_a21oi_1 _8121_ (.A1(_3118_),
    .A2(_3135_),
    .Y(_3148_),
    .B1(_3147_));
 sg13g2_nand2_2 _8122_ (.Y(_3149_),
    .A(_3091_),
    .B(_3148_));
 sg13g2_nand2_1 _8123_ (.Y(_3150_),
    .A(_2996_),
    .B(_3016_));
 sg13g2_nand2_1 _8124_ (.Y(_3151_),
    .A(_3150_),
    .B(net20));
 sg13g2_nand2_1 _8125_ (.Y(_3152_),
    .A(_3032_),
    .B(_3151_));
 sg13g2_nand2_1 _8126_ (.Y(_3153_),
    .A(_3030_),
    .B(_3024_));
 sg13g2_a21oi_1 _8127_ (.A1(_3014_),
    .A2(_3031_),
    .Y(_3154_),
    .B1(_3028_));
 sg13g2_a21oi_1 _8128_ (.A1(_3153_),
    .A2(_3154_),
    .Y(_3155_),
    .B1(_3089_));
 sg13g2_nand2_1 _8129_ (.Y(_3156_),
    .A(_3152_),
    .B(_3155_));
 sg13g2_nand2_1 _8130_ (.Y(_3157_),
    .A(_3103_),
    .B(_3031_));
 sg13g2_a21oi_1 _8131_ (.A1(_3070_),
    .A2(_3024_),
    .Y(_3158_),
    .B1(net18));
 sg13g2_a21oi_1 _8132_ (.A1(_3157_),
    .A2(_3158_),
    .Y(_3159_),
    .B1(_3039_));
 sg13g2_nand2_1 _8133_ (.Y(_3160_),
    .A(_3108_),
    .B(_3024_));
 sg13g2_nand2_1 _8134_ (.Y(_3161_),
    .A(_3114_),
    .B(_3031_));
 sg13g2_nand3_1 _8135_ (.B(_3161_),
    .C(_3027_),
    .A(_3160_),
    .Y(_3162_));
 sg13g2_nand2_1 _8136_ (.Y(_3163_),
    .A(_3159_),
    .B(_3162_));
 sg13g2_nor2b_1 _8137_ (.A(_3134_),
    .B_N(_3076_),
    .Y(_3164_));
 sg13g2_nand3_1 _8138_ (.B(_3163_),
    .C(_3164_),
    .A(_3156_),
    .Y(_3165_));
 sg13g2_o21ai_1 _8139_ (.B1(_3128_),
    .Y(_3166_),
    .A1(net16),
    .A2(net20));
 sg13g2_a22oi_1 _8140_ (.Y(_3167_),
    .B1(_3166_),
    .B2(_3131_),
    .A2(_3015_),
    .A1(net18));
 sg13g2_a21oi_1 _8141_ (.A1(net17),
    .A2(_3051_),
    .Y(_3168_),
    .B1(_2999_));
 sg13g2_o21ai_1 _8142_ (.B1(_3168_),
    .Y(_3169_),
    .A1(net17),
    .A2(_3043_));
 sg13g2_nand2_1 _8143_ (.Y(_3170_),
    .A(_3033_),
    .B(_2870_));
 sg13g2_nand3_1 _8144_ (.B(_3122_),
    .C(net20),
    .A(_3170_),
    .Y(_3171_));
 sg13g2_nand3_1 _8145_ (.B(_3171_),
    .C(_3101_),
    .A(_3169_),
    .Y(_3172_));
 sg13g2_nand2_1 _8146_ (.Y(_3173_),
    .A(_3120_),
    .B(_2998_));
 sg13g2_nand3_1 _8147_ (.B(net20),
    .C(_3123_),
    .A(_3122_),
    .Y(_3174_));
 sg13g2_nand3_1 _8148_ (.B(_3174_),
    .C(net16),
    .A(_3173_),
    .Y(_3175_));
 sg13g2_nand3_1 _8149_ (.B(_3175_),
    .C(net18),
    .A(_3172_),
    .Y(_3176_));
 sg13g2_nand2b_1 _8150_ (.Y(_3177_),
    .B(_3176_),
    .A_N(_3167_));
 sg13g2_nor2_1 _8151_ (.A(_3009_),
    .B(_2787_),
    .Y(_3178_));
 sg13g2_a21oi_1 _8152_ (.A1(_3177_),
    .A2(_3178_),
    .Y(_3179_),
    .B1(_3146_));
 sg13g2_a21oi_1 _8153_ (.A1(_4310_),
    .A2(_0942_),
    .Y(_3180_),
    .B1(_4370_));
 sg13g2_xnor2_1 _8154_ (.Y(_3181_),
    .A(_0034_),
    .B(_3180_));
 sg13g2_a21oi_1 _8155_ (.A1(_4310_),
    .A2(_0942_),
    .Y(_3182_),
    .B1(_4337_));
 sg13g2_xnor2_1 _8156_ (.Y(_3183_),
    .A(_0059_),
    .B(_3182_));
 sg13g2_nand2_1 _8157_ (.Y(_3184_),
    .A(_2973_),
    .B(_3183_));
 sg13g2_xor2_1 _8158_ (.B(_3184_),
    .A(_3181_),
    .X(_3185_));
 sg13g2_xnor2_1 _8159_ (.Y(_3186_),
    .A(_4341_),
    .B(_2819_));
 sg13g2_or2_1 _8160_ (.X(_3187_),
    .B(_2952_),
    .A(_0999_));
 sg13g2_a21oi_1 _8161_ (.A1(_0997_),
    .A2(_4383_),
    .Y(_3188_),
    .B1(_0996_));
 sg13g2_xnor2_1 _8162_ (.Y(_3189_),
    .A(_1018_),
    .B(_3188_));
 sg13g2_nand2_1 _8163_ (.Y(_3190_),
    .A(_3187_),
    .B(_3189_));
 sg13g2_xnor2_1 _8164_ (.Y(_3191_),
    .A(_3186_),
    .B(_3190_));
 sg13g2_nand2_1 _8165_ (.Y(_3192_),
    .A(_3191_),
    .B(_2855_));
 sg13g2_a21oi_1 _8166_ (.A1(_3192_),
    .A2(_2832_),
    .Y(_3193_),
    .B1(_2799_));
 sg13g2_o21ai_1 _8167_ (.B1(_3193_),
    .Y(_3194_),
    .A1(_2832_),
    .A2(_3185_));
 sg13g2_o21ai_1 _8168_ (.B1(_4288_),
    .Y(_3195_),
    .A1(_4461_),
    .A2(_2978_));
 sg13g2_nor2_1 _8169_ (.A(_3195_),
    .B(net22),
    .Y(_3196_));
 sg13g2_a21oi_1 _8170_ (.A1(\vgademo.plane_u[21] ),
    .A2(net22),
    .Y(_3197_),
    .B1(_3196_));
 sg13g2_xor2_1 _8171_ (.B(_3197_),
    .A(_3194_),
    .X(_3198_));
 sg13g2_nand2_1 _8172_ (.Y(_3199_),
    .A(_2992_),
    .B(_2986_));
 sg13g2_xor2_1 _8173_ (.B(_3187_),
    .A(_3189_),
    .X(_3200_));
 sg13g2_o21ai_1 _8174_ (.B1(_2824_),
    .Y(_3201_),
    .A1(_0939_),
    .A2(_3200_));
 sg13g2_nor2_1 _8175_ (.A(_3183_),
    .B(_2973_),
    .Y(_3202_));
 sg13g2_inv_1 _8176_ (.Y(_3203_),
    .A(_3184_));
 sg13g2_o21ai_1 _8177_ (.B1(_2833_),
    .Y(_3204_),
    .A1(_3202_),
    .A2(_3203_));
 sg13g2_nand3_1 _8178_ (.B(_2798_),
    .C(_3204_),
    .A(_3201_),
    .Y(_3205_));
 sg13g2_xnor2_1 _8179_ (.Y(_3206_),
    .A(_4442_),
    .B(_2978_));
 sg13g2_nor2_1 _8180_ (.A(_3206_),
    .B(net22),
    .Y(_3207_));
 sg13g2_a21oi_1 _8181_ (.A1(_1570_),
    .A2(net22),
    .Y(_3208_),
    .B1(_3207_));
 sg13g2_nor2_1 _8182_ (.A(_3205_),
    .B(_3208_),
    .Y(_3209_));
 sg13g2_nor2_1 _8183_ (.A(_3209_),
    .B(_2983_),
    .Y(_3210_));
 sg13g2_and2_1 _8184_ (.A(_3208_),
    .B(_3205_),
    .X(_3211_));
 sg13g2_a21oi_1 _8185_ (.A1(_3199_),
    .A2(_3210_),
    .Y(_3212_),
    .B1(_3211_));
 sg13g2_xnor2_1 _8186_ (.Y(_3213_),
    .A(_3198_),
    .B(_3212_));
 sg13g2_nor2_1 _8187_ (.A(_3209_),
    .B(_3211_),
    .Y(_3214_));
 sg13g2_nand2b_1 _8188_ (.Y(_3215_),
    .B(_2965_),
    .A_N(_2960_));
 sg13g2_nor2b_1 _8189_ (.A(_2983_),
    .B_N(_2959_),
    .Y(_3216_));
 sg13g2_a21oi_1 _8190_ (.A1(_3215_),
    .A2(_3216_),
    .Y(_3217_),
    .B1(_2985_));
 sg13g2_xor2_1 _8191_ (.B(_3217_),
    .A(_3214_),
    .X(_3218_));
 sg13g2_nand2_1 _8192_ (.Y(_3219_),
    .A(_3213_),
    .B(_3218_));
 sg13g2_a21oi_2 _8193_ (.B1(_3219_),
    .Y(_3220_),
    .A2(_3179_),
    .A1(_3165_));
 sg13g2_nand2_1 _8194_ (.Y(_3221_),
    .A(_3149_),
    .B(_3220_));
 sg13g2_nand2_1 _8195_ (.Y(_3222_),
    .A(_0599_),
    .B(_0889_));
 sg13g2_inv_1 _8196_ (.Y(_3223_),
    .A(_3222_));
 sg13g2_nor2_1 _8197_ (.A(net100),
    .B(_0889_),
    .Y(_3224_));
 sg13g2_inv_1 _8198_ (.Y(_3225_),
    .A(_0885_));
 sg13g2_a22oi_1 _8199_ (.Y(_3226_),
    .B1(_0660_),
    .B2(_0885_),
    .A2(_0881_),
    .A1(_0656_));
 sg13g2_inv_1 _8200_ (.Y(_3227_),
    .A(_0881_));
 sg13g2_inv_1 _8201_ (.Y(_3228_),
    .A(_0877_));
 sg13g2_nand2_1 _8202_ (.Y(_3229_),
    .A(_3228_),
    .B(_0590_));
 sg13g2_nor2_1 _8203_ (.A(_0590_),
    .B(_3228_),
    .Y(_3230_));
 sg13g2_a21oi_1 _8204_ (.A1(_2766_),
    .A2(_3229_),
    .Y(_3231_),
    .B1(_3230_));
 sg13g2_a21o_1 _8205_ (.A2(_3227_),
    .A1(_0588_),
    .B1(_3231_),
    .X(_3232_));
 sg13g2_a22oi_1 _8206_ (.Y(_3233_),
    .B1(_3226_),
    .B2(_3232_),
    .A2(_3225_),
    .A1(net119));
 sg13g2_o21ai_1 _8207_ (.B1(_3233_),
    .Y(_3234_),
    .A1(_3223_),
    .A2(_3224_));
 sg13g2_a22oi_1 _8208_ (.Y(_3235_),
    .B1(_0619_),
    .B2(_0889_),
    .A2(_0893_),
    .A1(_0553_));
 sg13g2_inv_1 _8209_ (.Y(_3236_),
    .A(_0893_));
 sg13g2_a22oi_1 _8210_ (.Y(_3237_),
    .B1(_0072_),
    .B2(_3137_),
    .A2(_3236_),
    .A1(_0554_));
 sg13g2_o21ai_1 _8211_ (.B1(_3237_),
    .Y(_3238_),
    .A1(_0072_),
    .A2(_3137_));
 sg13g2_a21o_1 _8212_ (.A2(_3235_),
    .A1(_3234_),
    .B1(_3238_),
    .X(_3239_));
 sg13g2_nor2_1 _8213_ (.A(_0611_),
    .B(_0554_),
    .Y(_3240_));
 sg13g2_inv_1 _8214_ (.Y(_3241_),
    .A(_3240_));
 sg13g2_a22oi_1 _8215_ (.Y(_3242_),
    .B1(net111),
    .B2(_3138_),
    .A2(_3241_),
    .A1(_0901_));
 sg13g2_nor2_1 _8216_ (.A(net100),
    .B(_0611_),
    .Y(_3243_));
 sg13g2_a21oi_2 _8217_ (.B1(_3243_),
    .Y(_3244_),
    .A2(net100),
    .A1(_3137_));
 sg13g2_xor2_1 _8218_ (.B(_3244_),
    .A(_0072_),
    .X(_3245_));
 sg13g2_nand2_1 _8219_ (.Y(_3246_),
    .A(net100),
    .B(_0553_));
 sg13g2_nand2_2 _8220_ (.Y(_3247_),
    .A(_0620_),
    .B(_3246_));
 sg13g2_xor2_1 _8221_ (.B(_3247_),
    .A(_0071_),
    .X(_3248_));
 sg13g2_nor2_1 _8222_ (.A(_3224_),
    .B(_3248_),
    .Y(_3249_));
 sg13g2_nand2b_1 _8223_ (.Y(_3250_),
    .B(_3222_),
    .A_N(_3233_));
 sg13g2_a22oi_1 _8224_ (.Y(_3251_),
    .B1(_3249_),
    .B2(_3250_),
    .A2(_3247_),
    .A1(_0893_));
 sg13g2_nand2_1 _8225_ (.Y(_3252_),
    .A(_3244_),
    .B(net111));
 sg13g2_o21ai_1 _8226_ (.B1(_3252_),
    .Y(_3253_),
    .A1(_3245_),
    .A2(_3251_));
 sg13g2_inv_1 _8227_ (.Y(_3254_),
    .A(_0901_));
 sg13g2_nor2_1 _8228_ (.A(_0611_),
    .B(_3246_),
    .Y(_3255_));
 sg13g2_nor2_1 _8229_ (.A(_3254_),
    .B(_3255_),
    .Y(_3256_));
 sg13g2_nor2_1 _8230_ (.A(_0901_),
    .B(_3241_),
    .Y(_3257_));
 sg13g2_a221oi_1 _8231_ (.B2(_3256_),
    .C1(_3257_),
    .B1(_3253_),
    .A1(_3239_),
    .Y(_3258_),
    .A2(_3242_));
 sg13g2_buf_1 _8232_ (.A(_3258_),
    .X(_3259_));
 sg13g2_nor2b_1 _8233_ (.A(_3221_),
    .B_N(_3259_),
    .Y(_3260_));
 sg13g2_buf_8 _8234_ (.A(_3260_),
    .X(_3261_));
 sg13g2_xor2_1 _8235_ (.B(net111),
    .A(net104),
    .X(_3262_));
 sg13g2_xnor2_1 _8236_ (.Y(_3263_),
    .A(net96),
    .B(_0889_));
 sg13g2_nand2_1 _8237_ (.Y(_3264_),
    .A(_0757_),
    .B(_0881_));
 sg13g2_xor2_1 _8238_ (.B(_0885_),
    .A(net107),
    .X(_3265_));
 sg13g2_nor2b_1 _8239_ (.A(_3264_),
    .B_N(_3265_),
    .Y(_3266_));
 sg13g2_a21oi_1 _8240_ (.A1(net107),
    .A2(_0885_),
    .Y(_3267_),
    .B1(_3266_));
 sg13g2_nand2_1 _8241_ (.Y(_3268_),
    .A(net96),
    .B(_0889_));
 sg13g2_o21ai_1 _8242_ (.B1(_3268_),
    .Y(_3269_),
    .A1(_3263_),
    .A2(_3267_));
 sg13g2_xor2_1 _8243_ (.B(_0893_),
    .A(net105),
    .X(_3270_));
 sg13g2_nand2_1 _8244_ (.Y(_3271_),
    .A(_3269_),
    .B(_3270_));
 sg13g2_o21ai_1 _8245_ (.B1(_3271_),
    .Y(_3272_),
    .A1(_4347_),
    .A2(_3236_));
 sg13g2_xor2_1 _8246_ (.B(_3272_),
    .A(_3262_),
    .X(_3273_));
 sg13g2_nor2_1 _8247_ (.A(_4578_),
    .B(\vgademo.plane_u[17] ),
    .Y(_3274_));
 sg13g2_nand2_1 _8248_ (.Y(_3275_),
    .A(_4578_),
    .B(\vgademo.plane_u[17] ));
 sg13g2_nor2b_1 _8249_ (.A(_3274_),
    .B_N(_3275_),
    .Y(_3276_));
 sg13g2_nor2_1 _8250_ (.A(_4503_),
    .B(\vgademo.plane_u[13] ),
    .Y(_3277_));
 sg13g2_nand2_1 _8251_ (.Y(_3278_),
    .A(_4533_),
    .B(\vgademo.plane_u[9] ));
 sg13g2_nor2_1 _8252_ (.A(_4540_),
    .B(_1224_),
    .Y(_3279_));
 sg13g2_nand2_1 _8253_ (.Y(_3280_),
    .A(_4540_),
    .B(_1224_));
 sg13g2_o21ai_1 _8254_ (.B1(_3280_),
    .Y(_3281_),
    .A1(_3278_),
    .A2(_3279_));
 sg13g2_nor2_1 _8255_ (.A(\vgademo.a_cos[6] ),
    .B(\vgademo.plane_u[11] ),
    .Y(_3282_));
 sg13g2_inv_1 _8256_ (.Y(_3283_),
    .A(_3282_));
 sg13g2_nand2_1 _8257_ (.Y(_3284_),
    .A(\vgademo.a_cos[6] ),
    .B(\vgademo.plane_u[11] ));
 sg13g2_inv_1 _8258_ (.Y(_3285_),
    .A(_3284_));
 sg13g2_a21oi_1 _8259_ (.A1(_3281_),
    .A2(_3283_),
    .Y(_3286_),
    .B1(_3285_));
 sg13g2_xor2_1 _8260_ (.B(_1396_),
    .A(_4507_),
    .X(_3287_));
 sg13g2_nor2b_1 _8261_ (.A(_3286_),
    .B_N(_3287_),
    .Y(_3288_));
 sg13g2_a21oi_1 _8262_ (.A1(_4507_),
    .A2(_1396_),
    .Y(_3289_),
    .B1(_3288_));
 sg13g2_nand2_1 _8263_ (.Y(_3290_),
    .A(_4503_),
    .B(\vgademo.plane_u[13] ));
 sg13g2_o21ai_1 _8264_ (.B1(_3290_),
    .Y(_3291_),
    .A1(_3277_),
    .A2(_3289_));
 sg13g2_xor2_1 _8265_ (.B(_1448_),
    .A(_4556_),
    .X(_3292_));
 sg13g2_nand2_1 _8266_ (.Y(_3293_),
    .A(_3291_),
    .B(_3292_));
 sg13g2_nand2_1 _8267_ (.Y(_3294_),
    .A(_4556_),
    .B(_1448_));
 sg13g2_nand2_1 _8268_ (.Y(_3295_),
    .A(_3293_),
    .B(_3294_));
 sg13g2_inv_1 _8269_ (.Y(_3296_),
    .A(_3295_));
 sg13g2_nand2_1 _8270_ (.Y(_3297_),
    .A(_4495_),
    .B(_1475_));
 sg13g2_nor2_1 _8271_ (.A(_4495_),
    .B(_1475_),
    .Y(_3298_));
 sg13g2_a21oi_1 _8272_ (.A1(_3296_),
    .A2(_3297_),
    .Y(_3299_),
    .B1(_3298_));
 sg13g2_inv_1 _8273_ (.Y(_3300_),
    .A(_3299_));
 sg13g2_nand2_1 _8274_ (.Y(_3301_),
    .A(_4563_),
    .B(\vgademo.plane_u[16] ));
 sg13g2_nor2_1 _8275_ (.A(_4563_),
    .B(\vgademo.plane_u[16] ),
    .Y(_3302_));
 sg13g2_a21oi_1 _8276_ (.A1(_3300_),
    .A2(_3301_),
    .Y(_3303_),
    .B1(_3302_));
 sg13g2_xor2_1 _8277_ (.B(_3303_),
    .A(_3276_),
    .X(_3304_));
 sg13g2_xor2_1 _8278_ (.B(_3304_),
    .A(_3273_),
    .X(_3305_));
 sg13g2_inv_1 _8279_ (.Y(_3306_),
    .A(_3305_));
 sg13g2_nand2_1 _8280_ (.Y(_3307_),
    .A(_3306_),
    .B(net88));
 sg13g2_nand2_1 _8281_ (.Y(_3308_),
    .A(_3305_),
    .B(_1661_));
 sg13g2_nor2b_1 _8282_ (.A(_3302_),
    .B_N(_3301_),
    .Y(_3309_));
 sg13g2_xor2_1 _8283_ (.B(_3299_),
    .A(_3309_),
    .X(_3310_));
 sg13g2_nand2_1 _8284_ (.Y(_3311_),
    .A(_3310_),
    .B(_0767_));
 sg13g2_xor2_1 _8285_ (.B(_3269_),
    .A(_3270_),
    .X(_3312_));
 sg13g2_inv_1 _8286_ (.Y(_3313_),
    .A(_3310_));
 sg13g2_o21ai_1 _8287_ (.B1(_0778_),
    .Y(_3314_),
    .A1(net79),
    .A2(_3312_));
 sg13g2_a221oi_1 _8288_ (.B2(net117),
    .C1(_3314_),
    .B1(_3313_),
    .A1(net79),
    .Y(_3315_),
    .A2(_3312_));
 sg13g2_nand4_1 _8289_ (.B(_3308_),
    .C(_3311_),
    .A(_3307_),
    .Y(_3316_),
    .D(_3315_));
 sg13g2_xor2_1 _8290_ (.B(_0901_),
    .A(net103),
    .X(_3317_));
 sg13g2_inv_1 _8291_ (.Y(_3318_),
    .A(net111));
 sg13g2_nand2_1 _8292_ (.Y(_3319_),
    .A(_3272_),
    .B(_3262_));
 sg13g2_o21ai_1 _8293_ (.B1(_3319_),
    .Y(_3320_),
    .A1(_4365_),
    .A2(_3318_));
 sg13g2_xor2_1 _8294_ (.B(_3320_),
    .A(_3317_),
    .X(_3321_));
 sg13g2_inv_1 _8295_ (.Y(_3322_),
    .A(_3321_));
 sg13g2_nor2_1 _8296_ (.A(_0381_),
    .B(\vgademo.plane_u[18] ),
    .Y(_3323_));
 sg13g2_nand2_1 _8297_ (.Y(_3324_),
    .A(_0381_),
    .B(\vgademo.plane_u[18] ));
 sg13g2_inv_1 _8298_ (.Y(_3325_),
    .A(_3324_));
 sg13g2_nor2_1 _8299_ (.A(_3323_),
    .B(_3325_),
    .Y(_3326_));
 sg13g2_inv_1 _8300_ (.Y(_3327_),
    .A(_3303_));
 sg13g2_o21ai_1 _8301_ (.B1(_3275_),
    .Y(_3328_),
    .A1(_3274_),
    .A2(_3327_));
 sg13g2_xnor2_1 _8302_ (.Y(_3329_),
    .A(_3326_),
    .B(_3328_));
 sg13g2_xnor2_1 _8303_ (.Y(_3330_),
    .A(_3322_),
    .B(_3329_));
 sg13g2_xnor2_1 _8304_ (.Y(_3331_),
    .A(net116),
    .B(_3330_));
 sg13g2_nor2_1 _8305_ (.A(_3316_),
    .B(_3331_),
    .Y(_3332_));
 sg13g2_buf_1 _8306_ (.A(_3332_),
    .X(_3333_));
 sg13g2_xnor2_1 _8307_ (.Y(_3334_),
    .A(net95),
    .B(_0398_));
 sg13g2_xor2_1 _8308_ (.B(\vgademo.plane_u[19] ),
    .A(_0866_),
    .X(_3335_));
 sg13g2_xnor2_1 _8309_ (.Y(_3336_),
    .A(_3334_),
    .B(_3335_));
 sg13g2_nand2_1 _8310_ (.Y(_3337_),
    .A(_3320_),
    .B(_3317_));
 sg13g2_o21ai_1 _8311_ (.B1(_3337_),
    .Y(_3338_),
    .A1(net106),
    .A2(_3254_));
 sg13g2_xnor2_1 _8312_ (.Y(_3339_),
    .A(_3336_),
    .B(_3338_));
 sg13g2_inv_1 _8313_ (.Y(_3340_),
    .A(_3323_));
 sg13g2_a21oi_1 _8314_ (.A1(_3328_),
    .A2(_3340_),
    .Y(_3341_),
    .B1(_3325_));
 sg13g2_xnor2_1 _8315_ (.Y(_3342_),
    .A(_3339_),
    .B(_3341_));
 sg13g2_inv_1 _8316_ (.Y(_3343_),
    .A(_3329_));
 sg13g2_inv_1 _8317_ (.Y(_3344_),
    .A(_3312_));
 sg13g2_nor2_1 _8318_ (.A(_3344_),
    .B(_3313_),
    .Y(_3345_));
 sg13g2_inv_1 _8319_ (.Y(_3346_),
    .A(_3345_));
 sg13g2_nor2_1 _8320_ (.A(_3346_),
    .B(_3306_),
    .Y(_3347_));
 sg13g2_a21oi_1 _8321_ (.A1(_3273_),
    .A2(_3304_),
    .Y(_3348_),
    .B1(_3347_));
 sg13g2_nor2_1 _8322_ (.A(_3330_),
    .B(_3348_),
    .Y(_3349_));
 sg13g2_a21oi_1 _8323_ (.A1(_3321_),
    .A2(_3343_),
    .Y(_3350_),
    .B1(_3349_));
 sg13g2_xnor2_1 _8324_ (.Y(_3351_),
    .A(_3342_),
    .B(_3350_));
 sg13g2_nor2_1 _8325_ (.A(net78),
    .B(_3351_),
    .Y(_3352_));
 sg13g2_nor2_1 _8326_ (.A(_3344_),
    .B(_3310_),
    .Y(_3353_));
 sg13g2_nor2_1 _8327_ (.A(_3312_),
    .B(_3313_),
    .Y(_3354_));
 sg13g2_nor2_1 _8328_ (.A(_3353_),
    .B(_3354_),
    .Y(_3355_));
 sg13g2_buf_2 _8329_ (.A(_3355_),
    .X(_3356_));
 sg13g2_nor3_1 _8330_ (.A(net97),
    .B(net88),
    .C(_3356_),
    .Y(_3357_));
 sg13g2_xnor2_1 _8331_ (.Y(_3358_),
    .A(_3346_),
    .B(_3305_));
 sg13g2_o21ai_1 _8332_ (.B1(net97),
    .Y(_3359_),
    .A1(net88),
    .A2(_3356_));
 sg13g2_o21ai_1 _8333_ (.B1(_3359_),
    .Y(_3360_),
    .A1(_3357_),
    .A2(_3358_));
 sg13g2_xor2_1 _8334_ (.B(_3348_),
    .A(_3330_),
    .X(_3361_));
 sg13g2_nand2_1 _8335_ (.Y(_3362_),
    .A(_3361_),
    .B(net77));
 sg13g2_nor2_1 _8336_ (.A(net77),
    .B(_3361_),
    .Y(_3363_));
 sg13g2_a221oi_1 _8337_ (.B2(net78),
    .C1(_3363_),
    .B1(_3351_),
    .A1(_3360_),
    .Y(_3364_),
    .A2(_3362_));
 sg13g2_nor3_2 _8338_ (.A(_1711_),
    .B(_3352_),
    .C(_3364_),
    .Y(_3365_));
 sg13g2_a21o_1 _8339_ (.A2(net26),
    .A1(_0080_),
    .B1(_3365_),
    .X(_3366_));
 sg13g2_inv_1 _8340_ (.Y(_3367_),
    .A(_3366_));
 sg13g2_inv_1 _8341_ (.Y(_3368_),
    .A(_3264_));
 sg13g2_nor3_1 _8342_ (.A(_3266_),
    .B(_3356_),
    .C(net26),
    .Y(_3369_));
 sg13g2_o21ai_1 _8343_ (.B1(_3369_),
    .Y(_3370_),
    .A1(_3368_),
    .A2(_3265_));
 sg13g2_nand2_1 _8344_ (.Y(_3371_),
    .A(_3367_),
    .B(_3370_));
 sg13g2_nand2_1 _8345_ (.Y(_3372_),
    .A(net14),
    .B(_3371_));
 sg13g2_nand3_1 _8346_ (.B(_3220_),
    .C(_3259_),
    .A(_3149_),
    .Y(_3373_));
 sg13g2_buf_2 _8347_ (.A(_3373_),
    .X(_3374_));
 sg13g2_buf_8 _8348_ (.A(_3374_),
    .X(_3375_));
 sg13g2_a21oi_1 _8349_ (.A1(_0075_),
    .A2(net26),
    .Y(_3376_),
    .B1(_3365_));
 sg13g2_inv_2 _8350_ (.Y(_3377_),
    .A(_3333_));
 sg13g2_inv_2 _8351_ (.Y(_3378_),
    .A(_3356_));
 sg13g2_nand3_1 _8352_ (.B(_0877_),
    .C(_3378_),
    .A(_3377_),
    .Y(_3379_));
 sg13g2_nand2_1 _8353_ (.Y(_3380_),
    .A(_3376_),
    .B(_3379_));
 sg13g2_nand2_1 _8354_ (.Y(_3381_),
    .A(net13),
    .B(_3380_));
 sg13g2_buf_1 _8355_ (.A(net22),
    .X(_3382_));
 sg13g2_nand3_1 _8356_ (.B(_3381_),
    .C(net21),
    .A(_3372_),
    .Y(_3383_));
 sg13g2_nor2_1 _8357_ (.A(_4456_),
    .B(_0591_),
    .Y(_3384_));
 sg13g2_nor2_1 _8358_ (.A(_2765_),
    .B(_3384_),
    .Y(_3385_));
 sg13g2_a21oi_1 _8359_ (.A1(_4456_),
    .A2(_0591_),
    .Y(_3386_),
    .B1(_3385_));
 sg13g2_nor2_1 _8360_ (.A(_0588_),
    .B(_0964_),
    .Y(_3387_));
 sg13g2_xnor2_1 _8361_ (.Y(_3388_),
    .A(_4458_),
    .B(net119));
 sg13g2_nand2_1 _8362_ (.Y(_3389_),
    .A(_0964_),
    .B(_0588_));
 sg13g2_nand3b_1 _8363_ (.B(_3388_),
    .C(_3389_),
    .Y(_3390_),
    .A_N(_3387_));
 sg13g2_nor2_1 _8364_ (.A(_0601_),
    .B(_4459_),
    .Y(_3391_));
 sg13g2_a21oi_1 _8365_ (.A1(_3388_),
    .A2(_3387_),
    .Y(_3392_),
    .B1(_3391_));
 sg13g2_o21ai_1 _8366_ (.B1(_3392_),
    .Y(_3393_),
    .A1(_3386_),
    .A2(_3390_));
 sg13g2_nand2_1 _8367_ (.Y(_3394_),
    .A(_4449_),
    .B(_0554_));
 sg13g2_nand2_1 _8368_ (.Y(_3395_),
    .A(_4448_),
    .B(_0553_));
 sg13g2_nor2_1 _8369_ (.A(net122),
    .B(net100),
    .Y(_3396_));
 sg13g2_nand2_1 _8370_ (.Y(_3397_),
    .A(net122),
    .B(net100));
 sg13g2_inv_1 _8371_ (.Y(_3398_),
    .A(_3397_));
 sg13g2_nor2_1 _8372_ (.A(_3396_),
    .B(_3398_),
    .Y(_3399_));
 sg13g2_inv_1 _8373_ (.Y(_3400_),
    .A(_3399_));
 sg13g2_nand4_1 _8374_ (.B(_3394_),
    .C(_3395_),
    .A(_3393_),
    .Y(_3401_),
    .D(_3400_));
 sg13g2_o21ai_1 _8375_ (.B1(_3395_),
    .Y(_3402_),
    .A1(_0599_),
    .A2(_4569_));
 sg13g2_a22oi_1 _8376_ (.Y(_3403_),
    .B1(_3394_),
    .B2(_3402_),
    .A2(_1033_),
    .A1(_3138_));
 sg13g2_xnor2_1 _8377_ (.Y(_3404_),
    .A(_1076_),
    .B(_3240_));
 sg13g2_a221oi_1 _8378_ (.B2(_3403_),
    .C1(_3404_),
    .B1(_3401_),
    .A1(_1031_),
    .Y(_3405_),
    .A2(_3137_));
 sg13g2_nor2b_1 _8379_ (.A(_3405_),
    .B_N(_2739_),
    .Y(_3406_));
 sg13g2_nand2_1 _8380_ (.Y(_3407_),
    .A(_3241_),
    .B(net121));
 sg13g2_nand2b_1 _8381_ (.Y(_3408_),
    .B(_0406_),
    .A_N(_3244_));
 sg13g2_o21ai_1 _8382_ (.B1(_1071_),
    .Y(_3409_),
    .A1(_1076_),
    .A2(_3255_));
 sg13g2_nand3_1 _8383_ (.B(_0040_),
    .C(_3409_),
    .A(_3408_),
    .Y(_3410_));
 sg13g2_nand2b_1 _8384_ (.Y(_3411_),
    .B(_3386_),
    .A_N(_3387_));
 sg13g2_nand4_1 _8385_ (.B(_3389_),
    .C(_3399_),
    .A(_3411_),
    .Y(_3412_),
    .D(_3388_));
 sg13g2_a21oi_1 _8386_ (.A1(_3399_),
    .A2(_3391_),
    .Y(_3413_),
    .B1(_3398_));
 sg13g2_xnor2_1 _8387_ (.Y(_3414_),
    .A(_2725_),
    .B(_3247_));
 sg13g2_a21oi_1 _8388_ (.A1(_3412_),
    .A2(_3413_),
    .Y(_3415_),
    .B1(_3414_));
 sg13g2_a22oi_1 _8389_ (.Y(_3416_),
    .B1(_4454_),
    .B2(_3244_),
    .A2(_3247_),
    .A1(_4448_));
 sg13g2_nor2b_1 _8390_ (.A(_3415_),
    .B_N(_3416_),
    .Y(_3417_));
 sg13g2_nand2_1 _8391_ (.Y(_3418_),
    .A(_3255_),
    .B(_1076_));
 sg13g2_a21oi_1 _8392_ (.A1(_3418_),
    .A2(_1073_),
    .Y(_3419_),
    .B1(_4447_));
 sg13g2_o21ai_1 _8393_ (.B1(_3419_),
    .Y(_3420_),
    .A1(_3410_),
    .A2(_3417_));
 sg13g2_a21oi_1 _8394_ (.A1(_3406_),
    .A2(_3407_),
    .Y(_3421_),
    .B1(_3420_));
 sg13g2_nor2b_2 _8395_ (.A(_3221_),
    .B_N(_3421_),
    .Y(_3422_));
 sg13g2_inv_4 _8396_ (.A(_3422_),
    .Y(_3423_));
 sg13g2_buf_8 _8397_ (.A(_3423_),
    .X(_3424_));
 sg13g2_nor2_1 _8398_ (.A(_4319_),
    .B(_4352_),
    .Y(_3425_));
 sg13g2_nor2_1 _8399_ (.A(_4447_),
    .B(net94),
    .Y(_3426_));
 sg13g2_nor2_1 _8400_ (.A(_0037_),
    .B(_3426_),
    .Y(_3427_));
 sg13g2_xor2_1 _8401_ (.B(net94),
    .A(_4447_),
    .X(_3428_));
 sg13g2_a21oi_1 _8402_ (.A1(_4451_),
    .A2(net83),
    .Y(_3429_),
    .B1(_3428_));
 sg13g2_inv_1 _8403_ (.Y(_3430_),
    .A(_3429_));
 sg13g2_nand3_1 _8404_ (.B(_4451_),
    .C(net83),
    .A(_3428_),
    .Y(_3431_));
 sg13g2_nand2_1 _8405_ (.Y(_3432_),
    .A(_3430_),
    .B(_3431_));
 sg13g2_xor2_1 _8406_ (.B(net95),
    .A(_4450_),
    .X(_3433_));
 sg13g2_nor3_1 _8407_ (.A(_0405_),
    .B(net106),
    .C(_3433_),
    .Y(_3434_));
 sg13g2_nor2_1 _8408_ (.A(_4446_),
    .B(net96),
    .Y(_3435_));
 sg13g2_xor2_1 _8409_ (.B(net105),
    .A(_4448_),
    .X(_3436_));
 sg13g2_o21ai_1 _8410_ (.B1(net107),
    .Y(_3437_),
    .A1(_4455_),
    .A2(_0757_));
 sg13g2_nand2_1 _8411_ (.Y(_3438_),
    .A(_4446_),
    .B(net96));
 sg13g2_inv_1 _8412_ (.Y(_3439_),
    .A(_3438_));
 sg13g2_nand3_1 _8413_ (.B(_4459_),
    .C(_0964_),
    .A(_0796_),
    .Y(_3440_));
 sg13g2_o21ai_1 _8414_ (.B1(_3440_),
    .Y(_3441_),
    .A1(_3435_),
    .A2(_3439_));
 sg13g2_o21ai_1 _8415_ (.B1(_3441_),
    .Y(_3442_),
    .A1(_4459_),
    .A2(_3437_));
 sg13g2_nand2_1 _8416_ (.Y(_3443_),
    .A(_3436_),
    .B(_3435_));
 sg13g2_nand2_1 _8417_ (.Y(_3444_),
    .A(_3442_),
    .B(_3443_));
 sg13g2_o21ai_1 _8418_ (.B1(_3444_),
    .Y(_3445_),
    .A1(_3435_),
    .A2(_3436_));
 sg13g2_nor2_1 _8419_ (.A(_4448_),
    .B(net105),
    .Y(_3446_));
 sg13g2_xnor2_1 _8420_ (.Y(_3447_),
    .A(_4454_),
    .B(net104));
 sg13g2_xnor2_1 _8421_ (.Y(_3448_),
    .A(_3446_),
    .B(_3447_));
 sg13g2_nor2b_1 _8422_ (.A(_3446_),
    .B_N(_3447_),
    .Y(_3449_));
 sg13g2_a21o_1 _8423_ (.A2(_3448_),
    .A1(_3445_),
    .B1(_3449_),
    .X(_3450_));
 sg13g2_nand2_1 _8424_ (.Y(_3451_),
    .A(_0406_),
    .B(_4365_));
 sg13g2_xor2_1 _8425_ (.B(net103),
    .A(_4453_),
    .X(_3452_));
 sg13g2_xor2_1 _8426_ (.B(_3452_),
    .A(_3451_),
    .X(_3453_));
 sg13g2_nand2_1 _8427_ (.Y(_3454_),
    .A(_3450_),
    .B(_3453_));
 sg13g2_nand2_1 _8428_ (.Y(_3455_),
    .A(_3452_),
    .B(_3451_));
 sg13g2_nand2_1 _8429_ (.Y(_3456_),
    .A(_3454_),
    .B(_3455_));
 sg13g2_inv_1 _8430_ (.Y(_3457_),
    .A(_3433_));
 sg13g2_a21oi_1 _8431_ (.A1(_4453_),
    .A2(net103),
    .Y(_3458_),
    .B1(_3457_));
 sg13g2_inv_1 _8432_ (.Y(_3459_),
    .A(_3458_));
 sg13g2_o21ai_1 _8433_ (.B1(_3459_),
    .Y(_3460_),
    .A1(_3434_),
    .A2(_3456_));
 sg13g2_o21ai_1 _8434_ (.B1(_3430_),
    .Y(_3461_),
    .A1(_3432_),
    .A2(_3460_));
 sg13g2_xnor2_1 _8435_ (.Y(_3462_),
    .A(_4312_),
    .B(_3426_));
 sg13g2_nand2_1 _8436_ (.Y(_3463_),
    .A(_3461_),
    .B(_3462_));
 sg13g2_inv_1 _8437_ (.Y(_3464_),
    .A(_3463_));
 sg13g2_a22oi_1 _8438_ (.Y(_3465_),
    .B1(_0060_),
    .B2(_3464_),
    .A2(_3427_),
    .A1(_4359_));
 sg13g2_xnor2_1 _8439_ (.Y(_3466_),
    .A(_3425_),
    .B(_3465_));
 sg13g2_buf_1 _8440_ (.A(_3466_),
    .X(_3467_));
 sg13g2_xnor2_1 _8441_ (.Y(_3468_),
    .A(_3448_),
    .B(_3445_));
 sg13g2_nor4_1 _8442_ (.A(_0813_),
    .B(_4364_),
    .C(_0760_),
    .D(_4339_),
    .Y(_3469_));
 sg13g2_nor2_1 _8443_ (.A(_4353_),
    .B(_3469_),
    .Y(_3470_));
 sg13g2_nor2_1 _8444_ (.A(_2791_),
    .B(_0797_),
    .Y(_3471_));
 sg13g2_nor2_1 _8445_ (.A(net94),
    .B(_0813_),
    .Y(_3472_));
 sg13g2_nand4_1 _8446_ (.B(_4379_),
    .C(_4326_),
    .A(_3471_),
    .Y(_3473_),
    .D(_3472_));
 sg13g2_nand2_1 _8447_ (.Y(_3474_),
    .A(_3473_),
    .B(_0758_));
 sg13g2_nor2_1 _8448_ (.A(_3470_),
    .B(_3474_),
    .Y(_3475_));
 sg13g2_nor2_1 _8449_ (.A(_3427_),
    .B(_3464_),
    .Y(_3476_));
 sg13g2_a21oi_1 _8450_ (.A1(_3476_),
    .A2(_4359_),
    .Y(_3477_),
    .B1(_4318_));
 sg13g2_xnor2_1 _8451_ (.Y(_3478_),
    .A(_0015_),
    .B(_3477_));
 sg13g2_inv_1 _8452_ (.Y(_3479_),
    .A(_3478_));
 sg13g2_nor2_1 _8453_ (.A(_3475_),
    .B(_3479_),
    .Y(_3480_));
 sg13g2_inv_1 _8454_ (.Y(_3481_),
    .A(_3480_));
 sg13g2_a21oi_1 _8455_ (.A1(_3467_),
    .A2(_3468_),
    .Y(_3482_),
    .B1(_3481_));
 sg13g2_nand2_1 _8456_ (.Y(_3483_),
    .A(net104),
    .B(net93));
 sg13g2_nand2_1 _8457_ (.Y(_3484_),
    .A(net103),
    .B(net115));
 sg13g2_nand2_1 _8458_ (.Y(_3485_),
    .A(_3483_),
    .B(_3484_));
 sg13g2_nand2_1 _8459_ (.Y(_3486_),
    .A(net104),
    .B(net115));
 sg13g2_nand2_1 _8460_ (.Y(_3487_),
    .A(net103),
    .B(net93));
 sg13g2_nor2_1 _8461_ (.A(_3486_),
    .B(_3487_),
    .Y(_3488_));
 sg13g2_a21oi_1 _8462_ (.A1(_3485_),
    .A2(\vgademo.linelfsr[9] ),
    .Y(_3489_),
    .B1(_3488_));
 sg13g2_nand2_1 _8463_ (.Y(_3490_),
    .A(net95),
    .B(_0829_));
 sg13g2_nand2_1 _8464_ (.Y(_3491_),
    .A(net95),
    .B(net115));
 sg13g2_nand2_1 _8465_ (.Y(_3492_),
    .A(_3487_),
    .B(_3491_));
 sg13g2_o21ai_1 _8466_ (.B1(_3492_),
    .Y(_3493_),
    .A1(_3484_),
    .A2(_3490_));
 sg13g2_xnor2_1 _8467_ (.Y(_3494_),
    .A(_0853_),
    .B(_3493_));
 sg13g2_nor2_1 _8468_ (.A(_3489_),
    .B(_3494_),
    .Y(_3495_));
 sg13g2_xnor2_1 _8469_ (.Y(_3496_),
    .A(_3489_),
    .B(_3494_));
 sg13g2_nor2_1 _8470_ (.A(_4341_),
    .B(_3496_),
    .Y(_3497_));
 sg13g2_nor2_1 _8471_ (.A(_3495_),
    .B(_3497_),
    .Y(_3498_));
 sg13g2_nor2_1 _8472_ (.A(_3484_),
    .B(_3490_),
    .Y(_3499_));
 sg13g2_a21oi_1 _8473_ (.A1(_3492_),
    .A2(\vgademo.linelfsr[10] ),
    .Y(_3500_),
    .B1(_3499_));
 sg13g2_nand2_1 _8474_ (.Y(_3501_),
    .A(net94),
    .B(net93));
 sg13g2_nor2_1 _8475_ (.A(_3491_),
    .B(_3501_),
    .Y(_3502_));
 sg13g2_o21ai_1 _8476_ (.B1(_3490_),
    .Y(_3503_),
    .A1(_4341_),
    .A2(_0827_));
 sg13g2_nand2b_1 _8477_ (.Y(_3504_),
    .B(_3503_),
    .A_N(_3502_));
 sg13g2_xnor2_1 _8478_ (.Y(_3505_),
    .A(_0836_),
    .B(_3504_));
 sg13g2_xnor2_1 _8479_ (.Y(_3506_),
    .A(_3500_),
    .B(_3505_));
 sg13g2_xnor2_1 _8480_ (.Y(_3507_),
    .A(_4335_),
    .B(_3506_));
 sg13g2_nor2_1 _8481_ (.A(_3498_),
    .B(_3507_),
    .Y(_3508_));
 sg13g2_nand2_1 _8482_ (.Y(_3509_),
    .A(_3507_),
    .B(_3498_));
 sg13g2_nor2b_1 _8483_ (.A(_3508_),
    .B_N(_3509_),
    .Y(_3510_));
 sg13g2_nand2_1 _8484_ (.Y(_3511_),
    .A(net105),
    .B(_0828_));
 sg13g2_nand2_1 _8485_ (.Y(_3512_),
    .A(_3511_),
    .B(_3486_));
 sg13g2_nand2_1 _8486_ (.Y(_3513_),
    .A(net105),
    .B(net115));
 sg13g2_nor2_1 _8487_ (.A(_3513_),
    .B(_3483_),
    .Y(_3514_));
 sg13g2_a21oi_1 _8488_ (.A1(_3512_),
    .A2(\vgademo.linelfsr[8] ),
    .Y(_3515_),
    .B1(_3514_));
 sg13g2_o21ai_1 _8489_ (.B1(_3485_),
    .Y(_3516_),
    .A1(_3486_),
    .A2(_3487_));
 sg13g2_xnor2_1 _8490_ (.Y(_3517_),
    .A(_0854_),
    .B(_3516_));
 sg13g2_nor2_1 _8491_ (.A(_3515_),
    .B(_3517_),
    .Y(_3518_));
 sg13g2_xnor2_1 _8492_ (.Y(_3519_),
    .A(_3515_),
    .B(_3517_));
 sg13g2_nor2_1 _8493_ (.A(net83),
    .B(_3519_),
    .Y(_3520_));
 sg13g2_nor2_1 _8494_ (.A(_3518_),
    .B(_3520_),
    .Y(_3521_));
 sg13g2_xnor2_1 _8495_ (.Y(_3522_),
    .A(_4341_),
    .B(_3496_));
 sg13g2_nor2_1 _8496_ (.A(_3521_),
    .B(_3522_),
    .Y(_3523_));
 sg13g2_nand2_1 _8497_ (.Y(_3524_),
    .A(net96),
    .B(_0828_));
 sg13g2_nand2_1 _8498_ (.Y(_3525_),
    .A(_3513_),
    .B(_3524_));
 sg13g2_nand2_1 _8499_ (.Y(_3526_),
    .A(net96),
    .B(net115));
 sg13g2_nor2_1 _8500_ (.A(_3511_),
    .B(_3526_),
    .Y(_3527_));
 sg13g2_a21oi_1 _8501_ (.A1(_3525_),
    .A2(\vgademo.linelfsr[7] ),
    .Y(_3528_),
    .B1(_3527_));
 sg13g2_o21ai_1 _8502_ (.B1(_3512_),
    .Y(_3529_),
    .A1(_3513_),
    .A2(_3483_));
 sg13g2_xnor2_1 _8503_ (.Y(_3530_),
    .A(_0849_),
    .B(_3529_));
 sg13g2_nor2_1 _8504_ (.A(_3528_),
    .B(_3530_),
    .Y(_3531_));
 sg13g2_xnor2_1 _8505_ (.Y(_3532_),
    .A(_3528_),
    .B(_3530_));
 sg13g2_nor2_1 _8506_ (.A(net106),
    .B(_3532_),
    .Y(_3533_));
 sg13g2_nor2_1 _8507_ (.A(_3531_),
    .B(_3533_),
    .Y(_3534_));
 sg13g2_xnor2_1 _8508_ (.Y(_3535_),
    .A(net83),
    .B(_3519_));
 sg13g2_nor2_1 _8509_ (.A(_3534_),
    .B(_3535_),
    .Y(_3536_));
 sg13g2_nand2_1 _8510_ (.Y(_3537_),
    .A(net107),
    .B(_0828_));
 sg13g2_nand2_1 _8511_ (.Y(_3538_),
    .A(_3526_),
    .B(_3537_));
 sg13g2_nand2_1 _8512_ (.Y(_3539_),
    .A(net107),
    .B(_0826_));
 sg13g2_nor2_1 _8513_ (.A(_3524_),
    .B(_3539_),
    .Y(_3540_));
 sg13g2_a21oi_1 _8514_ (.A1(_3538_),
    .A2(\vgademo.linelfsr[6] ),
    .Y(_3541_),
    .B1(_3540_));
 sg13g2_o21ai_1 _8515_ (.B1(_3525_),
    .Y(_3542_),
    .A1(_3511_),
    .A2(_3526_));
 sg13g2_xnor2_1 _8516_ (.Y(_3543_),
    .A(_0850_),
    .B(_3542_));
 sg13g2_nor2_1 _8517_ (.A(_3541_),
    .B(_3543_),
    .Y(_3544_));
 sg13g2_xnor2_1 _8518_ (.Y(_3545_),
    .A(_3541_),
    .B(_3543_));
 sg13g2_nor2_1 _8519_ (.A(_4365_),
    .B(_3545_),
    .Y(_3546_));
 sg13g2_nor2_1 _8520_ (.A(_3544_),
    .B(_3546_),
    .Y(_3547_));
 sg13g2_xnor2_1 _8521_ (.Y(_3548_),
    .A(net106),
    .B(_3532_));
 sg13g2_nor2_1 _8522_ (.A(_3547_),
    .B(_3548_),
    .Y(_3549_));
 sg13g2_nand2_1 _8523_ (.Y(_3550_),
    .A(_4324_),
    .B(_0826_));
 sg13g2_nor2_1 _8524_ (.A(_3537_),
    .B(_3550_),
    .Y(_3551_));
 sg13g2_nand2_1 _8525_ (.Y(_3552_),
    .A(_4324_),
    .B(_0828_));
 sg13g2_xnor2_1 _8526_ (.Y(_3553_),
    .A(_3539_),
    .B(_3552_));
 sg13g2_nor2_1 _8527_ (.A(_0847_),
    .B(_3553_),
    .Y(_3554_));
 sg13g2_nor2_1 _8528_ (.A(_3551_),
    .B(_3554_),
    .Y(_3555_));
 sg13g2_o21ai_1 _8529_ (.B1(_3538_),
    .Y(_3556_),
    .A1(_3524_),
    .A2(_3539_));
 sg13g2_xnor2_1 _8530_ (.Y(_3557_),
    .A(_0846_),
    .B(_3556_));
 sg13g2_nor2_1 _8531_ (.A(_3555_),
    .B(_3557_),
    .Y(_3558_));
 sg13g2_xnor2_1 _8532_ (.Y(_3559_),
    .A(_3555_),
    .B(_3557_));
 sg13g2_nor2_1 _8533_ (.A(_4347_),
    .B(_3559_),
    .Y(_3560_));
 sg13g2_nor2_1 _8534_ (.A(_3558_),
    .B(_3560_),
    .Y(_3561_));
 sg13g2_xnor2_1 _8535_ (.Y(_3562_),
    .A(_4365_),
    .B(_3545_));
 sg13g2_nor2_1 _8536_ (.A(_0845_),
    .B(_3550_),
    .Y(_3563_));
 sg13g2_nand2_1 _8537_ (.Y(_3564_),
    .A(_3550_),
    .B(_0845_));
 sg13g2_nor2b_1 _8538_ (.A(_3563_),
    .B_N(_3564_),
    .Y(_3565_));
 sg13g2_xnor2_1 _8539_ (.Y(_3566_),
    .A(_4323_),
    .B(_3565_));
 sg13g2_inv_1 _8540_ (.Y(_3567_),
    .A(_3566_));
 sg13g2_nor3_1 _8541_ (.A(_2875_),
    .B(_0841_),
    .C(_3567_),
    .Y(_3568_));
 sg13g2_inv_1 _8542_ (.Y(_3569_),
    .A(_3568_));
 sg13g2_a21oi_1 _8543_ (.A1(_3564_),
    .A2(net107),
    .Y(_3570_),
    .B1(_3563_));
 sg13g2_xnor2_1 _8544_ (.Y(_3571_),
    .A(_0847_),
    .B(_3553_));
 sg13g2_xnor2_1 _8545_ (.Y(_3572_),
    .A(_3570_),
    .B(_3571_));
 sg13g2_xnor2_1 _8546_ (.Y(_3573_),
    .A(_0942_),
    .B(_3572_));
 sg13g2_nor2_1 _8547_ (.A(_3569_),
    .B(_3573_),
    .Y(_3574_));
 sg13g2_inv_1 _8548_ (.Y(_3575_),
    .A(_3574_));
 sg13g2_nor2_1 _8549_ (.A(_3570_),
    .B(_3571_),
    .Y(_3576_));
 sg13g2_nor2_1 _8550_ (.A(_0942_),
    .B(_3572_),
    .Y(_3577_));
 sg13g2_nor2_1 _8551_ (.A(_3576_),
    .B(_3577_),
    .Y(_3578_));
 sg13g2_xnor2_1 _8552_ (.Y(_3579_),
    .A(_4347_),
    .B(_3559_));
 sg13g2_xnor2_1 _8553_ (.Y(_3580_),
    .A(_3578_),
    .B(_3579_));
 sg13g2_or2_1 _8554_ (.X(_3581_),
    .B(_3579_),
    .A(_3578_));
 sg13g2_o21ai_1 _8555_ (.B1(_3581_),
    .Y(_3582_),
    .A1(_3575_),
    .A2(_3580_));
 sg13g2_xor2_1 _8556_ (.B(_3562_),
    .A(_3561_),
    .X(_3583_));
 sg13g2_nand2_1 _8557_ (.Y(_3584_),
    .A(_3582_),
    .B(_3583_));
 sg13g2_o21ai_1 _8558_ (.B1(_3584_),
    .Y(_3585_),
    .A1(_3561_),
    .A2(_3562_));
 sg13g2_xor2_1 _8559_ (.B(_3548_),
    .A(_3547_),
    .X(_3586_));
 sg13g2_nand2_1 _8560_ (.Y(_3587_),
    .A(_3585_),
    .B(_3586_));
 sg13g2_nand2b_1 _8561_ (.Y(_3588_),
    .B(_3587_),
    .A_N(_3549_));
 sg13g2_xor2_1 _8562_ (.B(_3535_),
    .A(_3534_),
    .X(_3589_));
 sg13g2_nand2_1 _8563_ (.Y(_3590_),
    .A(_3588_),
    .B(_3589_));
 sg13g2_nand2b_1 _8564_ (.Y(_3591_),
    .B(_3590_),
    .A_N(_3536_));
 sg13g2_xor2_1 _8565_ (.B(_3522_),
    .A(_3521_),
    .X(_3592_));
 sg13g2_nand2_1 _8566_ (.Y(_3593_),
    .A(_3591_),
    .B(_3592_));
 sg13g2_nand2b_1 _8567_ (.Y(_3594_),
    .B(_3593_),
    .A_N(_3523_));
 sg13g2_xnor2_1 _8568_ (.Y(_3595_),
    .A(_3510_),
    .B(_3594_));
 sg13g2_inv_1 _8569_ (.Y(_3596_),
    .A(_3595_));
 sg13g2_xor2_1 _8570_ (.B(_3591_),
    .A(_3592_),
    .X(_3597_));
 sg13g2_inv_1 _8571_ (.Y(_3598_),
    .A(_3597_));
 sg13g2_xor2_1 _8572_ (.B(_3582_),
    .A(_3583_),
    .X(_3599_));
 sg13g2_buf_1 _8573_ (.A(_3599_),
    .X(_3600_));
 sg13g2_inv_1 _8574_ (.Y(_3601_),
    .A(_3600_));
 sg13g2_xnor2_1 _8575_ (.Y(_3602_),
    .A(_3569_),
    .B(_3573_));
 sg13g2_xor2_1 _8576_ (.B(\vgademo.linelfsr[3] ),
    .A(net99),
    .X(_3603_));
 sg13g2_inv_1 _8577_ (.Y(_3604_),
    .A(_3603_));
 sg13g2_nor2_1 _8578_ (.A(_3604_),
    .B(_3567_),
    .Y(_3605_));
 sg13g2_inv_1 _8579_ (.Y(_3606_),
    .A(_3605_));
 sg13g2_nand2_1 _8580_ (.Y(_3607_),
    .A(_3602_),
    .B(_3606_));
 sg13g2_nor2_1 _8581_ (.A(_3606_),
    .B(_3573_),
    .Y(_3608_));
 sg13g2_inv_1 _8582_ (.Y(_3609_),
    .A(_3608_));
 sg13g2_nand2_1 _8583_ (.Y(_3610_),
    .A(_3607_),
    .B(_3609_));
 sg13g2_o21ai_1 _8584_ (.B1(_3567_),
    .Y(_3611_),
    .A1(_2875_),
    .A2(_0841_));
 sg13g2_nand2_1 _8585_ (.Y(_3612_),
    .A(_3569_),
    .B(_3611_));
 sg13g2_nand2_1 _8586_ (.Y(_3613_),
    .A(_3612_),
    .B(_3604_));
 sg13g2_nand2_1 _8587_ (.Y(_3614_),
    .A(_3613_),
    .B(_3606_));
 sg13g2_xnor2_1 _8588_ (.Y(_3615_),
    .A(_1802_),
    .B(_3614_));
 sg13g2_nor2_1 _8589_ (.A(_1638_),
    .B(_3603_),
    .Y(_3616_));
 sg13g2_xnor2_1 _8590_ (.Y(_3617_),
    .A(_1638_),
    .B(_3603_));
 sg13g2_nor3_1 _8591_ (.A(\vgademo.audio_snare_frames[1] ),
    .B(_0840_),
    .C(_3617_),
    .Y(_3618_));
 sg13g2_nor2_1 _8592_ (.A(_3616_),
    .B(_3618_),
    .Y(_3619_));
 sg13g2_inv_1 _8593_ (.Y(_3620_),
    .A(_3619_));
 sg13g2_nor2_1 _8594_ (.A(_1636_),
    .B(_3614_),
    .Y(_3621_));
 sg13g2_a21oi_1 _8595_ (.A1(_3615_),
    .A2(_3620_),
    .Y(_3622_),
    .B1(_3621_));
 sg13g2_nor2_1 _8596_ (.A(_3610_),
    .B(_3622_),
    .Y(_3623_));
 sg13g2_xnor2_1 _8597_ (.Y(_3624_),
    .A(_3574_),
    .B(_3580_));
 sg13g2_buf_2 _8598_ (.A(_3624_),
    .X(_3625_));
 sg13g2_nand2_1 _8599_ (.Y(_3626_),
    .A(_3623_),
    .B(_3625_));
 sg13g2_nor2_1 _8600_ (.A(_3601_),
    .B(_3626_),
    .Y(_3627_));
 sg13g2_inv_1 _8601_ (.Y(_3628_),
    .A(_3627_));
 sg13g2_xor2_1 _8602_ (.B(_3585_),
    .A(_3586_),
    .X(_3629_));
 sg13g2_inv_1 _8603_ (.Y(_3630_),
    .A(_3629_));
 sg13g2_nor2_1 _8604_ (.A(_3628_),
    .B(_3630_),
    .Y(_3631_));
 sg13g2_inv_1 _8605_ (.Y(_3632_),
    .A(_3631_));
 sg13g2_xor2_1 _8606_ (.B(_3588_),
    .A(_3589_),
    .X(_3633_));
 sg13g2_inv_1 _8607_ (.Y(_3634_),
    .A(_3633_));
 sg13g2_nor2_2 _8608_ (.A(_3632_),
    .B(_3634_),
    .Y(_3635_));
 sg13g2_nor2b_1 _8609_ (.A(_3598_),
    .B_N(_3635_),
    .Y(_3636_));
 sg13g2_nand2_1 _8610_ (.Y(_3637_),
    .A(_3596_),
    .B(_3636_));
 sg13g2_inv_1 _8611_ (.Y(_3638_),
    .A(_3625_));
 sg13g2_nor2_1 _8612_ (.A(_3609_),
    .B(_3638_),
    .Y(_3639_));
 sg13g2_nand2_1 _8613_ (.Y(_3640_),
    .A(_3600_),
    .B(_3639_));
 sg13g2_nor2_1 _8614_ (.A(_3640_),
    .B(_3630_),
    .Y(_3641_));
 sg13g2_inv_1 _8615_ (.Y(_3642_),
    .A(_3641_));
 sg13g2_nor2_1 _8616_ (.A(_3642_),
    .B(_3634_),
    .Y(_3643_));
 sg13g2_inv_1 _8617_ (.Y(_3644_),
    .A(_3643_));
 sg13g2_nor2_1 _8618_ (.A(_3644_),
    .B(_3598_),
    .Y(_3645_));
 sg13g2_nand2_1 _8619_ (.Y(_3646_),
    .A(_3596_),
    .B(_3645_));
 sg13g2_a21oi_1 _8620_ (.A1(_3503_),
    .A2(\vgademo.linelfsr[11] ),
    .Y(_3647_),
    .B1(_3502_));
 sg13g2_xor2_1 _8621_ (.B(\vgademo.linelfsr[12] ),
    .A(_4317_),
    .X(_3648_));
 sg13g2_nand2_1 _8622_ (.Y(_3649_),
    .A(_4312_),
    .B(net115));
 sg13g2_xnor2_1 _8623_ (.Y(_3650_),
    .A(_3501_),
    .B(_3649_));
 sg13g2_xnor2_1 _8624_ (.Y(_3651_),
    .A(_3648_),
    .B(_3650_));
 sg13g2_xnor2_1 _8625_ (.Y(_3652_),
    .A(_3647_),
    .B(_3651_));
 sg13g2_nor2_1 _8626_ (.A(_3500_),
    .B(_3505_),
    .Y(_3653_));
 sg13g2_nor2_1 _8627_ (.A(_4335_),
    .B(_3506_),
    .Y(_3654_));
 sg13g2_nor2_1 _8628_ (.A(_3653_),
    .B(_3654_),
    .Y(_3655_));
 sg13g2_xnor2_1 _8629_ (.Y(_3656_),
    .A(_3652_),
    .B(_3655_));
 sg13g2_a21oi_1 _8630_ (.A1(_3594_),
    .A2(_3509_),
    .Y(_3657_),
    .B1(_3508_));
 sg13g2_xor2_1 _8631_ (.B(_3657_),
    .A(_3656_),
    .X(_3658_));
 sg13g2_xnor2_1 _8632_ (.Y(_3659_),
    .A(_3646_),
    .B(_3658_));
 sg13g2_xor2_1 _8633_ (.B(_3659_),
    .A(_3637_),
    .X(_3660_));
 sg13g2_xnor2_1 _8634_ (.Y(_3661_),
    .A(_4288_),
    .B(_3660_));
 sg13g2_nor4_1 _8635_ (.A(_3634_),
    .B(_3630_),
    .C(_3598_),
    .D(_3595_),
    .Y(_3662_));
 sg13g2_nor4_1 _8636_ (.A(_3612_),
    .B(_3602_),
    .C(_3638_),
    .D(_3601_),
    .Y(_3663_));
 sg13g2_nand3_1 _8637_ (.B(_3603_),
    .C(_3663_),
    .A(_3662_),
    .Y(_3664_));
 sg13g2_xnor2_1 _8638_ (.Y(_3665_),
    .A(_3644_),
    .B(_3597_));
 sg13g2_xnor2_1 _8639_ (.Y(_3666_),
    .A(_3642_),
    .B(_3633_));
 sg13g2_nand2_1 _8640_ (.Y(_3667_),
    .A(_3665_),
    .B(_3666_));
 sg13g2_xor2_1 _8641_ (.B(_3595_),
    .A(_3645_),
    .X(_3668_));
 sg13g2_nor3_1 _8642_ (.A(_3667_),
    .B(_3668_),
    .C(_3659_),
    .Y(_3669_));
 sg13g2_inv_1 _8643_ (.Y(_3670_),
    .A(_3640_));
 sg13g2_nand3_1 _8644_ (.B(_3609_),
    .C(_3607_),
    .A(_3625_),
    .Y(_3671_));
 sg13g2_nor2_1 _8645_ (.A(_3639_),
    .B(_3600_),
    .Y(_3672_));
 sg13g2_nor4_1 _8646_ (.A(_3670_),
    .B(_3671_),
    .C(_3672_),
    .D(_3630_),
    .Y(_3673_));
 sg13g2_nand3b_1 _8647_ (.B(_3669_),
    .C(_3673_),
    .Y(_3674_),
    .A_N(_3622_));
 sg13g2_o21ai_1 _8648_ (.B1(_3674_),
    .Y(_3675_),
    .A1(_3658_),
    .A2(_3664_));
 sg13g2_nor2_1 _8649_ (.A(_3661_),
    .B(_3675_),
    .Y(_3676_));
 sg13g2_xor2_1 _8650_ (.B(_3668_),
    .A(_3636_),
    .X(_3677_));
 sg13g2_xnor2_1 _8651_ (.Y(_3678_),
    .A(_4437_),
    .B(_3677_));
 sg13g2_inv_1 _8652_ (.Y(_3679_),
    .A(_3678_));
 sg13g2_nor2_1 _8653_ (.A(_3631_),
    .B(_3666_),
    .Y(_3680_));
 sg13g2_nor3_1 _8654_ (.A(_4281_),
    .B(_3635_),
    .C(_3680_),
    .Y(_3681_));
 sg13g2_xnor2_1 _8655_ (.Y(_3682_),
    .A(_3640_),
    .B(_3629_));
 sg13g2_xnor2_1 _8656_ (.Y(_3683_),
    .A(_3627_),
    .B(_3682_));
 sg13g2_nand2b_1 _8657_ (.Y(_3684_),
    .B(_4421_),
    .A_N(_3683_));
 sg13g2_inv_1 _8658_ (.Y(_3685_),
    .A(_4421_));
 sg13g2_a21oi_2 _8659_ (.B1(_3639_),
    .Y(_3686_),
    .A2(_3625_),
    .A1(_3623_));
 sg13g2_a21oi_1 _8660_ (.A1(_3686_),
    .A2(_3600_),
    .Y(_3687_),
    .B1(_4476_));
 sg13g2_o21ai_1 _8661_ (.B1(_3687_),
    .Y(_3688_),
    .A1(_3600_),
    .A2(_3686_));
 sg13g2_xor2_1 _8662_ (.B(_3622_),
    .A(_3610_),
    .X(_3689_));
 sg13g2_nor2_1 _8663_ (.A(_2810_),
    .B(_3689_),
    .Y(_3690_));
 sg13g2_nor3_1 _8664_ (.A(_3608_),
    .B(_3625_),
    .C(_3623_),
    .Y(_3691_));
 sg13g2_nand2b_1 _8665_ (.Y(_3692_),
    .B(_3686_),
    .A_N(_3691_));
 sg13g2_nand2_1 _8666_ (.Y(_3693_),
    .A(_3692_),
    .B(_4412_));
 sg13g2_nand2_1 _8667_ (.Y(_3694_),
    .A(_0840_),
    .B(net127));
 sg13g2_nor2_1 _8668_ (.A(net127),
    .B(_0840_),
    .Y(_3695_));
 sg13g2_a21oi_1 _8669_ (.A1(_3694_),
    .A2(_1758_),
    .Y(_3696_),
    .B1(_3695_));
 sg13g2_a21o_1 _8670_ (.A2(_3696_),
    .A1(net126),
    .B1(_3617_),
    .X(_3697_));
 sg13g2_inv_1 _8671_ (.Y(_3698_),
    .A(net126));
 sg13g2_nand2b_1 _8672_ (.Y(_3699_),
    .B(_3698_),
    .A_N(_3696_));
 sg13g2_a21oi_1 _8673_ (.A1(_3697_),
    .A2(_3699_),
    .Y(_3700_),
    .B1(_3618_));
 sg13g2_xnor2_1 _8674_ (.Y(_3701_),
    .A(_3619_),
    .B(_3615_));
 sg13g2_inv_1 _8675_ (.Y(_3702_),
    .A(_3701_));
 sg13g2_nor3_1 _8676_ (.A(_4405_),
    .B(_3700_),
    .C(_3702_),
    .Y(_3703_));
 sg13g2_nand2b_1 _8677_ (.Y(_3704_),
    .B(_4405_),
    .A_N(_3700_));
 sg13g2_a21oi_1 _8678_ (.A1(_4279_),
    .A2(_3704_),
    .Y(_3705_),
    .B1(_3701_));
 sg13g2_nand2_1 _8679_ (.Y(_3706_),
    .A(_3689_),
    .B(_2810_));
 sg13g2_o21ai_1 _8680_ (.B1(_3706_),
    .Y(_3707_),
    .A1(_3703_),
    .A2(_3705_));
 sg13g2_nand3b_1 _8681_ (.B(_3693_),
    .C(_3707_),
    .Y(_3708_),
    .A_N(_3690_));
 sg13g2_xnor2_1 _8682_ (.Y(_3709_),
    .A(_4419_),
    .B(_3600_));
 sg13g2_xnor2_1 _8683_ (.Y(_3710_),
    .A(_3686_),
    .B(_3709_));
 sg13g2_nand2b_1 _8684_ (.Y(_3711_),
    .B(_4411_),
    .A_N(_3692_));
 sg13g2_nand3_1 _8685_ (.B(_3710_),
    .C(_3711_),
    .A(_3708_),
    .Y(_3712_));
 sg13g2_a22oi_1 _8686_ (.Y(_3713_),
    .B1(_3688_),
    .B2(_3712_),
    .A2(_3683_),
    .A1(_3685_));
 sg13g2_a22oi_1 _8687_ (.Y(_3714_),
    .B1(_3684_),
    .B2(_3713_),
    .A2(_3683_),
    .A1(net124));
 sg13g2_o21ai_1 _8688_ (.B1(_4281_),
    .Y(_3715_),
    .A1(_3635_),
    .A2(_3680_));
 sg13g2_o21ai_1 _8689_ (.B1(_3715_),
    .Y(_3716_),
    .A1(_3681_),
    .A2(_3714_));
 sg13g2_xnor2_1 _8690_ (.Y(_3717_),
    .A(_3635_),
    .B(_3665_));
 sg13g2_xnor2_1 _8691_ (.Y(_3718_),
    .A(_0079_),
    .B(_3717_));
 sg13g2_nand4_1 _8692_ (.B(_3679_),
    .C(_3716_),
    .A(_3676_),
    .Y(_3719_),
    .D(_3718_));
 sg13g2_nand2_1 _8693_ (.Y(_3720_),
    .A(_3717_),
    .B(_4434_));
 sg13g2_nand2_1 _8694_ (.Y(_3721_),
    .A(_3677_),
    .B(_4289_));
 sg13g2_o21ai_1 _8695_ (.B1(_3721_),
    .Y(_3722_),
    .A1(_3720_),
    .A2(_3678_));
 sg13g2_nor3_1 _8696_ (.A(_4462_),
    .B(_3660_),
    .C(_3675_),
    .Y(_3723_));
 sg13g2_a21oi_1 _8697_ (.A1(_3676_),
    .A2(_3722_),
    .Y(_3724_),
    .B1(_3723_));
 sg13g2_nor2_1 _8698_ (.A(_3462_),
    .B(_3461_),
    .Y(_3725_));
 sg13g2_o21ai_1 _8699_ (.B1(_3467_),
    .Y(_3726_),
    .A1(_3464_),
    .A2(_3725_));
 sg13g2_xor2_1 _8700_ (.B(_3476_),
    .A(_0060_),
    .X(_3727_));
 sg13g2_xnor2_1 _8701_ (.Y(_3728_),
    .A(_3453_),
    .B(_3450_));
 sg13g2_nor2_1 _8702_ (.A(_3434_),
    .B(_3458_),
    .Y(_3729_));
 sg13g2_xnor2_1 _8703_ (.Y(_3730_),
    .A(_3729_),
    .B(_3456_));
 sg13g2_nor2_1 _8704_ (.A(_3728_),
    .B(_3730_),
    .Y(_3731_));
 sg13g2_xnor2_1 _8705_ (.Y(_3732_),
    .A(_3432_),
    .B(_3460_));
 sg13g2_nor2_1 _8706_ (.A(_3468_),
    .B(_3732_),
    .Y(_3733_));
 sg13g2_nand3b_1 _8707_ (.B(_3731_),
    .C(_3733_),
    .Y(_3734_),
    .A_N(_3727_));
 sg13g2_a21oi_1 _8708_ (.A1(_3734_),
    .A2(_3467_),
    .Y(_3735_),
    .B1(_3479_));
 sg13g2_nor2_1 _8709_ (.A(_4461_),
    .B(_3658_),
    .Y(_3736_));
 sg13g2_xnor2_1 _8710_ (.Y(_3737_),
    .A(_4442_),
    .B(_3658_));
 sg13g2_nor3_1 _8711_ (.A(_4437_),
    .B(_3595_),
    .C(_3737_),
    .Y(_3738_));
 sg13g2_nor2_1 _8712_ (.A(_4427_),
    .B(_3634_),
    .Y(_3739_));
 sg13g2_xnor2_1 _8713_ (.Y(_3740_),
    .A(_4434_),
    .B(_3597_));
 sg13g2_a22oi_1 _8714_ (.Y(_3741_),
    .B1(_3739_),
    .B2(_3740_),
    .A2(_3597_),
    .A1(_4399_));
 sg13g2_xnor2_1 _8715_ (.Y(_3742_),
    .A(_0057_),
    .B(_3595_));
 sg13g2_nor2b_1 _8716_ (.A(_3737_),
    .B_N(_3742_),
    .Y(_3743_));
 sg13g2_inv_1 _8717_ (.Y(_3744_),
    .A(_3743_));
 sg13g2_nor2_1 _8718_ (.A(_3741_),
    .B(_3744_),
    .Y(_3745_));
 sg13g2_nor3_1 _8719_ (.A(_3736_),
    .B(_3738_),
    .C(_3745_),
    .Y(_3746_));
 sg13g2_o21ai_1 _8720_ (.B1(_3740_),
    .Y(_3747_),
    .A1(_0056_),
    .A2(_3633_));
 sg13g2_nor3_1 _8721_ (.A(_3739_),
    .B(_3747_),
    .C(_3744_),
    .Y(_3748_));
 sg13g2_nor2_1 _8722_ (.A(_4419_),
    .B(_3601_),
    .Y(_3749_));
 sg13g2_xnor2_1 _8723_ (.Y(_3750_),
    .A(_3685_),
    .B(_3629_));
 sg13g2_nor2_1 _8724_ (.A(_4408_),
    .B(_3602_),
    .Y(_3751_));
 sg13g2_xnor2_1 _8725_ (.Y(_3752_),
    .A(_4411_),
    .B(_3625_));
 sg13g2_inv_1 _8726_ (.Y(_3753_),
    .A(_3752_));
 sg13g2_a22oi_1 _8727_ (.Y(_3754_),
    .B1(_3751_),
    .B2(_3753_),
    .A2(_3625_),
    .A1(_4417_));
 sg13g2_nand2_1 _8728_ (.Y(_3755_),
    .A(_3750_),
    .B(_3709_));
 sg13g2_nor2_1 _8729_ (.A(_3754_),
    .B(_3755_),
    .Y(_3756_));
 sg13g2_a221oi_1 _8730_ (.B2(_3750_),
    .C1(_3756_),
    .B1(_3749_),
    .A1(_4428_),
    .Y(_3757_),
    .A2(_3629_));
 sg13g2_nor2_1 _8731_ (.A(_3752_),
    .B(_3755_),
    .Y(_3758_));
 sg13g2_xnor2_1 _8732_ (.Y(_3759_),
    .A(_4405_),
    .B(_3612_));
 sg13g2_inv_1 _8733_ (.Y(_3760_),
    .A(_0066_));
 sg13g2_nor2_1 _8734_ (.A(_3760_),
    .B(_3604_),
    .Y(_3761_));
 sg13g2_inv_1 _8735_ (.Y(_3762_),
    .A(_3761_));
 sg13g2_nand2_1 _8736_ (.Y(_3763_),
    .A(_3604_),
    .B(_3760_));
 sg13g2_nand4_1 _8737_ (.B(_3694_),
    .C(_3762_),
    .A(_3759_),
    .Y(_3764_),
    .D(_3763_));
 sg13g2_nand3_1 _8738_ (.B(_4279_),
    .C(_3611_),
    .A(_3569_),
    .Y(_3765_));
 sg13g2_nand2_1 _8739_ (.Y(_3766_),
    .A(_3759_),
    .B(_3761_));
 sg13g2_nand3_1 _8740_ (.B(_3765_),
    .C(_3766_),
    .A(_3764_),
    .Y(_3767_));
 sg13g2_xnor2_1 _8741_ (.Y(_3768_),
    .A(_0052_),
    .B(_3602_));
 sg13g2_nand3_1 _8742_ (.B(_3767_),
    .C(_3768_),
    .A(_3758_),
    .Y(_3769_));
 sg13g2_nand2_1 _8743_ (.Y(_3770_),
    .A(_3757_),
    .B(_3769_));
 sg13g2_nand2_1 _8744_ (.Y(_3771_),
    .A(_3748_),
    .B(_3770_));
 sg13g2_nand2_1 _8745_ (.Y(_3772_),
    .A(_3746_),
    .B(_3771_));
 sg13g2_nor2_1 _8746_ (.A(_3695_),
    .B(_3764_),
    .Y(_3773_));
 sg13g2_nand4_1 _8747_ (.B(_3758_),
    .C(_3768_),
    .A(_3748_),
    .Y(_3774_),
    .D(_3773_));
 sg13g2_a22oi_1 _8748_ (.Y(_3775_),
    .B1(_3772_),
    .B2(_3774_),
    .A2(_3735_),
    .A1(_3726_));
 sg13g2_nand3_1 _8749_ (.B(_3724_),
    .C(_3775_),
    .A(_3719_),
    .Y(_3776_));
 sg13g2_buf_1 _8750_ (.A(_3776_),
    .X(_3777_));
 sg13g2_nand2_1 _8751_ (.Y(_3778_),
    .A(_3777_),
    .B(net23));
 sg13g2_inv_1 _8752_ (.Y(_3779_),
    .A(_3778_));
 sg13g2_nand2b_1 _8753_ (.Y(_3780_),
    .B(_3779_),
    .A_N(_3482_));
 sg13g2_nand3_1 _8754_ (.B(net11),
    .C(_3780_),
    .A(_3383_),
    .Y(_3781_));
 sg13g2_xor2_1 _8755_ (.B(_1979_),
    .A(net125),
    .X(_3782_));
 sg13g2_xor2_1 _8756_ (.B(_1981_),
    .A(net123),
    .X(_3783_));
 sg13g2_nor2_1 _8757_ (.A(\vgademo.scanline_audio_sample[6] ),
    .B(_4428_),
    .Y(_3784_));
 sg13g2_inv_1 _8758_ (.Y(_3785_),
    .A(_2005_));
 sg13g2_nor2_1 _8759_ (.A(_4285_),
    .B(_3785_),
    .Y(_3786_));
 sg13g2_inv_1 _8760_ (.Y(_3787_),
    .A(\vgademo.scanline_audio_sample[6] ));
 sg13g2_nor2_1 _8761_ (.A(net124),
    .B(_3787_),
    .Y(_3788_));
 sg13g2_nor3_1 _8762_ (.A(_3784_),
    .B(_3786_),
    .C(_3788_),
    .Y(_3789_));
 sg13g2_o21ai_1 _8763_ (.B1(_3789_),
    .Y(_3790_),
    .A1(_4476_),
    .A2(_2005_));
 sg13g2_nor3_1 _8764_ (.A(_3782_),
    .B(_3783_),
    .C(_3790_),
    .Y(_3791_));
 sg13g2_inv_1 _8765_ (.Y(_3792_),
    .A(\vgademo.scanline_audio_sample[1] ));
 sg13g2_nor2_1 _8766_ (.A(net126),
    .B(_3792_),
    .Y(_3793_));
 sg13g2_a21oi_1 _8767_ (.A1(net127),
    .A2(_1631_),
    .Y(_3794_),
    .B1(_3793_));
 sg13g2_o21ai_1 _8768_ (.B1(_3794_),
    .Y(_3795_),
    .A1(_3698_),
    .A2(\vgademo.scanline_audio_sample[1] ));
 sg13g2_nor2_1 _8769_ (.A(_4278_),
    .B(_1945_),
    .Y(_3796_));
 sg13g2_nor2_1 _8770_ (.A(_3793_),
    .B(_3796_),
    .Y(_3797_));
 sg13g2_nor2_1 _8771_ (.A(\vgademo.scanline_audio_sample[2] ),
    .B(_4279_),
    .Y(_3798_));
 sg13g2_a21oi_1 _8772_ (.A1(_3795_),
    .A2(_3797_),
    .Y(_3799_),
    .B1(_3798_));
 sg13g2_inv_1 _8773_ (.Y(_3800_),
    .A(_1979_));
 sg13g2_nor3_1 _8774_ (.A(net125),
    .B(_3800_),
    .C(_3783_),
    .Y(_3801_));
 sg13g2_a21oi_1 _8775_ (.A1(_4417_),
    .A2(_1981_),
    .Y(_3802_),
    .B1(_3801_));
 sg13g2_inv_1 _8776_ (.Y(_3803_),
    .A(_3784_));
 sg13g2_o21ai_1 _8777_ (.B1(_3803_),
    .Y(_3804_),
    .A1(_3786_),
    .A2(_3788_));
 sg13g2_o21ai_1 _8778_ (.B1(_3804_),
    .Y(_3805_),
    .A1(_3790_),
    .A2(_3802_));
 sg13g2_a21oi_1 _8779_ (.A1(_3791_),
    .A2(_3799_),
    .Y(_3806_),
    .B1(_3805_));
 sg13g2_nor2_1 _8780_ (.A(_3798_),
    .B(_3796_),
    .Y(_3807_));
 sg13g2_o21ai_1 _8781_ (.B1(_3807_),
    .Y(_3808_),
    .A1(net127),
    .A2(_1631_));
 sg13g2_nand3_1 _8782_ (.B(_4282_),
    .C(_4288_),
    .A(_4290_),
    .Y(_3809_));
 sg13g2_nor3_1 _8783_ (.A(_3808_),
    .B(_3809_),
    .C(_3795_),
    .Y(_3810_));
 sg13g2_nand2_1 _8784_ (.Y(_3811_),
    .A(_3791_),
    .B(_3810_));
 sg13g2_nor3_1 _8785_ (.A(_4281_),
    .B(_4461_),
    .C(_4291_),
    .Y(_3812_));
 sg13g2_nand3b_1 _8786_ (.B(_3811_),
    .C(_3812_),
    .Y(_3813_),
    .A_N(_3806_));
 sg13g2_buf_2 _8787_ (.A(_3813_),
    .X(_3814_));
 sg13g2_buf_1 _8788_ (.A(_3814_),
    .X(_3815_));
 sg13g2_xnor2_1 _8789_ (.Y(_3816_),
    .A(_4276_),
    .B(net99));
 sg13g2_nand3_1 _8790_ (.B(net47),
    .C(_3816_),
    .A(_3781_),
    .Y(_3817_));
 sg13g2_a21oi_1 _8791_ (.A1(_3467_),
    .A2(_3728_),
    .Y(_3818_),
    .B1(_3481_));
 sg13g2_inv_1 _8792_ (.Y(_3819_),
    .A(_3475_));
 sg13g2_nor2_1 _8793_ (.A(_4364_),
    .B(_3819_),
    .Y(_3820_));
 sg13g2_inv_1 _8794_ (.Y(_3821_),
    .A(_3820_));
 sg13g2_buf_8 _8795_ (.A(_3422_),
    .X(_3822_));
 sg13g2_a21oi_2 _8796_ (.B1(net12),
    .Y(_3823_),
    .A2(_3821_),
    .A1(_3779_));
 sg13g2_a21oi_1 _8797_ (.A1(net11),
    .A2(_3818_),
    .Y(_3824_),
    .B1(_3823_));
 sg13g2_nand2_1 _8798_ (.Y(_3825_),
    .A(_2875_),
    .B(_3227_));
 sg13g2_nand4_1 _8799_ (.B(_3264_),
    .C(_3378_),
    .A(_3377_),
    .Y(_3826_),
    .D(_3825_));
 sg13g2_a21oi_1 _8800_ (.A1(_0076_),
    .A2(net26),
    .Y(_3827_),
    .B1(_3365_));
 sg13g2_a21oi_1 _8801_ (.A1(_3826_),
    .A2(_3827_),
    .Y(_3828_),
    .B1(net14));
 sg13g2_inv_1 _8802_ (.Y(_3829_),
    .A(_3365_));
 sg13g2_nand2_1 _8803_ (.Y(_3830_),
    .A(net26),
    .B(_0074_));
 sg13g2_nand2_1 _8804_ (.Y(_3831_),
    .A(_3829_),
    .B(_3830_));
 sg13g2_inv_1 _8805_ (.Y(_3832_),
    .A(_3831_));
 sg13g2_xor2_1 _8806_ (.B(_3267_),
    .A(_3263_),
    .X(_3833_));
 sg13g2_nand3_1 _8807_ (.B(_3833_),
    .C(_3378_),
    .A(_3377_),
    .Y(_3834_));
 sg13g2_nand2_1 _8808_ (.Y(_3835_),
    .A(_3832_),
    .B(_3834_));
 sg13g2_nand2_1 _8809_ (.Y(_3836_),
    .A(net14),
    .B(_3835_));
 sg13g2_nand3b_1 _8810_ (.B(net21),
    .C(_3836_),
    .Y(_3837_),
    .A_N(_3828_));
 sg13g2_nand2b_1 _8811_ (.Y(_3838_),
    .B(_3837_),
    .A_N(_3824_));
 sg13g2_nand2_2 _8812_ (.Y(_3839_),
    .A(_3838_),
    .B(net47));
 sg13g2_nand2_1 _8813_ (.Y(_3840_),
    .A(_3781_),
    .B(net47));
 sg13g2_inv_1 _8814_ (.Y(_3841_),
    .A(_3816_));
 sg13g2_nand2_1 _8815_ (.Y(_3842_),
    .A(_3840_),
    .B(_3841_));
 sg13g2_inv_1 _8816_ (.Y(_3843_),
    .A(_3842_));
 sg13g2_a21oi_1 _8817_ (.A1(_3817_),
    .A2(_3839_),
    .Y(_3844_),
    .B1(_3843_));
 sg13g2_nor2_1 _8818_ (.A(_3332_),
    .B(_3365_),
    .Y(_3845_));
 sg13g2_nand2_1 _8819_ (.Y(_3846_),
    .A(_3378_),
    .B(_3273_));
 sg13g2_nand2_1 _8820_ (.Y(_3847_),
    .A(_3845_),
    .B(_3846_));
 sg13g2_nand2b_1 _8821_ (.Y(_3848_),
    .B(net14),
    .A_N(_3847_));
 sg13g2_nand2b_1 _8822_ (.Y(_3849_),
    .B(_3374_),
    .A_N(_3835_));
 sg13g2_nand3_1 _8823_ (.B(_3849_),
    .C(net21),
    .A(_3848_),
    .Y(_3850_));
 sg13g2_nand2_1 _8824_ (.Y(_3851_),
    .A(_3467_),
    .B(_3732_));
 sg13g2_nor2_1 _8825_ (.A(net22),
    .B(_3481_),
    .Y(_3852_));
 sg13g2_nand2_1 _8826_ (.Y(_3853_),
    .A(_3475_),
    .B(_0058_));
 sg13g2_a21oi_1 _8827_ (.A1(_3777_),
    .A2(_3853_),
    .Y(_3854_),
    .B1(net21));
 sg13g2_a21oi_1 _8828_ (.A1(_3851_),
    .A2(_3852_),
    .Y(_3855_),
    .B1(_3854_));
 sg13g2_nand2_1 _8829_ (.Y(_3856_),
    .A(_3850_),
    .B(_3855_));
 sg13g2_nand2_1 _8830_ (.Y(_3857_),
    .A(_3856_),
    .B(net11));
 sg13g2_xnor2_1 _8831_ (.Y(_3858_),
    .A(_2904_),
    .B(_2787_));
 sg13g2_xnor2_1 _8832_ (.Y(_3859_),
    .A(_2867_),
    .B(_3039_));
 sg13g2_nor2_1 _8833_ (.A(_2896_),
    .B(_3028_),
    .Y(_3860_));
 sg13g2_nand2b_1 _8834_ (.Y(_3861_),
    .B(_3860_),
    .A_N(_3859_));
 sg13g2_o21ai_1 _8835_ (.B1(_3861_),
    .Y(_3862_),
    .A1(_3039_),
    .A2(_2867_));
 sg13g2_xor2_1 _8836_ (.B(_3862_),
    .A(_3858_),
    .X(_3863_));
 sg13g2_xnor2_1 _8837_ (.Y(_3864_),
    .A(_3860_),
    .B(_3859_));
 sg13g2_nor2b_1 _8838_ (.A(_3863_),
    .B_N(_3864_),
    .Y(_3865_));
 sg13g2_inv_1 _8839_ (.Y(_3866_),
    .A(_3865_));
 sg13g2_inv_1 _8840_ (.Y(_3867_),
    .A(_3863_));
 sg13g2_nor2_1 _8841_ (.A(_3864_),
    .B(_3867_),
    .Y(_3868_));
 sg13g2_inv_1 _8842_ (.Y(_3869_),
    .A(_3868_));
 sg13g2_a21oi_1 _8843_ (.A1(_3866_),
    .A2(_3869_),
    .Y(_3870_),
    .B1(_3423_));
 sg13g2_xnor2_1 _8844_ (.Y(_3871_),
    .A(_2896_),
    .B(net18));
 sg13g2_inv_1 _8845_ (.Y(_3872_),
    .A(_3871_));
 sg13g2_nand2_1 _8846_ (.Y(_3873_),
    .A(_3870_),
    .B(_3872_));
 sg13g2_nand3_1 _8847_ (.B(_3814_),
    .C(_3873_),
    .A(_3857_),
    .Y(_3874_));
 sg13g2_buf_2 _8848_ (.A(_3874_),
    .X(_3875_));
 sg13g2_a21o_1 _8849_ (.A2(net26),
    .A1(_0073_),
    .B1(_3365_),
    .X(_3876_));
 sg13g2_inv_1 _8850_ (.Y(_3877_),
    .A(_3876_));
 sg13g2_nand2_1 _8851_ (.Y(_3878_),
    .A(_3377_),
    .B(_3353_));
 sg13g2_nand2_1 _8852_ (.Y(_3879_),
    .A(_3877_),
    .B(_3878_));
 sg13g2_nand2_1 _8853_ (.Y(_3880_),
    .A(net14),
    .B(_3879_));
 sg13g2_nand2_1 _8854_ (.Y(_3881_),
    .A(net13),
    .B(_3371_));
 sg13g2_nand3_1 _8855_ (.B(_3881_),
    .C(net21),
    .A(_3880_),
    .Y(_3882_));
 sg13g2_nor2_1 _8856_ (.A(_2853_),
    .B(_3819_),
    .Y(_3883_));
 sg13g2_nor2_1 _8857_ (.A(_3883_),
    .B(_3778_),
    .Y(_3884_));
 sg13g2_a21o_1 _8858_ (.A2(_3730_),
    .A1(_3467_),
    .B1(_3481_),
    .X(_3885_));
 sg13g2_a21oi_1 _8859_ (.A1(_3884_),
    .A2(_3885_),
    .Y(_3886_),
    .B1(net12));
 sg13g2_nand2_1 _8860_ (.Y(_3887_),
    .A(_3882_),
    .B(_3886_));
 sg13g2_inv_4 _8861_ (.A(_3814_),
    .Y(_3888_));
 sg13g2_a21oi_1 _8862_ (.A1(net12),
    .A2(_3867_),
    .Y(_3889_),
    .B1(net46));
 sg13g2_nand2_1 _8863_ (.Y(_3890_),
    .A(_3887_),
    .B(_3889_));
 sg13g2_xnor2_1 _8864_ (.Y(_3891_),
    .A(_0947_),
    .B(_3816_));
 sg13g2_inv_1 _8865_ (.Y(_3892_),
    .A(_3891_));
 sg13g2_nand2_1 _8866_ (.Y(_3893_),
    .A(_3890_),
    .B(_3892_));
 sg13g2_nand3_1 _8867_ (.B(_3889_),
    .C(_3891_),
    .A(_3887_),
    .Y(_3894_));
 sg13g2_nand2_1 _8868_ (.Y(_3895_),
    .A(_3893_),
    .B(_3894_));
 sg13g2_xor2_1 _8869_ (.B(_3895_),
    .A(_3875_),
    .X(_3896_));
 sg13g2_nor2_1 _8870_ (.A(_3844_),
    .B(_3896_),
    .Y(_3897_));
 sg13g2_nand2_1 _8871_ (.Y(_3898_),
    .A(_3842_),
    .B(_3817_));
 sg13g2_xor2_1 _8872_ (.B(_3898_),
    .A(_3839_),
    .X(_3899_));
 sg13g2_nand2_1 _8873_ (.Y(_3900_),
    .A(_3467_),
    .B(_3727_));
 sg13g2_nor2_1 _8874_ (.A(net23),
    .B(_3261_),
    .Y(_3901_));
 sg13g2_a22oi_1 _8875_ (.Y(_3902_),
    .B1(_3847_),
    .B2(_3901_),
    .A2(_3852_),
    .A1(_3900_));
 sg13g2_nor2_1 _8876_ (.A(_0806_),
    .B(_3819_),
    .Y(_3903_));
 sg13g2_inv_1 _8877_ (.Y(_3904_),
    .A(_3777_));
 sg13g2_o21ai_1 _8878_ (.B1(net23),
    .Y(_3905_),
    .A1(_3903_),
    .A2(_3904_));
 sg13g2_nand3_1 _8879_ (.B(net11),
    .C(_3905_),
    .A(_3902_),
    .Y(_3906_));
 sg13g2_nor2_1 _8880_ (.A(_3872_),
    .B(_3866_),
    .Y(_3907_));
 sg13g2_nor2_1 _8881_ (.A(_3907_),
    .B(_3423_),
    .Y(_3908_));
 sg13g2_nor2_1 _8882_ (.A(net46),
    .B(_3908_),
    .Y(_3909_));
 sg13g2_xnor2_1 _8883_ (.Y(_3910_),
    .A(_1981_),
    .B(_1979_));
 sg13g2_xnor2_1 _8884_ (.Y(_3911_),
    .A(_4411_),
    .B(_3910_));
 sg13g2_inv_1 _8885_ (.Y(_3912_),
    .A(_3911_));
 sg13g2_nand2_1 _8886_ (.Y(_3913_),
    .A(_3912_),
    .B(_3782_));
 sg13g2_inv_1 _8887_ (.Y(_3914_),
    .A(_3799_));
 sg13g2_nor2_1 _8888_ (.A(net125),
    .B(_1979_),
    .Y(_3915_));
 sg13g2_a22oi_1 _8889_ (.Y(_3916_),
    .B1(_3915_),
    .B2(_3912_),
    .A2(_3910_),
    .A1(_4417_));
 sg13g2_o21ai_1 _8890_ (.B1(_3916_),
    .Y(_3917_),
    .A1(_3913_),
    .A2(_3914_));
 sg13g2_nor2_1 _8891_ (.A(_1981_),
    .B(_1979_),
    .Y(_3918_));
 sg13g2_xnor2_1 _8892_ (.Y(_3919_),
    .A(_2005_),
    .B(_3918_));
 sg13g2_nor2_1 _8893_ (.A(_4419_),
    .B(_3919_),
    .Y(_3920_));
 sg13g2_nor2b_1 _8894_ (.A(_0054_),
    .B_N(_3919_),
    .Y(_3921_));
 sg13g2_nand2_1 _8895_ (.Y(_3922_),
    .A(_3918_),
    .B(_3785_));
 sg13g2_xnor2_1 _8896_ (.Y(_3923_),
    .A(_3787_),
    .B(_3922_));
 sg13g2_xnor2_1 _8897_ (.Y(_3924_),
    .A(_4421_),
    .B(_3923_));
 sg13g2_inv_1 _8898_ (.Y(_3925_),
    .A(_3924_));
 sg13g2_nor3_1 _8899_ (.A(_3920_),
    .B(_3921_),
    .C(_3925_),
    .Y(_3926_));
 sg13g2_nand2_1 _8900_ (.Y(_3927_),
    .A(_3924_),
    .B(_3920_));
 sg13g2_o21ai_1 _8901_ (.B1(_3927_),
    .Y(_3928_),
    .A1(net124),
    .A2(_3923_));
 sg13g2_a21oi_1 _8902_ (.A1(_3917_),
    .A2(_3926_),
    .Y(_3929_),
    .B1(_3928_));
 sg13g2_nand4_1 _8903_ (.B(_3782_),
    .C(_3810_),
    .A(_3926_),
    .Y(_3930_),
    .D(_3912_));
 sg13g2_nand3b_1 _8904_ (.B(_3812_),
    .C(_3930_),
    .Y(_3931_),
    .A_N(_3929_));
 sg13g2_nand2_2 _8905_ (.Y(_3932_),
    .A(_3931_),
    .B(net46));
 sg13g2_inv_1 _8906_ (.Y(_3933_),
    .A(_3932_));
 sg13g2_a21oi_1 _8907_ (.A1(_3906_),
    .A2(_3909_),
    .Y(_3934_),
    .B1(_3933_));
 sg13g2_buf_2 _8908_ (.A(_3934_),
    .X(_3935_));
 sg13g2_xor2_1 _8909_ (.B(net99),
    .A(_4278_),
    .X(_3936_));
 sg13g2_nand2_1 _8910_ (.Y(_3937_),
    .A(_3839_),
    .B(_3936_));
 sg13g2_nor2_1 _8911_ (.A(_3936_),
    .B(_3839_),
    .Y(_3938_));
 sg13g2_a21oi_1 _8912_ (.A1(_3935_),
    .A2(_3937_),
    .Y(_3939_),
    .B1(_3938_));
 sg13g2_nor2b_1 _8913_ (.A(_3899_),
    .B_N(_3939_),
    .Y(_3940_));
 sg13g2_nor2_1 _8914_ (.A(_3897_),
    .B(_3940_),
    .Y(_3941_));
 sg13g2_nand2_1 _8915_ (.Y(_3942_),
    .A(_3374_),
    .B(_3139_));
 sg13g2_nor2b_1 _8916_ (.A(_3942_),
    .B_N(_3879_),
    .Y(_3943_));
 sg13g2_nand2_1 _8917_ (.Y(_3944_),
    .A(_3475_),
    .B(_0802_));
 sg13g2_a21oi_1 _8918_ (.A1(_3777_),
    .A2(_3944_),
    .Y(_3945_),
    .B1(_3139_));
 sg13g2_nor2_1 _8919_ (.A(_3945_),
    .B(net12),
    .Y(_3946_));
 sg13g2_nand2_1 _8920_ (.Y(_3947_),
    .A(_3852_),
    .B(_3726_));
 sg13g2_nand2_1 _8921_ (.Y(_3948_),
    .A(_3946_),
    .B(_3947_));
 sg13g2_nor2_1 _8922_ (.A(_3943_),
    .B(_3948_),
    .Y(_3949_));
 sg13g2_o21ai_1 _8923_ (.B1(_3814_),
    .Y(_3950_),
    .A1(_3908_),
    .A2(_3949_));
 sg13g2_buf_2 _8924_ (.A(_3950_),
    .X(_3951_));
 sg13g2_inv_4 _8925_ (.A(_3875_),
    .Y(_3952_));
 sg13g2_xnor2_1 _8926_ (.Y(_3953_),
    .A(_4275_),
    .B(net99));
 sg13g2_nand2_1 _8927_ (.Y(_3954_),
    .A(_3952_),
    .B(_3953_));
 sg13g2_inv_1 _8928_ (.Y(_3955_),
    .A(_3953_));
 sg13g2_nand2_1 _8929_ (.Y(_3956_),
    .A(_3875_),
    .B(_3955_));
 sg13g2_nand2_1 _8930_ (.Y(_3957_),
    .A(_3954_),
    .B(_3956_));
 sg13g2_nand2b_1 _8931_ (.Y(_3958_),
    .B(_3957_),
    .A_N(_3951_));
 sg13g2_nand3_1 _8932_ (.B(_3956_),
    .C(_3951_),
    .A(_3954_),
    .Y(_3959_));
 sg13g2_inv_1 _8933_ (.Y(_3960_),
    .A(_3893_));
 sg13g2_a21oi_1 _8934_ (.A1(_3875_),
    .A2(_3894_),
    .Y(_3961_),
    .B1(_3960_));
 sg13g2_inv_1 _8935_ (.Y(_3962_),
    .A(_3961_));
 sg13g2_nand3_1 _8936_ (.B(_3959_),
    .C(_3962_),
    .A(_3958_),
    .Y(_3963_));
 sg13g2_nand2_1 _8937_ (.Y(_3964_),
    .A(_3896_),
    .B(_3844_));
 sg13g2_nand2_1 _8938_ (.Y(_3965_),
    .A(_3963_),
    .B(_3964_));
 sg13g2_nor2_1 _8939_ (.A(_3941_),
    .B(_3965_),
    .Y(_3966_));
 sg13g2_a21oi_1 _8940_ (.A1(_3958_),
    .A2(_3959_),
    .Y(_3967_),
    .B1(_3962_));
 sg13g2_xnor2_1 _8941_ (.Y(_3968_),
    .A(_0018_),
    .B(_3953_));
 sg13g2_inv_1 _8942_ (.Y(_3969_),
    .A(_3968_));
 sg13g2_nor2_1 _8943_ (.A(_3969_),
    .B(_3951_),
    .Y(_3970_));
 sg13g2_nand2_1 _8944_ (.Y(_3971_),
    .A(_3951_),
    .B(_3969_));
 sg13g2_nand2b_1 _8945_ (.Y(_3972_),
    .B(_3971_),
    .A_N(_3970_));
 sg13g2_xor2_1 _8946_ (.B(_3972_),
    .A(_3935_),
    .X(_3973_));
 sg13g2_inv_1 _8947_ (.Y(_3974_),
    .A(_3956_));
 sg13g2_a21oi_1 _8948_ (.A1(_3954_),
    .A2(_3951_),
    .Y(_3975_),
    .B1(_3974_));
 sg13g2_inv_1 _8949_ (.Y(_3976_),
    .A(_3975_));
 sg13g2_nand2_1 _8950_ (.Y(_3977_),
    .A(_3973_),
    .B(_3976_));
 sg13g2_xnor2_1 _8951_ (.Y(_3978_),
    .A(_3935_),
    .B(_3972_));
 sg13g2_nand2_1 _8952_ (.Y(_3979_),
    .A(_3978_),
    .B(_3975_));
 sg13g2_nand2_1 _8953_ (.Y(_3980_),
    .A(_3977_),
    .B(_3979_));
 sg13g2_nor2_1 _8954_ (.A(_3967_),
    .B(_3980_),
    .Y(_3981_));
 sg13g2_inv_1 _8955_ (.Y(_3982_),
    .A(_3979_));
 sg13g2_a21oi_1 _8956_ (.A1(_3963_),
    .A2(_3977_),
    .Y(_3983_),
    .B1(_3982_));
 sg13g2_a21oi_1 _8957_ (.A1(_3966_),
    .A2(_3981_),
    .Y(_3984_),
    .B1(_3983_));
 sg13g2_nand2b_1 _8958_ (.Y(_3985_),
    .B(_3963_),
    .A_N(_3897_));
 sg13g2_nor2b_1 _8959_ (.A(_3985_),
    .B_N(_3964_),
    .Y(_3986_));
 sg13g2_xor2_1 _8960_ (.B(_3899_),
    .A(_3939_),
    .X(_3987_));
 sg13g2_nor2b_1 _8961_ (.A(_3987_),
    .B_N(_3890_),
    .Y(_3988_));
 sg13g2_nand3_1 _8962_ (.B(_3988_),
    .C(_3981_),
    .A(_3986_),
    .Y(_3989_));
 sg13g2_nor2_1 _8963_ (.A(_3970_),
    .B(_3935_),
    .Y(_3990_));
 sg13g2_a21oi_1 _8964_ (.A1(_3935_),
    .A2(_3971_),
    .Y(_3991_),
    .B1(_3990_));
 sg13g2_inv_1 _8965_ (.Y(_3992_),
    .A(_3991_));
 sg13g2_a21oi_1 _8966_ (.A1(_3984_),
    .A2(_3989_),
    .Y(_3993_),
    .B1(_3992_));
 sg13g2_nand3_1 _8967_ (.B(_3989_),
    .C(_3992_),
    .A(_3984_),
    .Y(_3994_));
 sg13g2_nor4_1 _8968_ (.A(_4449_),
    .B(_0405_),
    .C(_0406_),
    .D(_2739_),
    .Y(_3995_));
 sg13g2_nand3b_1 _8969_ (.B(_1217_),
    .C(_2700_),
    .Y(_3996_),
    .A_N(_3995_));
 sg13g2_buf_1 _8970_ (.A(_3996_),
    .X(_3997_));
 sg13g2_inv_1 _8971_ (.Y(_3998_),
    .A(_3997_));
 sg13g2_nand2_1 _8972_ (.Y(_3999_),
    .A(_3994_),
    .B(_3998_));
 sg13g2_nor2_1 _8973_ (.A(_3993_),
    .B(_3999_),
    .Y(_0154_));
 sg13g2_or2_1 _8974_ (.X(_4000_),
    .B(_3988_),
    .A(_3940_));
 sg13g2_nand4_1 _8975_ (.B(_3981_),
    .C(_3986_),
    .A(_4000_),
    .Y(_4001_),
    .D(_3991_));
 sg13g2_a21oi_1 _8976_ (.A1(_3975_),
    .A2(_3970_),
    .Y(_4002_),
    .B1(_3935_));
 sg13g2_inv_1 _8977_ (.Y(_4003_),
    .A(_3985_));
 sg13g2_nor4_1 _8978_ (.A(_3967_),
    .B(_3992_),
    .C(_3980_),
    .D(_4003_),
    .Y(_4004_));
 sg13g2_nor2_1 _8979_ (.A(_4002_),
    .B(_4004_),
    .Y(_4005_));
 sg13g2_a21oi_1 _8980_ (.A1(_4001_),
    .A2(_4005_),
    .Y(_0155_),
    .B1(_3997_));
 sg13g2_o21ai_1 _8981_ (.B1(_3877_),
    .Y(_4006_),
    .A1(net26),
    .A2(_3846_));
 sg13g2_nand2_1 _8982_ (.Y(_4007_),
    .A(net14),
    .B(_4006_));
 sg13g2_nand2_1 _8983_ (.Y(_4008_),
    .A(_3367_),
    .B(_3834_));
 sg13g2_nand2_1 _8984_ (.Y(_4009_),
    .A(net13),
    .B(_4008_));
 sg13g2_nand3_1 _8985_ (.B(_4009_),
    .C(net21),
    .A(_4007_),
    .Y(_4010_));
 sg13g2_inv_1 _8986_ (.Y(_4011_),
    .A(_3884_));
 sg13g2_nand3_1 _8987_ (.B(net11),
    .C(_4011_),
    .A(_4010_),
    .Y(_4012_));
 sg13g2_nor2_1 _8988_ (.A(_3871_),
    .B(_3869_),
    .Y(_4013_));
 sg13g2_o21ai_1 _8989_ (.B1(net12),
    .Y(_4014_),
    .A1(_3907_),
    .A2(_4013_));
 sg13g2_nand2_1 _8990_ (.Y(_4015_),
    .A(_4012_),
    .B(_4014_));
 sg13g2_nand2_1 _8991_ (.Y(_4016_),
    .A(_3832_),
    .B(_3878_));
 sg13g2_nor2_1 _8992_ (.A(_4016_),
    .B(net14),
    .Y(_4017_));
 sg13g2_nor2_1 _8993_ (.A(_3322_),
    .B(_3356_),
    .Y(_4018_));
 sg13g2_inv_1 _8994_ (.Y(_4019_),
    .A(_4018_));
 sg13g2_a21oi_1 _8995_ (.A1(_3845_),
    .A2(_4019_),
    .Y(_4020_),
    .B1(net23));
 sg13g2_nor2_1 _8996_ (.A(_4020_),
    .B(_3901_),
    .Y(_4021_));
 sg13g2_inv_1 _8997_ (.Y(_4022_),
    .A(_3854_));
 sg13g2_o21ai_1 _8998_ (.B1(_4022_),
    .Y(_4023_),
    .A1(_4017_),
    .A2(_4021_));
 sg13g2_nor2_1 _8999_ (.A(net46),
    .B(_3870_),
    .Y(_4024_));
 sg13g2_inv_1 _9000_ (.Y(_4025_),
    .A(_4024_));
 sg13g2_a21oi_1 _9001_ (.A1(_4023_),
    .A2(net11),
    .Y(_4026_),
    .B1(_4025_));
 sg13g2_nand2b_1 _9002_ (.Y(_4027_),
    .B(_4026_),
    .A_N(_4015_));
 sg13g2_nand3_1 _9003_ (.B(net47),
    .C(_4014_),
    .A(_4012_),
    .Y(_4028_));
 sg13g2_nand2_1 _9004_ (.Y(_4029_),
    .A(_4023_),
    .B(net11));
 sg13g2_nand2_1 _9005_ (.Y(_4030_),
    .A(_4029_),
    .B(_4024_));
 sg13g2_nand2_1 _9006_ (.Y(_4031_),
    .A(_4028_),
    .B(_4030_));
 sg13g2_inv_1 _9007_ (.Y(_4032_),
    .A(_4031_));
 sg13g2_a21oi_1 _9008_ (.A1(_4027_),
    .A2(_3892_),
    .Y(_4033_),
    .B1(_4032_));
 sg13g2_inv_1 _9009_ (.Y(_4034_),
    .A(_4033_));
 sg13g2_nand2_1 _9010_ (.Y(_4035_),
    .A(_3901_),
    .B(_4006_));
 sg13g2_nand2_1 _9011_ (.Y(_4036_),
    .A(_4035_),
    .B(_3946_));
 sg13g2_inv_1 _9012_ (.Y(_4037_),
    .A(_3864_));
 sg13g2_a21oi_1 _9013_ (.A1(_3872_),
    .A2(_4037_),
    .Y(_4038_),
    .B1(_3867_));
 sg13g2_nor2_1 _9014_ (.A(_4038_),
    .B(_3424_),
    .Y(_4039_));
 sg13g2_nand2_1 _9015_ (.Y(_4040_),
    .A(_4039_),
    .B(_3866_));
 sg13g2_a21oi_2 _9016_ (.B1(net46),
    .Y(_4041_),
    .A2(_4040_),
    .A1(_4036_));
 sg13g2_inv_2 _9017_ (.Y(_4042_),
    .A(_4041_));
 sg13g2_nand2_1 _9018_ (.Y(_4043_),
    .A(_4030_),
    .B(_4042_));
 sg13g2_nand3_1 _9019_ (.B(_4024_),
    .C(_4041_),
    .A(_4029_),
    .Y(_4044_));
 sg13g2_nand3_1 _9020_ (.B(_4044_),
    .C(_3955_),
    .A(_4043_),
    .Y(_4045_));
 sg13g2_nand2_1 _9021_ (.Y(_4046_),
    .A(_4043_),
    .B(_4044_));
 sg13g2_nand2_1 _9022_ (.Y(_4047_),
    .A(_4046_),
    .B(_3953_));
 sg13g2_nand3_1 _9023_ (.B(_4045_),
    .C(_4047_),
    .A(_4034_),
    .Y(_4048_));
 sg13g2_nand2_1 _9024_ (.Y(_4049_),
    .A(_3375_),
    .B(_4020_));
 sg13g2_a21oi_1 _9025_ (.A1(_4049_),
    .A2(_3905_),
    .Y(_4050_),
    .B1(net12));
 sg13g2_o21ai_1 _9026_ (.B1(_3815_),
    .Y(_4051_),
    .A1(_4039_),
    .A2(_4050_));
 sg13g2_nand2_1 _9027_ (.Y(_4052_),
    .A(_4051_),
    .B(_3932_));
 sg13g2_nand2_1 _9028_ (.Y(_4053_),
    .A(_4052_),
    .B(_4042_));
 sg13g2_nand3_1 _9029_ (.B(_4041_),
    .C(_3932_),
    .A(_4051_),
    .Y(_4054_));
 sg13g2_nand2_1 _9030_ (.Y(_4055_),
    .A(_4053_),
    .B(_4054_));
 sg13g2_nand2_1 _9031_ (.Y(_4056_),
    .A(_4055_),
    .B(_3968_));
 sg13g2_nand3_1 _9032_ (.B(_4054_),
    .C(_3969_),
    .A(_4053_),
    .Y(_4057_));
 sg13g2_nand2_1 _9033_ (.Y(_4058_),
    .A(_4056_),
    .B(_4057_));
 sg13g2_nor2_1 _9034_ (.A(_4041_),
    .B(_4026_),
    .Y(_4059_));
 sg13g2_a21oi_1 _9035_ (.A1(_4044_),
    .A2(_3955_),
    .Y(_4060_),
    .B1(_4059_));
 sg13g2_nand2_1 _9036_ (.Y(_4061_),
    .A(_4058_),
    .B(_4060_));
 sg13g2_nor2b_1 _9037_ (.A(_4048_),
    .B_N(_4061_),
    .Y(_4062_));
 sg13g2_inv_1 _9038_ (.Y(_4063_),
    .A(_4060_));
 sg13g2_nand3_1 _9039_ (.B(_4056_),
    .C(_4057_),
    .A(_4063_),
    .Y(_4064_));
 sg13g2_buf_1 _9040_ (.A(_4064_),
    .X(_4065_));
 sg13g2_nand2b_1 _9041_ (.Y(_4066_),
    .B(_4065_),
    .A_N(_4062_));
 sg13g2_nand2_1 _9042_ (.Y(_4067_),
    .A(_4031_),
    .B(_4027_));
 sg13g2_nand2_1 _9043_ (.Y(_4068_),
    .A(_4067_),
    .B(_3891_));
 sg13g2_nand3_1 _9044_ (.B(_4027_),
    .C(_3892_),
    .A(_4031_),
    .Y(_4069_));
 sg13g2_nand2_1 _9045_ (.Y(_4070_),
    .A(_4068_),
    .B(_4069_));
 sg13g2_inv_1 _9046_ (.Y(_4071_),
    .A(_4016_));
 sg13g2_nand2_1 _9047_ (.Y(_4072_),
    .A(_3827_),
    .B(_3370_));
 sg13g2_a21oi_1 _9048_ (.A1(net13),
    .A2(_4072_),
    .Y(_4073_),
    .B1(net23));
 sg13g2_o21ai_1 _9049_ (.B1(_4073_),
    .Y(_4074_),
    .A1(net13),
    .A2(_4071_));
 sg13g2_nand2_1 _9050_ (.Y(_4075_),
    .A(_4074_),
    .B(_3823_));
 sg13g2_nand2_1 _9051_ (.Y(_4076_),
    .A(net14),
    .B(_4008_));
 sg13g2_nand2_1 _9052_ (.Y(_4077_),
    .A(_3376_),
    .B(_3826_));
 sg13g2_nand2_1 _9053_ (.Y(_4078_),
    .A(net13),
    .B(_4077_));
 sg13g2_nand3_1 _9054_ (.B(_4078_),
    .C(net21),
    .A(_4076_),
    .Y(_4079_));
 sg13g2_nor2_1 _9055_ (.A(_3779_),
    .B(net12),
    .Y(_4080_));
 sg13g2_nand2_1 _9056_ (.Y(_4081_),
    .A(_4079_),
    .B(_4080_));
 sg13g2_nand2_1 _9057_ (.Y(_4082_),
    .A(_4075_),
    .B(_4081_));
 sg13g2_nand2_1 _9058_ (.Y(_4083_),
    .A(_4075_),
    .B(net47));
 sg13g2_nand2_1 _9059_ (.Y(_4084_),
    .A(_4081_),
    .B(net47));
 sg13g2_nand2_1 _9060_ (.Y(_4085_),
    .A(_4083_),
    .B(_4084_));
 sg13g2_inv_1 _9061_ (.Y(_4086_),
    .A(_4085_));
 sg13g2_a21oi_1 _9062_ (.A1(_4015_),
    .A2(_4082_),
    .Y(_4087_),
    .B1(_4086_));
 sg13g2_nand2_1 _9063_ (.Y(_4088_),
    .A(_4070_),
    .B(_4087_));
 sg13g2_nand3_1 _9064_ (.B(_4065_),
    .C(_4061_),
    .A(_4088_),
    .Y(_4089_));
 sg13g2_nand2_1 _9065_ (.Y(_4090_),
    .A(_4047_),
    .B(_4045_));
 sg13g2_xnor2_1 _9066_ (.Y(_4091_),
    .A(_4034_),
    .B(_4090_));
 sg13g2_inv_1 _9067_ (.Y(_4092_),
    .A(_4087_));
 sg13g2_nand3_1 _9068_ (.B(_4069_),
    .C(_4092_),
    .A(_4068_),
    .Y(_4093_));
 sg13g2_inv_1 _9069_ (.Y(_4094_),
    .A(_4028_));
 sg13g2_nand2_1 _9070_ (.Y(_4095_),
    .A(_4085_),
    .B(_4082_));
 sg13g2_xnor2_1 _9071_ (.Y(_4096_),
    .A(_4094_),
    .B(_4095_));
 sg13g2_inv_1 _9072_ (.Y(_4097_),
    .A(_4083_));
 sg13g2_inv_1 _9073_ (.Y(_4098_),
    .A(_3936_));
 sg13g2_nand2_1 _9074_ (.Y(_4099_),
    .A(_4097_),
    .B(_4098_));
 sg13g2_nor2_1 _9075_ (.A(_4098_),
    .B(_4097_),
    .Y(_4100_));
 sg13g2_a21oi_1 _9076_ (.A1(_4099_),
    .A2(_4052_),
    .Y(_4101_),
    .B1(_4100_));
 sg13g2_inv_1 _9077_ (.Y(_4102_),
    .A(_4101_));
 sg13g2_nand2b_1 _9078_ (.Y(_4103_),
    .B(_4102_),
    .A_N(_4096_));
 sg13g2_nand2_1 _9079_ (.Y(_4104_),
    .A(_4093_),
    .B(_4103_));
 sg13g2_nand2_1 _9080_ (.Y(_4105_),
    .A(_4091_),
    .B(_4104_));
 sg13g2_nor2_1 _9081_ (.A(_4089_),
    .B(_4105_),
    .Y(_4106_));
 sg13g2_nor2_1 _9082_ (.A(_4066_),
    .B(_4106_),
    .Y(_4107_));
 sg13g2_nand2_1 _9083_ (.Y(_4108_),
    .A(_4088_),
    .B(_4093_));
 sg13g2_inv_2 _9084_ (.Y(_4109_),
    .A(_4091_));
 sg13g2_nor2_1 _9085_ (.A(_4108_),
    .B(_4109_),
    .Y(_4110_));
 sg13g2_nand2_1 _9086_ (.Y(_4111_),
    .A(_4065_),
    .B(_4061_));
 sg13g2_a21oi_1 _9087_ (.A1(_4096_),
    .A2(_4101_),
    .Y(_4112_),
    .B1(_3816_));
 sg13g2_nand2_1 _9088_ (.Y(_4113_),
    .A(_4112_),
    .B(_4103_));
 sg13g2_nor2_1 _9089_ (.A(_4111_),
    .B(_4113_),
    .Y(_4114_));
 sg13g2_nand2_1 _9090_ (.Y(_4115_),
    .A(_4110_),
    .B(_4114_));
 sg13g2_nand2_1 _9091_ (.Y(_4116_),
    .A(_4107_),
    .B(_4115_));
 sg13g2_a21oi_1 _9092_ (.A1(_3969_),
    .A2(_4042_),
    .Y(_4117_),
    .B1(_4052_));
 sg13g2_o21ai_1 _9093_ (.B1(_4052_),
    .Y(_4118_),
    .A1(_3969_),
    .A2(_4042_));
 sg13g2_nor2b_1 _9094_ (.A(_4117_),
    .B_N(_4118_),
    .Y(_4119_));
 sg13g2_inv_1 _9095_ (.Y(_4120_),
    .A(_4119_));
 sg13g2_nand2_1 _9096_ (.Y(_4121_),
    .A(_4116_),
    .B(_4120_));
 sg13g2_nand3_1 _9097_ (.B(_4115_),
    .C(_4119_),
    .A(_4107_),
    .Y(_4122_));
 sg13g2_a21oi_1 _9098_ (.A1(_4121_),
    .A2(_4122_),
    .Y(_0179_),
    .B1(_3997_));
 sg13g2_o21ai_1 _9099_ (.B1(_4048_),
    .Y(_4123_),
    .A1(_4093_),
    .A2(_4109_));
 sg13g2_nor2_1 _9100_ (.A(_4120_),
    .B(_4111_),
    .Y(_4124_));
 sg13g2_a21oi_1 _9101_ (.A1(_4065_),
    .A2(_4118_),
    .Y(_4125_),
    .B1(_4117_));
 sg13g2_a21oi_1 _9102_ (.A1(_4123_),
    .A2(_4124_),
    .Y(_4126_),
    .B1(_4125_));
 sg13g2_nand2_1 _9103_ (.Y(_4127_),
    .A(_4113_),
    .B(_4103_));
 sg13g2_nand3_1 _9104_ (.B(_4127_),
    .C(_4124_),
    .A(_4110_),
    .Y(_4128_));
 sg13g2_a21oi_1 _9105_ (.A1(_4126_),
    .A2(_4128_),
    .Y(_0180_),
    .B1(_3997_));
 sg13g2_nand2_1 _9106_ (.Y(_4129_),
    .A(_3378_),
    .B(_3304_));
 sg13g2_a21o_1 _9107_ (.A2(_4129_),
    .A1(_3845_),
    .B1(_2764_),
    .X(_4130_));
 sg13g2_nand2_1 _9108_ (.Y(_4131_),
    .A(_3942_),
    .B(_4130_));
 sg13g2_nor2b_1 _9109_ (.A(_3298_),
    .B_N(_3297_),
    .Y(_4132_));
 sg13g2_xnor2_1 _9110_ (.Y(_4133_),
    .A(_4132_),
    .B(_3295_));
 sg13g2_nor3_1 _9111_ (.A(_3356_),
    .B(_4133_),
    .C(net26),
    .Y(_4134_));
 sg13g2_nor2_1 _9112_ (.A(_4134_),
    .B(_3831_),
    .Y(_4135_));
 sg13g2_nand2_1 _9113_ (.Y(_4136_),
    .A(_3374_),
    .B(_4135_));
 sg13g2_nand2_1 _9114_ (.Y(_4137_),
    .A(_4131_),
    .B(_4136_));
 sg13g2_nand2_1 _9115_ (.Y(_4138_),
    .A(_4137_),
    .B(_4022_));
 sg13g2_nand2_1 _9116_ (.Y(_4139_),
    .A(_4138_),
    .B(net11));
 sg13g2_a21oi_1 _9117_ (.A1(net12),
    .A2(_3869_),
    .Y(_4140_),
    .B1(net46));
 sg13g2_nand2_1 _9118_ (.Y(_4141_),
    .A(_4139_),
    .B(_4140_));
 sg13g2_nand2_1 _9119_ (.Y(_4142_),
    .A(_3377_),
    .B(_3354_));
 sg13g2_a21oi_1 _9120_ (.A1(_3877_),
    .A2(_4142_),
    .Y(_4143_),
    .B1(_2764_));
 sg13g2_nand2_1 _9121_ (.Y(_4144_),
    .A(net13),
    .B(_4143_));
 sg13g2_nand2_1 _9122_ (.Y(_4145_),
    .A(_3946_),
    .B(_4144_));
 sg13g2_a21oi_1 _9123_ (.A1(_3863_),
    .A2(_3872_),
    .Y(_4146_),
    .B1(_3864_));
 sg13g2_a21oi_1 _9124_ (.A1(_3822_),
    .A2(_4146_),
    .Y(_4147_),
    .B1(net46));
 sg13g2_a21oi_1 _9125_ (.A1(_4145_),
    .A2(_4147_),
    .Y(_4148_),
    .B1(_3933_));
 sg13g2_inv_1 _9126_ (.Y(_4149_),
    .A(_4148_));
 sg13g2_nand2_1 _9127_ (.Y(_4150_),
    .A(_4141_),
    .B(_4149_));
 sg13g2_nand3_1 _9128_ (.B(_4140_),
    .C(_4148_),
    .A(_4139_),
    .Y(_4151_));
 sg13g2_nand2_1 _9129_ (.Y(_4152_),
    .A(_4150_),
    .B(_4151_));
 sg13g2_nand2_1 _9130_ (.Y(_4153_),
    .A(_4152_),
    .B(_3953_));
 sg13g2_nand3_1 _9131_ (.B(_4151_),
    .C(_3955_),
    .A(_4150_),
    .Y(_4154_));
 sg13g2_nand2_1 _9132_ (.Y(_4155_),
    .A(_4153_),
    .B(_4154_));
 sg13g2_or2_1 _9133_ (.X(_4156_),
    .B(_3291_),
    .A(_3292_));
 sg13g2_nand4_1 _9134_ (.B(_3293_),
    .C(_3378_),
    .A(_3377_),
    .Y(_4157_),
    .D(_4156_));
 sg13g2_nand2_1 _9135_ (.Y(_4158_),
    .A(_3367_),
    .B(_4157_));
 sg13g2_nand2_1 _9136_ (.Y(_4159_),
    .A(_3375_),
    .B(_4158_));
 sg13g2_nand2_1 _9137_ (.Y(_4160_),
    .A(_3877_),
    .B(_4142_));
 sg13g2_nand4_1 _9138_ (.B(_3220_),
    .C(_3259_),
    .A(_3149_),
    .Y(_4161_),
    .D(_4160_));
 sg13g2_nand3_1 _9139_ (.B(_4161_),
    .C(_3382_),
    .A(_4159_),
    .Y(_4162_));
 sg13g2_nand2_1 _9140_ (.Y(_4163_),
    .A(_4162_),
    .B(_4011_));
 sg13g2_nand2_1 _9141_ (.Y(_4164_),
    .A(_4163_),
    .B(_3424_));
 sg13g2_a21oi_1 _9142_ (.A1(_4164_),
    .A2(_3909_),
    .Y(_4165_),
    .B1(_3933_));
 sg13g2_inv_1 _9143_ (.Y(_4166_),
    .A(_4141_));
 sg13g2_nand2_1 _9144_ (.Y(_4167_),
    .A(_4165_),
    .B(_4166_));
 sg13g2_nand2_1 _9145_ (.Y(_4168_),
    .A(_4164_),
    .B(_3909_));
 sg13g2_nand2_1 _9146_ (.Y(_4169_),
    .A(_4168_),
    .B(_3932_));
 sg13g2_nand2_1 _9147_ (.Y(_4170_),
    .A(_4169_),
    .B(_4141_));
 sg13g2_inv_1 _9148_ (.Y(_4171_),
    .A(_4170_));
 sg13g2_a21oi_1 _9149_ (.A1(_4167_),
    .A2(_3892_),
    .Y(_4172_),
    .B1(_4171_));
 sg13g2_nor2_1 _9150_ (.A(_4155_),
    .B(_4172_),
    .Y(_4173_));
 sg13g2_nor2b_1 _9151_ (.A(_3277_),
    .B_N(_3290_),
    .Y(_4174_));
 sg13g2_xnor2_1 _9152_ (.Y(_4175_),
    .A(_4174_),
    .B(_3289_));
 sg13g2_nand3_1 _9153_ (.B(_3378_),
    .C(_4175_),
    .A(_3377_),
    .Y(_4176_));
 sg13g2_nand2_1 _9154_ (.Y(_4177_),
    .A(_3827_),
    .B(_4176_));
 sg13g2_nand2_1 _9155_ (.Y(_4178_),
    .A(net13),
    .B(_4177_));
 sg13g2_inv_1 _9156_ (.Y(_4179_),
    .A(_4135_));
 sg13g2_nand4_1 _9157_ (.B(_3220_),
    .C(_3259_),
    .A(_3149_),
    .Y(_4180_),
    .D(_4179_));
 sg13g2_nand3_1 _9158_ (.B(_4180_),
    .C(_3382_),
    .A(_4178_),
    .Y(_4181_));
 sg13g2_nand2_1 _9159_ (.Y(_4182_),
    .A(_4181_),
    .B(_3823_));
 sg13g2_nand2_1 _9160_ (.Y(_4183_),
    .A(_4182_),
    .B(_3815_));
 sg13g2_nor2b_1 _9161_ (.A(_3287_),
    .B_N(_3286_),
    .Y(_4184_));
 sg13g2_nor4_1 _9162_ (.A(_3288_),
    .B(_3356_),
    .C(_4184_),
    .D(_3333_),
    .Y(_4185_));
 sg13g2_nor2b_1 _9163_ (.A(_4185_),
    .B_N(_3376_),
    .Y(_4186_));
 sg13g2_nand2b_1 _9164_ (.Y(_4187_),
    .B(_3374_),
    .A_N(_4186_));
 sg13g2_nand4_1 _9165_ (.B(_3220_),
    .C(_3259_),
    .A(_3149_),
    .Y(_4188_),
    .D(_4158_));
 sg13g2_nand3_1 _9166_ (.B(_4188_),
    .C(net21),
    .A(_4187_),
    .Y(_4189_));
 sg13g2_nand2_1 _9167_ (.Y(_4190_),
    .A(_4189_),
    .B(_4080_));
 sg13g2_nor2b_1 _9168_ (.A(_4183_),
    .B_N(_4190_),
    .Y(_4191_));
 sg13g2_a21oi_2 _9169_ (.B1(net46),
    .Y(_4192_),
    .A2(_3823_),
    .A1(_4181_));
 sg13g2_a21oi_1 _9170_ (.A1(_4189_),
    .A2(_4080_),
    .Y(_4193_),
    .B1(_3888_));
 sg13g2_nor2_1 _9171_ (.A(_4192_),
    .B(_4193_),
    .Y(_4194_));
 sg13g2_nor2_1 _9172_ (.A(_4191_),
    .B(_4194_),
    .Y(_4195_));
 sg13g2_nand2_1 _9173_ (.Y(_4196_),
    .A(_4195_),
    .B(_4169_));
 sg13g2_nand2_1 _9174_ (.Y(_4197_),
    .A(_4190_),
    .B(net47));
 sg13g2_nand2_1 _9175_ (.Y(_4198_),
    .A(_4183_),
    .B(_4197_));
 sg13g2_nand2_1 _9176_ (.Y(_4199_),
    .A(_4192_),
    .B(_4190_));
 sg13g2_nand2_1 _9177_ (.Y(_4200_),
    .A(_4198_),
    .B(_4199_));
 sg13g2_nand2_1 _9178_ (.Y(_4201_),
    .A(_4200_),
    .B(_4165_));
 sg13g2_nand2_1 _9179_ (.Y(_4202_),
    .A(_4196_),
    .B(_4201_));
 sg13g2_o21ai_1 _9180_ (.B1(_3905_),
    .Y(_4203_),
    .A1(_4130_),
    .A2(_3261_));
 sg13g2_nand2_1 _9181_ (.Y(_4204_),
    .A(_4203_),
    .B(_3423_));
 sg13g2_o21ai_1 _9182_ (.B1(_3822_),
    .Y(_4205_),
    .A1(_3867_),
    .A2(_4037_));
 sg13g2_nand2_1 _9183_ (.Y(_4206_),
    .A(_4204_),
    .B(_4205_));
 sg13g2_nand2_1 _9184_ (.Y(_4207_),
    .A(_4206_),
    .B(_3814_));
 sg13g2_nand2_1 _9185_ (.Y(_4208_),
    .A(_4207_),
    .B(_3932_));
 sg13g2_nand2_1 _9186_ (.Y(_4209_),
    .A(_4192_),
    .B(_4098_));
 sg13g2_nor2_1 _9187_ (.A(_4098_),
    .B(_4192_),
    .Y(_4210_));
 sg13g2_a21oi_1 _9188_ (.A1(_4208_),
    .A2(_4209_),
    .Y(_4211_),
    .B1(_4210_));
 sg13g2_nand2_1 _9189_ (.Y(_4212_),
    .A(_4202_),
    .B(_4211_));
 sg13g2_nand2_1 _9190_ (.Y(_4213_),
    .A(_4212_),
    .B(_3841_));
 sg13g2_nor2_1 _9191_ (.A(_4173_),
    .B(_4213_),
    .Y(_4214_));
 sg13g2_nand2_1 _9192_ (.Y(_4215_),
    .A(_4167_),
    .B(_4170_));
 sg13g2_nand2_1 _9193_ (.Y(_4216_),
    .A(_4215_),
    .B(_3891_));
 sg13g2_nand3_1 _9194_ (.B(_4170_),
    .C(_3892_),
    .A(_4167_),
    .Y(_4217_));
 sg13g2_nand2_1 _9195_ (.Y(_4218_),
    .A(_4196_),
    .B(_4198_));
 sg13g2_nand3_1 _9196_ (.B(_4217_),
    .C(_4218_),
    .A(_4216_),
    .Y(_4219_));
 sg13g2_or2_1 _9197_ (.X(_4220_),
    .B(_4202_),
    .A(_4211_));
 sg13g2_buf_1 _9198_ (.A(_4220_),
    .X(_4221_));
 sg13g2_nand3_1 _9199_ (.B(_4219_),
    .C(_4221_),
    .A(_4214_),
    .Y(_4222_));
 sg13g2_nand2_1 _9200_ (.Y(_4223_),
    .A(_4219_),
    .B(_4221_));
 sg13g2_inv_1 _9201_ (.Y(_4224_),
    .A(_4173_));
 sg13g2_nand2_1 _9202_ (.Y(_4225_),
    .A(_4223_),
    .B(_4224_));
 sg13g2_nand2_1 _9203_ (.Y(_4226_),
    .A(_4222_),
    .B(_4225_));
 sg13g2_a21oi_1 _9204_ (.A1(_4216_),
    .A2(_4217_),
    .Y(_4227_),
    .B1(_4218_));
 sg13g2_inv_1 _9205_ (.Y(_4228_),
    .A(_4150_));
 sg13g2_a21oi_1 _9206_ (.A1(_4151_),
    .A2(_3955_),
    .Y(_4229_),
    .B1(_4228_));
 sg13g2_nand2_1 _9207_ (.Y(_4230_),
    .A(_4145_),
    .B(_4147_));
 sg13g2_inv_2 _9208_ (.Y(_4231_),
    .A(_4208_));
 sg13g2_nand2b_1 _9209_ (.Y(_4232_),
    .B(_4231_),
    .A_N(_4230_));
 sg13g2_nand3_1 _9210_ (.B(net47),
    .C(_4230_),
    .A(_4206_),
    .Y(_4233_));
 sg13g2_nand2_1 _9211_ (.Y(_4234_),
    .A(_4232_),
    .B(_4233_));
 sg13g2_nand2_1 _9212_ (.Y(_4235_),
    .A(_4234_),
    .B(_3969_));
 sg13g2_nand3_1 _9213_ (.B(_3968_),
    .C(_4233_),
    .A(_4232_),
    .Y(_4236_));
 sg13g2_nand2_1 _9214_ (.Y(_4237_),
    .A(_4235_),
    .B(_4236_));
 sg13g2_nand2b_1 _9215_ (.Y(_4238_),
    .B(_4237_),
    .A_N(_4229_));
 sg13g2_nand3_1 _9216_ (.B(_4236_),
    .C(_4229_),
    .A(_4235_),
    .Y(_4239_));
 sg13g2_nand2_1 _9217_ (.Y(_4240_),
    .A(_4238_),
    .B(_4239_));
 sg13g2_nand2_1 _9218_ (.Y(_4241_),
    .A(_4172_),
    .B(_4155_));
 sg13g2_nand2_1 _9219_ (.Y(_4242_),
    .A(_4240_),
    .B(_4241_));
 sg13g2_nor2_1 _9220_ (.A(_4227_),
    .B(_4242_),
    .Y(_4243_));
 sg13g2_nand2_1 _9221_ (.Y(_4244_),
    .A(_4226_),
    .B(_4243_));
 sg13g2_nor2_1 _9222_ (.A(_4229_),
    .B(_4237_),
    .Y(_4245_));
 sg13g2_a21oi_1 _9223_ (.A1(_4240_),
    .A2(_4173_),
    .Y(_4246_),
    .B1(_4245_));
 sg13g2_nand2_1 _9224_ (.Y(_4247_),
    .A(_4244_),
    .B(_4246_));
 sg13g2_a21oi_1 _9225_ (.A1(_3968_),
    .A2(_4148_),
    .Y(_4248_),
    .B1(_4231_));
 sg13g2_a21oi_1 _9226_ (.A1(_4235_),
    .A2(_4231_),
    .Y(_4249_),
    .B1(_4248_));
 sg13g2_nand2_1 _9227_ (.Y(_4250_),
    .A(_4247_),
    .B(_4249_));
 sg13g2_nand2_1 _9228_ (.Y(_4251_),
    .A(_4250_),
    .B(_3998_));
 sg13g2_nand3b_1 _9229_ (.B(_4244_),
    .C(_4246_),
    .Y(_4252_),
    .A_N(_4249_));
 sg13g2_nor2b_1 _9230_ (.A(_4251_),
    .B_N(_4252_),
    .Y(_0259_));
 sg13g2_nand2_1 _9231_ (.Y(_4253_),
    .A(_4219_),
    .B(_4224_));
 sg13g2_a21oi_1 _9232_ (.A1(_4221_),
    .A2(_4213_),
    .Y(_4254_),
    .B1(_4227_));
 sg13g2_nor2b_1 _9233_ (.A(_4242_),
    .B_N(_4249_),
    .Y(_4255_));
 sg13g2_o21ai_1 _9234_ (.B1(_4255_),
    .Y(_4256_),
    .A1(_4253_),
    .A2(_4254_));
 sg13g2_a21oi_1 _9235_ (.A1(_4245_),
    .A2(_4208_),
    .Y(_4257_),
    .B1(_4248_));
 sg13g2_a21oi_1 _9236_ (.A1(_4256_),
    .A2(_4257_),
    .Y(_0260_),
    .B1(_3997_));
 sg13g2_xor2_1 _9237_ (.B(\vgademo.soundtrack.sample_div[0] ),
    .A(\vgademo.soundtrack.sample_div[1] ),
    .X(\vgademo.soundtrack.sample_div_[1] ));
 sg13g2_xnor2_1 _9238_ (.Y(\vgademo.soundtrack.sample_div_[2] ),
    .A(\vgademo.soundtrack.sample_div[2] ),
    .B(_2018_));
 sg13g2_o21ai_1 _9239_ (.B1(_2016_),
    .Y(_4258_),
    .A1(_2017_),
    .A2(_2018_));
 sg13g2_nor2b_1 _9240_ (.A(_2019_),
    .B_N(_4258_),
    .Y(\vgademo.soundtrack.sample_div_[3] ));
 sg13g2_xor2_1 _9241_ (.B(_2019_),
    .A(\vgademo.soundtrack.sample_div[4] ),
    .X(\vgademo.soundtrack.sample_div_[4] ));
 sg13g2_xnor2_1 _9242_ (.Y(\vgademo.soundtrack.sample_div_[5] ),
    .A(\vgademo.soundtrack.sample_div[5] ),
    .B(_2020_));
 sg13g2_xor2_1 _9243_ (.B(_2021_),
    .A(\vgademo.soundtrack.sample_div[6] ),
    .X(\vgademo.soundtrack.sample_div_[6] ));
 sg13g2_xnor2_1 _9244_ (.Y(\vgademo.soundtrack.sample_div_[7] ),
    .A(\vgademo.soundtrack.sample_div[7] ),
    .B(_2022_));
 sg13g2_xor2_1 _9245_ (.B(_2023_),
    .A(\vgademo.soundtrack.sample_div[8] ),
    .X(\vgademo.soundtrack.sample_div_[8] ));
 sg13g2_xnor2_1 _9246_ (.Y(\vgademo.soundtrack.sample_div_[9] ),
    .A(\vgademo.soundtrack.sample_div[9] ),
    .B(_2024_));
 sg13g2_xnor2_1 _9247_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .A(\vgademo.soundtrack.sigma_delta_accum[0] ),
    .B(_2204_));
 sg13g2_xor2_1 _9248_ (.B(_2235_),
    .A(_2238_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[10] ));
 sg13g2_nor2_1 _9249_ (.A(_2243_),
    .B(_2241_),
    .Y(_4259_));
 sg13g2_inv_1 _9250_ (.Y(_4260_),
    .A(_2233_));
 sg13g2_nor2_1 _9251_ (.A(_4260_),
    .B(_2237_),
    .Y(_4261_));
 sg13g2_nor2_1 _9252_ (.A(_2234_),
    .B(_4260_),
    .Y(_4262_));
 sg13g2_nand3_1 _9253_ (.B(_2231_),
    .C(_4262_),
    .A(_2238_),
    .Y(_4263_));
 sg13g2_o21ai_1 _9254_ (.B1(_4263_),
    .Y(_4264_),
    .A1(_2236_),
    .A2(_4261_));
 sg13g2_xor2_1 _9255_ (.B(_4264_),
    .A(_4259_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[11] ));
 sg13g2_xor2_1 _9256_ (.B(_2244_),
    .A(_2246_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[12] ));
 sg13g2_nand2_1 _9257_ (.Y(_4265_),
    .A(_4264_),
    .B(_4259_));
 sg13g2_nor2_1 _9258_ (.A(_2241_),
    .B(_2182_),
    .Y(_4266_));
 sg13g2_a21oi_1 _9259_ (.A1(_4265_),
    .A2(_4266_),
    .Y(_4267_),
    .B1(_2245_));
 sg13g2_xnor2_1 _9260_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .A(_2187_),
    .B(_4267_));
 sg13g2_nor2_1 _9261_ (.A(_2252_),
    .B(_2180_),
    .Y(_4268_));
 sg13g2_xnor2_1 _9262_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .A(_4268_),
    .B(_2249_));
 sg13g2_nor2b_1 _9263_ (.A(_2177_),
    .B_N(_2251_),
    .Y(_4269_));
 sg13g2_nand2_1 _9264_ (.Y(_4270_),
    .A(_2250_),
    .B(_2253_));
 sg13g2_xnor2_1 _9265_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .A(_4269_),
    .B(_4270_));
 sg13g2_xnor2_1 _9266_ (.Y(_4271_),
    .A(_2202_),
    .B(_2201_));
 sg13g2_xnor2_1 _9267_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .A(_2205_),
    .B(_4271_));
 sg13g2_xor2_1 _9268_ (.B(_2209_),
    .A(_2207_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[2] ));
 sg13g2_xor2_1 _9269_ (.B(_2200_),
    .A(_2211_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[3] ));
 sg13g2_nand2b_1 _9270_ (.Y(_4272_),
    .B(_2216_),
    .A_N(_2217_));
 sg13g2_xnor2_1 _9271_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .A(_2213_),
    .B(_4272_));
 sg13g2_xnor2_1 _9272_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .A(_2197_),
    .B(_2218_));
 sg13g2_nor2b_1 _9273_ (.A(_2193_),
    .B_N(_2222_),
    .Y(_4273_));
 sg13g2_xor2_1 _9274_ (.B(_2220_),
    .A(_4273_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[6] ));
 sg13g2_nand2b_1 _9275_ (.Y(_4274_),
    .B(_2226_),
    .A_N(_2227_));
 sg13g2_xnor2_1 _9276_ (.Y(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .A(_2223_),
    .B(_4274_));
 sg13g2_xor2_1 _9277_ (.B(_2228_),
    .A(_2190_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[8] ));
 sg13g2_xor2_1 _9278_ (.B(_2231_),
    .A(_4262_),
    .X(\vgademo.soundtrack.sigma_delta_accum_[9] ));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _9288__167 (.L_HI(net167));
 sg13g2_buf_1 _9281_ (.A(net153),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9282_ (.A(net154),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9283_ (.A(net155),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9284_ (.A(net156),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9285_ (.A(net157),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9286_ (.A(net158),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9287_ (.A(net159),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9288_ (.A(net167),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9289_ (.A(net160),
    .X(uio_out[0]));
 sg13g2_buf_1 _9290_ (.A(net161),
    .X(uio_out[1]));
 sg13g2_buf_1 _9291_ (.A(net162),
    .X(uio_out[2]));
 sg13g2_buf_1 _9292_ (.A(net163),
    .X(uio_out[3]));
 sg13g2_buf_1 _9293_ (.A(net164),
    .X(uio_out[4]));
 sg13g2_buf_1 _9294_ (.A(net165),
    .X(uio_out[5]));
 sg13g2_buf_1 _9295_ (.A(net166),
    .X(uio_out[6]));
 sg13g2_buf_1 _9296_ (.A(audio),
    .X(net2));
 sg13g2_buf_1 _9297_ (.A(\vgademo.vsync ),
    .X(net6));
 sg13g2_buf_1 _9298_ (.A(hsync),
    .X(net10));
 sg13g2_dfrbp_1 \vgademo.a_cos[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net134),
    .D(_0112_),
    .Q_N(_4744_),
    .Q(\vgademo.a_cos[0] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net143),
    .D(_0113_),
    .Q_N(_4743_),
    .Q(\vgademo.a_cos[10] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net143),
    .D(_0114_),
    .Q_N(_4742_),
    .Q(\vgademo.a_cos[11] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net137),
    .D(_0115_),
    .Q_N(_4741_),
    .Q(\vgademo.a_cos[12] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[13]$_DFFE_PN1P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net137),
    .D(_0116_),
    .Q_N(\vgademo.a_cos[13] ),
    .Q(_0086_));
 sg13g2_dfrbp_1 \vgademo.a_cos[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net142),
    .D(_0117_),
    .Q_N(_4740_),
    .Q(\vgademo.a_cos[14] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net134),
    .D(_0118_),
    .Q_N(_4739_),
    .Q(\vgademo.a_cos[1] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net133),
    .D(_0119_),
    .Q_N(_4738_),
    .Q(\vgademo.a_cos[2] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net141),
    .D(_0120_),
    .Q_N(_4737_),
    .Q(\vgademo.a_cos[3] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net141),
    .D(_0121_),
    .Q_N(_4736_),
    .Q(\vgademo.a_cos[4] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net141),
    .D(_0122_),
    .Q_N(_4735_),
    .Q(\vgademo.a_cos[5] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net142),
    .D(_0123_),
    .Q_N(_4734_),
    .Q(\vgademo.a_cos[6] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net142),
    .D(_0124_),
    .Q_N(_4733_),
    .Q(\vgademo.a_cos[7] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net142),
    .D(_0125_),
    .Q_N(_4732_),
    .Q(\vgademo.a_cos[8] ));
 sg13g2_dfrbp_1 \vgademo.a_cos[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net142),
    .D(_0126_),
    .Q_N(_4731_),
    .Q(\vgademo.a_cos[9] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net141),
    .D(_0127_),
    .Q_N(_4730_),
    .Q(\vgademo.a_sin[0] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net141),
    .D(_0128_),
    .Q_N(_4729_),
    .Q(\vgademo.a_sin[10] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net141),
    .D(_0129_),
    .Q_N(_4728_),
    .Q(\vgademo.a_sin[11] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net133),
    .D(_0130_),
    .Q_N(_4727_),
    .Q(\vgademo.a_sin[12] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net133),
    .D(_0131_),
    .Q_N(_4726_),
    .Q(\vgademo.a_sin[13] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net142),
    .D(_0132_),
    .Q_N(_4725_),
    .Q(\vgademo.a_sin[14] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net141),
    .D(_0133_),
    .Q_N(_4724_),
    .Q(\vgademo.a_sin[1] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net142),
    .D(_0134_),
    .Q_N(_4723_),
    .Q(\vgademo.a_sin[2] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net144),
    .D(_0135_),
    .Q_N(_4722_),
    .Q(\vgademo.a_sin[3] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net144),
    .D(_0136_),
    .Q_N(_4721_),
    .Q(\vgademo.a_sin[4] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net134),
    .D(_0137_),
    .Q_N(_4720_),
    .Q(\vgademo.a_sin[5] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net135),
    .D(_0138_),
    .Q_N(_4719_),
    .Q(\vgademo.a_sin[6] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net135),
    .D(_0139_),
    .Q_N(_4718_),
    .Q(\vgademo.a_sin[7] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net133),
    .D(_0140_),
    .Q_N(_4717_),
    .Q(\vgademo.a_sin[8] ));
 sg13g2_dfrbp_1 \vgademo.a_sin[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net141),
    .D(_0141_),
    .Q_N(_4716_),
    .Q(\vgademo.a_sin[9] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[0]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net168),
    .D(_0142_),
    .Q_N(_4715_),
    .Q(\vgademo.b_cos[0] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[10]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net169),
    .D(_0143_),
    .Q_N(_4714_),
    .Q(\vgademo.b_cos[10] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net170),
    .D(_0144_),
    .Q_N(_4713_),
    .Q(\vgademo.b_cos[11] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[1]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net171),
    .D(_0145_),
    .Q_N(_4712_),
    .Q(\vgademo.b_cos[1] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[2]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net172),
    .D(_0146_),
    .Q_N(_4711_),
    .Q(\vgademo.b_cos[2] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net173),
    .D(_0147_),
    .Q_N(_4710_),
    .Q(\vgademo.b_cos[3] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[4]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net174),
    .D(_0148_),
    .Q_N(_4709_),
    .Q(\vgademo.b_cos[4] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[5]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net175),
    .D(_0149_),
    .Q_N(_4708_),
    .Q(\vgademo.b_cos[5] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net176),
    .D(_0150_),
    .Q_N(_4707_),
    .Q(\vgademo.b_cos[6] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net177),
    .D(_0151_),
    .Q_N(_4706_),
    .Q(\vgademo.b_cos[7] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[8]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net178),
    .D(_0152_),
    .Q_N(_4705_),
    .Q(\vgademo.b_cos[8] ));
 sg13g2_dfrbp_1 \vgademo.b_cos[9]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net179),
    .D(_0153_),
    .Q_N(_4704_),
    .Q(\vgademo.b_cos[9] ));
 sg13g2_dfrbp_1 \vgademo.b_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net180),
    .D(_0154_),
    .Q_N(_4703_),
    .Q(net9));
 sg13g2_dfrbp_1 \vgademo.b_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net181),
    .D(_0155_),
    .Q_N(_4702_),
    .Q(net5));
 sg13g2_dfrbp_1 \vgademo.b_sin[0]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net182),
    .D(_0156_),
    .Q_N(_4701_),
    .Q(\vgademo.b_sin[0] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net183),
    .D(_0157_),
    .Q_N(_4700_),
    .Q(\vgademo.b_sin[10] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[11]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net184),
    .D(_0158_),
    .Q_N(_4699_),
    .Q(\vgademo.b_sin[11] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[1]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net185),
    .D(_0159_),
    .Q_N(_4698_),
    .Q(\vgademo.b_sin[1] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net186),
    .D(_0160_),
    .Q_N(_4697_),
    .Q(\vgademo.b_sin[2] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[3]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net187),
    .D(_0161_),
    .Q_N(_4696_),
    .Q(\vgademo.b_sin[3] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net188),
    .D(_0162_),
    .Q_N(_4695_),
    .Q(\vgademo.b_sin[4] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[5]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net189),
    .D(_0163_),
    .Q_N(_4694_),
    .Q(\vgademo.b_sin[5] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[6]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net190),
    .D(_0164_),
    .Q_N(_4693_),
    .Q(\vgademo.b_sin[6] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net191),
    .D(_0165_),
    .Q_N(_4692_),
    .Q(\vgademo.b_sin[7] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[8]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net192),
    .D(_0166_),
    .Q_N(_4691_),
    .Q(\vgademo.b_sin[8] ));
 sg13g2_dfrbp_1 \vgademo.b_sin[9]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net193),
    .D(_0167_),
    .Q_N(_4690_),
    .Q(\vgademo.b_sin[9] ));
 sg13g2_dfrbp_1 \vgademo.frame[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net150),
    .D(_0168_),
    .Q_N(_0081_),
    .Q(\vgademo.a_scrolly[3] ));
 sg13g2_dfrbp_1 \vgademo.frame[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_0169_),
    .Q_N(_0015_),
    .Q(\vgademo.a_scrolly[13] ));
 sg13g2_dfrbp_1 \vgademo.frame[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net149),
    .D(_0170_),
    .Q_N(_0017_),
    .Q(\vgademo.a_scrolly[4] ));
 sg13g2_dfrbp_1 \vgademo.frame[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_0171_),
    .Q_N(_0058_),
    .Q(\vgademo.a_scrolly[5] ));
 sg13g2_dfrbp_1 \vgademo.frame[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net150),
    .D(_0172_),
    .Q_N(_0024_),
    .Q(\vgademo.a_scrolly[6] ));
 sg13g2_dfrbp_1 \vgademo.frame[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net150),
    .D(_0173_),
    .Q_N(_0014_),
    .Q(\vgademo.a_scrolly[7] ));
 sg13g2_dfrbp_1 \vgademo.frame[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net150),
    .D(_0174_),
    .Q_N(_0029_),
    .Q(\vgademo.a_scrolly[8] ));
 sg13g2_dfrbp_1 \vgademo.frame[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net150),
    .D(_0175_),
    .Q_N(_0059_),
    .Q(\vgademo.a_scrolly[9] ));
 sg13g2_dfrbp_1 \vgademo.frame[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net151),
    .D(_0176_),
    .Q_N(_0034_),
    .Q(\vgademo.a_scrolly[10] ));
 sg13g2_dfrbp_1 \vgademo.frame[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net151),
    .D(_0177_),
    .Q_N(_0037_),
    .Q(\vgademo.a_scrolly[11] ));
 sg13g2_dfrbp_1 \vgademo.frame[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net150),
    .D(_0178_),
    .Q_N(_0060_),
    .Q(\vgademo.a_scrolly[12] ));
 sg13g2_dfrbp_1 \vgademo.g_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net194),
    .D(_0179_),
    .Q_N(_4689_),
    .Q(net8));
 sg13g2_dfrbp_1 \vgademo.g_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net195),
    .D(_0180_),
    .Q_N(_4745_),
    .Q(net4));
 sg13g2_dfrbp_1 \vgademo.h_count[0]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net137),
    .D(_0000_),
    .Q_N(_4746_),
    .Q(\vgademo.h_count[0] ));
 sg13g2_dfrbp_1 \vgademo.h_count[10]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net143),
    .D(_0001_),
    .Q_N(_0078_),
    .Q(\vgademo.h_count[10] ));
 sg13g2_dfrbp_1 \vgademo.h_count[1]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net146),
    .D(_0002_),
    .Q_N(_0066_),
    .Q(\vgademo.h_count[1] ));
 sg13g2_dfrbp_1 \vgademo.h_count[2]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net138),
    .D(_0003_),
    .Q_N(_0051_),
    .Q(\vgademo.h_count[2] ));
 sg13g2_dfrbp_1 \vgademo.h_count[3]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net138),
    .D(_0004_),
    .Q_N(_0052_),
    .Q(\vgademo.h_count[3] ));
 sg13g2_dfrbp_1 \vgademo.h_count[4]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net138),
    .D(_0005_),
    .Q_N(_0053_),
    .Q(\vgademo.h_count[4] ));
 sg13g2_dfrbp_1 \vgademo.h_count[5]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net143),
    .D(_0006_),
    .Q_N(_0054_),
    .Q(\vgademo.h_count[5] ));
 sg13g2_dfrbp_1 \vgademo.h_count[6]$_DFF_PN0_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net143),
    .D(_0007_),
    .Q_N(_0055_),
    .Q(\vgademo.h_count[6] ));
 sg13g2_dfrbp_1 \vgademo.h_count[7]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net143),
    .D(_0008_),
    .Q_N(_0056_),
    .Q(\vgademo.h_count[7] ));
 sg13g2_dfrbp_1 \vgademo.h_count[8]$_DFF_PN0_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net143),
    .D(_0009_),
    .Q_N(_0079_),
    .Q(\vgademo.h_count[8] ));
 sg13g2_dfrbp_1 \vgademo.h_count[9]$_DFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0010_),
    .Q_N(_0057_),
    .Q(\vgademo.h_count[9] ));
 sg13g2_dfrbp_1 \vgademo.hsync$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net196),
    .D(_0011_),
    .Q_N(_4688_),
    .Q(hsync));
 sg13g2_dfrbp_1 \vgademo.linelfsr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net197),
    .D(_0181_),
    .Q_N(_4687_),
    .Q(\vgademo.linelfsr[0] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net198),
    .D(_0182_),
    .Q_N(_4686_),
    .Q(\vgademo.linelfsr[10] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[11]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net199),
    .D(_0183_),
    .Q_N(_4685_),
    .Q(\vgademo.linelfsr[11] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[12]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net200),
    .D(_0184_),
    .Q_N(_4684_),
    .Q(\vgademo.linelfsr[12] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[1]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net201),
    .D(_0185_),
    .Q_N(_4683_),
    .Q(\vgademo.linelfsr[1] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net202),
    .D(_0186_),
    .Q_N(_4682_),
    .Q(\vgademo.linelfsr[2] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[3]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net203),
    .D(_0187_),
    .Q_N(_4681_),
    .Q(\vgademo.linelfsr[3] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[4]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net204),
    .D(_0188_),
    .Q_N(_4680_),
    .Q(\vgademo.linelfsr[4] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[5]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net205),
    .D(_0189_),
    .Q_N(_4679_),
    .Q(\vgademo.linelfsr[5] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[6]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net206),
    .D(_0190_),
    .Q_N(_4678_),
    .Q(\vgademo.linelfsr[6] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[7]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net207),
    .D(_0191_),
    .Q_N(_4677_),
    .Q(\vgademo.linelfsr[7] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net208),
    .D(_0192_),
    .Q_N(_4676_),
    .Q(\vgademo.linelfsr[8] ));
 sg13g2_dfrbp_1 \vgademo.linelfsr[9]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net209),
    .D(_0193_),
    .Q_N(_4675_),
    .Q(\vgademo.linelfsr[9] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[0]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net210),
    .D(_0194_),
    .Q_N(_4674_),
    .Q(\vgademo.plane_du[0] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[10]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net211),
    .D(_0195_),
    .Q_N(_4673_),
    .Q(\vgademo.plane_du[10] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net212),
    .D(_0196_),
    .Q_N(_4672_),
    .Q(\vgademo.plane_du[1] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[2]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net213),
    .D(_0197_),
    .Q_N(_4671_),
    .Q(\vgademo.plane_du[2] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[3]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net214),
    .D(_0198_),
    .Q_N(_0068_),
    .Q(\vgademo.plane_du[3] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[4]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net215),
    .D(_0199_),
    .Q_N(_0067_),
    .Q(\vgademo.plane_du[4] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net216),
    .D(_0200_),
    .Q_N(_0069_),
    .Q(\vgademo.plane_du[5] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[6]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net217),
    .D(_0201_),
    .Q_N(_0070_),
    .Q(\vgademo.plane_du[6] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net218),
    .D(_0202_),
    .Q_N(_0071_),
    .Q(\vgademo.plane_du[7] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[8]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net219),
    .D(_0203_),
    .Q_N(_0072_),
    .Q(\vgademo.plane_du[8] ));
 sg13g2_dfrbp_1 \vgademo.plane_du[9]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net220),
    .D(_0204_),
    .Q_N(_4670_),
    .Q(\vgademo.plane_du[9] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[16]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net221),
    .D(_0013_),
    .Q_N(_0026_),
    .Q(\vgademo.plane_dx_div.d[16] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[17]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net222),
    .D(_0205_),
    .Q_N(_0019_),
    .Q(\vgademo.plane_dx_div.d[17] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[18]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net223),
    .D(_0206_),
    .Q_N(_0022_),
    .Q(\vgademo.plane_dx_div.d[18] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[19]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net224),
    .D(_0207_),
    .Q_N(_0025_),
    .Q(\vgademo.plane_dx_div.d[19] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[20]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net225),
    .D(_0208_),
    .Q_N(_0028_),
    .Q(\vgademo.plane_dx_div.d[20] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[21]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net226),
    .D(_0209_),
    .Q_N(_0030_),
    .Q(\vgademo.plane_dx_div.d[21] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[22]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net227),
    .D(_0210_),
    .Q_N(_0033_),
    .Q(\vgademo.plane_dx_div.d[22] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[23]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net228),
    .D(_0211_),
    .Q_N(_0035_),
    .Q(\vgademo.plane_dx_div.d[23] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.d[24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net229),
    .D(_0212_),
    .Q_N(_0039_),
    .Q(\vgademo.plane_dx_div.d[24] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.i[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net230),
    .D(_0213_),
    .Q_N(_0082_),
    .Q(\vgademo.plane_dx_div.i[0] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.i[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net231),
    .D(_0214_),
    .Q_N(_4669_),
    .Q(\vgademo.plane_dx_div.i[1] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.i[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net232),
    .D(_0215_),
    .Q_N(_4668_),
    .Q(\vgademo.plane_dx_div.i[2] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.i[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net233),
    .D(_0216_),
    .Q_N(_4667_),
    .Q(\vgademo.plane_dx_div.i[3] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[0]$_SDFFE_PP1P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net234),
    .D(_0217_),
    .Q_N(_4666_),
    .Q(\vgademo.plane_dx[1] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net235),
    .D(_0218_),
    .Q_N(_4665_),
    .Q(\vgademo.plane_dx[2] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net236),
    .D(_0219_),
    .Q_N(_4664_),
    .Q(\vgademo.plane_dx_div.q[2] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net237),
    .D(_0220_),
    .Q_N(_4663_),
    .Q(\vgademo.plane_dx_div.q[3] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net238),
    .D(_0221_),
    .Q_N(_4662_),
    .Q(\vgademo.plane_dx_div.q[4] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net239),
    .D(_0222_),
    .Q_N(_4661_),
    .Q(\vgademo.plane_dx_div.q[5] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net240),
    .D(_0223_),
    .Q_N(_4660_),
    .Q(\vgademo.plane_dx_div.q[6] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net241),
    .D(_0224_),
    .Q_N(_4659_),
    .Q(\vgademo.plane_dx_div.q[7] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net242),
    .D(_0225_),
    .Q_N(_4658_),
    .Q(\vgademo.plane_dx_div.q[8] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.q[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net243),
    .D(_0226_),
    .Q_N(_4657_),
    .Q(\vgademo.plane_dx_div.q[9] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[16]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net244),
    .D(_0227_),
    .Q_N(_4656_),
    .Q(\vgademo.plane_dx_div.r[16] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[17]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net245),
    .D(_0228_),
    .Q_N(_4655_),
    .Q(\vgademo.plane_dx_div.r[17] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[18]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net246),
    .D(_0229_),
    .Q_N(_4654_),
    .Q(\vgademo.plane_dx_div.r[18] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[19]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net247),
    .D(_0230_),
    .Q_N(_4653_),
    .Q(\vgademo.plane_dx_div.r[19] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[20]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net248),
    .D(_0231_),
    .Q_N(_4652_),
    .Q(\vgademo.plane_dx_div.r[20] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[21]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net249),
    .D(_0232_),
    .Q_N(_4651_),
    .Q(\vgademo.plane_dx_div.r[21] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[22]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net250),
    .D(_0233_),
    .Q_N(_4650_),
    .Q(\vgademo.plane_dx_div.r[22] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[23]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net251),
    .D(_0234_),
    .Q_N(_4649_),
    .Q(\vgademo.plane_dx_div.r[23] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[24]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net252),
    .D(_0235_),
    .Q_N(_4648_),
    .Q(\vgademo.plane_dx_div.r[24] ));
 sg13g2_dfrbp_1 \vgademo.plane_dx_div.r[25]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net253),
    .D(_0236_),
    .Q_N(\vgademo.plane_dx[0] ),
    .Q(\vgademo.plane_dx_div.r[25] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net254),
    .D(_0237_),
    .Q_N(_4647_),
    .Q(\vgademo.plane_u[0] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net255),
    .D(_0238_),
    .Q_N(_4646_),
    .Q(\vgademo.plane_u[10] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[11]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net256),
    .D(_0239_),
    .Q_N(_0041_),
    .Q(\vgademo.plane_u[11] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[12]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net257),
    .D(_0240_),
    .Q_N(_0042_),
    .Q(\vgademo.plane_u[12] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[13]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net258),
    .D(_0241_),
    .Q_N(_0043_),
    .Q(\vgademo.plane_u[13] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[14]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net259),
    .D(_0242_),
    .Q_N(_0044_),
    .Q(\vgademo.plane_u[14] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[15]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net260),
    .D(_0243_),
    .Q_N(_0045_),
    .Q(\vgademo.plane_u[15] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net261),
    .D(_0244_),
    .Q_N(_0046_),
    .Q(\vgademo.plane_u[16] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[17]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net262),
    .D(_0245_),
    .Q_N(_0047_),
    .Q(\vgademo.plane_u[17] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[18]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net263),
    .D(_0246_),
    .Q_N(_0048_),
    .Q(\vgademo.plane_u[18] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[19]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net264),
    .D(_0247_),
    .Q_N(_0049_),
    .Q(\vgademo.plane_u[19] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[1]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net265),
    .D(_0248_),
    .Q_N(_4645_),
    .Q(\vgademo.plane_u[1] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[20]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net266),
    .D(_0249_),
    .Q_N(_0050_),
    .Q(\vgademo.plane_u[20] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[21]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net267),
    .D(_0250_),
    .Q_N(_4644_),
    .Q(\vgademo.plane_u[21] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net268),
    .D(_0251_),
    .Q_N(_4643_),
    .Q(\vgademo.plane_u[2] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[3]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net269),
    .D(_0252_),
    .Q_N(_4642_),
    .Q(\vgademo.plane_u[3] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net270),
    .D(_0253_),
    .Q_N(_4641_),
    .Q(\vgademo.plane_u[4] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net271),
    .D(_0254_),
    .Q_N(_4640_),
    .Q(\vgademo.plane_u[5] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[6]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net272),
    .D(_0255_),
    .Q_N(_4639_),
    .Q(\vgademo.plane_u[6] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[7]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net273),
    .D(_0256_),
    .Q_N(_4638_),
    .Q(\vgademo.plane_u[7] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[8]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net274),
    .D(_0257_),
    .Q_N(_4637_),
    .Q(\vgademo.plane_u[8] ));
 sg13g2_dfrbp_1 \vgademo.plane_u[9]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net275),
    .D(_0258_),
    .Q_N(_4636_),
    .Q(\vgademo.plane_u[9] ));
 sg13g2_dfrbp_1 \vgademo.r_out[0]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net276),
    .D(_0259_),
    .Q_N(_4635_),
    .Q(net7));
 sg13g2_dfrbp_1 \vgademo.r_out[1]$_SDFF_PN0_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net277),
    .D(_0260_),
    .Q_N(_4634_),
    .Q(net3));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[0]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net278),
    .D(_0261_),
    .Q_N(_4633_),
    .Q(\vgademo.scanline_audio_sample[0] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net279),
    .D(_0262_),
    .Q_N(_4632_),
    .Q(\vgademo.scanline_audio_sample[1] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[2]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net280),
    .D(_0263_),
    .Q_N(_4631_),
    .Q(\vgademo.scanline_audio_sample[2] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[3]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net281),
    .D(_0264_),
    .Q_N(_4630_),
    .Q(\vgademo.scanline_audio_sample[3] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[4]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net282),
    .D(_0265_),
    .Q_N(_4629_),
    .Q(\vgademo.scanline_audio_sample[4] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net283),
    .D(_0266_),
    .Q_N(_4628_),
    .Q(\vgademo.scanline_audio_sample[5] ));
 sg13g2_dfrbp_1 \vgademo.scanline_audio_sample[6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net284),
    .D(_0267_),
    .Q_N(_4627_),
    .Q(\vgademo.scanline_audio_sample[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.beat_div[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0268_),
    .Q_N(_0075_),
    .Q(\vgademo.audio_beat_out[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.beat_div[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0269_),
    .Q_N(_0076_),
    .Q(\vgademo.audio_beat_out[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.beat_div[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net145),
    .D(_0270_),
    .Q_N(_0080_),
    .Q(\vgademo.audio_beat_out[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.beat_div[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0271_),
    .Q_N(_0074_),
    .Q(\vgademo.audio_beat_out[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.beat_div[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net146),
    .D(_0272_),
    .Q_N(_0073_),
    .Q(\vgademo.audio_beat_out[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.kick_frames[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0273_),
    .Q_N(_0077_),
    .Q(\vgademo.audio_kick_frames[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.kick_frames[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0274_),
    .Q_N(_0016_),
    .Q(\vgademo.audio_kick_frames[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.kick_frames[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net146),
    .D(_0275_),
    .Q_N(_4626_),
    .Q(\vgademo.audio_kick_frames[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net128),
    .D(_0276_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[0] ),
    .Q(_0087_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[10]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(_0277_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[10] ),
    .Q(_0088_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[11]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(_0278_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[11] ),
    .Q(_0089_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[12]$_DFFE_PN1P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(_0279_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[12] ),
    .Q(_0090_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net128),
    .D(_0280_),
    .Q_N(_0085_),
    .Q(\vgademo.soundtrack.noise_lfsr[13] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net128),
    .D(_0281_),
    .Q_N(_4625_),
    .Q(\vgademo.soundtrack.noise_lfsr[14] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net128),
    .D(_0282_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[1] ),
    .Q(_0091_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net131),
    .D(_0283_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[2] ),
    .Q(_0092_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(_0284_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[3] ),
    .Q(_0093_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(_0285_),
    .Q_N(_0063_),
    .Q(\vgademo.soundtrack.noise_lfsr[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net132),
    .D(_0286_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[5] ),
    .Q(_0094_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net132),
    .D(_0287_),
    .Q_N(_0084_),
    .Q(\vgademo.soundtrack.noise_lfsr[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net130),
    .D(_0288_),
    .Q_N(\vgademo.soundtrack.noise_lfsr[7] ),
    .Q(_0095_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net132),
    .D(_0289_),
    .Q_N(_0083_),
    .Q(\vgademo.soundtrack.noise_lfsr[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_lfsr[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(_0290_),
    .Q_N(_4624_),
    .Q(\vgademo.soundtrack.noise_lfsr[9] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_vol[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net134),
    .D(_0291_),
    .Q_N(\vgademo.audio_snare_frames[0] ),
    .Q(_0096_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_vol[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net134),
    .D(_0292_),
    .Q_N(\vgademo.audio_snare_frames[1] ),
    .Q(_0097_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_vol[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net138),
    .D(_0293_),
    .Q_N(\vgademo.audio_snare_frames[2] ),
    .Q(_0098_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.noise_vol[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net134),
    .D(_0294_),
    .Q_N(\vgademo.audio_snare_frames[3] ),
    .Q(_0099_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.out$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net285),
    .D(_0295_),
    .Q_N(_4623_),
    .Q(audio));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net286),
    .D(_0296_),
    .Q_N(_4622_),
    .Q(\vgademo.soundtrack.pulse_osc_p[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[10]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net287),
    .D(_0297_),
    .Q_N(_4621_),
    .Q(\vgademo.soundtrack.pulse_osc_p[10] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[11]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net288),
    .D(_0298_),
    .Q_N(_4620_),
    .Q(\vgademo.soundtrack.pulse_osc_p[11] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[12]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net289),
    .D(_0299_),
    .Q_N(_0062_),
    .Q(\vgademo.soundtrack.pulse_osc_p[12] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net290),
    .D(_0300_),
    .Q_N(_0061_),
    .Q(\vgademo.soundtrack.pulse_osc_p[13] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[1]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net291),
    .D(_0301_),
    .Q_N(_4619_),
    .Q(\vgademo.soundtrack.pulse_osc_p[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net292),
    .D(_0302_),
    .Q_N(_4618_),
    .Q(\vgademo.soundtrack.pulse_osc_p[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net293),
    .D(_0303_),
    .Q_N(_4617_),
    .Q(\vgademo.soundtrack.pulse_osc_p[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net294),
    .D(_0304_),
    .Q_N(_4616_),
    .Q(\vgademo.soundtrack.pulse_osc_p[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[5]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net295),
    .D(_0305_),
    .Q_N(_4615_),
    .Q(\vgademo.soundtrack.pulse_osc_p[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net296),
    .D(_0306_),
    .Q_N(_4614_),
    .Q(\vgademo.soundtrack.pulse_osc_p[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net297),
    .D(_0307_),
    .Q_N(_4613_),
    .Q(\vgademo.soundtrack.pulse_osc_p[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[8]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net298),
    .D(_0308_),
    .Q_N(_0064_),
    .Q(\vgademo.soundtrack.pulse_osc_p[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_osc_p[9]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net299),
    .D(_0309_),
    .Q_N(_4612_),
    .Q(\vgademo.soundtrack.pulse_osc_p[9] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_vol[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0310_),
    .Q_N(\vgademo.soundtrack.pulse_vol[0] ),
    .Q(_0100_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_vol[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0311_),
    .Q_N(\vgademo.soundtrack.pulse_vol[1] ),
    .Q(_0101_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_vol[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0312_),
    .Q_N(\vgademo.soundtrack.pulse_vol[2] ),
    .Q(_0102_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.pulse_vol[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net139),
    .D(_0313_),
    .Q_N(\vgademo.soundtrack.pulse_vol[3] ),
    .Q(_0103_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[0]$_DFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net131),
    .D(\vgademo.soundtrack.sample_div_[0] ),
    .Q_N(\vgademo.soundtrack.sample_div_[0] ),
    .Q(\vgademo.soundtrack.sample_div[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[1]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net129),
    .D(\vgademo.soundtrack.sample_div_[1] ),
    .Q_N(_4747_),
    .Q(\vgademo.soundtrack.sample_div[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[2]$_DFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net129),
    .D(\vgademo.soundtrack.sample_div_[2] ),
    .Q_N(_4748_),
    .Q(\vgademo.soundtrack.sample_div[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[3]$_DFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net128),
    .D(\vgademo.soundtrack.sample_div_[3] ),
    .Q_N(_4749_),
    .Q(\vgademo.soundtrack.sample_div[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[4]$_DFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net128),
    .D(\vgademo.soundtrack.sample_div_[4] ),
    .Q_N(_4750_),
    .Q(\vgademo.soundtrack.sample_div[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[5]$_DFF_PN0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net128),
    .D(\vgademo.soundtrack.sample_div_[5] ),
    .Q_N(_4751_),
    .Q(\vgademo.soundtrack.sample_div[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[6]$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net128),
    .D(\vgademo.soundtrack.sample_div_[6] ),
    .Q_N(_4752_),
    .Q(\vgademo.soundtrack.sample_div[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[7]$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net130),
    .D(\vgademo.soundtrack.sample_div_[7] ),
    .Q_N(_4753_),
    .Q(\vgademo.soundtrack.sample_div[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[8]$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net132),
    .D(\vgademo.soundtrack.sample_div_[8] ),
    .Q_N(_4754_),
    .Q(\vgademo.soundtrack.sample_div[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sample_div[9]$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net132),
    .D(\vgademo.soundtrack.sample_div_[9] ),
    .Q_N(_4755_),
    .Q(\vgademo.soundtrack.sample_div[9] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[0]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net139),
    .D(\vgademo.soundtrack.sigma_delta_accum_[0] ),
    .Q_N(_4756_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[10]$_DFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net135),
    .D(\vgademo.soundtrack.sigma_delta_accum_[10] ),
    .Q_N(_4757_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[10] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[11]$_DFF_PN0_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net137),
    .D(\vgademo.soundtrack.sigma_delta_accum_[11] ),
    .Q_N(_4758_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[11] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[12]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net137),
    .D(\vgademo.soundtrack.sigma_delta_accum_[12] ),
    .Q_N(_4759_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[12] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[13]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net137),
    .D(\vgademo.soundtrack.sigma_delta_accum_[13] ),
    .Q_N(_4760_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[13] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[14]$_DFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net138),
    .D(\vgademo.soundtrack.sigma_delta_accum_[14] ),
    .Q_N(_4761_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[14] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[15]$_DFF_PN0_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net138),
    .D(\vgademo.soundtrack.sigma_delta_accum_[15] ),
    .Q_N(_4762_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[15] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[1]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net139),
    .D(\vgademo.soundtrack.sigma_delta_accum_[1] ),
    .Q_N(_4763_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[2]$_DFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net139),
    .D(\vgademo.soundtrack.sigma_delta_accum_[2] ),
    .Q_N(_4764_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[3]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net139),
    .D(\vgademo.soundtrack.sigma_delta_accum_[3] ),
    .Q_N(_4765_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[4]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net131),
    .D(\vgademo.soundtrack.sigma_delta_accum_[4] ),
    .Q_N(_4766_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[5]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net131),
    .D(\vgademo.soundtrack.sigma_delta_accum_[5] ),
    .Q_N(_4767_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[6]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net131),
    .D(\vgademo.soundtrack.sigma_delta_accum_[6] ),
    .Q_N(_4768_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[7]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net131),
    .D(\vgademo.soundtrack.sigma_delta_accum_[7] ),
    .Q_N(_4769_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[8]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net137),
    .D(\vgademo.soundtrack.sigma_delta_accum_[8] ),
    .Q_N(_4770_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.sigma_delta_accum[9]$_DFF_PN0_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net134),
    .D(\vgademo.soundtrack.sigma_delta_accum_[9] ),
    .Q_N(_4611_),
    .Q(\vgademo.soundtrack.sigma_delta_accum[9] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net147),
    .D(_0314_),
    .Q_N(\vgademo.audio_songpos[0] ),
    .Q(_0104_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0315_),
    .Q_N(\vgademo.audio_songpos[1] ),
    .Q(_0105_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[2]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0316_),
    .Q_N(\vgademo.audio_songpos[2] ),
    .Q(_0106_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0317_),
    .Q_N(\vgademo.audio_songpos[3] ),
    .Q(_0107_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[4]$_DFFE_PN1P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net148),
    .D(_0318_),
    .Q_N(\vgademo.audio_songpos[4] ),
    .Q(_0108_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[5]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0319_),
    .Q_N(\vgademo.audio_songpos[5] ),
    .Q(_0109_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[6]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0320_),
    .Q_N(\vgademo.audio_songpos[6] ),
    .Q(_0110_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.songpos[7]$_DFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net148),
    .D(_0321_),
    .Q_N(\vgademo.audio_songpos[7] ),
    .Q(_0111_));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net132),
    .D(_0322_),
    .Q_N(\vgademo.soundtrack.tick_div_[0] ),
    .Q(\vgademo.soundtrack.tick_div[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net132),
    .D(_0323_),
    .Q_N(_4610_),
    .Q(\vgademo.soundtrack.tick_div[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net133),
    .D(_0324_),
    .Q_N(_4609_),
    .Q(\vgademo.soundtrack.tick_div[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net133),
    .D(_0325_),
    .Q_N(_4608_),
    .Q(\vgademo.soundtrack.tick_div[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net132),
    .D(_0326_),
    .Q_N(_4607_),
    .Q(\vgademo.soundtrack.tick_div[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net133),
    .D(_0327_),
    .Q_N(_4606_),
    .Q(\vgademo.soundtrack.tick_div[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net135),
    .D(_0328_),
    .Q_N(_4605_),
    .Q(\vgademo.soundtrack.tick_div[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tick_div[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net134),
    .D(_0329_),
    .Q_N(_4604_),
    .Q(\vgademo.soundtrack.tick_div[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net145),
    .D(_0330_),
    .Q_N(_4603_),
    .Q(\vgademo.soundtrack.tri_osc_i[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net147),
    .D(_0331_),
    .Q_N(_4602_),
    .Q(\vgademo.soundtrack.tri_osc_i[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net147),
    .D(_0332_),
    .Q_N(_4601_),
    .Q(\vgademo.soundtrack.tri_osc_i[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0333_),
    .Q_N(_4600_),
    .Q(\vgademo.soundtrack.tri_osc_i[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net145),
    .D(_0334_),
    .Q_N(_4599_),
    .Q(\vgademo.soundtrack.tri_osc_i[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net145),
    .D(_0335_),
    .Q_N(_4598_),
    .Q(\vgademo.soundtrack.tri_osc_i[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0336_),
    .Q_N(_4597_),
    .Q(\vgademo.soundtrack.tri_osc_i[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0337_),
    .Q_N(_4596_),
    .Q(\vgademo.soundtrack.tri_osc_i[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_i[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net145),
    .D(_0338_),
    .Q_N(_4595_),
    .Q(\vgademo.soundtrack.tri_osc_i[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[0]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net300),
    .D(_0339_),
    .Q_N(_4594_),
    .Q(\vgademo.soundtrack.tri_osc_p[0] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[10]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net301),
    .D(_0340_),
    .Q_N(_4593_),
    .Q(\vgademo.soundtrack.tri_osc_p[10] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net302),
    .D(_0341_),
    .Q_N(_4592_),
    .Q(\vgademo.soundtrack.tri_osc_p[11] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[12]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net303),
    .D(_0342_),
    .Q_N(_4591_),
    .Q(\vgademo.soundtrack.tri_osc_p[12] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[13]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net304),
    .D(_0343_),
    .Q_N(_4590_),
    .Q(\vgademo.soundtrack.tri_osc_p[13] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[14]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net305),
    .D(_0344_),
    .Q_N(_4589_),
    .Q(\vgademo.soundtrack.tri_osc_p[14] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net306),
    .D(_0345_),
    .Q_N(_4588_),
    .Q(\vgademo.soundtrack.tri_osc_p[15] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[1]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net307),
    .D(_0346_),
    .Q_N(_4587_),
    .Q(\vgademo.soundtrack.tri_osc_p[1] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[2]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net308),
    .D(_0347_),
    .Q_N(_4586_),
    .Q(\vgademo.soundtrack.tri_osc_p[2] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[3]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net309),
    .D(_0348_),
    .Q_N(_4585_),
    .Q(\vgademo.soundtrack.tri_osc_p[3] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[4]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net310),
    .D(_0349_),
    .Q_N(_4584_),
    .Q(\vgademo.soundtrack.tri_osc_p[4] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[5]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net311),
    .D(_0350_),
    .Q_N(_4583_),
    .Q(\vgademo.soundtrack.tri_osc_p[5] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net312),
    .D(_0351_),
    .Q_N(_4582_),
    .Q(\vgademo.soundtrack.tri_osc_p[6] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[7]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net313),
    .D(_0352_),
    .Q_N(_4581_),
    .Q(\vgademo.soundtrack.tri_osc_p[7] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[8]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net314),
    .D(_0353_),
    .Q_N(_4580_),
    .Q(\vgademo.soundtrack.tri_osc_p[8] ));
 sg13g2_dfrbp_1 \vgademo.soundtrack.tri_osc_p[9]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net315),
    .D(_0354_),
    .Q_N(_0065_),
    .Q(\vgademo.soundtrack.tri_osc_p[9] ));
 sg13g2_dfrbp_1 \vgademo.v_count[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0355_),
    .Q_N(_0018_),
    .Q(\vgademo.bayer_j[0] ));
 sg13g2_dfrbp_1 \vgademo.v_count[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0356_),
    .Q_N(_0021_),
    .Q(\vgademo.bayer_j[1] ));
 sg13g2_dfrbp_1 \vgademo.v_count[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0357_),
    .Q_N(_0020_),
    .Q(\vgademo.v_count[2] ));
 sg13g2_dfrbp_1 \vgademo.v_count[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0358_),
    .Q_N(_0023_),
    .Q(\vgademo.v_count[3] ));
 sg13g2_dfrbp_1 \vgademo.v_count[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0359_),
    .Q_N(_0027_),
    .Q(\vgademo.v_count[4] ));
 sg13g2_dfrbp_1 \vgademo.v_count[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net151),
    .D(_0360_),
    .Q_N(_0032_),
    .Q(\vgademo.v_count[5] ));
 sg13g2_dfrbp_1 \vgademo.v_count[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net151),
    .D(_0361_),
    .Q_N(_0031_),
    .Q(\vgademo.v_count[6] ));
 sg13g2_dfrbp_1 \vgademo.v_count[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net144),
    .D(_0362_),
    .Q_N(_0038_),
    .Q(\vgademo.v_count[7] ));
 sg13g2_dfrbp_1 \vgademo.v_count[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net149),
    .D(_0363_),
    .Q_N(_0036_),
    .Q(\vgademo.v_count[8] ));
 sg13g2_dfrbp_1 \vgademo.v_count[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net149),
    .D(_0364_),
    .Q_N(_0040_),
    .Q(\vgademo.v_count[9] ));
 sg13g2_dfrbp_1 \vgademo.vsync$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net316),
    .D(_0012_),
    .Q_N(_4579_),
    .Q(\vgademo.vsync ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[7]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_3424_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_3822_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_3375_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_3261_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_2943_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_2967_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_2928_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_3027_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2894_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_3000_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_3382_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_3139_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_2764_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_2756_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0403_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_3333_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2755_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0671_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2481_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2406_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1354_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1227_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2412_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2407_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2348_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1226_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1220_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1089_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0837_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1088_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0730_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0643_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0637_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0608_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0559_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_3888_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_3815_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2130_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2129_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1100_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0905_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0640_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0634_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0556_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0550_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0542_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0537_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2049_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0953_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0785_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0555_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0545_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0541_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0411_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0939_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0870_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0862_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0861_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_0437_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0421_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_4576_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_4575_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_4404_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2493_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2060_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2045_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2142_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2103_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_2087_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1740_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1701_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1133_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1018_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0777_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1734_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1730_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1729_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1690_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1683_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1639_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1637_),
    .X(net91));
 sg13g2_buf_4 fanout92 (.X(net92),
    .A(_1633_));
 sg13g2_buf_2 fanout93 (.A(_0829_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_0818_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0813_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0787_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0772_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0764_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0757_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_0599_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_0579_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_4500_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_4382_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_4348_),
    .X(net104));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_4346_));
 sg13g2_buf_2 fanout106 (.A(_4337_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_4332_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1658_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1643_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_0899_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0897_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0875_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_0872_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_0864_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_0826_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_0768_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_0766_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_0765_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_0601_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0560_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_4453_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_4446_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_4284_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_4283_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_4277_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_4276_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_4275_),
    .X(net127));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net130));
 sg13g2_buf_2 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net131));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(net140));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(net136));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net136));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net136));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net140),
    .X(net136));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net140));
 sg13g2_buf_2 fanout138 (.A(net140),
    .X(net138));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net140));
 sg13g2_buf_1 fanout140 (.A(net152),
    .X(net140));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(net142));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(net144));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(net144));
 sg13g2_buf_2 fanout144 (.A(net152),
    .X(net144));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net147));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(net147));
 sg13g2_buf_2 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(net152));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(net151));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(net151));
 sg13g2_buf_2 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_1 fanout152 (.A(net1),
    .X(net152));
 sg13g2_tielo _9281__153 (.L_LO(net153));
 sg13g2_tielo _9282__154 (.L_LO(net154));
 sg13g2_tielo _9283__155 (.L_LO(net155));
 sg13g2_tielo _9284__156 (.L_LO(net156));
 sg13g2_tielo _9285__157 (.L_LO(net157));
 sg13g2_tielo _9286__158 (.L_LO(net158));
 sg13g2_tielo _9287__159 (.L_LO(net159));
 sg13g2_tielo _9289__160 (.L_LO(net160));
 sg13g2_tielo _9290__161 (.L_LO(net161));
 sg13g2_tielo _9291__162 (.L_LO(net162));
 sg13g2_tielo _9292__163 (.L_LO(net163));
 sg13g2_tielo _9293__164 (.L_LO(net164));
 sg13g2_tielo _9294__165 (.L_LO(net165));
 sg13g2_tielo _9295__166 (.L_LO(net166));
 sg13g2_tiehi \vgademo.b_cos[0]$_DFFE_PP__168  (.L_HI(net168));
 sg13g2_tiehi \vgademo.b_cos[10]$_DFFE_PP__169  (.L_HI(net169));
 sg13g2_tiehi \vgademo.b_cos[11]$_DFFE_PP__170  (.L_HI(net170));
 sg13g2_tiehi \vgademo.b_cos[1]$_DFFE_PP__171  (.L_HI(net171));
 sg13g2_tiehi \vgademo.b_cos[2]$_DFFE_PP__172  (.L_HI(net172));
 sg13g2_tiehi \vgademo.b_cos[3]$_DFFE_PP__173  (.L_HI(net173));
 sg13g2_tiehi \vgademo.b_cos[4]$_DFFE_PP__174  (.L_HI(net174));
 sg13g2_tiehi \vgademo.b_cos[5]$_DFFE_PP__175  (.L_HI(net175));
 sg13g2_tiehi \vgademo.b_cos[6]$_DFFE_PP__176  (.L_HI(net176));
 sg13g2_tiehi \vgademo.b_cos[7]$_DFFE_PP__177  (.L_HI(net177));
 sg13g2_tiehi \vgademo.b_cos[8]$_DFFE_PP__178  (.L_HI(net178));
 sg13g2_tiehi \vgademo.b_cos[9]$_DFFE_PP__179  (.L_HI(net179));
 sg13g2_tiehi \vgademo.b_out[0]$_SDFF_PN0__180  (.L_HI(net180));
 sg13g2_tiehi \vgademo.b_out[1]$_SDFF_PN0__181  (.L_HI(net181));
 sg13g2_tiehi \vgademo.b_sin[0]$_DFFE_PP__182  (.L_HI(net182));
 sg13g2_tiehi \vgademo.b_sin[10]$_DFFE_PP__183  (.L_HI(net183));
 sg13g2_tiehi \vgademo.b_sin[11]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \vgademo.b_sin[1]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \vgademo.b_sin[2]$_DFFE_PP__186  (.L_HI(net186));
 sg13g2_tiehi \vgademo.b_sin[3]$_DFFE_PP__187  (.L_HI(net187));
 sg13g2_tiehi \vgademo.b_sin[4]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \vgademo.b_sin[5]$_DFFE_PP__189  (.L_HI(net189));
 sg13g2_tiehi \vgademo.b_sin[6]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \vgademo.b_sin[7]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \vgademo.b_sin[8]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \vgademo.b_sin[9]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \vgademo.g_out[0]$_SDFF_PN0__194  (.L_HI(net194));
 sg13g2_tiehi \vgademo.g_out[1]$_SDFF_PN0__195  (.L_HI(net195));
 sg13g2_tiehi \vgademo.hsync$_DFF_P__196  (.L_HI(net196));
 sg13g2_tiehi \vgademo.linelfsr[0]$_SDFFCE_PN0P__197  (.L_HI(net197));
 sg13g2_tiehi \vgademo.linelfsr[10]$_SDFFCE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \vgademo.linelfsr[11]$_SDFFCE_PN1P__199  (.L_HI(net199));
 sg13g2_tiehi \vgademo.linelfsr[12]$_SDFFCE_PN1P__200  (.L_HI(net200));
 sg13g2_tiehi \vgademo.linelfsr[1]$_SDFFCE_PN1P__201  (.L_HI(net201));
 sg13g2_tiehi \vgademo.linelfsr[2]$_SDFFCE_PN0P__202  (.L_HI(net202));
 sg13g2_tiehi \vgademo.linelfsr[3]$_SDFFCE_PN1P__203  (.L_HI(net203));
 sg13g2_tiehi \vgademo.linelfsr[4]$_SDFFCE_PN1P__204  (.L_HI(net204));
 sg13g2_tiehi \vgademo.linelfsr[5]$_SDFFCE_PN1P__205  (.L_HI(net205));
 sg13g2_tiehi \vgademo.linelfsr[6]$_SDFFCE_PN1P__206  (.L_HI(net206));
 sg13g2_tiehi \vgademo.linelfsr[7]$_SDFFCE_PN1P__207  (.L_HI(net207));
 sg13g2_tiehi \vgademo.linelfsr[8]$_SDFFCE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \vgademo.linelfsr[9]$_SDFFCE_PN1P__209  (.L_HI(net209));
 sg13g2_tiehi \vgademo.plane_du[0]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \vgademo.plane_du[10]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \vgademo.plane_du[1]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \vgademo.plane_du[2]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \vgademo.plane_du[3]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \vgademo.plane_du[4]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \vgademo.plane_du[5]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \vgademo.plane_du[6]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \vgademo.plane_du[7]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \vgademo.plane_du[8]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \vgademo.plane_du[9]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \vgademo.plane_dx_div.d[16]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \vgademo.plane_dx_div.d[17]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \vgademo.plane_dx_div.d[18]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \vgademo.plane_dx_div.d[19]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \vgademo.plane_dx_div.d[20]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \vgademo.plane_dx_div.d[21]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \vgademo.plane_dx_div.d[22]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \vgademo.plane_dx_div.d[23]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \vgademo.plane_dx_div.d[24]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \vgademo.plane_dx_div.i[0]$_SDFFE_PP1P__230  (.L_HI(net230));
 sg13g2_tiehi \vgademo.plane_dx_div.i[1]$_SDFFE_PP0P__231  (.L_HI(net231));
 sg13g2_tiehi \vgademo.plane_dx_div.i[2]$_SDFFE_PP0P__232  (.L_HI(net232));
 sg13g2_tiehi \vgademo.plane_dx_div.i[3]$_SDFFE_PP0P__233  (.L_HI(net233));
 sg13g2_tiehi \vgademo.plane_dx_div.q[0]$_SDFFE_PP1P__234  (.L_HI(net234));
 sg13g2_tiehi \vgademo.plane_dx_div.q[1]$_SDFFE_PP0P__235  (.L_HI(net235));
 sg13g2_tiehi \vgademo.plane_dx_div.q[2]$_SDFFE_PP0P__236  (.L_HI(net236));
 sg13g2_tiehi \vgademo.plane_dx_div.q[3]$_SDFFE_PP0P__237  (.L_HI(net237));
 sg13g2_tiehi \vgademo.plane_dx_div.q[4]$_SDFFE_PP0P__238  (.L_HI(net238));
 sg13g2_tiehi \vgademo.plane_dx_div.q[5]$_SDFFE_PP0P__239  (.L_HI(net239));
 sg13g2_tiehi \vgademo.plane_dx_div.q[6]$_SDFFE_PP0P__240  (.L_HI(net240));
 sg13g2_tiehi \vgademo.plane_dx_div.q[7]$_SDFFE_PP0P__241  (.L_HI(net241));
 sg13g2_tiehi \vgademo.plane_dx_div.q[8]$_SDFFE_PP0P__242  (.L_HI(net242));
 sg13g2_tiehi \vgademo.plane_dx_div.q[9]$_SDFFE_PP0P__243  (.L_HI(net243));
 sg13g2_tiehi \vgademo.plane_dx_div.r[16]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \vgademo.plane_dx_div.r[17]$_DFFE_PP__245  (.L_HI(net245));
 sg13g2_tiehi \vgademo.plane_dx_div.r[18]$_DFFE_PP__246  (.L_HI(net246));
 sg13g2_tiehi \vgademo.plane_dx_div.r[19]$_DFFE_PP__247  (.L_HI(net247));
 sg13g2_tiehi \vgademo.plane_dx_div.r[20]$_DFFE_PP__248  (.L_HI(net248));
 sg13g2_tiehi \vgademo.plane_dx_div.r[21]$_DFFE_PP__249  (.L_HI(net249));
 sg13g2_tiehi \vgademo.plane_dx_div.r[22]$_DFFE_PP__250  (.L_HI(net250));
 sg13g2_tiehi \vgademo.plane_dx_div.r[23]$_DFFE_PP__251  (.L_HI(net251));
 sg13g2_tiehi \vgademo.plane_dx_div.r[24]$_DFFE_PP__252  (.L_HI(net252));
 sg13g2_tiehi \vgademo.plane_dx_div.r[25]$_DFFE_PP__253  (.L_HI(net253));
 sg13g2_tiehi \vgademo.plane_u[0]$_SDFFCE_PP0P__254  (.L_HI(net254));
 sg13g2_tiehi \vgademo.plane_u[10]$_DFFE_PP__255  (.L_HI(net255));
 sg13g2_tiehi \vgademo.plane_u[11]$_DFFE_PP__256  (.L_HI(net256));
 sg13g2_tiehi \vgademo.plane_u[12]$_DFFE_PP__257  (.L_HI(net257));
 sg13g2_tiehi \vgademo.plane_u[13]$_DFFE_PP__258  (.L_HI(net258));
 sg13g2_tiehi \vgademo.plane_u[14]$_DFFE_PP__259  (.L_HI(net259));
 sg13g2_tiehi \vgademo.plane_u[15]$_DFFE_PP__260  (.L_HI(net260));
 sg13g2_tiehi \vgademo.plane_u[16]$_DFFE_PP__261  (.L_HI(net261));
 sg13g2_tiehi \vgademo.plane_u[17]$_DFFE_PP__262  (.L_HI(net262));
 sg13g2_tiehi \vgademo.plane_u[18]$_DFFE_PP__263  (.L_HI(net263));
 sg13g2_tiehi \vgademo.plane_u[19]$_DFFE_PP__264  (.L_HI(net264));
 sg13g2_tiehi \vgademo.plane_u[1]$_DFFE_PP__265  (.L_HI(net265));
 sg13g2_tiehi \vgademo.plane_u[20]$_DFFE_PP__266  (.L_HI(net266));
 sg13g2_tiehi \vgademo.plane_u[21]$_DFFE_PP__267  (.L_HI(net267));
 sg13g2_tiehi \vgademo.plane_u[2]$_DFFE_PP__268  (.L_HI(net268));
 sg13g2_tiehi \vgademo.plane_u[3]$_DFFE_PP__269  (.L_HI(net269));
 sg13g2_tiehi \vgademo.plane_u[4]$_DFFE_PP__270  (.L_HI(net270));
 sg13g2_tiehi \vgademo.plane_u[5]$_DFFE_PP__271  (.L_HI(net271));
 sg13g2_tiehi \vgademo.plane_u[6]$_DFFE_PP__272  (.L_HI(net272));
 sg13g2_tiehi \vgademo.plane_u[7]$_DFFE_PP__273  (.L_HI(net273));
 sg13g2_tiehi \vgademo.plane_u[8]$_DFFE_PP__274  (.L_HI(net274));
 sg13g2_tiehi \vgademo.plane_u[9]$_DFFE_PP__275  (.L_HI(net275));
 sg13g2_tiehi \vgademo.r_out[0]$_SDFF_PN0__276  (.L_HI(net276));
 sg13g2_tiehi \vgademo.r_out[1]$_SDFF_PN0__277  (.L_HI(net277));
 sg13g2_tiehi \vgademo.scanline_audio_sample[0]$_DFFE_PP__278  (.L_HI(net278));
 sg13g2_tiehi \vgademo.scanline_audio_sample[1]$_DFFE_PP__279  (.L_HI(net279));
 sg13g2_tiehi \vgademo.scanline_audio_sample[2]$_DFFE_PP__280  (.L_HI(net280));
 sg13g2_tiehi \vgademo.scanline_audio_sample[3]$_DFFE_PP__281  (.L_HI(net281));
 sg13g2_tiehi \vgademo.scanline_audio_sample[4]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \vgademo.scanline_audio_sample[5]$_DFFE_PP__283  (.L_HI(net283));
 sg13g2_tiehi \vgademo.scanline_audio_sample[6]$_DFFE_PP__284  (.L_HI(net284));
 sg13g2_tiehi \vgademo.soundtrack.out$_DFFE_PP__285  (.L_HI(net285));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[0]$_DFFE_PP__286  (.L_HI(net286));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[10]$_DFFE_PP__287  (.L_HI(net287));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[11]$_DFFE_PP__288  (.L_HI(net288));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[12]$_DFFE_PP__289  (.L_HI(net289));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[13]$_DFFE_PP__290  (.L_HI(net290));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[1]$_DFFE_PP__291  (.L_HI(net291));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[2]$_DFFE_PP__292  (.L_HI(net292));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[3]$_DFFE_PP__293  (.L_HI(net293));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[4]$_DFFE_PP__294  (.L_HI(net294));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[5]$_DFFE_PP__295  (.L_HI(net295));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[6]$_DFFE_PP__296  (.L_HI(net296));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[7]$_DFFE_PP__297  (.L_HI(net297));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[8]$_DFFE_PP__298  (.L_HI(net298));
 sg13g2_tiehi \vgademo.soundtrack.pulse_osc_p[9]$_DFFE_PP__299  (.L_HI(net299));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[0]$_DFFE_PP__300  (.L_HI(net300));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[10]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[11]$_DFFE_PP__302  (.L_HI(net302));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[12]$_DFFE_PP__303  (.L_HI(net303));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[13]$_DFFE_PP__304  (.L_HI(net304));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[14]$_DFFE_PP__305  (.L_HI(net305));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[15]$_DFFE_PP__306  (.L_HI(net306));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[1]$_DFFE_PP__307  (.L_HI(net307));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[2]$_DFFE_PP__308  (.L_HI(net308));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[3]$_DFFE_PP__309  (.L_HI(net309));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[4]$_DFFE_PP__310  (.L_HI(net310));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[5]$_DFFE_PP__311  (.L_HI(net311));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[6]$_DFFE_PP__312  (.L_HI(net312));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[7]$_DFFE_PP__313  (.L_HI(net313));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[8]$_DFFE_PP__314  (.L_HI(net314));
 sg13g2_tiehi \vgademo.soundtrack.tri_osc_p[9]$_DFFE_PP__315  (.L_HI(net315));
 sg13g2_tiehi \vgademo.vsync$_DFF_P__316  (.L_HI(net316));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_2 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_2 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_2 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_2 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_2 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload3 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_2 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_41_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_35_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_leaf_26_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_27_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_buf_16 clkload12 (.A(clknet_leaf_25_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_leaf_10_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_13_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_21_clk));
 sg13g2_inv_1 clkload18 (.A(clknet_leaf_34_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_14_clk));
 sg13g2_buf_16 clkload20 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_17_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0011_));
 sg13g2_antennanp ANTENNA_2 (.A(_0012_));
 sg13g2_antennanp ANTENNA_3 (.A(_0011_));
 sg13g2_antennanp ANTENNA_4 (.A(_0012_));
 sg13g2_antennanp ANTENNA_5 (.A(_0011_));
 sg13g2_antennanp ANTENNA_6 (.A(_0012_));
 sg13g2_antennanp ANTENNA_7 (.A(_0011_));
 sg13g2_antennanp ANTENNA_8 (.A(_0012_));
 sg13g2_antennanp ANTENNA_9 (.A(_0011_));
 sg13g2_antennanp ANTENNA_10 (.A(_0012_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_4 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_26 ();
 sg13g2_fill_2 FILLER_0_33 ();
 sg13g2_fill_1 FILLER_0_35 ();
 sg13g2_fill_1 FILLER_0_48 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_117 ();
 sg13g2_decap_8 FILLER_0_124 ();
 sg13g2_decap_8 FILLER_0_131 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_4 FILLER_0_166 ();
 sg13g2_fill_1 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_4 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_145 ();
 sg13g2_decap_8 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_184 ();
 sg13g2_decap_8 FILLER_1_228 ();
 sg13g2_decap_8 FILLER_1_235 ();
 sg13g2_fill_2 FILLER_1_242 ();
 sg13g2_fill_1 FILLER_1_252 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_8 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_1_412 ();
 sg13g2_decap_8 FILLER_1_419 ();
 sg13g2_decap_4 FILLER_1_426 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_4 FILLER_2_83 ();
 sg13g2_fill_1 FILLER_2_87 ();
 sg13g2_decap_4 FILLER_2_100 ();
 sg13g2_decap_4 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_124 ();
 sg13g2_fill_1 FILLER_2_129 ();
 sg13g2_decap_8 FILLER_2_136 ();
 sg13g2_decap_8 FILLER_2_143 ();
 sg13g2_decap_8 FILLER_2_150 ();
 sg13g2_decap_4 FILLER_2_157 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_174 ();
 sg13g2_fill_1 FILLER_2_184 ();
 sg13g2_fill_2 FILLER_2_193 ();
 sg13g2_fill_2 FILLER_2_200 ();
 sg13g2_fill_2 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_213 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_fill_1 FILLER_2_267 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_fill_2 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_26 ();
 sg13g2_fill_1 FILLER_3_33 ();
 sg13g2_fill_1 FILLER_3_43 ();
 sg13g2_fill_2 FILLER_3_52 ();
 sg13g2_decap_4 FILLER_3_120 ();
 sg13g2_fill_2 FILLER_3_128 ();
 sg13g2_fill_2 FILLER_3_164 ();
 sg13g2_fill_1 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_208 ();
 sg13g2_fill_1 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_289 ();
 sg13g2_fill_2 FILLER_3_317 ();
 sg13g2_fill_2 FILLER_3_323 ();
 sg13g2_fill_1 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_419 ();
 sg13g2_decap_4 FILLER_3_426 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_83 ();
 sg13g2_fill_2 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_118 ();
 sg13g2_fill_2 FILLER_4_129 ();
 sg13g2_fill_1 FILLER_4_162 ();
 sg13g2_fill_2 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_217 ();
 sg13g2_decap_4 FILLER_4_242 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_fill_2 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_290 ();
 sg13g2_fill_2 FILLER_4_332 ();
 sg13g2_fill_2 FILLER_4_361 ();
 sg13g2_fill_1 FILLER_4_371 ();
 sg13g2_fill_1 FILLER_4_391 ();
 sg13g2_fill_2 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_7 ();
 sg13g2_fill_2 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_fill_2 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_202 ();
 sg13g2_decap_4 FILLER_5_212 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_220 ();
 sg13g2_decap_4 FILLER_5_225 ();
 sg13g2_fill_2 FILLER_5_229 ();
 sg13g2_fill_1 FILLER_5_315 ();
 sg13g2_fill_2 FILLER_5_327 ();
 sg13g2_fill_1 FILLER_5_344 ();
 sg13g2_fill_1 FILLER_5_350 ();
 sg13g2_fill_1 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_416 ();
 sg13g2_decap_8 FILLER_5_423 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_115 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_255 ();
 sg13g2_fill_2 FILLER_6_294 ();
 sg13g2_fill_1 FILLER_6_313 ();
 sg13g2_fill_1 FILLER_6_352 ();
 sg13g2_fill_2 FILLER_6_357 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_fill_1 FILLER_6_371 ();
 sg13g2_fill_1 FILLER_6_393 ();
 sg13g2_fill_1 FILLER_6_398 ();
 sg13g2_fill_2 FILLER_6_404 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_fill_2 FILLER_7_121 ();
 sg13g2_decap_4 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_153 ();
 sg13g2_fill_1 FILLER_7_159 ();
 sg13g2_fill_2 FILLER_7_164 ();
 sg13g2_fill_1 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_176 ();
 sg13g2_decap_4 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_fill_1 FILLER_7_211 ();
 sg13g2_fill_1 FILLER_7_233 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_fill_1 FILLER_7_244 ();
 sg13g2_fill_2 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_265 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_326 ();
 sg13g2_fill_2 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_413 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_decap_4 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_25 ();
 sg13g2_fill_1 FILLER_8_73 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_128 ();
 sg13g2_fill_2 FILLER_8_132 ();
 sg13g2_fill_1 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_322 ();
 sg13g2_fill_2 FILLER_8_387 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_9 ();
 sg13g2_fill_1 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_68 ();
 sg13g2_fill_1 FILLER_9_82 ();
 sg13g2_fill_1 FILLER_9_87 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_decap_4 FILLER_9_286 ();
 sg13g2_fill_1 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_295 ();
 sg13g2_fill_1 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_304 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_1 FILLER_9_316 ();
 sg13g2_fill_1 FILLER_9_385 ();
 sg13g2_fill_2 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_fill_1 FILLER_9_416 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_85 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_fill_2 FILLER_10_183 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_224 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_decap_4 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_fill_2 FILLER_10_320 ();
 sg13g2_fill_1 FILLER_10_330 ();
 sg13g2_fill_1 FILLER_10_341 ();
 sg13g2_fill_1 FILLER_10_347 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_decap_8 FILLER_11_48 ();
 sg13g2_fill_2 FILLER_11_55 ();
 sg13g2_fill_2 FILLER_11_103 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_fill_2 FILLER_11_230 ();
 sg13g2_fill_1 FILLER_11_232 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_306 ();
 sg13g2_fill_2 FILLER_11_337 ();
 sg13g2_fill_1 FILLER_11_344 ();
 sg13g2_fill_1 FILLER_11_394 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_55 ();
 sg13g2_fill_2 FILLER_12_74 ();
 sg13g2_fill_1 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_186 ();
 sg13g2_fill_1 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_fill_1 FILLER_12_274 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_fill_2 FILLER_12_324 ();
 sg13g2_fill_2 FILLER_12_374 ();
 sg13g2_fill_2 FILLER_12_410 ();
 sg13g2_fill_1 FILLER_12_421 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_14 ();
 sg13g2_fill_2 FILLER_13_24 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_decap_4 FILLER_13_102 ();
 sg13g2_fill_1 FILLER_13_110 ();
 sg13g2_decap_4 FILLER_13_114 ();
 sg13g2_decap_8 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_239 ();
 sg13g2_fill_1 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_305 ();
 sg13g2_fill_2 FILLER_13_384 ();
 sg13g2_fill_2 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_14_26 ();
 sg13g2_fill_2 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_95 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_124 ();
 sg13g2_fill_1 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_211 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_fill_1 FILLER_14_226 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_2 FILLER_14_340 ();
 sg13g2_fill_1 FILLER_14_369 ();
 sg13g2_fill_1 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_12 ();
 sg13g2_fill_1 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_fill_1 FILLER_15_69 ();
 sg13g2_fill_2 FILLER_15_75 ();
 sg13g2_fill_2 FILLER_15_85 ();
 sg13g2_fill_1 FILLER_15_87 ();
 sg13g2_fill_1 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_273 ();
 sg13g2_fill_1 FILLER_15_415 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_1 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_fill_2 FILLER_16_22 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_101 ();
 sg13g2_decap_8 FILLER_16_132 ();
 sg13g2_decap_4 FILLER_16_139 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_190 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_259 ();
 sg13g2_fill_2 FILLER_16_284 ();
 sg13g2_fill_2 FILLER_16_312 ();
 sg13g2_fill_1 FILLER_16_318 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_16_423 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_2 FILLER_17_10 ();
 sg13g2_fill_2 FILLER_17_23 ();
 sg13g2_fill_2 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_99 ();
 sg13g2_fill_2 FILLER_17_114 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_196 ();
 sg13g2_fill_2 FILLER_17_202 ();
 sg13g2_fill_1 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_fill_1 FILLER_17_397 ();
 sg13g2_fill_2 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_18_39 ();
 sg13g2_fill_2 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_70 ();
 sg13g2_fill_1 FILLER_18_72 ();
 sg13g2_fill_2 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_96 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_1 FILLER_18_125 ();
 sg13g2_fill_2 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_decap_4 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_198 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_339 ();
 sg13g2_fill_2 FILLER_18_345 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_2 FILLER_18_409 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_13 ();
 sg13g2_fill_2 FILLER_19_30 ();
 sg13g2_fill_2 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_2 FILLER_19_170 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_308 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_373 ();
 sg13g2_fill_1 FILLER_19_395 ();
 sg13g2_fill_2 FILLER_19_410 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_1 FILLER_20_247 ();
 sg13g2_fill_1 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_317 ();
 sg13g2_fill_1 FILLER_20_358 ();
 sg13g2_fill_2 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_379 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_6 ();
 sg13g2_fill_2 FILLER_21_20 ();
 sg13g2_fill_1 FILLER_21_22 ();
 sg13g2_fill_1 FILLER_21_40 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_71 ();
 sg13g2_fill_1 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_87 ();
 sg13g2_fill_2 FILLER_21_97 ();
 sg13g2_fill_2 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_108 ();
 sg13g2_fill_2 FILLER_21_148 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_236 ();
 sg13g2_decap_4 FILLER_21_242 ();
 sg13g2_decap_4 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_255 ();
 sg13g2_fill_1 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_405 ();
 sg13g2_fill_1 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_58 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_fill_2 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_165 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_176 ();
 sg13g2_fill_1 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_229 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_fill_1 FILLER_22_235 ();
 sg13g2_fill_1 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_396 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_22 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_72 ();
 sg13g2_fill_1 FILLER_23_74 ();
 sg13g2_fill_1 FILLER_23_79 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_127 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_246 ();
 sg13g2_fill_1 FILLER_23_248 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_412 ();
 sg13g2_fill_1 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_49 ();
 sg13g2_fill_1 FILLER_24_61 ();
 sg13g2_fill_2 FILLER_24_94 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_135 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_24_377 ();
 sg13g2_fill_1 FILLER_24_423 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_10 ();
 sg13g2_fill_1 FILLER_25_12 ();
 sg13g2_fill_1 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_1 FILLER_25_39 ();
 sg13g2_fill_1 FILLER_25_45 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_fill_1 FILLER_25_64 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_decap_4 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_218 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_229 ();
 sg13g2_decap_4 FILLER_25_238 ();
 sg13g2_fill_2 FILLER_25_242 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_286 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_2 FILLER_25_313 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_38 ();
 sg13g2_decap_8 FILLER_26_48 ();
 sg13g2_fill_1 FILLER_26_55 ();
 sg13g2_fill_1 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_146 ();
 sg13g2_fill_2 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_217 ();
 sg13g2_fill_1 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_241 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_1 FILLER_26_377 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_26_422 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_fill_1 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_53 ();
 sg13g2_fill_1 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_66 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_192 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_115 ();
 sg13g2_fill_1 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_217 ();
 sg13g2_decap_4 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_decap_8 FILLER_28_240 ();
 sg13g2_fill_1 FILLER_28_251 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_267 ();
 sg13g2_decap_4 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_decap_4 FILLER_29_26 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_fill_1 FILLER_29_87 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_114 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_135 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_1 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_fill_2 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_373 ();
 sg13g2_fill_1 FILLER_29_378 ();
 sg13g2_fill_1 FILLER_29_384 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_98 ();
 sg13g2_fill_1 FILLER_30_108 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_1 FILLER_30_178 ();
 sg13g2_fill_2 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_229 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_241 ();
 sg13g2_fill_1 FILLER_30_243 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_292 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_341 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_48 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_151 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_2 FILLER_31_251 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_402 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_50 ();
 sg13g2_fill_1 FILLER_32_97 ();
 sg13g2_fill_1 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_decap_4 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_360 ();
 sg13g2_fill_2 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_2 FILLER_32_421 ();
 sg13g2_fill_2 FILLER_32_428 ();
 sg13g2_fill_1 FILLER_33_17 ();
 sg13g2_fill_1 FILLER_33_70 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_1 FILLER_33_81 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_103 ();
 sg13g2_fill_2 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_fill_1 FILLER_33_198 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_2 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_390 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_fill_1 FILLER_34_39 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_decap_8 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_85 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_114 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_2 FILLER_34_196 ();
 sg13g2_fill_1 FILLER_34_198 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_256 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_412 ();
 sg13g2_decap_4 FILLER_34_421 ();
 sg13g2_fill_1 FILLER_34_425 ();
 sg13g2_fill_1 FILLER_35_34 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_2 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_51 ();
 sg13g2_fill_2 FILLER_36_94 ();
 sg13g2_fill_1 FILLER_36_96 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_153 ();
 sg13g2_fill_1 FILLER_36_175 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_2 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_325 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_fill_2 FILLER_36_372 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_37_31 ();
 sg13g2_fill_2 FILLER_37_88 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_182 ();
 sg13g2_fill_2 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_fill_1 FILLER_37_220 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_1 FILLER_37_357 ();
 sg13g2_fill_2 FILLER_37_366 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_fill_1 FILLER_38_19 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_64 ();
 sg13g2_decap_4 FILLER_38_91 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_fill_1 FILLER_38_145 ();
 sg13g2_fill_1 FILLER_38_162 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_2 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_383 ();
 sg13g2_fill_1 FILLER_38_394 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_15 ();
 sg13g2_fill_1 FILLER_39_28 ();
 sg13g2_fill_1 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_43 ();
 sg13g2_fill_2 FILLER_39_83 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_230 ();
 sg13g2_fill_1 FILLER_39_257 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_2 FILLER_39_269 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_358 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_1 FILLER_39_373 ();
 sg13g2_fill_2 FILLER_39_378 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_409 ();
 sg13g2_decap_4 FILLER_39_423 ();
 sg13g2_fill_2 FILLER_40_26 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_60 ();
 sg13g2_fill_1 FILLER_40_123 ();
 sg13g2_decap_4 FILLER_40_149 ();
 sg13g2_fill_1 FILLER_40_153 ();
 sg13g2_fill_2 FILLER_40_165 ();
 sg13g2_fill_1 FILLER_40_167 ();
 sg13g2_fill_1 FILLER_40_172 ();
 sg13g2_fill_1 FILLER_40_177 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_fill_1 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_190 ();
 sg13g2_fill_1 FILLER_40_195 ();
 sg13g2_fill_2 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_228 ();
 sg13g2_decap_8 FILLER_40_244 ();
 sg13g2_fill_2 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_258 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_273 ();
 sg13g2_fill_1 FILLER_40_278 ();
 sg13g2_fill_2 FILLER_40_284 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_fill_1 FILLER_40_308 ();
 sg13g2_fill_1 FILLER_40_320 ();
 sg13g2_fill_2 FILLER_40_325 ();
 sg13g2_fill_2 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_fill_2 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_fill_1 FILLER_41_82 ();
 sg13g2_decap_8 FILLER_41_92 ();
 sg13g2_decap_4 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_decap_4 FILLER_41_112 ();
 sg13g2_fill_1 FILLER_41_127 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_144 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_168 ();
 sg13g2_fill_1 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_181 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_245 ();
 sg13g2_fill_2 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_264 ();
 sg13g2_fill_2 FILLER_41_287 ();
 sg13g2_fill_1 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_307 ();
 sg13g2_fill_1 FILLER_41_309 ();
 sg13g2_fill_2 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_fill_1 FILLER_41_335 ();
 sg13g2_fill_2 FILLER_41_340 ();
 sg13g2_fill_2 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_2 FILLER_42_19 ();
 sg13g2_fill_1 FILLER_42_26 ();
 sg13g2_fill_1 FILLER_42_31 ();
 sg13g2_fill_1 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_52 ();
 sg13g2_decap_4 FILLER_42_58 ();
 sg13g2_decap_4 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_fill_1 FILLER_42_85 ();
 sg13g2_decap_4 FILLER_42_91 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_147 ();
 sg13g2_fill_2 FILLER_42_157 ();
 sg13g2_fill_1 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_178 ();
 sg13g2_decap_8 FILLER_42_212 ();
 sg13g2_fill_2 FILLER_42_219 ();
 sg13g2_fill_1 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_1 FILLER_42_281 ();
 sg13g2_fill_1 FILLER_42_372 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_2 FILLER_43_59 ();
 sg13g2_fill_1 FILLER_43_91 ();
 sg13g2_fill_2 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_fill_2 FILLER_43_146 ();
 sg13g2_fill_1 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_159 ();
 sg13g2_fill_2 FILLER_43_181 ();
 sg13g2_fill_1 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_204 ();
 sg13g2_decap_8 FILLER_43_239 ();
 sg13g2_fill_2 FILLER_43_246 ();
 sg13g2_fill_2 FILLER_43_269 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_fill_1 FILLER_43_288 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_324 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_decap_8 FILLER_43_335 ();
 sg13g2_fill_2 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_356 ();
 sg13g2_decap_4 FILLER_43_362 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_44_5 ();
 sg13g2_fill_1 FILLER_44_11 ();
 sg13g2_fill_2 FILLER_44_34 ();
 sg13g2_fill_2 FILLER_44_50 ();
 sg13g2_fill_1 FILLER_44_137 ();
 sg13g2_fill_1 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_159 ();
 sg13g2_fill_1 FILLER_44_164 ();
 sg13g2_fill_1 FILLER_44_179 ();
 sg13g2_fill_1 FILLER_44_188 ();
 sg13g2_fill_2 FILLER_44_193 ();
 sg13g2_fill_1 FILLER_44_202 ();
 sg13g2_fill_1 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_269 ();
 sg13g2_fill_1 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_280 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_fill_2 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_317 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_369 ();
 sg13g2_fill_1 FILLER_44_406 ();
 sg13g2_fill_2 FILLER_44_415 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_2 FILLER_45_15 ();
 sg13g2_fill_1 FILLER_45_21 ();
 sg13g2_fill_1 FILLER_45_26 ();
 sg13g2_fill_1 FILLER_45_37 ();
 sg13g2_fill_2 FILLER_45_46 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_fill_1 FILLER_45_112 ();
 sg13g2_fill_1 FILLER_45_144 ();
 sg13g2_fill_1 FILLER_45_161 ();
 sg13g2_fill_1 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_172 ();
 sg13g2_fill_1 FILLER_45_186 ();
 sg13g2_fill_2 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_218 ();
 sg13g2_fill_1 FILLER_45_237 ();
 sg13g2_fill_1 FILLER_45_245 ();
 sg13g2_fill_1 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_263 ();
 sg13g2_fill_1 FILLER_45_288 ();
 sg13g2_fill_1 FILLER_45_293 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_decap_4 FILLER_45_345 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_1 FILLER_45_388 ();
 sg13g2_fill_1 FILLER_45_398 ();
 sg13g2_fill_1 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_79 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_2 FILLER_46_86 ();
 sg13g2_fill_1 FILLER_46_88 ();
 sg13g2_decap_4 FILLER_46_94 ();
 sg13g2_fill_1 FILLER_46_98 ();
 sg13g2_fill_2 FILLER_46_105 ();
 sg13g2_decap_4 FILLER_46_110 ();
 sg13g2_fill_2 FILLER_46_119 ();
 sg13g2_decap_4 FILLER_46_125 ();
 sg13g2_fill_2 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_201 ();
 sg13g2_decap_4 FILLER_46_205 ();
 sg13g2_fill_2 FILLER_46_209 ();
 sg13g2_decap_4 FILLER_46_219 ();
 sg13g2_decap_8 FILLER_46_233 ();
 sg13g2_decap_4 FILLER_46_240 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_fill_2 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_306 ();
 sg13g2_fill_2 FILLER_46_312 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_fill_1 FILLER_46_327 ();
 sg13g2_fill_1 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_359 ();
 sg13g2_fill_1 FILLER_46_365 ();
 sg13g2_fill_2 FILLER_47_4 ();
 sg13g2_fill_1 FILLER_47_37 ();
 sg13g2_fill_1 FILLER_47_43 ();
 sg13g2_fill_1 FILLER_47_50 ();
 sg13g2_fill_1 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_127 ();
 sg13g2_fill_1 FILLER_47_134 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_146 ();
 sg13g2_fill_1 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_187 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_fill_2 FILLER_47_230 ();
 sg13g2_fill_1 FILLER_47_265 ();
 sg13g2_decap_4 FILLER_47_275 ();
 sg13g2_fill_2 FILLER_47_279 ();
 sg13g2_decap_8 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_293 ();
 sg13g2_fill_2 FILLER_47_303 ();
 sg13g2_fill_1 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_fill_1 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_355 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_fill_2 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_13 ();
 sg13g2_fill_1 FILLER_48_15 ();
 sg13g2_fill_2 FILLER_48_20 ();
 sg13g2_fill_1 FILLER_48_22 ();
 sg13g2_decap_4 FILLER_48_27 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_1 FILLER_48_52 ();
 sg13g2_fill_2 FILLER_48_80 ();
 sg13g2_fill_1 FILLER_48_82 ();
 sg13g2_fill_1 FILLER_48_95 ();
 sg13g2_fill_2 FILLER_48_100 ();
 sg13g2_fill_2 FILLER_48_136 ();
 sg13g2_fill_1 FILLER_48_172 ();
 sg13g2_fill_1 FILLER_48_181 ();
 sg13g2_fill_1 FILLER_48_186 ();
 sg13g2_decap_4 FILLER_48_211 ();
 sg13g2_fill_1 FILLER_48_223 ();
 sg13g2_decap_8 FILLER_48_232 ();
 sg13g2_decap_4 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_243 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_1 FILLER_48_252 ();
 sg13g2_fill_2 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_259 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_295 ();
 sg13g2_fill_2 FILLER_48_304 ();
 sg13g2_decap_4 FILLER_48_341 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_fill_1 FILLER_48_355 ();
 sg13g2_fill_1 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_27 ();
 sg13g2_fill_1 FILLER_49_33 ();
 sg13g2_fill_2 FILLER_49_39 ();
 sg13g2_fill_2 FILLER_49_61 ();
 sg13g2_fill_2 FILLER_49_85 ();
 sg13g2_fill_1 FILLER_49_91 ();
 sg13g2_fill_1 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_1 FILLER_49_185 ();
 sg13g2_fill_2 FILLER_49_194 ();
 sg13g2_fill_2 FILLER_49_208 ();
 sg13g2_fill_1 FILLER_49_218 ();
 sg13g2_fill_1 FILLER_49_227 ();
 sg13g2_decap_4 FILLER_49_232 ();
 sg13g2_fill_2 FILLER_49_236 ();
 sg13g2_fill_1 FILLER_49_250 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_333 ();
 sg13g2_fill_1 FILLER_49_335 ();
 sg13g2_fill_2 FILLER_49_340 ();
 sg13g2_fill_1 FILLER_49_347 ();
 sg13g2_fill_1 FILLER_49_352 ();
 sg13g2_fill_1 FILLER_49_358 ();
 sg13g2_fill_1 FILLER_49_366 ();
 sg13g2_fill_1 FILLER_49_375 ();
 sg13g2_fill_1 FILLER_49_391 ();
 sg13g2_fill_1 FILLER_49_421 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_50_57 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_fill_2 FILLER_50_222 ();
 sg13g2_fill_2 FILLER_50_252 ();
 sg13g2_fill_2 FILLER_50_267 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_fill_2 FILLER_50_313 ();
 sg13g2_fill_2 FILLER_50_331 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_fill_1 FILLER_50_361 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_50_421 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_fill_2 FILLER_51_34 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_51 ();
 sg13g2_fill_1 FILLER_51_61 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_85 ();
 sg13g2_fill_2 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_131 ();
 sg13g2_fill_1 FILLER_51_158 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_fill_2 FILLER_51_195 ();
 sg13g2_fill_2 FILLER_51_229 ();
 sg13g2_fill_2 FILLER_51_235 ();
 sg13g2_fill_1 FILLER_51_241 ();
 sg13g2_fill_2 FILLER_51_254 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_283 ();
 sg13g2_fill_1 FILLER_51_293 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_313 ();
 sg13g2_fill_1 FILLER_51_318 ();
 sg13g2_fill_2 FILLER_51_324 ();
 sg13g2_fill_1 FILLER_51_326 ();
 sg13g2_fill_1 FILLER_51_355 ();
 sg13g2_fill_1 FILLER_51_360 ();
 sg13g2_fill_1 FILLER_51_371 ();
 sg13g2_fill_2 FILLER_51_383 ();
 sg13g2_fill_1 FILLER_51_389 ();
 sg13g2_fill_1 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_52_22 ();
 sg13g2_fill_2 FILLER_52_34 ();
 sg13g2_fill_1 FILLER_52_81 ();
 sg13g2_fill_1 FILLER_52_96 ();
 sg13g2_fill_2 FILLER_52_102 ();
 sg13g2_fill_1 FILLER_52_151 ();
 sg13g2_fill_1 FILLER_52_156 ();
 sg13g2_fill_1 FILLER_52_186 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_fill_1 FILLER_52_215 ();
 sg13g2_decap_8 FILLER_52_233 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_fill_1 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_260 ();
 sg13g2_fill_2 FILLER_52_269 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_fill_1 FILLER_52_327 ();
 sg13g2_fill_1 FILLER_52_338 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_fill_1 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_365 ();
 sg13g2_fill_1 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_39 ();
 sg13g2_fill_1 FILLER_53_65 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_fill_1 FILLER_53_75 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_fill_1 FILLER_53_210 ();
 sg13g2_fill_2 FILLER_53_216 ();
 sg13g2_decap_4 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_262 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_272 ();
 sg13g2_fill_1 FILLER_53_281 ();
 sg13g2_fill_2 FILLER_53_290 ();
 sg13g2_fill_2 FILLER_53_311 ();
 sg13g2_fill_1 FILLER_53_313 ();
 sg13g2_decap_4 FILLER_53_322 ();
 sg13g2_fill_2 FILLER_53_326 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_2 FILLER_53_359 ();
 sg13g2_decap_4 FILLER_53_366 ();
 sg13g2_fill_1 FILLER_53_370 ();
 sg13g2_decap_4 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_131 ();
 sg13g2_fill_1 FILLER_54_224 ();
 sg13g2_fill_2 FILLER_54_229 ();
 sg13g2_fill_1 FILLER_54_231 ();
 sg13g2_fill_2 FILLER_54_240 ();
 sg13g2_fill_1 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_282 ();
 sg13g2_fill_1 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_316 ();
 sg13g2_fill_2 FILLER_54_336 ();
 sg13g2_fill_1 FILLER_54_342 ();
 sg13g2_fill_1 FILLER_54_351 ();
 sg13g2_decap_4 FILLER_54_362 ();
 sg13g2_fill_1 FILLER_54_403 ();
 sg13g2_fill_1 FILLER_54_412 ();
 sg13g2_fill_2 FILLER_54_417 ();
 sg13g2_fill_2 FILLER_54_427 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_2 ();
 sg13g2_fill_2 FILLER_55_11 ();
 sg13g2_fill_1 FILLER_55_13 ();
 sg13g2_fill_1 FILLER_55_90 ();
 sg13g2_fill_1 FILLER_55_96 ();
 sg13g2_fill_1 FILLER_55_128 ();
 sg13g2_decap_4 FILLER_55_199 ();
 sg13g2_fill_2 FILLER_55_203 ();
 sg13g2_fill_2 FILLER_55_208 ();
 sg13g2_decap_4 FILLER_55_214 ();
 sg13g2_fill_1 FILLER_55_222 ();
 sg13g2_decap_4 FILLER_55_229 ();
 sg13g2_fill_1 FILLER_55_258 ();
 sg13g2_fill_1 FILLER_55_288 ();
 sg13g2_fill_1 FILLER_55_293 ();
 sg13g2_fill_1 FILLER_55_299 ();
 sg13g2_fill_1 FILLER_55_312 ();
 sg13g2_fill_1 FILLER_55_319 ();
 sg13g2_decap_8 FILLER_55_335 ();
 sg13g2_fill_2 FILLER_55_342 ();
 sg13g2_decap_4 FILLER_55_357 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_fill_2 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_fill_1 FILLER_56_47 ();
 sg13g2_fill_2 FILLER_56_86 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_fill_1 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_214 ();
 sg13g2_fill_2 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_317 ();
 sg13g2_fill_1 FILLER_56_319 ();
 sg13g2_fill_2 FILLER_56_342 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_fill_2 FILLER_56_400 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_fill_1 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_fill_1 FILLER_57_64 ();
 sg13g2_fill_2 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_126 ();
 sg13g2_fill_1 FILLER_57_197 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_211 ();
 sg13g2_decap_4 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_312 ();
 sg13g2_fill_1 FILLER_57_314 ();
 sg13g2_decap_4 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_370 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_fill_1 FILLER_58_12 ();
 sg13g2_fill_1 FILLER_58_64 ();
 sg13g2_fill_2 FILLER_58_73 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_fill_1 FILLER_58_193 ();
 sg13g2_fill_1 FILLER_58_205 ();
 sg13g2_fill_1 FILLER_58_214 ();
 sg13g2_fill_1 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_224 ();
 sg13g2_fill_2 FILLER_58_230 ();
 sg13g2_fill_2 FILLER_58_237 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_2 FILLER_58_275 ();
 sg13g2_fill_2 FILLER_58_302 ();
 sg13g2_fill_1 FILLER_58_304 ();
 sg13g2_fill_2 FILLER_58_326 ();
 sg13g2_fill_1 FILLER_58_332 ();
 sg13g2_fill_2 FILLER_58_341 ();
 sg13g2_decap_4 FILLER_58_348 ();
 sg13g2_fill_2 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_fill_2 FILLER_58_377 ();
 sg13g2_fill_1 FILLER_58_389 ();
 sg13g2_fill_1 FILLER_58_393 ();
 sg13g2_fill_1 FILLER_58_412 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_59_35 ();
 sg13g2_fill_2 FILLER_59_48 ();
 sg13g2_fill_2 FILLER_59_65 ();
 sg13g2_fill_1 FILLER_59_72 ();
 sg13g2_fill_2 FILLER_59_123 ();
 sg13g2_fill_1 FILLER_59_125 ();
 sg13g2_fill_2 FILLER_59_143 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_fill_1 FILLER_59_213 ();
 sg13g2_fill_2 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_229 ();
 sg13g2_fill_2 FILLER_59_235 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_246 ();
 sg13g2_fill_2 FILLER_59_267 ();
 sg13g2_decap_8 FILLER_59_282 ();
 sg13g2_decap_8 FILLER_59_289 ();
 sg13g2_decap_8 FILLER_59_296 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_fill_1 FILLER_59_315 ();
 sg13g2_fill_1 FILLER_59_321 ();
 sg13g2_fill_1 FILLER_59_326 ();
 sg13g2_fill_1 FILLER_59_335 ();
 sg13g2_fill_2 FILLER_59_340 ();
 sg13g2_fill_2 FILLER_59_350 ();
 sg13g2_fill_1 FILLER_59_352 ();
 sg13g2_fill_1 FILLER_59_359 ();
 sg13g2_fill_2 FILLER_59_363 ();
 sg13g2_fill_1 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_422 ();
 sg13g2_fill_2 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_fill_2 FILLER_60_23 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_156 ();
 sg13g2_fill_1 FILLER_60_171 ();
 sg13g2_fill_2 FILLER_60_181 ();
 sg13g2_fill_1 FILLER_60_207 ();
 sg13g2_fill_2 FILLER_60_221 ();
 sg13g2_fill_1 FILLER_60_233 ();
 sg13g2_fill_2 FILLER_60_238 ();
 sg13g2_fill_1 FILLER_60_240 ();
 sg13g2_fill_1 FILLER_60_248 ();
 sg13g2_decap_4 FILLER_60_271 ();
 sg13g2_fill_2 FILLER_60_322 ();
 sg13g2_fill_1 FILLER_60_324 ();
 sg13g2_decap_4 FILLER_60_329 ();
 sg13g2_fill_2 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_1 FILLER_60_350 ();
 sg13g2_fill_1 FILLER_60_355 ();
 sg13g2_fill_2 FILLER_60_361 ();
 sg13g2_fill_1 FILLER_60_367 ();
 sg13g2_fill_2 FILLER_60_376 ();
 sg13g2_decap_4 FILLER_60_382 ();
 sg13g2_fill_1 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_60_419 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_fill_2 FILLER_61_26 ();
 sg13g2_fill_2 FILLER_61_85 ();
 sg13g2_fill_2 FILLER_61_104 ();
 sg13g2_fill_2 FILLER_61_135 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_183 ();
 sg13g2_fill_2 FILLER_61_222 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_fill_2 FILLER_61_229 ();
 sg13g2_fill_1 FILLER_61_235 ();
 sg13g2_fill_2 FILLER_61_241 ();
 sg13g2_fill_1 FILLER_61_248 ();
 sg13g2_fill_2 FILLER_61_288 ();
 sg13g2_fill_2 FILLER_61_307 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_fill_1 FILLER_61_318 ();
 sg13g2_fill_1 FILLER_61_324 ();
 sg13g2_fill_1 FILLER_61_331 ();
 sg13g2_fill_2 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_349 ();
 sg13g2_fill_1 FILLER_61_354 ();
 sg13g2_fill_1 FILLER_61_360 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_1 FILLER_61_377 ();
 sg13g2_decap_4 FILLER_61_383 ();
 sg13g2_fill_1 FILLER_61_387 ();
 sg13g2_fill_2 FILLER_61_419 ();
 sg13g2_fill_1 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_62_82 ();
 sg13g2_fill_1 FILLER_62_97 ();
 sg13g2_fill_1 FILLER_62_101 ();
 sg13g2_fill_1 FILLER_62_107 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_fill_2 FILLER_62_138 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_153 ();
 sg13g2_fill_1 FILLER_62_155 ();
 sg13g2_fill_1 FILLER_62_163 ();
 sg13g2_fill_2 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_177 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_1 FILLER_62_188 ();
 sg13g2_fill_1 FILLER_62_202 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_1 FILLER_62_284 ();
 sg13g2_fill_1 FILLER_62_289 ();
 sg13g2_fill_1 FILLER_62_317 ();
 sg13g2_fill_2 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_338 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_346 ();
 sg13g2_fill_2 FILLER_62_355 ();
 sg13g2_fill_1 FILLER_62_357 ();
 sg13g2_fill_2 FILLER_62_402 ();
 sg13g2_fill_1 FILLER_63_30 ();
 sg13g2_fill_2 FILLER_63_70 ();
 sg13g2_fill_1 FILLER_63_133 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_decap_4 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_180 ();
 sg13g2_fill_1 FILLER_63_185 ();
 sg13g2_fill_1 FILLER_63_190 ();
 sg13g2_fill_2 FILLER_63_202 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_1 FILLER_63_215 ();
 sg13g2_fill_1 FILLER_63_221 ();
 sg13g2_fill_1 FILLER_63_227 ();
 sg13g2_decap_4 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_264 ();
 sg13g2_fill_2 FILLER_63_279 ();
 sg13g2_fill_1 FILLER_63_281 ();
 sg13g2_fill_2 FILLER_63_289 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_1 FILLER_63_315 ();
 sg13g2_fill_1 FILLER_63_382 ();
 sg13g2_fill_2 FILLER_63_397 ();
 sg13g2_fill_1 FILLER_64_16 ();
 sg13g2_fill_1 FILLER_64_66 ();
 sg13g2_fill_1 FILLER_64_76 ();
 sg13g2_fill_1 FILLER_64_101 ();
 sg13g2_decap_8 FILLER_64_121 ();
 sg13g2_fill_1 FILLER_64_128 ();
 sg13g2_fill_2 FILLER_64_145 ();
 sg13g2_decap_4 FILLER_64_152 ();
 sg13g2_fill_2 FILLER_64_156 ();
 sg13g2_fill_1 FILLER_64_193 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_fill_1 FILLER_64_203 ();
 sg13g2_fill_2 FILLER_64_225 ();
 sg13g2_fill_1 FILLER_64_232 ();
 sg13g2_fill_1 FILLER_64_238 ();
 sg13g2_fill_1 FILLER_64_255 ();
 sg13g2_fill_2 FILLER_64_267 ();
 sg13g2_fill_1 FILLER_64_281 ();
 sg13g2_fill_2 FILLER_64_309 ();
 sg13g2_fill_2 FILLER_64_316 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_decap_4 FILLER_64_337 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_1 FILLER_64_352 ();
 sg13g2_fill_1 FILLER_64_357 ();
 sg13g2_fill_1 FILLER_64_363 ();
 sg13g2_fill_1 FILLER_64_368 ();
 sg13g2_fill_1 FILLER_64_374 ();
 sg13g2_fill_1 FILLER_64_383 ();
 sg13g2_fill_1 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_fill_1 FILLER_65_60 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_109 ();
 sg13g2_fill_2 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_141 ();
 sg13g2_fill_1 FILLER_65_150 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_fill_2 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_204 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_219 ();
 sg13g2_fill_2 FILLER_65_225 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_2 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_275 ();
 sg13g2_fill_2 FILLER_65_307 ();
 sg13g2_fill_1 FILLER_65_323 ();
 sg13g2_fill_2 FILLER_65_343 ();
 sg13g2_fill_1 FILLER_65_350 ();
 sg13g2_fill_1 FILLER_65_359 ();
 sg13g2_fill_2 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_402 ();
 sg13g2_fill_1 FILLER_66_5 ();
 sg13g2_fill_1 FILLER_66_11 ();
 sg13g2_fill_1 FILLER_66_20 ();
 sg13g2_fill_1 FILLER_66_25 ();
 sg13g2_fill_2 FILLER_66_67 ();
 sg13g2_fill_2 FILLER_66_117 ();
 sg13g2_fill_1 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_150 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_2 FILLER_66_164 ();
 sg13g2_fill_2 FILLER_66_170 ();
 sg13g2_fill_1 FILLER_66_181 ();
 sg13g2_fill_1 FILLER_66_240 ();
 sg13g2_decap_8 FILLER_66_256 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_2 FILLER_66_290 ();
 sg13g2_fill_1 FILLER_66_292 ();
 sg13g2_fill_1 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_decap_4 FILLER_66_309 ();
 sg13g2_fill_1 FILLER_66_321 ();
 sg13g2_fill_1 FILLER_66_334 ();
 sg13g2_fill_2 FILLER_66_346 ();
 sg13g2_fill_1 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_397 ();
 sg13g2_fill_2 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_410 ();
 sg13g2_decap_4 FILLER_66_419 ();
 sg13g2_fill_2 FILLER_66_423 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_fill_1 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_53 ();
 sg13g2_fill_1 FILLER_67_59 ();
 sg13g2_fill_2 FILLER_67_68 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_fill_1 FILLER_67_179 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_decap_4 FILLER_67_194 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_224 ();
 sg13g2_fill_2 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_232 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_fill_1 FILLER_67_259 ();
 sg13g2_decap_4 FILLER_67_278 ();
 sg13g2_decap_4 FILLER_67_306 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_1 FILLER_67_333 ();
 sg13g2_fill_1 FILLER_67_337 ();
 sg13g2_fill_1 FILLER_67_343 ();
 sg13g2_fill_2 FILLER_67_348 ();
 sg13g2_decap_8 FILLER_67_356 ();
 sg13g2_decap_8 FILLER_67_363 ();
 sg13g2_fill_2 FILLER_67_370 ();
 sg13g2_fill_1 FILLER_67_372 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_fill_2 FILLER_67_393 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_67_400 ();
 sg13g2_fill_1 FILLER_67_405 ();
 sg13g2_fill_1 FILLER_67_414 ();
 sg13g2_fill_1 FILLER_67_423 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_26 ();
 sg13g2_fill_1 FILLER_68_52 ();
 sg13g2_fill_2 FILLER_68_61 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_fill_1 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_150 ();
 sg13g2_fill_1 FILLER_68_167 ();
 sg13g2_fill_1 FILLER_68_184 ();
 sg13g2_decap_4 FILLER_68_198 ();
 sg13g2_fill_2 FILLER_68_202 ();
 sg13g2_fill_1 FILLER_68_208 ();
 sg13g2_fill_2 FILLER_68_213 ();
 sg13g2_fill_2 FILLER_68_220 ();
 sg13g2_fill_2 FILLER_68_227 ();
 sg13g2_decap_4 FILLER_68_234 ();
 sg13g2_fill_1 FILLER_68_245 ();
 sg13g2_fill_2 FILLER_68_250 ();
 sg13g2_fill_2 FILLER_68_255 ();
 sg13g2_fill_2 FILLER_68_262 ();
 sg13g2_fill_1 FILLER_68_270 ();
 sg13g2_fill_1 FILLER_68_299 ();
 sg13g2_fill_1 FILLER_68_306 ();
 sg13g2_fill_1 FILLER_68_311 ();
 sg13g2_decap_4 FILLER_68_317 ();
 sg13g2_fill_2 FILLER_68_329 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_fill_2 FILLER_68_356 ();
 sg13g2_fill_1 FILLER_68_358 ();
 sg13g2_fill_2 FILLER_68_376 ();
 sg13g2_fill_2 FILLER_68_386 ();
 sg13g2_fill_2 FILLER_68_409 ();
 sg13g2_decap_8 FILLER_68_423 ();
 sg13g2_fill_1 FILLER_69_46 ();
 sg13g2_fill_1 FILLER_69_97 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_decap_8 FILLER_69_134 ();
 sg13g2_fill_1 FILLER_69_216 ();
 sg13g2_fill_2 FILLER_69_221 ();
 sg13g2_fill_1 FILLER_69_223 ();
 sg13g2_fill_1 FILLER_69_244 ();
 sg13g2_fill_1 FILLER_69_325 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_fill_1 FILLER_69_336 ();
 sg13g2_fill_2 FILLER_69_355 ();
 sg13g2_fill_1 FILLER_69_357 ();
 sg13g2_fill_1 FILLER_69_411 ();
 sg13g2_fill_1 FILLER_70_34 ();
 sg13g2_fill_2 FILLER_70_42 ();
 sg13g2_fill_1 FILLER_70_71 ();
 sg13g2_fill_1 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_102 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_1 FILLER_70_116 ();
 sg13g2_fill_2 FILLER_70_121 ();
 sg13g2_fill_2 FILLER_70_144 ();
 sg13g2_decap_4 FILLER_70_150 ();
 sg13g2_decap_4 FILLER_70_159 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_fill_1 FILLER_70_169 ();
 sg13g2_decap_4 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_224 ();
 sg13g2_fill_1 FILLER_70_231 ();
 sg13g2_fill_1 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_262 ();
 sg13g2_fill_2 FILLER_70_280 ();
 sg13g2_fill_2 FILLER_70_306 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_2 FILLER_70_356 ();
 sg13g2_fill_1 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_367 ();
 sg13g2_fill_1 FILLER_70_374 ();
 sg13g2_fill_1 FILLER_70_380 ();
 sg13g2_fill_2 FILLER_70_409 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_fill_1 FILLER_71_47 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_76 ();
 sg13g2_fill_1 FILLER_71_80 ();
 sg13g2_fill_1 FILLER_71_91 ();
 sg13g2_fill_1 FILLER_71_109 ();
 sg13g2_fill_1 FILLER_71_145 ();
 sg13g2_fill_1 FILLER_71_151 ();
 sg13g2_fill_1 FILLER_71_156 ();
 sg13g2_fill_1 FILLER_71_161 ();
 sg13g2_fill_1 FILLER_71_167 ();
 sg13g2_fill_1 FILLER_71_171 ();
 sg13g2_fill_2 FILLER_71_185 ();
 sg13g2_decap_8 FILLER_71_237 ();
 sg13g2_fill_2 FILLER_71_244 ();
 sg13g2_fill_1 FILLER_71_246 ();
 sg13g2_fill_2 FILLER_71_256 ();
 sg13g2_fill_2 FILLER_71_264 ();
 sg13g2_fill_1 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_283 ();
 sg13g2_fill_1 FILLER_71_315 ();
 sg13g2_fill_1 FILLER_71_320 ();
 sg13g2_fill_1 FILLER_71_329 ();
 sg13g2_fill_1 FILLER_71_334 ();
 sg13g2_fill_1 FILLER_71_343 ();
 sg13g2_fill_1 FILLER_71_357 ();
 sg13g2_decap_4 FILLER_71_366 ();
 sg13g2_fill_1 FILLER_71_381 ();
 sg13g2_fill_1 FILLER_71_386 ();
 sg13g2_fill_1 FILLER_71_391 ();
 sg13g2_fill_1 FILLER_71_397 ();
 sg13g2_fill_1 FILLER_71_415 ();
 sg13g2_fill_1 FILLER_71_424 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_72_18 ();
 sg13g2_fill_1 FILLER_72_68 ();
 sg13g2_fill_1 FILLER_72_113 ();
 sg13g2_fill_2 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_1 FILLER_72_226 ();
 sg13g2_decap_4 FILLER_72_266 ();
 sg13g2_fill_1 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_296 ();
 sg13g2_decap_4 FILLER_72_344 ();
 sg13g2_fill_2 FILLER_72_366 ();
 sg13g2_fill_1 FILLER_72_386 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_fill_2 FILLER_72_417 ();
 sg13g2_fill_1 FILLER_72_419 ();
 sg13g2_decap_4 FILLER_72_424 ();
 sg13g2_fill_2 FILLER_72_428 ();
 sg13g2_fill_2 FILLER_73_29 ();
 sg13g2_fill_2 FILLER_73_134 ();
 sg13g2_fill_2 FILLER_73_155 ();
 sg13g2_fill_1 FILLER_73_162 ();
 sg13g2_fill_1 FILLER_73_180 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_fill_2 FILLER_73_200 ();
 sg13g2_fill_2 FILLER_73_211 ();
 sg13g2_fill_2 FILLER_73_221 ();
 sg13g2_fill_1 FILLER_73_223 ();
 sg13g2_decap_4 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_237 ();
 sg13g2_decap_8 FILLER_73_247 ();
 sg13g2_fill_2 FILLER_73_268 ();
 sg13g2_fill_1 FILLER_73_275 ();
 sg13g2_fill_1 FILLER_73_284 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_1 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_326 ();
 sg13g2_fill_1 FILLER_73_332 ();
 sg13g2_decap_4 FILLER_73_342 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_fill_2 FILLER_73_356 ();
 sg13g2_decap_4 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_366 ();
 sg13g2_fill_2 FILLER_73_380 ();
 sg13g2_fill_1 FILLER_73_387 ();
 sg13g2_fill_2 FILLER_73_392 ();
 sg13g2_decap_4 FILLER_73_424 ();
 sg13g2_fill_2 FILLER_73_428 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_19 ();
 sg13g2_fill_1 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_114 ();
 sg13g2_fill_2 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_168 ();
 sg13g2_fill_2 FILLER_74_175 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_fill_2 FILLER_74_223 ();
 sg13g2_fill_1 FILLER_74_225 ();
 sg13g2_fill_2 FILLER_74_230 ();
 sg13g2_fill_1 FILLER_74_334 ();
 sg13g2_fill_2 FILLER_74_338 ();
 sg13g2_fill_1 FILLER_74_340 ();
 sg13g2_fill_1 FILLER_74_346 ();
 sg13g2_fill_2 FILLER_74_352 ();
 sg13g2_fill_1 FILLER_74_415 ();
 sg13g2_fill_1 FILLER_74_420 ();
 sg13g2_decap_4 FILLER_74_426 ();
 sg13g2_fill_2 FILLER_75_19 ();
 sg13g2_fill_2 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_49 ();
 sg13g2_fill_1 FILLER_75_67 ();
 sg13g2_fill_1 FILLER_75_73 ();
 sg13g2_fill_1 FILLER_75_79 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_93 ();
 sg13g2_fill_1 FILLER_75_138 ();
 sg13g2_fill_1 FILLER_75_144 ();
 sg13g2_fill_1 FILLER_75_150 ();
 sg13g2_fill_2 FILLER_75_179 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_223 ();
 sg13g2_fill_2 FILLER_75_260 ();
 sg13g2_fill_1 FILLER_75_262 ();
 sg13g2_fill_2 FILLER_75_267 ();
 sg13g2_fill_1 FILLER_75_278 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_288 ();
 sg13g2_fill_1 FILLER_75_297 ();
 sg13g2_fill_1 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_307 ();
 sg13g2_fill_1 FILLER_75_313 ();
 sg13g2_fill_1 FILLER_75_320 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_336 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_2 FILLER_75_347 ();
 sg13g2_fill_1 FILLER_75_369 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_2 FILLER_75_394 ();
 sg13g2_fill_1 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_75_424 ();
 sg13g2_fill_1 FILLER_76_76 ();
 sg13g2_fill_2 FILLER_76_82 ();
 sg13g2_fill_1 FILLER_76_88 ();
 sg13g2_fill_1 FILLER_76_140 ();
 sg13g2_fill_2 FILLER_76_145 ();
 sg13g2_fill_1 FILLER_76_177 ();
 sg13g2_fill_1 FILLER_76_181 ();
 sg13g2_fill_1 FILLER_76_189 ();
 sg13g2_fill_1 FILLER_76_203 ();
 sg13g2_fill_2 FILLER_76_213 ();
 sg13g2_fill_1 FILLER_76_220 ();
 sg13g2_fill_1 FILLER_76_225 ();
 sg13g2_fill_2 FILLER_76_231 ();
 sg13g2_fill_1 FILLER_76_238 ();
 sg13g2_fill_1 FILLER_76_248 ();
 sg13g2_fill_2 FILLER_76_278 ();
 sg13g2_fill_2 FILLER_76_288 ();
 sg13g2_fill_1 FILLER_76_295 ();
 sg13g2_fill_1 FILLER_76_304 ();
 sg13g2_fill_1 FILLER_76_331 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_fill_1 FILLER_76_359 ();
 sg13g2_fill_1 FILLER_76_392 ();
 sg13g2_fill_2 FILLER_76_397 ();
 sg13g2_fill_2 FILLER_76_408 ();
 sg13g2_fill_1 FILLER_76_410 ();
 sg13g2_fill_1 FILLER_76_424 ();
 sg13g2_fill_1 FILLER_77_30 ();
 sg13g2_fill_1 FILLER_77_35 ();
 sg13g2_fill_2 FILLER_77_102 ();
 sg13g2_fill_1 FILLER_77_108 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_fill_1 FILLER_77_118 ();
 sg13g2_fill_1 FILLER_77_127 ();
 sg13g2_fill_1 FILLER_77_140 ();
 sg13g2_fill_1 FILLER_77_145 ();
 sg13g2_fill_1 FILLER_77_154 ();
 sg13g2_fill_2 FILLER_77_202 ();
 sg13g2_fill_1 FILLER_77_208 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_298 ();
 sg13g2_fill_2 FILLER_77_304 ();
 sg13g2_fill_1 FILLER_77_338 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_fill_1 FILLER_77_354 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_fill_1 FILLER_77_365 ();
 sg13g2_fill_1 FILLER_77_370 ();
 sg13g2_fill_1 FILLER_77_390 ();
 sg13g2_fill_1 FILLER_77_395 ();
 sg13g2_fill_2 FILLER_77_406 ();
 sg13g2_fill_1 FILLER_77_413 ();
 sg13g2_fill_2 FILLER_78_26 ();
 sg13g2_fill_2 FILLER_78_169 ();
 sg13g2_fill_1 FILLER_78_179 ();
 sg13g2_fill_2 FILLER_78_184 ();
 sg13g2_fill_1 FILLER_78_203 ();
 sg13g2_fill_1 FILLER_78_237 ();
 sg13g2_fill_1 FILLER_78_242 ();
 sg13g2_fill_1 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_253 ();
 sg13g2_fill_2 FILLER_78_263 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_1 FILLER_78_359 ();
 sg13g2_fill_2 FILLER_78_373 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_fill_2 FILLER_79_9 ();
 sg13g2_fill_1 FILLER_79_32 ();
 sg13g2_fill_2 FILLER_79_182 ();
 sg13g2_fill_2 FILLER_79_223 ();
 sg13g2_fill_1 FILLER_79_355 ();
 sg13g2_fill_2 FILLER_79_371 ();
 sg13g2_fill_2 FILLER_79_411 ();
 sg13g2_fill_1 FILLER_79_413 ();
 sg13g2_fill_2 FILLER_79_422 ();
 sg13g2_fill_1 FILLER_79_424 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_fill_2 FILLER_80_94 ();
 sg13g2_fill_1 FILLER_80_112 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_fill_2 FILLER_80_259 ();
 sg13g2_fill_1 FILLER_80_265 ();
 sg13g2_fill_1 FILLER_80_271 ();
 sg13g2_fill_1 FILLER_80_276 ();
 sg13g2_fill_1 FILLER_80_338 ();
 sg13g2_fill_2 FILLER_80_352 ();
 sg13g2_fill_1 FILLER_80_365 ();
 sg13g2_fill_2 FILLER_80_370 ();
 sg13g2_fill_2 FILLER_80_376 ();
 sg13g2_fill_1 FILLER_80_378 ();
 sg13g2_fill_1 FILLER_80_388 ();
 sg13g2_fill_2 FILLER_80_397 ();
 sg13g2_fill_1 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_422 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
