module tt_um_meiniKi_ttihp_fazyrv_exotiny (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire _4704_;
 wire _4705_;
 wire _4706_;
 wire _4707_;
 wire _4708_;
 wire _4709_;
 wire _4710_;
 wire _4711_;
 wire _4712_;
 wire _4713_;
 wire _4714_;
 wire _4715_;
 wire _4716_;
 wire _4717_;
 wire _4718_;
 wire _4719_;
 wire _4720_;
 wire _4721_;
 wire _4722_;
 wire _4723_;
 wire _4724_;
 wire _4725_;
 wire _4726_;
 wire _4727_;
 wire _4728_;
 wire _4729_;
 wire _4730_;
 wire _4731_;
 wire _4732_;
 wire _4733_;
 wire _4734_;
 wire _4735_;
 wire _4736_;
 wire _4737_;
 wire _4738_;
 wire _4739_;
 wire _4740_;
 wire _4741_;
 wire _4742_;
 wire _4743_;
 wire _4744_;
 wire _4745_;
 wire _4746_;
 wire _4747_;
 wire _4748_;
 wire _4749_;
 wire _4750_;
 wire _4751_;
 wire _4752_;
 wire _4753_;
 wire _4754_;
 wire _4755_;
 wire _4756_;
 wire _4757_;
 wire _4758_;
 wire _4759_;
 wire _4760_;
 wire _4761_;
 wire _4762_;
 wire _4763_;
 wire _4764_;
 wire _4765_;
 wire _4766_;
 wire _4767_;
 wire _4768_;
 wire _4769_;
 wire _4770_;
 wire _4771_;
 wire _4772_;
 wire _4773_;
 wire _4774_;
 wire _4775_;
 wire _4776_;
 wire _4777_;
 wire _4778_;
 wire _4779_;
 wire _4780_;
 wire _4781_;
 wire _4782_;
 wire _4783_;
 wire _4784_;
 wire _4785_;
 wire _4786_;
 wire _4787_;
 wire _4788_;
 wire _4789_;
 wire _4790_;
 wire _4791_;
 wire _4792_;
 wire _4793_;
 wire _4794_;
 wire _4795_;
 wire _4796_;
 wire _4797_;
 wire _4798_;
 wire _4799_;
 wire _4800_;
 wire _4801_;
 wire _4802_;
 wire _4803_;
 wire _4804_;
 wire _4805_;
 wire _4806_;
 wire _4807_;
 wire _4808_;
 wire _4809_;
 wire _4810_;
 wire _4811_;
 wire _4812_;
 wire _4813_;
 wire _4814_;
 wire _4815_;
 wire _4816_;
 wire _4817_;
 wire _4818_;
 wire _4819_;
 wire _4820_;
 wire _4821_;
 wire _4822_;
 wire _4823_;
 wire _4824_;
 wire _4825_;
 wire _4826_;
 wire _4827_;
 wire _4828_;
 wire _4829_;
 wire _4830_;
 wire _4831_;
 wire _4832_;
 wire _4833_;
 wire _4834_;
 wire _4835_;
 wire _4836_;
 wire _4837_;
 wire _4838_;
 wire _4839_;
 wire _4840_;
 wire _4841_;
 wire _4842_;
 wire _4843_;
 wire _4844_;
 wire _4845_;
 wire _4846_;
 wire _4847_;
 wire _4848_;
 wire _4849_;
 wire _4850_;
 wire _4851_;
 wire _4852_;
 wire _4853_;
 wire _4854_;
 wire _4855_;
 wire _4856_;
 wire _4857_;
 wire _4858_;
 wire _4859_;
 wire _4860_;
 wire _4861_;
 wire _4862_;
 wire _4863_;
 wire _4864_;
 wire _4865_;
 wire _4866_;
 wire _4867_;
 wire _4868_;
 wire _4869_;
 wire _4870_;
 wire _4871_;
 wire _4872_;
 wire _4873_;
 wire _4874_;
 wire _4875_;
 wire _4876_;
 wire _4877_;
 wire _4878_;
 wire _4879_;
 wire _4880_;
 wire _4881_;
 wire _4882_;
 wire _4883_;
 wire _4884_;
 wire _4885_;
 wire _4886_;
 wire _4887_;
 wire _4888_;
 wire _4889_;
 wire _4890_;
 wire _4891_;
 wire _4892_;
 wire _4893_;
 wire _4894_;
 wire _4895_;
 wire _4896_;
 wire _4897_;
 wire _4898_;
 wire _4899_;
 wire _4900_;
 wire _4901_;
 wire _4902_;
 wire _4903_;
 wire _4904_;
 wire _4905_;
 wire _4906_;
 wire _4907_;
 wire _4908_;
 wire _4909_;
 wire _4910_;
 wire _4911_;
 wire _4912_;
 wire _4913_;
 wire _4914_;
 wire _4915_;
 wire _4916_;
 wire _4917_;
 wire _4918_;
 wire _4919_;
 wire _4920_;
 wire _4921_;
 wire _4922_;
 wire _4923_;
 wire _4924_;
 wire _4925_;
 wire _4926_;
 wire _4927_;
 wire _4928_;
 wire _4929_;
 wire _4930_;
 wire _4931_;
 wire _4932_;
 wire _4933_;
 wire _4934_;
 wire _4935_;
 wire _4936_;
 wire _4937_;
 wire _4938_;
 wire _4939_;
 wire _4940_;
 wire _4941_;
 wire _4942_;
 wire _4943_;
 wire _4944_;
 wire _4945_;
 wire _4946_;
 wire _4947_;
 wire _4948_;
 wire _4949_;
 wire _4950_;
 wire _4951_;
 wire _4952_;
 wire _4953_;
 wire _4954_;
 wire _4955_;
 wire _4956_;
 wire _4957_;
 wire _4958_;
 wire _4959_;
 wire _4960_;
 wire _4961_;
 wire _4962_;
 wire _4963_;
 wire _4964_;
 wire _4965_;
 wire _4966_;
 wire _4967_;
 wire _4968_;
 wire _4969_;
 wire _4970_;
 wire _4971_;
 wire _4972_;
 wire _4973_;
 wire _4974_;
 wire _4975_;
 wire _4976_;
 wire _4977_;
 wire _4978_;
 wire _4979_;
 wire _4980_;
 wire _4981_;
 wire _4982_;
 wire _4983_;
 wire _4984_;
 wire _4985_;
 wire _4986_;
 wire _4987_;
 wire _4988_;
 wire _4989_;
 wire _4990_;
 wire _4991_;
 wire _4992_;
 wire _4993_;
 wire _4994_;
 wire _4995_;
 wire _4996_;
 wire _4997_;
 wire _4998_;
 wire _4999_;
 wire _5000_;
 wire _5001_;
 wire _5002_;
 wire _5003_;
 wire _5004_;
 wire _5005_;
 wire _5006_;
 wire _5007_;
 wire _5008_;
 wire _5009_;
 wire _5010_;
 wire _5011_;
 wire _5012_;
 wire _5013_;
 wire _5014_;
 wire _5015_;
 wire _5016_;
 wire _5017_;
 wire _5018_;
 wire _5019_;
 wire _5020_;
 wire _5021_;
 wire _5022_;
 wire _5023_;
 wire _5024_;
 wire _5025_;
 wire _5026_;
 wire _5027_;
 wire _5028_;
 wire _5029_;
 wire _5030_;
 wire _5031_;
 wire _5032_;
 wire _5033_;
 wire _5034_;
 wire _5035_;
 wire _5036_;
 wire _5037_;
 wire _5038_;
 wire _5039_;
 wire _5040_;
 wire _5041_;
 wire _5042_;
 wire _5043_;
 wire _5044_;
 wire _5045_;
 wire _5046_;
 wire _5047_;
 wire _5048_;
 wire _5049_;
 wire _5050_;
 wire _5051_;
 wire _5052_;
 wire _5053_;
 wire _5054_;
 wire _5055_;
 wire _5056_;
 wire _5057_;
 wire _5058_;
 wire _5059_;
 wire _5060_;
 wire _5061_;
 wire _5062_;
 wire _5063_;
 wire _5064_;
 wire _5065_;
 wire _5066_;
 wire _5067_;
 wire _5068_;
 wire _5069_;
 wire _5070_;
 wire _5071_;
 wire _5072_;
 wire _5073_;
 wire _5074_;
 wire _5075_;
 wire _5076_;
 wire _5077_;
 wire _5078_;
 wire _5079_;
 wire _5080_;
 wire _5081_;
 wire _5082_;
 wire _5083_;
 wire _5084_;
 wire _5085_;
 wire _5086_;
 wire _5087_;
 wire _5088_;
 wire _5089_;
 wire _5090_;
 wire _5091_;
 wire _5092_;
 wire _5093_;
 wire _5094_;
 wire _5095_;
 wire _5096_;
 wire _5097_;
 wire _5098_;
 wire _5099_;
 wire _5100_;
 wire _5101_;
 wire _5102_;
 wire _5103_;
 wire _5104_;
 wire _5105_;
 wire _5106_;
 wire _5107_;
 wire _5108_;
 wire _5109_;
 wire _5110_;
 wire _5111_;
 wire _5112_;
 wire _5113_;
 wire _5114_;
 wire _5115_;
 wire _5116_;
 wire _5117_;
 wire _5118_;
 wire _5119_;
 wire _5120_;
 wire _5121_;
 wire _5122_;
 wire _5123_;
 wire _5124_;
 wire _5125_;
 wire _5126_;
 wire _5127_;
 wire _5128_;
 wire _5129_;
 wire _5130_;
 wire _5131_;
 wire _5132_;
 wire _5133_;
 wire _5134_;
 wire _5135_;
 wire _5136_;
 wire _5137_;
 wire _5138_;
 wire _5139_;
 wire _5140_;
 wire _5141_;
 wire _5142_;
 wire _5143_;
 wire _5144_;
 wire _5145_;
 wire _5146_;
 wire _5147_;
 wire _5148_;
 wire _5149_;
 wire _5150_;
 wire _5151_;
 wire _5152_;
 wire _5153_;
 wire _5154_;
 wire _5155_;
 wire _5156_;
 wire _5157_;
 wire _5158_;
 wire _5159_;
 wire _5160_;
 wire _5161_;
 wire _5162_;
 wire _5163_;
 wire _5164_;
 wire _5165_;
 wire _5166_;
 wire _5167_;
 wire _5168_;
 wire _5169_;
 wire _5170_;
 wire _5171_;
 wire _5172_;
 wire _5173_;
 wire _5174_;
 wire _5175_;
 wire _5176_;
 wire _5177_;
 wire _5178_;
 wire _5179_;
 wire _5180_;
 wire _5181_;
 wire _5182_;
 wire _5183_;
 wire _5184_;
 wire _5185_;
 wire _5186_;
 wire _5187_;
 wire _5188_;
 wire _5189_;
 wire _5190_;
 wire _5191_;
 wire _5192_;
 wire _5193_;
 wire _5194_;
 wire _5195_;
 wire _5196_;
 wire _5197_;
 wire _5198_;
 wire _5199_;
 wire _5200_;
 wire _5201_;
 wire _5202_;
 wire _5203_;
 wire _5204_;
 wire _5205_;
 wire _5206_;
 wire _5207_;
 wire _5208_;
 wire _5209_;
 wire _5210_;
 wire _5211_;
 wire _5212_;
 wire _5213_;
 wire _5214_;
 wire _5215_;
 wire _5216_;
 wire _5217_;
 wire _5218_;
 wire _5219_;
 wire _5220_;
 wire _5221_;
 wire _5222_;
 wire _5223_;
 wire _5224_;
 wire _5225_;
 wire _5226_;
 wire _5227_;
 wire _5228_;
 wire _5229_;
 wire _5230_;
 wire _5231_;
 wire _5232_;
 wire _5233_;
 wire _5234_;
 wire _5235_;
 wire _5236_;
 wire _5237_;
 wire _5238_;
 wire _5239_;
 wire _5240_;
 wire _5241_;
 wire _5242_;
 wire _5243_;
 wire _5244_;
 wire _5245_;
 wire _5246_;
 wire _5247_;
 wire _5248_;
 wire _5249_;
 wire _5250_;
 wire _5251_;
 wire _5252_;
 wire _5253_;
 wire _5254_;
 wire _5255_;
 wire _5256_;
 wire _5257_;
 wire _5258_;
 wire _5259_;
 wire _5260_;
 wire _5261_;
 wire _5262_;
 wire _5263_;
 wire _5264_;
 wire _5265_;
 wire _5266_;
 wire _5267_;
 wire _5268_;
 wire _5269_;
 wire _5270_;
 wire _5271_;
 wire _5272_;
 wire _5273_;
 wire _5274_;
 wire _5275_;
 wire _5276_;
 wire _5277_;
 wire _5278_;
 wire _5279_;
 wire _5280_;
 wire _5281_;
 wire _5282_;
 wire _5283_;
 wire _5284_;
 wire _5285_;
 wire _5286_;
 wire _5287_;
 wire _5288_;
 wire _5289_;
 wire _5290_;
 wire _5291_;
 wire _5292_;
 wire _5293_;
 wire _5294_;
 wire _5295_;
 wire _5296_;
 wire _5297_;
 wire _5298_;
 wire _5299_;
 wire _5300_;
 wire _5301_;
 wire _5302_;
 wire _5303_;
 wire _5304_;
 wire _5305_;
 wire _5306_;
 wire _5307_;
 wire _5308_;
 wire _5309_;
 wire _5310_;
 wire _5311_;
 wire _5312_;
 wire _5313_;
 wire _5314_;
 wire _5315_;
 wire _5316_;
 wire _5317_;
 wire _5318_;
 wire _5319_;
 wire _5320_;
 wire _5321_;
 wire _5322_;
 wire _5323_;
 wire _5324_;
 wire _5325_;
 wire _5326_;
 wire _5327_;
 wire _5328_;
 wire _5329_;
 wire _5330_;
 wire _5331_;
 wire _5332_;
 wire _5333_;
 wire _5334_;
 wire _5335_;
 wire _5336_;
 wire _5337_;
 wire _5338_;
 wire _5339_;
 wire _5340_;
 wire _5341_;
 wire _5342_;
 wire _5343_;
 wire _5344_;
 wire _5345_;
 wire _5346_;
 wire _5347_;
 wire _5348_;
 wire _5349_;
 wire _5350_;
 wire _5351_;
 wire _5352_;
 wire _5353_;
 wire _5354_;
 wire _5355_;
 wire _5356_;
 wire _5357_;
 wire _5358_;
 wire _5359_;
 wire _5360_;
 wire _5361_;
 wire _5362_;
 wire _5363_;
 wire _5364_;
 wire _5365_;
 wire _5366_;
 wire _5367_;
 wire _5368_;
 wire _5369_;
 wire _5370_;
 wire _5371_;
 wire _5372_;
 wire _5373_;
 wire _5374_;
 wire _5375_;
 wire _5376_;
 wire _5377_;
 wire _5378_;
 wire _5379_;
 wire _5380_;
 wire _5381_;
 wire _5382_;
 wire _5383_;
 wire _5384_;
 wire _5385_;
 wire _5386_;
 wire _5387_;
 wire _5388_;
 wire _5389_;
 wire _5390_;
 wire _5391_;
 wire _5392_;
 wire _5393_;
 wire _5394_;
 wire net1646;
 wire net340;
 wire cs_ram_n;
 wire cs_rom_n;
 wire \i_exotiny._0000_ ;
 wire \i_exotiny._0001_ ;
 wire \i_exotiny._0002_ ;
 wire \i_exotiny._0003_ ;
 wire \i_exotiny._0004_ ;
 wire \i_exotiny._0005_ ;
 wire \i_exotiny._0006_ ;
 wire \i_exotiny._0007_ ;
 wire \i_exotiny._0008_ ;
 wire \i_exotiny._0009_ ;
 wire \i_exotiny._0010_ ;
 wire \i_exotiny._0011_ ;
 wire \i_exotiny._0012_ ;
 wire \i_exotiny._0013_ ;
 wire \i_exotiny._0014_ ;
 wire \i_exotiny._0015_ ;
 wire \i_exotiny._0062_ ;
 wire \i_exotiny._0063_ ;
 wire \i_exotiny._0064_ ;
 wire \i_exotiny._0065_ ;
 wire \i_exotiny._0066_ ;
 wire \i_exotiny._0067_ ;
 wire \i_exotiny._0068_ ;
 wire \i_exotiny._0069_ ;
 wire \i_exotiny._0070_ ;
 wire \i_exotiny._0071_ ;
 wire \i_exotiny._0072_ ;
 wire \i_exotiny._0073_ ;
 wire \i_exotiny._0074_ ;
 wire \i_exotiny._0075_ ;
 wire \i_exotiny._0076_ ;
 wire \i_exotiny._0077_ ;
 wire \i_exotiny._0078_ ;
 wire \i_exotiny._0079_ ;
 wire \i_exotiny._0080_ ;
 wire \i_exotiny._0081_ ;
 wire \i_exotiny._0082_ ;
 wire \i_exotiny._0083_ ;
 wire \i_exotiny._0084_ ;
 wire \i_exotiny._0085_ ;
 wire \i_exotiny._2356_[0] ;
 wire \i_exotiny._2358_[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_ack ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_shft ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_two ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_msb ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.ex_cmp_tmp ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[11] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[31] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[9] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[12] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[15] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[16] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ld_sext_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_w_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.genblk1[3].i_fazyrv_fadd_x.c_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.imem_stb_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.c_o ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[28] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[7] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[8] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[10] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[16] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[17] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[9] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ;
 wire \i_exotiny.i_wb_qspi_mem.cnt_r[0] ;
 wire \i_exotiny.i_wb_qspi_mem.cnt_r[1] ;
 wire \i_exotiny.i_wb_qspi_mem.cnt_r[2] ;
 wire \i_exotiny.i_wb_qspi_mem.crm_r ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[0] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[1] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[2] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[3] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[4] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[5] ;
 wire \i_exotiny.i_wb_qspi_mem.state_r_reg[6] ;
 wire \i_exotiny.i_wb_qspi_mem.wb_mem_ack_o ;
 wire \i_exotiny.i_wb_regs.spi_auto_cs_o ;
 wire \i_exotiny.i_wb_regs.spi_cpol_o ;
 wire \i_exotiny.i_wb_regs.spi_presc_o[0] ;
 wire \i_exotiny.i_wb_regs.spi_presc_o[1] ;
 wire \i_exotiny.i_wb_regs.spi_presc_o[2] ;
 wire \i_exotiny.i_wb_regs.spi_presc_o[3] ;
 wire \i_exotiny.i_wb_regs.spi_rdy_i ;
 wire \i_exotiny.i_wb_regs.spi_size_o[0] ;
 wire \i_exotiny.i_wb_regs.spi_size_o[1] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[0] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[1] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[2] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[3] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[4] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[5] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[6] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[0] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[1] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[2] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[3] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[4] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[5] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_n[6] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[0] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[1] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[2] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[3] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[4] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[5] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[6] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[0] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[10] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[11] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[12] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[13] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[14] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[15] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[16] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[17] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[18] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[19] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[1] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[20] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[21] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[22] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[23] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[24] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[25] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[26] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[27] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[28] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[29] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[2] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[30] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[31] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[3] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[4] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[5] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[6] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[7] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[8] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[9] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[0] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[10] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[11] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[12] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[13] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[14] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[15] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[16] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[17] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[18] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[19] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[1] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[20] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[21] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[22] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[23] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[24] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[25] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[26] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[27] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[28] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[29] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[2] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[30] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[3] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[4] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[5] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[6] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[7] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[8] ;
 wire \i_exotiny.i_wb_spi.dat_tx_r_reg[9] ;
 wire \i_exotiny.i_wb_spi.state_r_reg[1] ;
 wire clknet_leaf_0_clk;
 wire \i_exotiny.spi_sck_o ;
 wire \i_exotiny.spi_sdo_o ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_buf_1 _5397_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_shft ),
    .X(_1367_));
 sg13g2_buf_1 _5398_ (.A(_1367_),
    .X(_1368_));
 sg13g2_buf_1 _5399_ (.A(net319),
    .X(_1369_));
 sg13g2_buf_2 _5400_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[6] ),
    .X(_1370_));
 sg13g2_buf_8 _5401_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[6] ),
    .X(_1371_));
 sg13g2_inv_1 _5402_ (.Y(_1372_),
    .A(net337));
 sg13g2_buf_2 _5403_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[5] ),
    .X(_1373_));
 sg13g2_buf_1 _5404_ (.A(_0090_),
    .X(_1374_));
 sg13g2_nor2b_1 _5405_ (.A(_1373_),
    .B_N(net336),
    .Y(_1375_));
 sg13g2_buf_8 _5406_ (.A(_1375_),
    .X(_1376_));
 sg13g2_buf_1 _5407_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ld_sext_o ),
    .X(_1377_));
 sg13g2_buf_8 _5408_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_w_o ),
    .X(_1378_));
 sg13g2_o21ai_1 _5409_ (.B1(_1378_),
    .Y(_1379_),
    .A1(net335),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o ));
 sg13g2_buf_1 _5410_ (.A(_1379_),
    .X(_1380_));
 sg13g2_and3_1 _5411_ (.X(_1381_),
    .A(_1372_),
    .B(_1376_),
    .C(_1380_));
 sg13g2_buf_1 _5412_ (.A(_1381_),
    .X(_1382_));
 sg13g2_buf_1 _5413_ (.A(net248),
    .X(_1383_));
 sg13g2_nor2_1 _5414_ (.A(_1370_),
    .B(net230),
    .Y(_1384_));
 sg13g2_nand2_1 _5415_ (.Y(_1385_),
    .A(_1367_),
    .B(_0044_));
 sg13g2_o21ai_1 _5416_ (.B1(_1385_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[0] ),
    .A1(net290),
    .A2(_1384_));
 sg13g2_buf_1 _5417_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[11] ),
    .X(_1386_));
 sg13g2_buf_2 _5418_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ),
    .X(_1387_));
 sg13g2_buf_1 _5419_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.imem_stb_o ),
    .X(_1388_));
 sg13g2_buf_1 _5420_ (.A(_1388_),
    .X(_1389_));
 sg13g2_buf_1 _5421_ (.A(net318),
    .X(_1390_));
 sg13g2_buf_1 _5422_ (.A(\i_exotiny.i_wb_qspi_mem.wb_mem_ack_o ),
    .X(_1391_));
 sg13g2_nand2_1 _5423_ (.Y(_1392_),
    .A(_1390_),
    .B(_1391_));
 sg13g2_buf_2 _5424_ (.A(_1392_),
    .X(_1393_));
 sg13g2_buf_1 _5425_ (.A(_1393_),
    .X(_1394_));
 sg13g2_mux2_1 _5426_ (.A0(_1386_),
    .A1(_1387_),
    .S(net229),
    .X(_1114_));
 sg13g2_mux2_1 _5427_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .S(_1394_),
    .X(_1115_));
 sg13g2_mux2_1 _5428_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .S(net229),
    .X(_1116_));
 sg13g2_mux2_1 _5429_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .S(net229),
    .X(_1117_));
 sg13g2_mux2_1 _5430_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .S(net229),
    .X(_1118_));
 sg13g2_buf_1 _5431_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[0] ),
    .X(_1395_));
 sg13g2_buf_1 _5432_ (.A(_1395_),
    .X(_1396_));
 sg13g2_inv_2 _5433_ (.Y(_1397_),
    .A(net317));
 sg13g2_and2_1 _5434_ (.A(net318),
    .B(_1391_),
    .X(_1398_));
 sg13g2_buf_2 _5435_ (.A(_1398_),
    .X(_1399_));
 sg13g2_buf_1 _5436_ (.A(_1399_),
    .X(_1400_));
 sg13g2_buf_1 _5437_ (.A(_1400_),
    .X(_1401_));
 sg13g2_buf_1 _5438_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[15] ),
    .X(_1402_));
 sg13g2_buf_1 _5439_ (.A(_1399_),
    .X(_1403_));
 sg13g2_nand2_1 _5440_ (.Y(_1404_),
    .A(_1402_),
    .B(net246));
 sg13g2_o21ai_1 _5441_ (.B1(_1404_),
    .Y(_1119_),
    .A1(_1397_),
    .A2(net228));
 sg13g2_buf_1 _5442_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[1] ),
    .X(_1405_));
 sg13g2_buf_1 _5443_ (.A(net334),
    .X(_1406_));
 sg13g2_inv_2 _5444_ (.Y(_1407_),
    .A(net316));
 sg13g2_buf_1 _5445_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[16] ),
    .X(_1408_));
 sg13g2_nand2_1 _5446_ (.Y(_1409_),
    .A(_1408_),
    .B(net246));
 sg13g2_o21ai_1 _5447_ (.B1(_1409_),
    .Y(_1120_),
    .A1(_1407_),
    .A2(net228));
 sg13g2_buf_1 _5448_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[2] ),
    .X(_1410_));
 sg13g2_buf_1 _5449_ (.A(_1410_),
    .X(_1411_));
 sg13g2_buf_1 _5450_ (.A(net315),
    .X(_1412_));
 sg13g2_buf_1 _5451_ (.A(net288),
    .X(_1413_));
 sg13g2_mux2_1 _5452_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ),
    .A1(net265),
    .S(_1394_),
    .X(_1121_));
 sg13g2_buf_2 _5453_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[3] ),
    .X(_1414_));
 sg13g2_buf_1 _5454_ (.A(_1414_),
    .X(_1415_));
 sg13g2_inv_1 _5455_ (.Y(_1416_),
    .A(_1415_));
 sg13g2_nand2_1 _5456_ (.Y(_1417_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ),
    .B(net246));
 sg13g2_o21ai_1 _5457_ (.B1(_1417_),
    .Y(_1122_),
    .A1(net287),
    .A2(net228));
 sg13g2_buf_1 _5458_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[4] ),
    .X(_1418_));
 sg13g2_inv_1 _5459_ (.Y(_1419_),
    .A(_1418_));
 sg13g2_nand2_1 _5460_ (.Y(_1420_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ),
    .B(net246));
 sg13g2_o21ai_1 _5461_ (.B1(_1420_),
    .Y(_1123_),
    .A1(net313),
    .A2(net228));
 sg13g2_buf_1 _5462_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[0] ),
    .X(_1421_));
 sg13g2_buf_1 _5463_ (.A(_1421_),
    .X(_1422_));
 sg13g2_buf_1 _5464_ (.A(net312),
    .X(_1423_));
 sg13g2_buf_1 _5465_ (.A(net286),
    .X(_1424_));
 sg13g2_mux2_1 _5466_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ),
    .A1(net264),
    .S(net229),
    .X(_1124_));
 sg13g2_buf_1 _5467_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[1] ),
    .X(_1425_));
 sg13g2_buf_1 _5468_ (.A(_1425_),
    .X(_1426_));
 sg13g2_buf_1 _5469_ (.A(net311),
    .X(_1427_));
 sg13g2_inv_2 _5470_ (.Y(_1428_),
    .A(net285));
 sg13g2_nand2_1 _5471_ (.Y(_1429_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ),
    .B(net246));
 sg13g2_o21ai_1 _5472_ (.B1(_1429_),
    .Y(_1125_),
    .A1(_1428_),
    .A2(net228));
 sg13g2_buf_2 _5473_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[2] ),
    .X(_1430_));
 sg13g2_inv_1 _5474_ (.Y(_1431_),
    .A(_1430_));
 sg13g2_buf_1 _5475_ (.A(_1431_),
    .X(_1432_));
 sg13g2_nand2_1 _5476_ (.Y(_1433_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ),
    .B(net246));
 sg13g2_o21ai_1 _5477_ (.B1(_1433_),
    .Y(_1126_),
    .A1(_1432_),
    .A2(net228));
 sg13g2_buf_1 _5478_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[3] ),
    .X(_1434_));
 sg13g2_buf_1 _5479_ (.A(_1434_),
    .X(_1435_));
 sg13g2_inv_1 _5480_ (.Y(_1436_),
    .A(net310));
 sg13g2_nand2_1 _5481_ (.Y(_1437_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ),
    .B(_1403_));
 sg13g2_o21ai_1 _5482_ (.B1(_1437_),
    .Y(_1127_),
    .A1(net283),
    .A2(_1401_));
 sg13g2_buf_1 _5483_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[4] ),
    .X(_1438_));
 sg13g2_inv_2 _5484_ (.Y(_1439_),
    .A(net333));
 sg13g2_nand2_1 _5485_ (.Y(_1440_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ),
    .B(_1403_));
 sg13g2_o21ai_1 _5486_ (.B1(_1440_),
    .Y(_1128_),
    .A1(_1439_),
    .A2(_1401_));
 sg13g2_buf_1 _5487_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4] ),
    .X(_1441_));
 sg13g2_inv_2 _5488_ (.Y(_1442_),
    .A(net332));
 sg13g2_buf_2 _5489_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[1] ),
    .X(_1443_));
 sg13g2_buf_2 _5490_ (.A(_0091_),
    .X(_1444_));
 sg13g2_buf_1 _5491_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[2] ),
    .X(_1445_));
 sg13g2_buf_1 _5492_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o ),
    .X(_1446_));
 sg13g2_nand2b_1 _5493_ (.Y(_1447_),
    .B(net331),
    .A_N(net336));
 sg13g2_or2_1 _5494_ (.X(_1448_),
    .B(net337),
    .A(_1378_));
 sg13g2_buf_2 _5495_ (.A(_1448_),
    .X(_1449_));
 sg13g2_nor4_2 _5496_ (.A(_1444_),
    .B(_1445_),
    .C(_1447_),
    .Y(_1450_),
    .D(_1449_));
 sg13g2_buf_8 _5497_ (.A(_1378_),
    .X(_1451_));
 sg13g2_nor2_2 _5498_ (.A(net309),
    .B(net337),
    .Y(_1452_));
 sg13g2_buf_2 _5499_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[3] ),
    .X(_1453_));
 sg13g2_nor2_2 _5500_ (.A(_1373_),
    .B(_1453_),
    .Y(_1454_));
 sg13g2_and2_1 _5501_ (.A(_1452_),
    .B(_1454_),
    .X(_1455_));
 sg13g2_buf_2 _5502_ (.A(_0025_),
    .X(_1456_));
 sg13g2_inv_1 _5503_ (.Y(_1457_),
    .A(_1456_));
 sg13g2_nor2_1 _5504_ (.A(_1457_),
    .B(_1447_),
    .Y(_1458_));
 sg13g2_nand2_1 _5505_ (.Y(_1459_),
    .A(_1455_),
    .B(_1458_));
 sg13g2_nand2b_1 _5506_ (.Y(_1460_),
    .B(_1459_),
    .A_N(_1450_));
 sg13g2_buf_1 _5507_ (.A(_1460_),
    .X(_1461_));
 sg13g2_inv_1 _5508_ (.Y(_1462_),
    .A(_1391_));
 sg13g2_nor2b_1 _5509_ (.A(_1388_),
    .B_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29] ),
    .Y(_1463_));
 sg13g2_a21o_1 _5510_ (.A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ),
    .A1(net318),
    .B1(_1463_),
    .X(_1464_));
 sg13g2_buf_2 _5511_ (.A(_1464_),
    .X(_1465_));
 sg13g2_mux2_1 _5512_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30] ),
    .S(_1388_),
    .X(_1466_));
 sg13g2_buf_1 _5513_ (.A(_1466_),
    .X(_1467_));
 sg13g2_nor2_1 _5514_ (.A(_1465_),
    .B(_1467_),
    .Y(_1468_));
 sg13g2_buf_1 _5515_ (.A(_0089_),
    .X(_1469_));
 sg13g2_a21oi_2 _5516_ (.B1(_1469_),
    .Y(_1470_),
    .A2(_1468_),
    .A1(_1462_));
 sg13g2_nor3_1 _5517_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ),
    .C(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ),
    .Y(_1471_));
 sg13g2_xnor2_1 _5518_ (.Y(_1472_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ),
    .B(_1471_));
 sg13g2_nor2_1 _5519_ (.A(_1385_),
    .B(_1472_),
    .Y(_1473_));
 sg13g2_buf_1 _5520_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ),
    .X(_1474_));
 sg13g2_buf_1 _5521_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .X(_1475_));
 sg13g2_nand2_1 _5522_ (.Y(_1476_),
    .A(_1474_),
    .B(_1475_));
 sg13g2_buf_1 _5523_ (.A(_0029_),
    .X(_1477_));
 sg13g2_inv_1 _5524_ (.Y(_1478_),
    .A(net330));
 sg13g2_nand2b_1 _5525_ (.Y(_1479_),
    .B(_1478_),
    .A_N(_1476_));
 sg13g2_buf_1 _5526_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_two ),
    .X(_1480_));
 sg13g2_buf_1 _5527_ (.A(_1480_),
    .X(_1481_));
 sg13g2_nor2_1 _5528_ (.A(net308),
    .B(_1443_),
    .Y(_1482_));
 sg13g2_buf_2 _5529_ (.A(_1482_),
    .X(_1483_));
 sg13g2_nor2_1 _5530_ (.A(_1479_),
    .B(_1483_),
    .Y(_1484_));
 sg13g2_buf_1 _5531_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_ack ),
    .X(_1485_));
 sg13g2_or2_1 _5532_ (.X(_1486_),
    .B(_1443_),
    .A(net308));
 sg13g2_buf_2 _5533_ (.A(_1486_),
    .X(_1487_));
 sg13g2_nor3_1 _5534_ (.A(net329),
    .B(net319),
    .C(_1487_),
    .Y(_1488_));
 sg13g2_or4_1 _5535_ (.A(_1470_),
    .B(_1473_),
    .C(_1484_),
    .D(_1488_),
    .X(_1489_));
 sg13g2_buf_1 _5536_ (.A(_1489_),
    .X(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_msb ));
 sg13g2_nand2_1 _5537_ (.Y(_1490_),
    .A(net175),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_msb ));
 sg13g2_nand2_1 _5538_ (.Y(_1491_),
    .A(_1443_),
    .B(_1490_));
 sg13g2_buf_1 _5539_ (.A(_1491_),
    .X(_1492_));
 sg13g2_buf_1 _5540_ (.A(_1492_),
    .X(_1493_));
 sg13g2_buf_1 _5541_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[0] ),
    .X(_1494_));
 sg13g2_buf_1 _5542_ (.A(_1494_),
    .X(_1495_));
 sg13g2_buf_1 _5543_ (.A(_1492_),
    .X(_1496_));
 sg13g2_nand2_1 _5544_ (.Y(_1497_),
    .A(net307),
    .B(net74));
 sg13g2_o21ai_1 _5545_ (.B1(_1497_),
    .Y(_1132_),
    .A1(_1442_),
    .A2(net75));
 sg13g2_buf_1 _5546_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5] ),
    .X(_1498_));
 sg13g2_inv_1 _5547_ (.Y(_1499_),
    .A(net328));
 sg13g2_buf_1 _5548_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[1] ),
    .X(_1500_));
 sg13g2_nand2_1 _5549_ (.Y(_1501_),
    .A(net327),
    .B(net74));
 sg13g2_o21ai_1 _5550_ (.B1(_1501_),
    .Y(_1133_),
    .A1(_1499_),
    .A2(net75));
 sg13g2_buf_1 _5551_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[9] ),
    .X(_1502_));
 sg13g2_buf_1 _5552_ (.A(rst_n),
    .X(_1503_));
 sg13g2_buf_1 _5553_ (.A(_1503_),
    .X(_1504_));
 sg13g2_nand2_1 _5554_ (.Y(_1505_),
    .A(net326),
    .B(_1393_));
 sg13g2_buf_1 _5555_ (.A(_1505_),
    .X(_1506_));
 sg13g2_buf_1 _5556_ (.A(_1506_),
    .X(_1507_));
 sg13g2_mux2_1 _5557_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29] ),
    .A1(_1502_),
    .S(net100),
    .X(_1138_));
 sg13g2_buf_2 _5558_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[2] ),
    .X(_1508_));
 sg13g2_mux2_1 _5559_ (.A0(_1445_),
    .A1(_1508_),
    .S(net100),
    .X(_1139_));
 sg13g2_mux2_1 _5560_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ),
    .S(net100),
    .X(_1140_));
 sg13g2_buf_1 _5561_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[3] ),
    .X(_1509_));
 sg13g2_mux2_1 _5562_ (.A0(_1453_),
    .A1(_1509_),
    .S(net100),
    .X(_1141_));
 sg13g2_buf_2 _5563_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[4] ),
    .X(_1510_));
 sg13g2_inv_1 _5564_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_buf_2 _5565_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[4] ),
    .X(_1512_));
 sg13g2_nand2_1 _5566_ (.Y(_1513_),
    .A(_1512_),
    .B(_1506_));
 sg13g2_o21ai_1 _5567_ (.B1(_1513_),
    .Y(_1142_),
    .A1(_1511_),
    .A2(_1507_));
 sg13g2_buf_1 _5568_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[5] ),
    .X(_1514_));
 sg13g2_mux2_1 _5569_ (.A0(_1373_),
    .A1(_1514_),
    .S(net100),
    .X(_1143_));
 sg13g2_buf_1 _5570_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[6] ),
    .X(_1515_));
 sg13g2_nand2_1 _5571_ (.Y(_1516_),
    .A(_1515_),
    .B(_1506_));
 sg13g2_o21ai_1 _5572_ (.B1(_1516_),
    .Y(_1144_),
    .A1(_1372_),
    .A2(net100));
 sg13g2_nor2b_1 _5573_ (.A(_1377_),
    .B_N(net309),
    .Y(_1517_));
 sg13g2_nand2b_1 _5574_ (.Y(_1518_),
    .B(net337),
    .A_N(_1510_));
 sg13g2_nor3_2 _5575_ (.A(_1453_),
    .B(_1517_),
    .C(_1518_),
    .Y(_1519_));
 sg13g2_and2_1 _5576_ (.A(_1456_),
    .B(_1519_),
    .X(_1520_));
 sg13g2_buf_1 _5577_ (.A(_1520_),
    .X(_1521_));
 sg13g2_a21oi_1 _5578_ (.A1(_1443_),
    .A2(_1521_),
    .Y(_1522_),
    .B1(_1483_));
 sg13g2_nor2_1 _5579_ (.A(_1399_),
    .B(_1522_),
    .Y(_1523_));
 sg13g2_buf_1 _5580_ (.A(_1523_),
    .X(_1524_));
 sg13g2_buf_1 _5581_ (.A(_1524_),
    .X(_1525_));
 sg13g2_buf_1 _5582_ (.A(_1393_),
    .X(_1526_));
 sg13g2_inv_1 _5583_ (.Y(_1527_),
    .A(_0108_));
 sg13g2_inv_1 _5584_ (.Y(_1528_),
    .A(_1514_));
 sg13g2_nand2b_1 _5585_ (.Y(_1529_),
    .B(net325),
    .A_N(_1512_));
 sg13g2_nand2_1 _5586_ (.Y(_1530_),
    .A(_1528_),
    .B(_1529_));
 sg13g2_inv_1 _5587_ (.Y(_1531_),
    .A(_1509_));
 sg13g2_nand2_1 _5588_ (.Y(_1532_),
    .A(_1512_),
    .B(_1514_));
 sg13g2_nand4_1 _5589_ (.B(_1531_),
    .C(net325),
    .A(_1508_),
    .Y(_1533_),
    .D(_1532_));
 sg13g2_o21ai_1 _5590_ (.B1(_1533_),
    .Y(_1534_),
    .A1(_1508_),
    .A2(_1530_));
 sg13g2_nor4_1 _5591_ (.A(_1508_),
    .B(net325),
    .C(_1512_),
    .D(_1528_),
    .Y(_1535_));
 sg13g2_a22oi_1 _5592_ (.Y(_1536_),
    .B1(_1535_),
    .B2(_1386_),
    .A2(_1534_),
    .A1(_1527_));
 sg13g2_nor2_1 _5593_ (.A(_1526_),
    .B(_1536_),
    .Y(_1537_));
 sg13g2_a21oi_1 _5594_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4] ),
    .A2(net229),
    .Y(_1538_),
    .B1(_1537_));
 sg13g2_buf_1 _5595_ (.A(_1524_),
    .X(_1539_));
 sg13g2_nand2_1 _5596_ (.Y(_1540_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .B(net91));
 sg13g2_o21ai_1 _5597_ (.B1(_1540_),
    .Y(_1145_),
    .A1(net92),
    .A2(_1538_));
 sg13g2_nor2_1 _5598_ (.A(_1508_),
    .B(_1512_),
    .Y(_1541_));
 sg13g2_o21ai_1 _5599_ (.B1(_1541_),
    .Y(_1542_),
    .A1(net325),
    .A2(_1514_));
 sg13g2_buf_1 _5600_ (.A(_1542_),
    .X(_1543_));
 sg13g2_inv_2 _5601_ (.Y(_1544_),
    .A(_1508_));
 sg13g2_o21ai_1 _5602_ (.B1(_1532_),
    .Y(_1545_),
    .A1(_1544_),
    .A2(net325));
 sg13g2_a22oi_1 _5603_ (.Y(_1546_),
    .B1(_1545_),
    .B2(_1531_),
    .A2(_1530_),
    .A1(_1544_));
 sg13g2_buf_1 _5604_ (.A(_1546_),
    .X(_1547_));
 sg13g2_nand2b_1 _5605_ (.Y(_1548_),
    .B(_1547_),
    .A_N(_0020_));
 sg13g2_o21ai_1 _5606_ (.B1(_1548_),
    .Y(_1549_),
    .A1(_0105_),
    .A2(_1543_));
 sg13g2_buf_1 _5607_ (.A(_1393_),
    .X(_1550_));
 sg13g2_and2_1 _5608_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5] ),
    .B(_1550_),
    .X(_1551_));
 sg13g2_a21oi_1 _5609_ (.A1(net247),
    .A2(_1549_),
    .Y(_1552_),
    .B1(_1551_));
 sg13g2_nand2_1 _5610_ (.Y(_1553_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .B(net91));
 sg13g2_o21ai_1 _5611_ (.B1(_1553_),
    .Y(_1146_),
    .A1(net92),
    .A2(_1552_));
 sg13g2_inv_1 _5612_ (.Y(_1554_),
    .A(_1543_));
 sg13g2_nor3_2 _5613_ (.A(_1544_),
    .B(_1509_),
    .C(net325),
    .Y(_1555_));
 sg13g2_buf_1 _5614_ (.A(_1555_),
    .X(_1556_));
 sg13g2_a221oi_1 _5615_ (.B2(_0019_),
    .C1(_1556_),
    .B1(_1554_),
    .A1(_0018_),
    .Y(_1557_),
    .A2(_1547_));
 sg13g2_and2_1 _5616_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6] ),
    .B(_1550_),
    .X(_1558_));
 sg13g2_a21oi_1 _5617_ (.A1(net247),
    .A2(_1557_),
    .Y(_1559_),
    .B1(_1558_));
 sg13g2_buf_1 _5618_ (.A(_1524_),
    .X(_1560_));
 sg13g2_nand2_1 _5619_ (.Y(_1561_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .B(_1560_));
 sg13g2_o21ai_1 _5620_ (.B1(_1561_),
    .Y(_1147_),
    .A1(_1525_),
    .A2(_1559_));
 sg13g2_nand2b_1 _5621_ (.Y(_1562_),
    .B(_1547_),
    .A_N(_0016_));
 sg13g2_o21ai_1 _5622_ (.B1(_1562_),
    .Y(_1563_),
    .A1(_0017_),
    .A2(_1543_));
 sg13g2_and2_1 _5623_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7] ),
    .B(_1393_),
    .X(_1564_));
 sg13g2_a21oi_1 _5624_ (.A1(net247),
    .A2(_1563_),
    .Y(_1565_),
    .B1(_1564_));
 sg13g2_nand2_1 _5625_ (.Y(_1566_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .B(net90));
 sg13g2_o21ai_1 _5626_ (.B1(_1566_),
    .Y(_1148_),
    .A1(_1525_),
    .A2(_1565_));
 sg13g2_buf_1 _5627_ (.A(_1393_),
    .X(_1567_));
 sg13g2_nand2b_1 _5628_ (.Y(_1568_),
    .B(_1543_),
    .A_N(_1547_));
 sg13g2_buf_2 _5629_ (.A(_1568_),
    .X(_1569_));
 sg13g2_nor2_1 _5630_ (.A(_0010_),
    .B(net227),
    .Y(_1570_));
 sg13g2_a22oi_1 _5631_ (.Y(_1571_),
    .B1(_1569_),
    .B2(_1570_),
    .A2(net225),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14] ));
 sg13g2_nand2_1 _5632_ (.Y(_1572_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10] ),
    .B(_1560_));
 sg13g2_o21ai_1 _5633_ (.B1(_1572_),
    .Y(_1149_),
    .A1(net92),
    .A2(_1571_));
 sg13g2_nor2_1 _5634_ (.A(_0009_),
    .B(_1545_),
    .Y(_1573_));
 sg13g2_mux2_1 _5635_ (.A0(_1527_),
    .A1(_1573_),
    .S(_1531_),
    .X(_1574_));
 sg13g2_mux2_1 _5636_ (.A0(_1386_),
    .A1(_1573_),
    .S(_1529_),
    .X(_1575_));
 sg13g2_mux2_1 _5637_ (.A0(_1574_),
    .A1(_1575_),
    .S(_1544_),
    .X(_1576_));
 sg13g2_and2_1 _5638_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15] ),
    .B(_1393_),
    .X(_1577_));
 sg13g2_a21oi_1 _5639_ (.A1(net247),
    .A2(_1576_),
    .Y(_1578_),
    .B1(_1577_));
 sg13g2_nand2_1 _5640_ (.Y(_1579_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11] ),
    .B(net90));
 sg13g2_o21ai_1 _5641_ (.B1(_1579_),
    .Y(_1150_),
    .A1(net92),
    .A2(_1578_));
 sg13g2_buf_1 _5642_ (.A(_1524_),
    .X(_1580_));
 sg13g2_nor2_1 _5643_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16] ),
    .B(net247),
    .Y(_1581_));
 sg13g2_buf_2 _5644_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[12] ),
    .X(_1582_));
 sg13g2_a21oi_1 _5645_ (.A1(_1531_),
    .A2(net325),
    .Y(_1583_),
    .B1(_1544_));
 sg13g2_buf_1 _5646_ (.A(_1583_),
    .X(_1584_));
 sg13g2_buf_1 _5647_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[31] ),
    .X(_1585_));
 sg13g2_nand2_1 _5648_ (.Y(_1586_),
    .A(_1585_),
    .B(_1532_));
 sg13g2_o21ai_1 _5649_ (.B1(_1399_),
    .Y(_1587_),
    .A1(_1584_),
    .A2(_1586_));
 sg13g2_buf_2 _5650_ (.A(_1587_),
    .X(_1588_));
 sg13g2_a21oi_1 _5651_ (.A1(_1582_),
    .A2(net262),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_nor3_1 _5652_ (.A(net89),
    .B(_1581_),
    .C(_1589_),
    .Y(_1590_));
 sg13g2_a21o_1 _5653_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12] ),
    .B1(_1590_),
    .X(_1151_));
 sg13g2_nor2_1 _5654_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17] ),
    .B(_1400_),
    .Y(_1591_));
 sg13g2_a21oi_1 _5655_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ),
    .A2(net262),
    .Y(_1592_),
    .B1(_1588_));
 sg13g2_nor3_1 _5656_ (.A(_1580_),
    .B(_1591_),
    .C(_1592_),
    .Y(_1593_));
 sg13g2_a21o_1 _5657_ (.A2(_1539_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13] ),
    .B1(_1593_),
    .X(_1152_));
 sg13g2_nor2_1 _5658_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18] ),
    .B(net247),
    .Y(_1594_));
 sg13g2_a21oi_1 _5659_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ),
    .A2(net262),
    .Y(_1595_),
    .B1(_1588_));
 sg13g2_nor3_1 _5660_ (.A(net89),
    .B(_1594_),
    .C(_1595_),
    .Y(_1596_));
 sg13g2_a21o_1 _5661_ (.A2(_1539_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14] ),
    .B1(_1596_),
    .X(_1153_));
 sg13g2_nor2_1 _5662_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19] ),
    .B(net247),
    .Y(_1597_));
 sg13g2_a21oi_1 _5663_ (.A1(_1402_),
    .A2(net262),
    .Y(_1598_),
    .B1(_1588_));
 sg13g2_nor3_1 _5664_ (.A(net89),
    .B(_1597_),
    .C(_1598_),
    .Y(_1599_));
 sg13g2_a21o_1 _5665_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15] ),
    .B1(_1599_),
    .X(_1154_));
 sg13g2_nor2_1 _5666_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20] ),
    .B(_1399_),
    .Y(_1600_));
 sg13g2_a21oi_1 _5667_ (.A1(_1408_),
    .A2(net262),
    .Y(_1601_),
    .B1(_1588_));
 sg13g2_nor3_1 _5668_ (.A(net89),
    .B(_1600_),
    .C(_1601_),
    .Y(_1602_));
 sg13g2_a21o_1 _5669_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16] ),
    .B1(_1602_),
    .X(_1155_));
 sg13g2_nor2_1 _5670_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21] ),
    .B(_1399_),
    .Y(_1603_));
 sg13g2_a21oi_1 _5671_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ),
    .A2(net262),
    .Y(_1604_),
    .B1(_1588_));
 sg13g2_nor3_1 _5672_ (.A(net89),
    .B(_1603_),
    .C(_1604_),
    .Y(_1605_));
 sg13g2_a21o_1 _5673_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17] ),
    .B1(_1605_),
    .X(_1156_));
 sg13g2_nor2_1 _5674_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22] ),
    .B(_1399_),
    .Y(_1606_));
 sg13g2_a21oi_1 _5675_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ),
    .A2(net262),
    .Y(_1607_),
    .B1(_1588_));
 sg13g2_nor3_1 _5676_ (.A(net89),
    .B(_1606_),
    .C(_1607_),
    .Y(_1608_));
 sg13g2_a21o_1 _5677_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18] ),
    .B1(_1608_),
    .X(_1157_));
 sg13g2_nor2_1 _5678_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23] ),
    .B(_1399_),
    .Y(_1609_));
 sg13g2_a21oi_1 _5679_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ),
    .A2(net262),
    .Y(_1610_),
    .B1(_1588_));
 sg13g2_nor3_1 _5680_ (.A(net89),
    .B(_1609_),
    .C(_1610_),
    .Y(_1611_));
 sg13g2_a21o_1 _5681_ (.A2(net91),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19] ),
    .B1(_1611_),
    .X(_1158_));
 sg13g2_and2_1 _5682_ (.A(_1585_),
    .B(_1569_),
    .X(_1612_));
 sg13g2_buf_1 _5683_ (.A(_1612_),
    .X(_1613_));
 sg13g2_a21oi_1 _5684_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ),
    .A2(net263),
    .Y(_1614_),
    .B1(net98));
 sg13g2_nor2_1 _5685_ (.A(net226),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_a21oi_1 _5686_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24] ),
    .A2(net229),
    .Y(_1616_),
    .B1(_1615_));
 sg13g2_nand2_1 _5687_ (.Y(_1617_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20] ),
    .B(net90));
 sg13g2_o21ai_1 _5688_ (.B1(_1617_),
    .Y(_1159_),
    .A1(net92),
    .A2(_1616_));
 sg13g2_a21oi_1 _5689_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ),
    .A2(net263),
    .Y(_1618_),
    .B1(net98));
 sg13g2_nor2_1 _5690_ (.A(net226),
    .B(_1618_),
    .Y(_1619_));
 sg13g2_a21oi_1 _5691_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25] ),
    .A2(net225),
    .Y(_1620_),
    .B1(_1619_));
 sg13g2_nand2_1 _5692_ (.Y(_1621_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21] ),
    .B(net90));
 sg13g2_o21ai_1 _5693_ (.B1(_1621_),
    .Y(_1160_),
    .A1(net92),
    .A2(_1620_));
 sg13g2_a21oi_1 _5694_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ),
    .A2(net263),
    .Y(_1622_),
    .B1(net98));
 sg13g2_nor2_1 _5695_ (.A(net226),
    .B(_1622_),
    .Y(_1623_));
 sg13g2_a21oi_1 _5696_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26] ),
    .A2(net225),
    .Y(_1624_),
    .B1(_1623_));
 sg13g2_nand2_1 _5697_ (.Y(_1625_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22] ),
    .B(net90));
 sg13g2_o21ai_1 _5698_ (.B1(_1625_),
    .Y(_1161_),
    .A1(net92),
    .A2(_1624_));
 sg13g2_a21oi_1 _5699_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ),
    .A2(net263),
    .Y(_1626_),
    .B1(net98));
 sg13g2_nor2_1 _5700_ (.A(net226),
    .B(_1626_),
    .Y(_1627_));
 sg13g2_a21oi_1 _5701_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27] ),
    .A2(net225),
    .Y(_1628_),
    .B1(_1627_));
 sg13g2_nand2_1 _5702_ (.Y(_1629_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23] ),
    .B(net90));
 sg13g2_o21ai_1 _5703_ (.B1(_1629_),
    .Y(_1162_),
    .A1(net92),
    .A2(_1628_));
 sg13g2_buf_1 _5704_ (.A(_1524_),
    .X(_1630_));
 sg13g2_a21oi_1 _5705_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ),
    .A2(net263),
    .Y(_1631_),
    .B1(_1613_));
 sg13g2_nor2_1 _5706_ (.A(net226),
    .B(_1631_),
    .Y(_1632_));
 sg13g2_a21oi_1 _5707_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28] ),
    .A2(_1567_),
    .Y(_1633_),
    .B1(_1632_));
 sg13g2_nand2_1 _5708_ (.Y(_1634_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24] ),
    .B(net90));
 sg13g2_o21ai_1 _5709_ (.B1(_1634_),
    .Y(_1163_),
    .A1(_1630_),
    .A2(_1633_));
 sg13g2_a21oi_1 _5710_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5] ),
    .A2(_1555_),
    .Y(_1635_),
    .B1(net98));
 sg13g2_nor2_1 _5711_ (.A(net226),
    .B(_1635_),
    .Y(_1636_));
 sg13g2_a21oi_1 _5712_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29] ),
    .A2(_1567_),
    .Y(_1637_),
    .B1(_1636_));
 sg13g2_nand2_1 _5713_ (.Y(_1638_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25] ),
    .B(net90));
 sg13g2_o21ai_1 _5714_ (.B1(_1638_),
    .Y(_1164_),
    .A1(net88),
    .A2(_1637_));
 sg13g2_a21oi_1 _5715_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6] ),
    .A2(_1555_),
    .Y(_1639_),
    .B1(net98));
 sg13g2_nor2_1 _5716_ (.A(net226),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_a21oi_1 _5717_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30] ),
    .A2(net225),
    .Y(_1641_),
    .B1(_1640_));
 sg13g2_buf_1 _5718_ (.A(_1524_),
    .X(_1642_));
 sg13g2_nand2_1 _5719_ (.Y(_1643_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26] ),
    .B(net87));
 sg13g2_o21ai_1 _5720_ (.B1(_1643_),
    .Y(_1165_),
    .A1(net88),
    .A2(_1641_));
 sg13g2_a21oi_1 _5721_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7] ),
    .A2(_1555_),
    .Y(_1644_),
    .B1(net98));
 sg13g2_nor2_1 _5722_ (.A(net226),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_a21oi_1 _5723_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31] ),
    .A2(net225),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_nand2_1 _5724_ (.Y(_1647_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27] ),
    .B(net87));
 sg13g2_o21ai_1 _5725_ (.B1(_1647_),
    .Y(_1166_),
    .A1(_1630_),
    .A2(_1646_));
 sg13g2_or2_1 _5726_ (.X(_1648_),
    .B(net98),
    .A(_1524_));
 sg13g2_buf_1 _5727_ (.A(_1648_),
    .X(_1649_));
 sg13g2_a21oi_1 _5728_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8] ),
    .A2(net263),
    .Y(_1650_),
    .B1(_1649_));
 sg13g2_a21oi_1 _5729_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28] ),
    .A2(_1642_),
    .Y(_1651_),
    .B1(net228));
 sg13g2_nor2_1 _5730_ (.A(_1650_),
    .B(_1651_),
    .Y(_1167_));
 sg13g2_a21oi_1 _5731_ (.A1(_1502_),
    .A2(net263),
    .Y(_1652_),
    .B1(_1649_));
 sg13g2_a21oi_1 _5732_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29] ),
    .A2(_1580_),
    .Y(_1653_),
    .B1(net228));
 sg13g2_nor2_1 _5733_ (.A(_1652_),
    .B(_1653_),
    .Y(_1168_));
 sg13g2_a21oi_1 _5734_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ),
    .A2(net263),
    .Y(_1654_),
    .B1(_1649_));
 sg13g2_a21oi_1 _5735_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30] ),
    .A2(net89),
    .Y(_1655_),
    .B1(net246));
 sg13g2_nor2_1 _5736_ (.A(_1654_),
    .B(_1655_),
    .Y(_1169_));
 sg13g2_nor2_1 _5737_ (.A(_1556_),
    .B(_1569_),
    .Y(_1656_));
 sg13g2_nand2_1 _5738_ (.Y(_1657_),
    .A(_1585_),
    .B(net246));
 sg13g2_nand2_1 _5739_ (.Y(_1658_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31] ),
    .B(_1642_));
 sg13g2_o21ai_1 _5740_ (.B1(_1658_),
    .Y(_1170_),
    .A1(_1656_),
    .A2(_1657_));
 sg13g2_inv_1 _5741_ (.Y(_1659_),
    .A(_0000_));
 sg13g2_nand2_1 _5742_ (.Y(_1660_),
    .A(_1659_),
    .B(_1547_));
 sg13g2_o21ai_1 _5743_ (.B1(_1660_),
    .Y(_1661_),
    .A1(_0015_),
    .A2(_1543_));
 sg13g2_and2_1 _5744_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8] ),
    .B(_1393_),
    .X(_1662_));
 sg13g2_a21oi_1 _5745_ (.A1(net247),
    .A2(_1661_),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nand2_1 _5746_ (.Y(_1664_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4] ),
    .B(net87));
 sg13g2_o21ai_1 _5747_ (.B1(_1664_),
    .Y(_1171_),
    .A1(net88),
    .A2(_1663_));
 sg13g2_nor2_1 _5748_ (.A(_0014_),
    .B(net227),
    .Y(_1665_));
 sg13g2_a22oi_1 _5749_ (.Y(_1666_),
    .B1(_1569_),
    .B2(_1665_),
    .A2(net225),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9] ));
 sg13g2_nand2_1 _5750_ (.Y(_1667_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5] ),
    .B(net87));
 sg13g2_o21ai_1 _5751_ (.B1(_1667_),
    .Y(_1172_),
    .A1(net88),
    .A2(_1666_));
 sg13g2_nor2_1 _5752_ (.A(_0013_),
    .B(net227),
    .Y(_1668_));
 sg13g2_a22oi_1 _5753_ (.Y(_1669_),
    .B1(_1569_),
    .B2(_1668_),
    .A2(net225),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10] ));
 sg13g2_nand2_1 _5754_ (.Y(_1670_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6] ),
    .B(net87));
 sg13g2_o21ai_1 _5755_ (.B1(_1670_),
    .Y(_1173_),
    .A1(net88),
    .A2(_1669_));
 sg13g2_nor2_1 _5756_ (.A(_0012_),
    .B(net227),
    .Y(_1671_));
 sg13g2_a22oi_1 _5757_ (.Y(_1672_),
    .B1(_1569_),
    .B2(_1671_),
    .A2(net227),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11] ));
 sg13g2_nand2_1 _5758_ (.Y(_1673_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7] ),
    .B(net87));
 sg13g2_o21ai_1 _5759_ (.B1(_1673_),
    .Y(_1174_),
    .A1(net88),
    .A2(_1672_));
 sg13g2_nor2_1 _5760_ (.A(_0114_),
    .B(net227),
    .Y(_1674_));
 sg13g2_a22oi_1 _5761_ (.Y(_1675_),
    .B1(_1569_),
    .B2(_1674_),
    .A2(net227),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12] ));
 sg13g2_nand2_1 _5762_ (.Y(_1676_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8] ),
    .B(net87));
 sg13g2_o21ai_1 _5763_ (.B1(_1676_),
    .Y(_1175_),
    .A1(net88),
    .A2(_1675_));
 sg13g2_nor2_1 _5764_ (.A(_0011_),
    .B(_1526_),
    .Y(_1677_));
 sg13g2_a22oi_1 _5765_ (.Y(_1678_),
    .B1(_1569_),
    .B2(_1677_),
    .A2(net227),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13] ));
 sg13g2_nand2_1 _5766_ (.Y(_1679_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9] ),
    .B(net87));
 sg13g2_o21ai_1 _5767_ (.B1(_1679_),
    .Y(_1176_),
    .A1(net88),
    .A2(_1678_));
 sg13g2_inv_1 _5768_ (.Y(_1680_),
    .A(net335));
 sg13g2_nand2_1 _5769_ (.Y(_1681_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ),
    .B(_1506_));
 sg13g2_o21ai_1 _5770_ (.B1(_1681_),
    .Y(_1181_),
    .A1(_1680_),
    .A2(net100));
 sg13g2_inv_2 _5771_ (.Y(_1682_),
    .A(net331));
 sg13g2_nand2_1 _5772_ (.Y(_1683_),
    .A(_1582_),
    .B(_1506_));
 sg13g2_o21ai_1 _5773_ (.B1(_1683_),
    .Y(_1182_),
    .A1(_1682_),
    .A2(net100));
 sg13g2_mux2_1 _5774_ (.A0(net309),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ),
    .S(_1507_),
    .X(_1183_));
 sg13g2_mux2_1 _5775_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10] ),
    .S(net75),
    .X(_1216_));
 sg13g2_mux2_1 _5776_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11] ),
    .S(net75),
    .X(_1217_));
 sg13g2_buf_1 _5777_ (.A(_1492_),
    .X(_1684_));
 sg13g2_mux2_1 _5778_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12] ),
    .S(net73),
    .X(_1218_));
 sg13g2_mux2_1 _5779_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13] ),
    .S(net73),
    .X(_1219_));
 sg13g2_mux2_1 _5780_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14] ),
    .S(net73),
    .X(_1220_));
 sg13g2_mux2_1 _5781_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15] ),
    .S(net73),
    .X(_1221_));
 sg13g2_mux2_1 _5782_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16] ),
    .S(net73),
    .X(_1222_));
 sg13g2_mux2_1 _5783_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17] ),
    .S(net73),
    .X(_1223_));
 sg13g2_mux2_1 _5784_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18] ),
    .S(net73),
    .X(_1224_));
 sg13g2_mux2_1 _5785_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19] ),
    .S(net73),
    .X(_1225_));
 sg13g2_mux2_1 _5786_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20] ),
    .S(_1684_),
    .X(_1226_));
 sg13g2_mux2_1 _5787_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21] ),
    .S(_1684_),
    .X(_1227_));
 sg13g2_buf_1 _5788_ (.A(_1492_),
    .X(_1685_));
 sg13g2_mux2_1 _5789_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22] ),
    .S(net72),
    .X(_1228_));
 sg13g2_mux2_1 _5790_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23] ),
    .S(net72),
    .X(_1229_));
 sg13g2_mux2_1 _5791_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24] ),
    .S(net72),
    .X(_1230_));
 sg13g2_mux2_1 _5792_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25] ),
    .S(net72),
    .X(_1231_));
 sg13g2_mux2_1 _5793_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26] ),
    .S(net72),
    .X(_1232_));
 sg13g2_mux2_1 _5794_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27] ),
    .S(net72),
    .X(_1233_));
 sg13g2_buf_1 _5795_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ),
    .X(_1686_));
 sg13g2_nand2b_1 _5796_ (.Y(_1687_),
    .B(_1510_),
    .A_N(_1444_));
 sg13g2_buf_1 _5797_ (.A(_0022_),
    .X(_1688_));
 sg13g2_nand2b_1 _5798_ (.Y(_1689_),
    .B(net324),
    .A_N(net336));
 sg13g2_or2_1 _5799_ (.X(_1690_),
    .B(net337),
    .A(net335));
 sg13g2_buf_1 _5800_ (.A(_1690_),
    .X(_1691_));
 sg13g2_a21o_1 _5801_ (.A2(_1689_),
    .A1(_1687_),
    .B1(_1691_),
    .X(_1692_));
 sg13g2_buf_1 _5802_ (.A(_1692_),
    .X(_1693_));
 sg13g2_buf_1 _5803_ (.A(net245),
    .X(_1694_));
 sg13g2_nand2_1 _5804_ (.Y(_1695_),
    .A(net328),
    .B(net224));
 sg13g2_or3_1 _5805_ (.A(net335),
    .B(net337),
    .C(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5] ),
    .X(_1696_));
 sg13g2_a21oi_1 _5806_ (.A1(_1687_),
    .A2(_1689_),
    .Y(_1697_),
    .B1(_1696_));
 sg13g2_o21ai_1 _5807_ (.B1(net332),
    .Y(_1698_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3] ),
    .A2(_1697_));
 sg13g2_a21o_1 _5808_ (.A2(_1698_),
    .A1(_1695_),
    .B1(net230),
    .X(_1699_));
 sg13g2_nor2_1 _5809_ (.A(_1499_),
    .B(net248),
    .Y(_1700_));
 sg13g2_inv_1 _5810_ (.Y(_1701_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2] ));
 sg13g2_a21oi_1 _5811_ (.A1(_1687_),
    .A2(_1689_),
    .Y(_1702_),
    .B1(_1691_));
 sg13g2_buf_1 _5812_ (.A(_1702_),
    .X(_1703_));
 sg13g2_nor2_1 _5813_ (.A(_1701_),
    .B(net244),
    .Y(_1704_));
 sg13g2_nand3_1 _5814_ (.B(_1376_),
    .C(_1380_),
    .A(_1372_),
    .Y(_1705_));
 sg13g2_buf_2 _5815_ (.A(_1705_),
    .X(_1706_));
 sg13g2_nand2_1 _5816_ (.Y(_1707_),
    .A(net332),
    .B(_1706_));
 sg13g2_o21ai_1 _5817_ (.B1(_1707_),
    .Y(_1708_),
    .A1(_1700_),
    .A2(_1704_));
 sg13g2_buf_2 _5818_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[2] ),
    .X(_1709_));
 sg13g2_buf_1 _5819_ (.A(_1703_),
    .X(_1710_));
 sg13g2_nand2_1 _5820_ (.Y(_1711_),
    .A(net328),
    .B(_1706_));
 sg13g2_nand3_1 _5821_ (.B(net223),
    .C(_1711_),
    .A(_1709_),
    .Y(_1712_));
 sg13g2_nand4_1 _5822_ (.B(_1699_),
    .C(_1708_),
    .A(net308),
    .Y(_1713_),
    .D(_1712_));
 sg13g2_inv_1 _5823_ (.Y(_1714_),
    .A(_1480_));
 sg13g2_inv_1 _5824_ (.Y(_1715_),
    .A(_1709_));
 sg13g2_nand2b_1 _5825_ (.Y(_1716_),
    .B(net336),
    .A_N(_1373_));
 sg13g2_buf_1 _5826_ (.A(_1716_),
    .X(_1717_));
 sg13g2_nor2_1 _5827_ (.A(net337),
    .B(_1717_),
    .Y(_1718_));
 sg13g2_xnor2_1 _5828_ (.Y(_1719_),
    .A(net328),
    .B(net244));
 sg13g2_a221oi_1 _5829_ (.B2(_1441_),
    .C1(net306),
    .B1(_1719_),
    .A1(_1718_),
    .Y(_1720_),
    .A2(_1380_));
 sg13g2_buf_1 _5830_ (.A(_1720_),
    .X(_1721_));
 sg13g2_or2_1 _5831_ (.X(_1722_),
    .B(net328),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4] ));
 sg13g2_a21oi_1 _5832_ (.A1(_1706_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(net224));
 sg13g2_buf_2 _5833_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[1] ),
    .X(_1724_));
 sg13g2_inv_1 _5834_ (.Y(_1725_),
    .A(_1724_));
 sg13g2_nor2_1 _5835_ (.A(net332),
    .B(_1499_),
    .Y(_1726_));
 sg13g2_buf_2 _5836_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[0] ),
    .X(_1727_));
 sg13g2_inv_1 _5837_ (.Y(_1728_),
    .A(_1727_));
 sg13g2_a22oi_1 _5838_ (.Y(_1729_),
    .B1(_1726_),
    .B2(_1728_),
    .A2(_1725_),
    .A1(net332));
 sg13g2_a21oi_1 _5839_ (.A1(_1709_),
    .A2(_1723_),
    .Y(_1730_),
    .B1(_1729_));
 sg13g2_a221oi_1 _5840_ (.B2(_1730_),
    .C1(net328),
    .B1(_1721_),
    .A1(net306),
    .Y(_1731_),
    .A2(_1715_));
 sg13g2_buf_1 _5841_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[1] ),
    .X(_1732_));
 sg13g2_o21ai_1 _5842_ (.B1(net332),
    .Y(_1733_),
    .A1(_1732_),
    .A2(_1697_));
 sg13g2_a21o_1 _5843_ (.A2(_1733_),
    .A1(_1695_),
    .B1(net230),
    .X(_1734_));
 sg13g2_and2_1 _5844_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0] ),
    .B(_1694_),
    .X(_1735_));
 sg13g2_o21ai_1 _5845_ (.B1(_1707_),
    .Y(_1736_),
    .A1(_1700_),
    .A2(_1735_));
 sg13g2_nand3_1 _5846_ (.B(net223),
    .C(_1711_),
    .A(_1727_),
    .Y(_1737_));
 sg13g2_nand4_1 _5847_ (.B(_1734_),
    .C(_1736_),
    .A(net308),
    .Y(_1738_),
    .D(_1737_));
 sg13g2_inv_1 _5848_ (.Y(_1739_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3] ));
 sg13g2_a22oi_1 _5849_ (.Y(_1740_),
    .B1(_1726_),
    .B2(_1701_),
    .A2(_1739_),
    .A1(net332));
 sg13g2_a21oi_1 _5850_ (.A1(_1727_),
    .A2(_1723_),
    .Y(_1741_),
    .B1(_1740_));
 sg13g2_a221oi_1 _5851_ (.B2(_1741_),
    .C1(_1499_),
    .B1(_1721_),
    .A1(net306),
    .Y(_1742_),
    .A2(_1728_));
 sg13g2_a22oi_1 _5852_ (.Y(_1743_),
    .B1(_1738_),
    .B2(_1742_),
    .A2(_1731_),
    .A1(_1713_));
 sg13g2_nor2_2 _5853_ (.A(net335),
    .B(_1371_),
    .Y(_1744_));
 sg13g2_nand2_1 _5854_ (.Y(_1745_),
    .A(_1687_),
    .B(_1689_));
 sg13g2_nand4_1 _5855_ (.B(_1682_),
    .C(_1376_),
    .A(_1372_),
    .Y(_1746_),
    .D(_1517_));
 sg13g2_o21ai_1 _5856_ (.B1(_0110_),
    .Y(_1747_),
    .A1(_1717_),
    .A2(_1449_));
 sg13g2_a221oi_1 _5857_ (.B2(_1747_),
    .C1(_1478_),
    .B1(_1746_),
    .A1(_1744_),
    .Y(_1748_),
    .A2(_1745_));
 sg13g2_and4_1 _5858_ (.A(_1478_),
    .B(net245),
    .C(_1746_),
    .D(_1747_),
    .X(_1749_));
 sg13g2_buf_1 _5859_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[8] ),
    .X(_1750_));
 sg13g2_inv_1 _5860_ (.Y(_1751_),
    .A(_1750_));
 sg13g2_nand2_1 _5861_ (.Y(_1752_),
    .A(_1751_),
    .B(_1478_));
 sg13g2_nand2_1 _5862_ (.Y(_1753_),
    .A(_1750_),
    .B(net330));
 sg13g2_a21oi_1 _5863_ (.A1(_1752_),
    .A2(_1753_),
    .Y(_1754_),
    .B1(net245));
 sg13g2_or3_1 _5864_ (.A(_1748_),
    .B(_1749_),
    .C(_1754_),
    .X(_1755_));
 sg13g2_buf_1 _5865_ (.A(_1755_),
    .X(_1756_));
 sg13g2_buf_1 _5866_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[7] ),
    .X(_1757_));
 sg13g2_nand2b_1 _5867_ (.Y(_1758_),
    .B(net309),
    .A_N(net335));
 sg13g2_nand2b_1 _5868_ (.Y(_1759_),
    .B(net331),
    .A_N(net309));
 sg13g2_o21ai_1 _5869_ (.B1(_1759_),
    .Y(_1760_),
    .A1(net331),
    .A2(_1758_));
 sg13g2_a21o_1 _5870_ (.A2(_1760_),
    .A1(_1718_),
    .B1(net244),
    .X(_1761_));
 sg13g2_nor3_1 _5871_ (.A(net331),
    .B(_1717_),
    .C(_1449_),
    .Y(_1762_));
 sg13g2_nor2_1 _5872_ (.A(net323),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_buf_1 _5873_ (.A(_0030_),
    .X(_1764_));
 sg13g2_a221oi_1 _5874_ (.B2(net245),
    .C1(net322),
    .B1(_1763_),
    .A1(net323),
    .Y(_1765_),
    .A2(_1761_));
 sg13g2_buf_1 _5875_ (.A(_1765_),
    .X(_1766_));
 sg13g2_inv_1 _5876_ (.Y(_1767_),
    .A(net322));
 sg13g2_nand3_1 _5877_ (.B(_1376_),
    .C(_1452_),
    .A(_1682_),
    .Y(_1768_));
 sg13g2_a21oi_1 _5878_ (.A1(net245),
    .A2(_1768_),
    .Y(_1769_),
    .B1(net323));
 sg13g2_inv_1 _5879_ (.Y(_1770_),
    .A(net323));
 sg13g2_a221oi_1 _5880_ (.B2(_1718_),
    .C1(_1770_),
    .B1(_1760_),
    .A1(_1744_),
    .Y(_1771_),
    .A2(_1745_));
 sg13g2_buf_1 _5881_ (.A(_1771_),
    .X(_1772_));
 sg13g2_nor3_2 _5882_ (.A(_1767_),
    .B(_1769_),
    .C(_1772_),
    .Y(_1773_));
 sg13g2_nor2_1 _5883_ (.A(net248),
    .B(net244),
    .Y(_1774_));
 sg13g2_buf_1 _5884_ (.A(_0031_),
    .X(_1775_));
 sg13g2_inv_1 _5885_ (.Y(_1776_),
    .A(\i_exotiny._2356_[0] ));
 sg13g2_nor2_1 _5886_ (.A(_1775_),
    .B(_1776_),
    .Y(_1777_));
 sg13g2_inv_1 _5887_ (.Y(_1778_),
    .A(_1370_));
 sg13g2_a21oi_1 _5888_ (.A1(_1778_),
    .A2(net244),
    .Y(_1779_),
    .B1(\i_exotiny._2356_[0] ));
 sg13g2_nand3b_1 _5889_ (.B(_1706_),
    .C(net245),
    .Y(_1780_),
    .A_N(_1775_));
 sg13g2_nor3_1 _5890_ (.A(_1370_),
    .B(_1776_),
    .C(net245),
    .Y(_1781_));
 sg13g2_a221oi_1 _5891_ (.B2(_1780_),
    .C1(_1781_),
    .B1(_1779_),
    .A1(_1774_),
    .Y(_1782_),
    .A2(_1777_));
 sg13g2_buf_1 _5892_ (.A(_1782_),
    .X(_1783_));
 sg13g2_nor4_2 _5893_ (.A(_1756_),
    .B(_1766_),
    .C(_1773_),
    .Y(_1784_),
    .D(_1783_));
 sg13g2_buf_8 _5894_ (.A(_1784_),
    .X(_1785_));
 sg13g2_nand2_1 _5895_ (.Y(_1786_),
    .A(_1510_),
    .B(_0037_));
 sg13g2_o21ai_1 _5896_ (.B1(_1786_),
    .Y(_1787_),
    .A1(_1680_),
    .A2(_1510_));
 sg13g2_nor2_1 _5897_ (.A(_1707_),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_nand2_1 _5898_ (.Y(_1789_),
    .A(_1785_),
    .B(_1788_));
 sg13g2_nor2_1 _5899_ (.A(_0036_),
    .B(_1722_),
    .Y(_1790_));
 sg13g2_nor3_1 _5900_ (.A(_0007_),
    .B(net332),
    .C(_1499_),
    .Y(_1791_));
 sg13g2_buf_1 _5901_ (.A(_1706_),
    .X(_1792_));
 sg13g2_a22oi_1 _5902_ (.Y(_1793_),
    .B1(_1791_),
    .B2(net222),
    .A2(_1790_),
    .A1(net224));
 sg13g2_nand3b_1 _5903_ (.B(net248),
    .C(net224),
    .Y(_1794_),
    .A_N(_0036_));
 sg13g2_a21o_1 _5904_ (.A2(_1794_),
    .A1(_1793_),
    .B1(net306),
    .X(_1795_));
 sg13g2_inv_1 _5905_ (.Y(_1796_),
    .A(_0006_));
 sg13g2_buf_1 _5906_ (.A(_1441_),
    .X(_1797_));
 sg13g2_nand4_1 _5907_ (.B(net305),
    .C(net308),
    .A(_1796_),
    .Y(_1798_),
    .D(_1706_));
 sg13g2_or4_1 _5908_ (.A(_0008_),
    .B(_1442_),
    .C(net306),
    .D(net248),
    .X(_1799_));
 sg13g2_mux2_1 _5909_ (.A0(_1798_),
    .A1(_1799_),
    .S(_1719_),
    .X(_1800_));
 sg13g2_o21ai_1 _5910_ (.B1(net223),
    .Y(_1801_),
    .A1(_1442_),
    .A2(_1383_));
 sg13g2_a21o_1 _5911_ (.A2(_1801_),
    .A1(_1481_),
    .B1(_0004_),
    .X(_1802_));
 sg13g2_nand4_1 _5912_ (.B(_1795_),
    .C(_1800_),
    .A(_1711_),
    .Y(_1803_),
    .D(_1802_));
 sg13g2_nand2_1 _5913_ (.Y(_1804_),
    .A(net328),
    .B(_1725_));
 sg13g2_o21ai_1 _5914_ (.B1(_1442_),
    .Y(_1805_),
    .A1(_1481_),
    .A2(_1804_));
 sg13g2_a21oi_1 _5915_ (.A1(net222),
    .A2(_1805_),
    .Y(_1806_),
    .B1(_1787_));
 sg13g2_nand3_1 _5916_ (.B(_1727_),
    .C(net222),
    .A(net305),
    .Y(_1807_));
 sg13g2_nand3_1 _5917_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2] ),
    .C(_1706_),
    .A(net305),
    .Y(_1808_));
 sg13g2_mux2_1 _5918_ (.A0(_1807_),
    .A1(_1808_),
    .S(_1719_),
    .X(_1809_));
 sg13g2_o21ai_1 _5919_ (.B1(net328),
    .Y(_1810_),
    .A1(_1739_),
    .A2(net248));
 sg13g2_inv_1 _5920_ (.Y(_1811_),
    .A(_1732_));
 sg13g2_nand3_1 _5921_ (.B(_1811_),
    .C(_1694_),
    .A(_1499_),
    .Y(_1812_));
 sg13g2_nand3_1 _5922_ (.B(_1810_),
    .C(_1812_),
    .A(_1442_),
    .Y(_1813_));
 sg13g2_nand4_1 _5923_ (.B(_1700_),
    .C(_1809_),
    .A(net308),
    .Y(_1814_),
    .D(_1813_));
 sg13g2_nand4_1 _5924_ (.B(_1803_),
    .C(_1806_),
    .A(_1785_),
    .Y(_1815_),
    .D(_1814_));
 sg13g2_o21ai_1 _5925_ (.B1(_1815_),
    .Y(_1816_),
    .A1(_1743_),
    .A2(_1789_));
 sg13g2_buf_8 _5926_ (.A(_1816_),
    .X(_1817_));
 sg13g2_nand3_1 _5927_ (.B(_1746_),
    .C(_1747_),
    .A(_1693_),
    .Y(_1818_));
 sg13g2_buf_2 _5928_ (.A(_1818_),
    .X(_1819_));
 sg13g2_o21ai_1 _5929_ (.B1(_1819_),
    .Y(_1820_),
    .A1(_1750_),
    .A2(net224));
 sg13g2_inv_1 _5930_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_or3_1 _5931_ (.A(_1766_),
    .B(_1773_),
    .C(_1783_),
    .X(_1822_));
 sg13g2_buf_2 _5932_ (.A(_1822_),
    .X(_1823_));
 sg13g2_buf_1 _5933_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ),
    .X(_1824_));
 sg13g2_a21oi_1 _5934_ (.A1(_1751_),
    .A2(net244),
    .Y(_1825_),
    .B1(_1824_));
 sg13g2_nand2_1 _5935_ (.Y(_1826_),
    .A(_1819_),
    .B(_1825_));
 sg13g2_nand3_1 _5936_ (.B(_1474_),
    .C(net223),
    .A(_1778_),
    .Y(_1827_));
 sg13g2_inv_1 _5937_ (.Y(_1828_),
    .A(_1474_));
 sg13g2_or4_1 _5938_ (.A(_1775_),
    .B(_1828_),
    .C(net248),
    .D(net244),
    .X(_1829_));
 sg13g2_nor3_1 _5939_ (.A(net323),
    .B(net223),
    .C(_1762_),
    .Y(_1830_));
 sg13g2_a221oi_1 _5940_ (.B2(_1829_),
    .C1(_1830_),
    .B1(_1827_),
    .A1(net323),
    .Y(_1831_),
    .A2(_1761_));
 sg13g2_nor3_1 _5941_ (.A(_1370_),
    .B(_1828_),
    .C(net245),
    .Y(_1832_));
 sg13g2_nor4_1 _5942_ (.A(_1775_),
    .B(_1828_),
    .C(_1382_),
    .D(net244),
    .Y(_1833_));
 sg13g2_or4_1 _5943_ (.A(_1769_),
    .B(_1772_),
    .C(_1832_),
    .D(_1833_),
    .X(_1834_));
 sg13g2_buf_1 _5944_ (.A(_1834_),
    .X(_1835_));
 sg13g2_a21oi_1 _5945_ (.A1(_1819_),
    .A2(_1825_),
    .Y(_1836_),
    .B1(net322));
 sg13g2_a22oi_1 _5946_ (.Y(_1837_),
    .B1(_1835_),
    .B2(_1836_),
    .A2(_1831_),
    .A1(_1826_));
 sg13g2_nand4_1 _5947_ (.B(_1821_),
    .C(_1823_),
    .A(_1478_),
    .Y(_1838_),
    .D(_1837_));
 sg13g2_nor2_1 _5948_ (.A(net305),
    .B(_1498_),
    .Y(_1839_));
 sg13g2_nor2_1 _5949_ (.A(net230),
    .B(_1839_),
    .Y(_1840_));
 sg13g2_and2_1 _5950_ (.A(_1819_),
    .B(_1825_),
    .X(_1841_));
 sg13g2_buf_1 _5951_ (.A(_1841_),
    .X(_1842_));
 sg13g2_buf_1 _5952_ (.A(net224),
    .X(_1843_));
 sg13g2_a221oi_1 _5953_ (.B2(net330),
    .C1(net174),
    .B1(_1842_),
    .A1(_1785_),
    .Y(_1844_),
    .A2(_1840_));
 sg13g2_nand4_1 _5954_ (.B(_1820_),
    .C(_1823_),
    .A(net330),
    .Y(_1845_),
    .D(_1837_));
 sg13g2_and3_1 _5955_ (.X(_1846_),
    .A(_1838_),
    .B(_1844_),
    .C(_1845_));
 sg13g2_nor2_1 _5956_ (.A(_1769_),
    .B(_1772_),
    .Y(_1847_));
 sg13g2_o21ai_1 _5957_ (.B1(_1776_),
    .Y(_1848_),
    .A1(_1832_),
    .A2(_1833_));
 sg13g2_o21ai_1 _5958_ (.B1(net322),
    .Y(_1849_),
    .A1(_1847_),
    .A2(_1848_));
 sg13g2_buf_1 _5959_ (.A(_1849_),
    .X(_1850_));
 sg13g2_a21oi_1 _5960_ (.A1(_1847_),
    .A2(_1848_),
    .Y(_1851_),
    .B1(_1842_));
 sg13g2_nor3_1 _5961_ (.A(_1748_),
    .B(_1749_),
    .C(_1754_),
    .Y(_1852_));
 sg13g2_o21ai_1 _5962_ (.B1(net224),
    .Y(_1853_),
    .A1(_1852_),
    .A2(_1842_));
 sg13g2_a21oi_1 _5963_ (.A1(_1850_),
    .A2(_1851_),
    .Y(_1854_),
    .B1(_1853_));
 sg13g2_or2_1 _5964_ (.X(_1855_),
    .B(_1854_),
    .A(net319));
 sg13g2_or4_1 _5965_ (.A(_1686_),
    .B(_1817_),
    .C(_1846_),
    .D(_1855_),
    .X(_1856_));
 sg13g2_nor2b_1 _5966_ (.A(_1510_),
    .B_N(net337),
    .Y(_1857_));
 sg13g2_a22oi_1 _5967_ (.Y(_1858_),
    .B1(_1857_),
    .B2(_1457_),
    .A2(_1452_),
    .A1(_1376_));
 sg13g2_nand2_1 _5968_ (.Y(_1859_),
    .A(net309),
    .B(net331));
 sg13g2_nand3_1 _5969_ (.B(_1744_),
    .C(_1859_),
    .A(_1511_),
    .Y(_1860_));
 sg13g2_nor2_1 _5970_ (.A(_1480_),
    .B(_1367_),
    .Y(_1861_));
 sg13g2_nand2_1 _5971_ (.Y(_1862_),
    .A(_0103_),
    .B(_1861_));
 sg13g2_buf_2 _5972_ (.A(_1862_),
    .X(_1863_));
 sg13g2_a21o_1 _5973_ (.A2(_1860_),
    .A1(_1858_),
    .B1(_1863_),
    .X(_1864_));
 sg13g2_nor2b_1 _5974_ (.A(_0026_),
    .B_N(_1510_),
    .Y(_1865_));
 sg13g2_nor2_2 _5975_ (.A(_1451_),
    .B(net335),
    .Y(_1866_));
 sg13g2_nand4_1 _5976_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29] ),
    .C(_1865_),
    .A(_1682_),
    .Y(_1867_),
    .D(_1866_));
 sg13g2_nor2_2 _5977_ (.A(_1371_),
    .B(net336),
    .Y(_1868_));
 sg13g2_nand3_1 _5978_ (.B(_1454_),
    .C(_1868_),
    .A(_1445_),
    .Y(_1869_));
 sg13g2_and2_1 _5979_ (.A(_1867_),
    .B(_1869_),
    .X(_1870_));
 sg13g2_buf_1 _5980_ (.A(_1870_),
    .X(_1871_));
 sg13g2_and2_1 _5981_ (.A(_1445_),
    .B(_1868_),
    .X(_1872_));
 sg13g2_and4_1 _5982_ (.A(_1456_),
    .B(_1454_),
    .C(_1868_),
    .D(_1759_),
    .X(_1873_));
 sg13g2_a21oi_1 _5983_ (.A1(_1373_),
    .A2(_1872_),
    .Y(_1874_),
    .B1(_1873_));
 sg13g2_and4_1 _5984_ (.A(_0103_),
    .B(_1452_),
    .C(_1454_),
    .D(_1861_),
    .X(_1875_));
 sg13g2_a21oi_1 _5985_ (.A1(_1519_),
    .A2(_1863_),
    .Y(_1876_),
    .B1(_1875_));
 sg13g2_and4_1 _5986_ (.A(_1864_),
    .B(_1871_),
    .C(_1874_),
    .D(_1876_),
    .X(_1877_));
 sg13g2_buf_2 _5987_ (.A(_1877_),
    .X(_1878_));
 sg13g2_nor2_1 _5988_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .B(_1878_),
    .Y(_1879_));
 sg13g2_o21ai_1 _5989_ (.B1(_1863_),
    .Y(_1880_),
    .A1(net248),
    .A2(_1450_));
 sg13g2_and2_1 _5990_ (.A(_1459_),
    .B(_1880_),
    .X(_1881_));
 sg13g2_buf_1 _5991_ (.A(_1881_),
    .X(_1882_));
 sg13g2_nor2b_1 _5992_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0] ),
    .B_N(net319),
    .Y(_1883_));
 sg13g2_nor3_1 _5993_ (.A(_1879_),
    .B(_1882_),
    .C(_1883_),
    .Y(_1884_));
 sg13g2_a22oi_1 _5994_ (.Y(_1885_),
    .B1(_1721_),
    .B2(_1741_),
    .A2(_1728_),
    .A1(net306));
 sg13g2_a21oi_1 _5995_ (.A1(_1738_),
    .A2(_1885_),
    .Y(_1886_),
    .B1(_1368_));
 sg13g2_nand4_1 _5996_ (.B(_1844_),
    .C(_1845_),
    .A(_1838_),
    .Y(_1887_),
    .D(_1886_));
 sg13g2_nand2_1 _5997_ (.Y(_1888_),
    .A(_1854_),
    .B(_1886_));
 sg13g2_and3_1 _5998_ (.X(_1889_),
    .A(_1884_),
    .B(_1887_),
    .C(_1888_));
 sg13g2_buf_2 _5999_ (.A(_1430_),
    .X(_1890_));
 sg13g2_buf_1 _6000_ (.A(net304),
    .X(_1891_));
 sg13g2_nand2_1 _6001_ (.Y(_1892_),
    .A(net311),
    .B(_1422_));
 sg13g2_nor2_1 _6002_ (.A(net333),
    .B(_1892_),
    .Y(_1893_));
 sg13g2_buf_2 _6003_ (.A(_1893_),
    .X(_1894_));
 sg13g2_buf_1 _6004_ (.A(_0027_),
    .X(_1895_));
 sg13g2_buf_1 _6005_ (.A(_1895_),
    .X(_1896_));
 sg13g2_nand2b_1 _6006_ (.Y(_1897_),
    .B(_1421_),
    .A_N(_1425_));
 sg13g2_buf_1 _6007_ (.A(_1897_),
    .X(_1898_));
 sg13g2_nor2_1 _6008_ (.A(net303),
    .B(_1898_),
    .Y(_1899_));
 sg13g2_buf_2 _6009_ (.A(_1899_),
    .X(_1900_));
 sg13g2_a22oi_1 _6010_ (.Y(_1901_),
    .B1(_1900_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ),
    .A2(_1894_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0] ));
 sg13g2_nor2_1 _6011_ (.A(_1428_),
    .B(net286),
    .Y(_1902_));
 sg13g2_inv_1 _6012_ (.Y(_1903_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0] ));
 sg13g2_nand2_1 _6013_ (.Y(_1904_),
    .A(net286),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0] ));
 sg13g2_o21ai_1 _6014_ (.B1(_1904_),
    .Y(_1905_),
    .A1(net264),
    .A2(_1903_));
 sg13g2_a22oi_1 _6015_ (.Y(_1906_),
    .B1(_1905_),
    .B2(_1428_),
    .A2(_1902_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0] ));
 sg13g2_nand3b_1 _6016_ (.B(net282),
    .C(_1439_),
    .Y(_1907_),
    .A_N(_1906_));
 sg13g2_o21ai_1 _6017_ (.B1(_1907_),
    .Y(_1908_),
    .A1(net282),
    .A2(_1901_));
 sg13g2_nand2b_1 _6018_ (.Y(_1909_),
    .B(_1430_),
    .A_N(net303));
 sg13g2_nor2b_1 _6019_ (.A(net310),
    .B_N(net311),
    .Y(_1910_));
 sg13g2_nor2b_1 _6020_ (.A(net311),
    .B_N(_1435_),
    .Y(_1911_));
 sg13g2_a22oi_1 _6021_ (.Y(_1912_),
    .B1(_1911_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ),
    .A2(_1910_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ));
 sg13g2_buf_1 _6022_ (.A(_1435_),
    .X(_1913_));
 sg13g2_buf_1 _6023_ (.A(net281),
    .X(_1914_));
 sg13g2_buf_1 _6024_ (.A(net285),
    .X(_1915_));
 sg13g2_nand2_1 _6025_ (.Y(_1916_),
    .A(net260),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ));
 sg13g2_nand3_1 _6026_ (.B(_1428_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ),
    .A(net304),
    .Y(_1917_));
 sg13g2_o21ai_1 _6027_ (.B1(_1917_),
    .Y(_1918_),
    .A1(net282),
    .A2(_1916_));
 sg13g2_nand3_1 _6028_ (.B(_1439_),
    .C(_1918_),
    .A(net261),
    .Y(_1919_));
 sg13g2_o21ai_1 _6029_ (.B1(_1919_),
    .Y(_1920_),
    .A1(_1909_),
    .A2(_1912_));
 sg13g2_buf_1 _6030_ (.A(net333),
    .X(_1921_));
 sg13g2_inv_1 _6031_ (.Y(_1922_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0] ));
 sg13g2_nor4_1 _6032_ (.A(net283),
    .B(net302),
    .C(_1922_),
    .D(_1892_),
    .Y(_1923_));
 sg13g2_buf_1 _6033_ (.A(net303),
    .X(_1924_));
 sg13g2_inv_1 _6034_ (.Y(_1925_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0] ));
 sg13g2_nor4_1 _6035_ (.A(net281),
    .B(net280),
    .C(_1925_),
    .D(_1898_),
    .Y(_1926_));
 sg13g2_o21ai_1 _6036_ (.B1(_1891_),
    .Y(_1927_),
    .A1(_1923_),
    .A2(_1926_));
 sg13g2_and2_1 _6037_ (.A(net310),
    .B(_1430_),
    .X(_1928_));
 sg13g2_buf_2 _6038_ (.A(_1928_),
    .X(_1929_));
 sg13g2_nor3_1 _6039_ (.A(net311),
    .B(net312),
    .C(_1895_),
    .Y(_1930_));
 sg13g2_and2_1 _6040_ (.A(_1929_),
    .B(_1930_),
    .X(_1931_));
 sg13g2_buf_1 _6041_ (.A(_1931_),
    .X(_1932_));
 sg13g2_nand2b_1 _6042_ (.Y(_1933_),
    .B(_1426_),
    .A_N(net312));
 sg13g2_buf_1 _6043_ (.A(_1933_),
    .X(_1934_));
 sg13g2_nor2_1 _6044_ (.A(net280),
    .B(_1934_),
    .Y(_1935_));
 sg13g2_mux4_1 _6045_ (.S0(_1890_),
    .A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0] ),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0] ),
    .A3(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0] ),
    .S1(_1913_),
    .X(_1936_));
 sg13g2_a22oi_1 _6046_ (.Y(_1937_),
    .B1(_1935_),
    .B2(_1936_),
    .A2(_1932_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0] ));
 sg13g2_nand2_1 _6047_ (.Y(_1938_),
    .A(_1927_),
    .B(_1937_));
 sg13g2_a221oi_1 _6048_ (.B2(_1424_),
    .C1(_1938_),
    .B1(_1920_),
    .A1(net283),
    .Y(_1939_),
    .A2(_1908_));
 sg13g2_nor2_1 _6049_ (.A(_1434_),
    .B(_1430_),
    .Y(_1940_));
 sg13g2_buf_2 _6050_ (.A(_1940_),
    .X(_1941_));
 sg13g2_nor2b_1 _6051_ (.A(net311),
    .B_N(net312),
    .Y(_1942_));
 sg13g2_a22oi_1 _6052_ (.Y(_1943_),
    .B1(_1902_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0] ),
    .A2(_1942_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ));
 sg13g2_nor2_1 _6053_ (.A(net280),
    .B(_1892_),
    .Y(_1944_));
 sg13g2_nand2_1 _6054_ (.Y(_1945_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0] ),
    .B(_1944_));
 sg13g2_o21ai_1 _6055_ (.B1(_1945_),
    .Y(_1946_),
    .A1(net302),
    .A2(_1943_));
 sg13g2_nor3_1 _6056_ (.A(net310),
    .B(_1427_),
    .C(net286),
    .Y(_1947_));
 sg13g2_nand2_1 _6057_ (.Y(_1948_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0] ),
    .B(_1947_));
 sg13g2_and2_1 _6058_ (.A(_1425_),
    .B(_1421_),
    .X(_1949_));
 sg13g2_buf_2 _6059_ (.A(_1949_),
    .X(_1950_));
 sg13g2_nand3_1 _6060_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0] ),
    .C(_1950_),
    .A(net281),
    .Y(_1951_));
 sg13g2_a21oi_1 _6061_ (.A1(_1948_),
    .A2(_1951_),
    .Y(_1952_),
    .B1(_1909_));
 sg13g2_a21o_1 _6062_ (.A2(_1946_),
    .A1(_1941_),
    .B1(_1952_),
    .X(_1953_));
 sg13g2_nor2_2 _6063_ (.A(net333),
    .B(_1934_),
    .Y(_1954_));
 sg13g2_nor3_2 _6064_ (.A(net311),
    .B(net312),
    .C(net333),
    .Y(_1955_));
 sg13g2_a22oi_1 _6065_ (.Y(_1956_),
    .B1(_1955_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0] ),
    .A2(_1954_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0] ));
 sg13g2_nand3_1 _6066_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0] ),
    .C(_1954_),
    .A(net284),
    .Y(_1957_));
 sg13g2_o21ai_1 _6067_ (.B1(_1957_),
    .Y(_1958_),
    .A1(net284),
    .A2(_1956_));
 sg13g2_and2_1 _6068_ (.A(net261),
    .B(_1958_),
    .X(_1959_));
 sg13g2_inv_1 _6069_ (.Y(_1960_),
    .A(_1895_));
 sg13g2_a22oi_1 _6070_ (.Y(_1961_),
    .B1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0] ),
    .B2(_1439_),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0] ),
    .A1(_1960_));
 sg13g2_nor2_2 _6071_ (.A(net311),
    .B(net312),
    .Y(_1962_));
 sg13g2_nor2_1 _6072_ (.A(net283),
    .B(net304),
    .Y(_1963_));
 sg13g2_nand2_1 _6073_ (.Y(_1964_),
    .A(_1962_),
    .B(_1963_));
 sg13g2_nor2_1 _6074_ (.A(net281),
    .B(net284),
    .Y(_1965_));
 sg13g2_nand3_1 _6075_ (.B(_1894_),
    .C(_1965_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0] ),
    .Y(_1966_));
 sg13g2_o21ai_1 _6076_ (.B1(_1966_),
    .Y(_1967_),
    .A1(_1961_),
    .A2(_1964_));
 sg13g2_nor3_1 _6077_ (.A(net283),
    .B(net302),
    .C(_1898_),
    .Y(_1968_));
 sg13g2_mux2_1 _6078_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0] ),
    .S(net285),
    .X(_1969_));
 sg13g2_nand3_1 _6079_ (.B(net264),
    .C(_1969_),
    .A(net281),
    .Y(_1970_));
 sg13g2_nand2_1 _6080_ (.Y(_1971_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0] ),
    .B(_1947_));
 sg13g2_nand2_1 _6081_ (.Y(_1972_),
    .A(_1970_),
    .B(_1971_));
 sg13g2_a22oi_1 _6082_ (.Y(_1973_),
    .B1(_1972_),
    .B2(_1960_),
    .A2(_1968_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0] ));
 sg13g2_nor2_1 _6083_ (.A(net282),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_nor4_1 _6084_ (.A(_1953_),
    .B(_1959_),
    .C(_1967_),
    .D(_1974_),
    .Y(_1975_));
 sg13g2_a21oi_1 _6085_ (.A1(_1962_),
    .A2(_1941_),
    .Y(_1976_),
    .B1(net333));
 sg13g2_nand2b_1 _6086_ (.Y(_1977_),
    .B(net303),
    .A_N(_1976_));
 sg13g2_nand3_1 _6087_ (.B(_1880_),
    .C(_1977_),
    .A(_1459_),
    .Y(_1978_));
 sg13g2_buf_1 _6088_ (.A(_1978_),
    .X(_1979_));
 sg13g2_a21oi_1 _6089_ (.A1(_1939_),
    .A2(_1975_),
    .Y(_1980_),
    .B1(_1979_));
 sg13g2_mux2_1 _6090_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .A1(_1980_),
    .S(_1878_),
    .X(_1981_));
 sg13g2_a21oi_2 _6091_ (.B1(_1981_),
    .Y(_1982_),
    .A2(_1889_),
    .A1(_1856_));
 sg13g2_nor2_1 _6092_ (.A(_1444_),
    .B(_1446_),
    .Y(_1983_));
 sg13g2_nand4_1 _6093_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30] ),
    .C(_1868_),
    .A(_1456_),
    .Y(_1984_),
    .D(_1983_));
 sg13g2_buf_1 _6094_ (.A(_1984_),
    .X(_1985_));
 sg13g2_buf_1 _6095_ (.A(_1985_),
    .X(_1986_));
 sg13g2_nor3_1 _6096_ (.A(net335),
    .B(_1372_),
    .C(net336),
    .Y(_1987_));
 sg13g2_nor3_1 _6097_ (.A(_1450_),
    .B(_1455_),
    .C(_1987_),
    .Y(_1988_));
 sg13g2_nor2_1 _6098_ (.A(_1863_),
    .B(_1988_),
    .Y(_1989_));
 sg13g2_nor2_1 _6099_ (.A(_1456_),
    .B(_1518_),
    .Y(_1990_));
 sg13g2_nand2_1 _6100_ (.Y(_1991_),
    .A(_1863_),
    .B(_1990_));
 sg13g2_nor2b_1 _6101_ (.A(_1989_),
    .B_N(_1991_),
    .Y(_1992_));
 sg13g2_buf_2 _6102_ (.A(_1992_),
    .X(_1993_));
 sg13g2_buf_1 _6103_ (.A(_1993_),
    .X(_1994_));
 sg13g2_nand2_1 _6104_ (.Y(_1995_),
    .A(net243),
    .B(net97));
 sg13g2_nand4_1 _6105_ (.B(_1871_),
    .C(_1874_),
    .A(_1864_),
    .Y(_1996_),
    .D(_1876_));
 sg13g2_buf_2 _6106_ (.A(_1996_),
    .X(_1997_));
 sg13g2_inv_1 _6107_ (.Y(_1998_),
    .A(_1879_));
 sg13g2_o21ai_1 _6108_ (.B1(_1998_),
    .Y(_1999_),
    .A1(_1997_),
    .A2(_1980_));
 sg13g2_o21ai_1 _6109_ (.B1(_1991_),
    .Y(_2000_),
    .A1(_1863_),
    .A2(_1988_));
 sg13g2_buf_1 _6110_ (.A(_2000_),
    .X(_2001_));
 sg13g2_nor2_1 _6111_ (.A(_1985_),
    .B(net173),
    .Y(_2002_));
 sg13g2_nor2_1 _6112_ (.A(_1985_),
    .B(_1993_),
    .Y(_2003_));
 sg13g2_buf_1 _6113_ (.A(_1418_),
    .X(_2004_));
 sg13g2_and2_1 _6114_ (.A(net334),
    .B(_1395_),
    .X(_2005_));
 sg13g2_buf_1 _6115_ (.A(_2005_),
    .X(_2006_));
 sg13g2_nor2_2 _6116_ (.A(net334),
    .B(net317),
    .Y(_2007_));
 sg13g2_a22oi_1 _6117_ (.Y(_2008_),
    .B1(_2007_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0] ),
    .A2(_2006_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0] ));
 sg13g2_buf_1 _6118_ (.A(_0038_),
    .X(_2009_));
 sg13g2_buf_1 _6119_ (.A(_2009_),
    .X(_2010_));
 sg13g2_mux2_1 _6120_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ),
    .S(_1396_),
    .X(_2011_));
 sg13g2_a22oi_1 _6121_ (.Y(_2012_),
    .B1(_2011_),
    .B2(net316),
    .A2(_2007_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0] ));
 sg13g2_or2_1 _6122_ (.X(_2013_),
    .B(_2012_),
    .A(net300));
 sg13g2_o21ai_1 _6123_ (.B1(_2013_),
    .Y(_2014_),
    .A1(net301),
    .A2(_2008_));
 sg13g2_inv_1 _6124_ (.Y(_2015_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0] ));
 sg13g2_nor2_1 _6125_ (.A(net288),
    .B(_2015_),
    .Y(_2016_));
 sg13g2_nor3_1 _6126_ (.A(net316),
    .B(net317),
    .C(_2009_),
    .Y(_2017_));
 sg13g2_buf_1 _6127_ (.A(net314),
    .X(_2018_));
 sg13g2_buf_1 _6128_ (.A(net279),
    .X(_2019_));
 sg13g2_a221oi_1 _6129_ (.B2(_2017_),
    .C1(net259),
    .B1(_2016_),
    .A1(_1413_),
    .Y(_2020_),
    .A2(_2014_));
 sg13g2_inv_2 _6130_ (.Y(_2021_),
    .A(_2009_));
 sg13g2_a221oi_1 _6131_ (.B2(net313),
    .C1(net317),
    .B1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0] ),
    .A1(_2021_),
    .Y(_2022_),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0] ));
 sg13g2_a221oi_1 _6132_ (.B2(net313),
    .C1(_1397_),
    .B1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0] ),
    .A1(_2021_),
    .Y(_2023_),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0] ));
 sg13g2_nor3_1 _6133_ (.A(_1407_),
    .B(_2022_),
    .C(_2023_),
    .Y(_2024_));
 sg13g2_nor2b_1 _6134_ (.A(net334),
    .B_N(_1395_),
    .Y(_2025_));
 sg13g2_buf_2 _6135_ (.A(_2025_),
    .X(_2026_));
 sg13g2_and3_1 _6136_ (.X(_2027_),
    .A(net313),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ),
    .C(_2026_));
 sg13g2_o21ai_1 _6137_ (.B1(_1412_),
    .Y(_2028_),
    .A1(_2024_),
    .A2(_2027_));
 sg13g2_nor2b_1 _6138_ (.A(_1410_),
    .B_N(net334),
    .Y(_2029_));
 sg13g2_buf_1 _6139_ (.A(_2029_),
    .X(_2030_));
 sg13g2_nor2b_1 _6140_ (.A(_2009_),
    .B_N(_1395_),
    .Y(_2031_));
 sg13g2_buf_2 _6141_ (.A(_2031_),
    .X(_2032_));
 sg13g2_nand3_1 _6142_ (.B(_2030_),
    .C(_2032_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0] ),
    .Y(_2033_));
 sg13g2_nor2_1 _6143_ (.A(_1395_),
    .B(_1418_),
    .Y(_2034_));
 sg13g2_buf_2 _6144_ (.A(_2034_),
    .X(_2035_));
 sg13g2_nor2_2 _6145_ (.A(_1410_),
    .B(net334),
    .Y(_2036_));
 sg13g2_nand3_1 _6146_ (.B(_2035_),
    .C(_2036_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0] ),
    .Y(_2037_));
 sg13g2_nor2_1 _6147_ (.A(net317),
    .B(_2009_),
    .Y(_2038_));
 sg13g2_buf_2 _6148_ (.A(_2038_),
    .X(_2039_));
 sg13g2_nor2b_1 _6149_ (.A(_1405_),
    .B_N(_1410_),
    .Y(_2040_));
 sg13g2_buf_1 _6150_ (.A(_2040_),
    .X(_2041_));
 sg13g2_nand3_1 _6151_ (.B(_2039_),
    .C(_2041_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0] ),
    .Y(_2042_));
 sg13g2_nand3_1 _6152_ (.B(_2037_),
    .C(_2042_),
    .A(_2033_),
    .Y(_2043_));
 sg13g2_nor2b_1 _6153_ (.A(net317),
    .B_N(net334),
    .Y(_2044_));
 sg13g2_a22oi_1 _6154_ (.Y(_2045_),
    .B1(_2044_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0] ),
    .A2(_2026_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0] ));
 sg13g2_nor3_1 _6155_ (.A(net315),
    .B(net301),
    .C(_2045_),
    .Y(_2046_));
 sg13g2_nor2_1 _6156_ (.A(_2043_),
    .B(_2046_),
    .Y(_2047_));
 sg13g2_and3_1 _6157_ (.X(_2048_),
    .A(net259),
    .B(_2028_),
    .C(_2047_));
 sg13g2_a22oi_1 _6158_ (.Y(_2049_),
    .B1(_2044_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0] ),
    .A2(_2026_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ));
 sg13g2_or4_1 _6159_ (.A(net314),
    .B(net315),
    .C(net301),
    .D(_2049_),
    .X(_2050_));
 sg13g2_nor2_1 _6160_ (.A(_1414_),
    .B(_1418_),
    .Y(_2051_));
 sg13g2_nand4_1 _6161_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0] ),
    .C(_2026_),
    .A(net315),
    .Y(_2052_),
    .D(_2051_));
 sg13g2_nor2b_1 _6162_ (.A(net315),
    .B_N(_1414_),
    .Y(_2053_));
 sg13g2_nand3_1 _6163_ (.B(_2017_),
    .C(_2053_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0] ),
    .Y(_2054_));
 sg13g2_mux2_1 _6164_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ),
    .S(_1414_),
    .X(_2055_));
 sg13g2_and3_1 _6165_ (.X(_2056_),
    .A(_2021_),
    .B(_2026_),
    .C(_2055_));
 sg13g2_nor2_1 _6166_ (.A(_1414_),
    .B(_1410_),
    .Y(_2057_));
 sg13g2_and3_1 _6167_ (.X(_2058_),
    .A(net313),
    .B(_2006_),
    .C(_2057_));
 sg13g2_buf_1 _6168_ (.A(_2058_),
    .X(_2059_));
 sg13g2_a22oi_1 _6169_ (.Y(_2060_),
    .B1(_2059_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0] ),
    .A2(_2056_),
    .A1(net315));
 sg13g2_nand4_1 _6170_ (.B(_2052_),
    .C(_2054_),
    .A(_2050_),
    .Y(_2061_),
    .D(_2060_));
 sg13g2_nor2b_1 _6171_ (.A(net314),
    .B_N(net316),
    .Y(_2062_));
 sg13g2_nor2b_1 _6172_ (.A(net334),
    .B_N(_1414_),
    .Y(_2063_));
 sg13g2_buf_1 _6173_ (.A(_2063_),
    .X(_2064_));
 sg13g2_a22oi_1 _6174_ (.Y(_2065_),
    .B1(_2064_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0] ),
    .A2(_2062_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0] ));
 sg13g2_nand2_1 _6175_ (.Y(_2066_),
    .A(net288),
    .B(_2035_));
 sg13g2_buf_1 _6176_ (.A(_2039_),
    .X(_2067_));
 sg13g2_inv_1 _6177_ (.Y(_2068_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0] ));
 sg13g2_nand2_1 _6178_ (.Y(_2069_),
    .A(net314),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0] ));
 sg13g2_o21ai_1 _6179_ (.B1(_2069_),
    .Y(_2070_),
    .A1(net314),
    .A2(_2068_));
 sg13g2_nand3_1 _6180_ (.B(net242),
    .C(_2070_),
    .A(_2030_),
    .Y(_2071_));
 sg13g2_o21ai_1 _6181_ (.B1(_2071_),
    .Y(_2072_),
    .A1(_2065_),
    .A2(_2066_));
 sg13g2_nand2_1 _6182_ (.Y(_2073_),
    .A(_1445_),
    .B(_1857_));
 sg13g2_o21ai_1 _6183_ (.B1(_1869_),
    .Y(_2074_),
    .A1(net324),
    .A2(_2073_));
 sg13g2_o21ai_1 _6184_ (.B1(_1863_),
    .Y(_2075_),
    .A1(_1519_),
    .A2(_1990_));
 sg13g2_nand2b_1 _6185_ (.Y(_2076_),
    .B(_2075_),
    .A_N(_2074_));
 sg13g2_buf_2 _6186_ (.A(_2076_),
    .X(_2077_));
 sg13g2_buf_1 _6187_ (.A(_1406_),
    .X(_2078_));
 sg13g2_nand2b_1 _6188_ (.Y(_2079_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ),
    .A_N(_2009_));
 sg13g2_nand3b_1 _6189_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ),
    .C(net316),
    .Y(_2080_),
    .A_N(_1418_));
 sg13g2_o21ai_1 _6190_ (.B1(_2080_),
    .Y(_2081_),
    .A1(net278),
    .A2(_2079_));
 sg13g2_mux2_1 _6191_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0] ),
    .S(net316),
    .X(_2082_));
 sg13g2_nor2_1 _6192_ (.A(net314),
    .B(net300),
    .Y(_2083_));
 sg13g2_a22oi_1 _6193_ (.Y(_2084_),
    .B1(_2082_),
    .B2(_2083_),
    .A2(_2081_),
    .A1(net279));
 sg13g2_nand2b_1 _6194_ (.Y(_2085_),
    .B(net317),
    .A_N(net315));
 sg13g2_buf_1 _6195_ (.A(_2085_),
    .X(_2086_));
 sg13g2_nor2_1 _6196_ (.A(_2084_),
    .B(_2086_),
    .Y(_2087_));
 sg13g2_nor4_1 _6197_ (.A(_2061_),
    .B(_2072_),
    .C(_2077_),
    .D(_2087_),
    .Y(_2088_));
 sg13g2_o21ai_1 _6198_ (.B1(_2088_),
    .Y(_2089_),
    .A1(_2020_),
    .A2(_2048_));
 sg13g2_buf_1 _6199_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .X(_2090_));
 sg13g2_nand2b_1 _6200_ (.Y(_2091_),
    .B(_2077_),
    .A_N(_2090_));
 sg13g2_nand2_1 _6201_ (.Y(_2092_),
    .A(_2089_),
    .B(_2091_));
 sg13g2_buf_2 _6202_ (.A(_2092_),
    .X(_2093_));
 sg13g2_and4_1 _6203_ (.A(_1456_),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30] ),
    .C(_1868_),
    .D(_1983_),
    .X(_2094_));
 sg13g2_buf_2 _6204_ (.A(_2094_),
    .X(_2095_));
 sg13g2_nor2_1 _6205_ (.A(_2095_),
    .B(_1993_),
    .Y(_2096_));
 sg13g2_nor2b_1 _6206_ (.A(_2093_),
    .B_N(_2096_),
    .Y(_2097_));
 sg13g2_a221oi_1 _6207_ (.B2(_2093_),
    .C1(_2097_),
    .B1(_2003_),
    .A1(_1999_),
    .Y(_2098_),
    .A2(_2002_));
 sg13g2_o21ai_1 _6208_ (.B1(_2098_),
    .Y(_2099_),
    .A1(_1982_),
    .A2(_1995_));
 sg13g2_a21o_1 _6209_ (.A2(_1889_),
    .A1(_1856_),
    .B1(_1981_),
    .X(_2100_));
 sg13g2_nand2_1 _6210_ (.Y(_2101_),
    .A(_1456_),
    .B(_1519_));
 sg13g2_and2_1 _6211_ (.A(_1864_),
    .B(_1871_),
    .X(_2102_));
 sg13g2_inv_1 _6212_ (.Y(_2103_),
    .A(_1454_));
 sg13g2_nand2_1 _6213_ (.Y(_2104_),
    .A(_1456_),
    .B(_1868_));
 sg13g2_a21oi_1 _6214_ (.A1(_1444_),
    .A2(_2103_),
    .Y(_2105_),
    .B1(_2104_));
 sg13g2_nand2_1 _6215_ (.Y(_2106_),
    .A(_2105_),
    .B(_1759_));
 sg13g2_and3_1 _6216_ (.X(_2107_),
    .A(_2101_),
    .B(_2102_),
    .C(_2106_));
 sg13g2_buf_1 _6217_ (.A(_2107_),
    .X(_2108_));
 sg13g2_buf_1 _6218_ (.A(_2108_),
    .X(_2109_));
 sg13g2_nor2_1 _6219_ (.A(_1993_),
    .B(net86),
    .Y(_2110_));
 sg13g2_nor2_1 _6220_ (.A(net173),
    .B(_2108_),
    .Y(_2111_));
 sg13g2_nor2b_1 _6221_ (.A(_2093_),
    .B_N(_2111_),
    .Y(_2112_));
 sg13g2_a21o_1 _6222_ (.A2(_2110_),
    .A1(_2100_),
    .B1(_2112_),
    .X(_2113_));
 sg13g2_buf_1 _6223_ (.A(_2113_),
    .X(_2114_));
 sg13g2_nand2_1 _6224_ (.Y(_2115_),
    .A(_2099_),
    .B(_2114_));
 sg13g2_inv_1 _6225_ (.Y(_2116_),
    .A(_1444_));
 sg13g2_o21ai_1 _6226_ (.B1(_1452_),
    .Y(_2117_),
    .A1(_2116_),
    .A2(net324));
 sg13g2_nor2_1 _6227_ (.A(_1374_),
    .B(_2117_),
    .Y(_2118_));
 sg13g2_nor2_1 _6228_ (.A(_1717_),
    .B(_1449_),
    .Y(_2119_));
 sg13g2_buf_1 _6229_ (.A(net308),
    .X(_2120_));
 sg13g2_inv_1 _6230_ (.Y(_2121_),
    .A(_0103_));
 sg13g2_nor3_1 _6231_ (.A(net277),
    .B(net290),
    .C(_2121_),
    .Y(_2122_));
 sg13g2_a21oi_1 _6232_ (.A1(_2119_),
    .A2(_2122_),
    .Y(_2123_),
    .B1(net223));
 sg13g2_nor3_1 _6233_ (.A(_1446_),
    .B(_1717_),
    .C(_1691_),
    .Y(_2124_));
 sg13g2_nor2_1 _6234_ (.A(_1460_),
    .B(_2124_),
    .Y(_2125_));
 sg13g2_o21ai_1 _6235_ (.B1(_1872_),
    .Y(_2126_),
    .A1(_1373_),
    .A2(_1454_));
 sg13g2_nor2_1 _6236_ (.A(net309),
    .B(net331),
    .Y(_2127_));
 sg13g2_buf_2 _6237_ (.A(_2127_),
    .X(_2128_));
 sg13g2_nor2b_1 _6238_ (.A(_2128_),
    .B_N(_1865_),
    .Y(_2129_));
 sg13g2_a22oi_1 _6239_ (.Y(_2130_),
    .B1(_2129_),
    .B2(_1680_),
    .A2(_1863_),
    .A1(_2119_));
 sg13g2_and3_1 _6240_ (.X(_2131_),
    .A(_2125_),
    .B(_2126_),
    .C(_2130_));
 sg13g2_buf_1 _6241_ (.A(_2131_),
    .X(_2132_));
 sg13g2_a21oi_1 _6242_ (.A1(net324),
    .A2(_1453_),
    .Y(_2133_),
    .B1(_2073_));
 sg13g2_and4_1 _6243_ (.A(_2116_),
    .B(net336),
    .C(_1744_),
    .D(_1859_),
    .X(_2134_));
 sg13g2_buf_1 _6244_ (.A(_2134_),
    .X(_2135_));
 sg13g2_nor3_1 _6245_ (.A(_1521_),
    .B(_2133_),
    .C(_2135_),
    .Y(_2136_));
 sg13g2_and4_1 _6246_ (.A(_1867_),
    .B(_2123_),
    .C(_2132_),
    .D(_2136_),
    .X(_2137_));
 sg13g2_buf_1 _6247_ (.A(_2137_),
    .X(_2138_));
 sg13g2_nand2b_1 _6248_ (.Y(_2139_),
    .B(_2138_),
    .A_N(_2118_));
 sg13g2_nand2b_1 _6249_ (.Y(_2140_),
    .B(_2105_),
    .A_N(_1859_));
 sg13g2_and2_1 _6250_ (.A(_2138_),
    .B(_2140_),
    .X(_2141_));
 sg13g2_buf_1 _6251_ (.A(_2141_),
    .X(_2142_));
 sg13g2_mux2_1 _6252_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ),
    .A1(_2095_),
    .S(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb ),
    .X(_2143_));
 sg13g2_buf_2 _6253_ (.A(_2143_),
    .X(_2144_));
 sg13g2_nor2_1 _6254_ (.A(_2138_),
    .B(_2144_),
    .Y(_2145_));
 sg13g2_nor2_1 _6255_ (.A(_2142_),
    .B(_2145_),
    .Y(_2146_));
 sg13g2_nand4_1 _6256_ (.B(_2123_),
    .C(_2132_),
    .A(_1867_),
    .Y(_2147_),
    .D(_2136_));
 sg13g2_buf_1 _6257_ (.A(_2147_),
    .X(_2148_));
 sg13g2_nand2_1 _6258_ (.Y(_2149_),
    .A(_2148_),
    .B(_2144_));
 sg13g2_xnor2_1 _6259_ (.Y(_2150_),
    .A(_2099_),
    .B(_2114_));
 sg13g2_mux2_1 _6260_ (.A0(_2146_),
    .A1(_2149_),
    .S(_2150_),
    .X(_2151_));
 sg13g2_o21ai_1 _6261_ (.B1(_2151_),
    .Y(_2152_),
    .A1(_2115_),
    .A2(_2139_));
 sg13g2_buf_1 _6262_ (.A(_2152_),
    .X(_2153_));
 sg13g2_nand2_1 _6263_ (.Y(_2154_),
    .A(net175),
    .B(_1982_));
 sg13g2_o21ai_1 _6264_ (.B1(_2154_),
    .Y(_2155_),
    .A1(net175),
    .A2(_2153_));
 sg13g2_nand2_1 _6265_ (.Y(_2156_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28] ),
    .B(net74));
 sg13g2_o21ai_1 _6266_ (.B1(_2156_),
    .Y(_1234_),
    .A1(net75),
    .A2(_2155_));
 sg13g2_nor2_1 _6267_ (.A(_1997_),
    .B(_1979_),
    .Y(_2157_));
 sg13g2_a221oi_1 _6268_ (.B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ),
    .C1(net304),
    .B1(_1900_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ),
    .Y(_2158_),
    .A2(_1894_));
 sg13g2_a21oi_1 _6269_ (.A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ),
    .A2(_1894_),
    .Y(_2159_),
    .B1(_1431_));
 sg13g2_nor3_1 _6270_ (.A(net281),
    .B(_2158_),
    .C(_2159_),
    .Y(_2160_));
 sg13g2_nor2b_1 _6271_ (.A(_1896_),
    .B_N(net286),
    .Y(_2161_));
 sg13g2_mux2_1 _6272_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ),
    .S(net285),
    .X(_2162_));
 sg13g2_a22oi_1 _6273_ (.Y(_2163_),
    .B1(_2161_),
    .B2(_2162_),
    .A2(_1955_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ));
 sg13g2_mux2_1 _6274_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ),
    .S(net312),
    .X(_2164_));
 sg13g2_a21oi_1 _6275_ (.A1(net312),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ),
    .Y(_2165_),
    .B1(net285));
 sg13g2_nor2_1 _6276_ (.A(net302),
    .B(_2165_),
    .Y(_2166_));
 sg13g2_o21ai_1 _6277_ (.B1(_2166_),
    .Y(_2167_),
    .A1(_1428_),
    .A2(_2164_));
 sg13g2_nand2_1 _6278_ (.Y(_2168_),
    .A(net310),
    .B(net284));
 sg13g2_a21oi_1 _6279_ (.A1(_2163_),
    .A2(_2167_),
    .Y(_2169_),
    .B1(_2168_));
 sg13g2_nand2_1 _6280_ (.Y(_2170_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ),
    .B(_1955_));
 sg13g2_nand3_1 _6281_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ),
    .C(_1942_),
    .A(_1960_),
    .Y(_2171_));
 sg13g2_nand3_1 _6282_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ),
    .C(_1942_),
    .A(_1439_),
    .Y(_2172_));
 sg13g2_nor2b_1 _6283_ (.A(net303),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ),
    .Y(_2173_));
 sg13g2_a22oi_1 _6284_ (.Y(_2174_),
    .B1(_2173_),
    .B2(_1950_),
    .A2(_1930_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ));
 sg13g2_and4_1 _6285_ (.A(_2170_),
    .B(_2171_),
    .C(_2172_),
    .D(_2174_),
    .X(_2175_));
 sg13g2_nor2_1 _6286_ (.A(_1438_),
    .B(_1898_),
    .Y(_2176_));
 sg13g2_nand2b_1 _6287_ (.Y(_2177_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ),
    .A_N(net333));
 sg13g2_o21ai_1 _6288_ (.B1(_2177_),
    .Y(_2178_),
    .A1(_1896_),
    .A2(_0039_));
 sg13g2_a22oi_1 _6289_ (.Y(_2179_),
    .B1(_2178_),
    .B2(_1950_),
    .A2(_2176_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ));
 sg13g2_a21oi_1 _6290_ (.A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ),
    .A2(_1900_),
    .Y(_2180_),
    .B1(net283));
 sg13g2_a221oi_1 _6291_ (.B2(_2180_),
    .C1(net284),
    .B1(_2179_),
    .A1(net283),
    .Y(_2181_),
    .A2(_2175_));
 sg13g2_inv_1 _6292_ (.Y(_2182_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1] ));
 sg13g2_or2_1 _6293_ (.X(_2183_),
    .B(_1430_),
    .A(_1434_));
 sg13g2_buf_1 _6294_ (.A(_2183_),
    .X(_2184_));
 sg13g2_nand3_1 _6295_ (.B(_1430_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ),
    .A(net310),
    .Y(_2185_));
 sg13g2_o21ai_1 _6296_ (.B1(_2185_),
    .Y(_2186_),
    .A1(_2182_),
    .A2(_2184_));
 sg13g2_and2_1 _6297_ (.A(net286),
    .B(_1941_),
    .X(_2187_));
 sg13g2_nand2b_1 _6298_ (.Y(_2188_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ),
    .A_N(net333));
 sg13g2_nand3b_1 _6299_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ),
    .C(net285),
    .Y(_2189_),
    .A_N(net303));
 sg13g2_o21ai_1 _6300_ (.B1(_2189_),
    .Y(_2190_),
    .A1(net285),
    .A2(_2188_));
 sg13g2_a22oi_1 _6301_ (.Y(_2191_),
    .B1(_2187_),
    .B2(_2190_),
    .A2(_2186_),
    .A1(_1954_));
 sg13g2_a22oi_1 _6302_ (.Y(_2192_),
    .B1(_1929_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ),
    .A2(_1941_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ));
 sg13g2_nand2b_1 _6303_ (.Y(_2193_),
    .B(_1930_),
    .A_N(_2192_));
 sg13g2_a22oi_1 _6304_ (.Y(_2194_),
    .B1(_1911_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ),
    .A2(_1910_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ));
 sg13g2_nor2_2 _6305_ (.A(net286),
    .B(_1921_),
    .Y(_2195_));
 sg13g2_nand3b_1 _6306_ (.B(_2195_),
    .C(net304),
    .Y(_2196_),
    .A_N(_2194_));
 sg13g2_nor4_1 _6307_ (.A(net283),
    .B(_1430_),
    .C(_1422_),
    .D(net303),
    .Y(_2197_));
 sg13g2_mux2_1 _6308_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ),
    .S(_1426_),
    .X(_2198_));
 sg13g2_mux2_1 _6309_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ),
    .S(net310),
    .X(_2199_));
 sg13g2_nor2_1 _6310_ (.A(_1909_),
    .B(_1934_),
    .Y(_2200_));
 sg13g2_inv_1 _6311_ (.Y(_2201_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ));
 sg13g2_nor4_1 _6312_ (.A(net303),
    .B(_2201_),
    .C(_2184_),
    .D(_1934_),
    .Y(_2202_));
 sg13g2_a221oi_1 _6313_ (.B2(_2200_),
    .C1(_2202_),
    .B1(_2199_),
    .A1(_2197_),
    .Y(_2203_),
    .A2(_2198_));
 sg13g2_nand4_1 _6314_ (.B(_2193_),
    .C(_2196_),
    .A(_2191_),
    .Y(_2204_),
    .D(_2203_));
 sg13g2_or4_1 _6315_ (.A(_2160_),
    .B(_2169_),
    .C(_2181_),
    .D(_2204_),
    .X(_2205_));
 sg13g2_a22oi_1 _6316_ (.Y(_2206_),
    .B1(_2157_),
    .B2(_2205_),
    .A2(_1997_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ));
 sg13g2_nand2_1 _6317_ (.Y(_2207_),
    .A(_1785_),
    .B(_1711_));
 sg13g2_or4_1 _6318_ (.A(net330),
    .B(_1766_),
    .C(_1773_),
    .D(_1783_),
    .X(_2208_));
 sg13g2_a22oi_1 _6319_ (.Y(_2209_),
    .B1(_1842_),
    .B2(_2208_),
    .A2(_1785_),
    .A1(_1442_));
 sg13g2_o21ai_1 _6320_ (.B1(_1835_),
    .Y(_2210_),
    .A1(_1767_),
    .A2(_1831_));
 sg13g2_nand3_1 _6321_ (.B(_1823_),
    .C(_2210_),
    .A(_1852_),
    .Y(_2211_));
 sg13g2_nand4_1 _6322_ (.B(_2207_),
    .C(_2209_),
    .A(net174),
    .Y(_2212_),
    .D(_2211_));
 sg13g2_a221oi_1 _6323_ (.B2(_1851_),
    .C1(net224),
    .B1(_1850_),
    .A1(_1756_),
    .Y(_2213_),
    .A2(_1826_));
 sg13g2_nand2_1 _6324_ (.Y(_2214_),
    .A(_2207_),
    .B(_2213_));
 sg13g2_and3_1 _6325_ (.X(_2215_),
    .A(_2206_),
    .B(_2212_),
    .C(_2214_));
 sg13g2_buf_1 _6326_ (.A(_2215_),
    .X(_2216_));
 sg13g2_nand2b_1 _6327_ (.Y(_2217_),
    .B(_2206_),
    .A_N(_1686_));
 sg13g2_a21oi_1 _6328_ (.A1(_1367_),
    .A2(_1811_),
    .Y(_2218_),
    .B1(_1882_));
 sg13g2_o21ai_1 _6329_ (.B1(_2218_),
    .Y(_2219_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .A2(_1878_));
 sg13g2_buf_1 _6330_ (.A(_2219_),
    .X(_2220_));
 sg13g2_nand2_1 _6331_ (.Y(_2221_),
    .A(_2206_),
    .B(_2220_));
 sg13g2_o21ai_1 _6332_ (.B1(_2221_),
    .Y(_2222_),
    .A1(_1817_),
    .A2(_2217_));
 sg13g2_buf_1 _6333_ (.A(_2222_),
    .X(_2223_));
 sg13g2_inv_1 _6334_ (.Y(_2224_),
    .A(_2220_));
 sg13g2_o21ai_1 _6335_ (.B1(net223),
    .Y(_2225_),
    .A1(net230),
    .A2(_1839_));
 sg13g2_a21oi_1 _6336_ (.A1(net308),
    .A2(_2225_),
    .Y(_2226_),
    .B1(_1724_));
 sg13g2_o21ai_1 _6337_ (.B1(_1383_),
    .Y(_2227_),
    .A1(_1732_),
    .A2(_1710_));
 sg13g2_nand4_1 _6338_ (.B(_1809_),
    .C(_1813_),
    .A(net277),
    .Y(_2228_),
    .D(_2227_));
 sg13g2_nand2b_1 _6339_ (.Y(_2229_),
    .B(_2228_),
    .A_N(_2226_));
 sg13g2_nor3_1 _6340_ (.A(_2213_),
    .B(_2220_),
    .C(_2229_),
    .Y(_2230_));
 sg13g2_nand3_1 _6341_ (.B(_2209_),
    .C(_2211_),
    .A(net174),
    .Y(_2231_));
 sg13g2_nor3_1 _6342_ (.A(_2207_),
    .B(_2220_),
    .C(_2229_),
    .Y(_2232_));
 sg13g2_a221oi_1 _6343_ (.B2(_2231_),
    .C1(_2232_),
    .B1(_2230_),
    .A1(net319),
    .Y(_2233_),
    .A2(_2224_));
 sg13g2_o21ai_1 _6344_ (.B1(_2233_),
    .Y(_2234_),
    .A1(_2216_),
    .A2(_2223_));
 sg13g2_buf_2 _6345_ (.A(_2234_),
    .X(_2235_));
 sg13g2_inv_1 _6346_ (.Y(_2236_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ));
 sg13g2_nand3_1 _6347_ (.B(_1397_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ),
    .A(net315),
    .Y(_2237_));
 sg13g2_o21ai_1 _6348_ (.B1(_2237_),
    .Y(_2238_),
    .A1(_2236_),
    .A2(_2086_));
 sg13g2_nand3_1 _6349_ (.B(net313),
    .C(_2238_),
    .A(_1407_),
    .Y(_2239_));
 sg13g2_nand2_1 _6350_ (.Y(_2240_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ),
    .B(_2039_));
 sg13g2_nor2b_2 _6351_ (.A(net301),
    .B_N(_1396_),
    .Y(_2241_));
 sg13g2_a22oi_1 _6352_ (.Y(_2242_),
    .B1(_2241_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ),
    .A2(_2032_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ));
 sg13g2_nand3_1 _6353_ (.B(_2240_),
    .C(_2242_),
    .A(_1407_),
    .Y(_2243_));
 sg13g2_buf_1 _6354_ (.A(_2078_),
    .X(_2244_));
 sg13g2_nand2_1 _6355_ (.Y(_2245_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ),
    .B(_2241_));
 sg13g2_a22oi_1 _6356_ (.Y(_2246_),
    .B1(_2039_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ),
    .A2(_2035_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ));
 sg13g2_nand3_1 _6357_ (.B(_2245_),
    .C(_2246_),
    .A(net258),
    .Y(_2247_));
 sg13g2_nand3_1 _6358_ (.B(_2243_),
    .C(_2247_),
    .A(net265),
    .Y(_2248_));
 sg13g2_and2_1 _6359_ (.A(_2021_),
    .B(_2026_),
    .X(_2249_));
 sg13g2_mux2_1 _6360_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ),
    .S(net278),
    .X(_2250_));
 sg13g2_a22oi_1 _6361_ (.Y(_2251_),
    .B1(_2250_),
    .B2(net242),
    .A2(_2249_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ));
 sg13g2_or2_1 _6362_ (.X(_2252_),
    .B(_2251_),
    .A(net265));
 sg13g2_nand4_1 _6363_ (.B(_2239_),
    .C(_2248_),
    .A(net287),
    .Y(_2253_),
    .D(_2252_));
 sg13g2_nand2b_1 _6364_ (.Y(_2254_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ),
    .A_N(_1418_));
 sg13g2_o21ai_1 _6365_ (.B1(_2254_),
    .Y(_2255_),
    .A1(net300),
    .A2(_0039_));
 sg13g2_nor2b_1 _6366_ (.A(net300),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ),
    .Y(_2256_));
 sg13g2_nor2b_1 _6367_ (.A(net300),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ),
    .Y(_2257_));
 sg13g2_nor2b_1 _6368_ (.A(_1418_),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ),
    .Y(_2258_));
 sg13g2_a21o_1 _6369_ (.A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ),
    .A1(_2021_),
    .B1(_2258_),
    .X(_2259_));
 sg13g2_mux4_1 _6370_ (.S0(_1397_),
    .A0(_2255_),
    .A1(_2256_),
    .A2(_2257_),
    .A3(_2259_),
    .S1(_1407_),
    .X(_2260_));
 sg13g2_a22oi_1 _6371_ (.Y(_2261_),
    .B1(_2044_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ),
    .A2(_2026_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ));
 sg13g2_o21ai_1 _6372_ (.B1(net288),
    .Y(_2262_),
    .A1(net301),
    .A2(_2261_));
 sg13g2_nand3_1 _6373_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ),
    .C(_2035_),
    .A(net258),
    .Y(_2263_));
 sg13g2_mux2_1 _6374_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ),
    .S(net316),
    .X(_2264_));
 sg13g2_mux2_1 _6375_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ),
    .S(_1406_),
    .X(_2265_));
 sg13g2_a22oi_1 _6376_ (.Y(_2266_),
    .B1(_2265_),
    .B2(_2032_),
    .A2(_2264_),
    .A1(_2241_));
 sg13g2_nand3b_1 _6377_ (.B(_2263_),
    .C(_2266_),
    .Y(_2267_),
    .A_N(net288));
 sg13g2_o21ai_1 _6378_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_2260_),
    .A2(_2262_));
 sg13g2_nand2_1 _6379_ (.Y(_2269_),
    .A(net259),
    .B(_2268_));
 sg13g2_buf_1 _6380_ (.A(net317),
    .X(_2270_));
 sg13g2_a22oi_1 _6381_ (.Y(_2271_),
    .B1(_2064_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ),
    .A2(_2062_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1] ));
 sg13g2_or4_1 _6382_ (.A(net265),
    .B(net276),
    .C(net301),
    .D(_2271_),
    .X(_2272_));
 sg13g2_mux2_1 _6383_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ),
    .S(net288),
    .X(_2273_));
 sg13g2_nand3_1 _6384_ (.B(_2083_),
    .C(_2273_),
    .A(_2006_),
    .Y(_2274_));
 sg13g2_mux2_1 _6385_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ),
    .S(_2244_),
    .X(_2275_));
 sg13g2_nand3_1 _6386_ (.B(_2053_),
    .C(_2275_),
    .A(_2067_),
    .Y(_2276_));
 sg13g2_nand3_1 _6387_ (.B(_2274_),
    .C(_2276_),
    .A(_2272_),
    .Y(_2277_));
 sg13g2_a221oi_1 _6388_ (.B2(_2269_),
    .C1(_2277_),
    .B1(_2253_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ),
    .Y(_2278_),
    .A2(_2059_));
 sg13g2_nand2_1 _6389_ (.Y(_2279_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .B(_2077_));
 sg13g2_o21ai_1 _6390_ (.B1(_2279_),
    .Y(_2280_),
    .A1(_2077_),
    .A2(_2278_));
 sg13g2_buf_2 _6391_ (.A(_2280_),
    .X(_2281_));
 sg13g2_a22oi_1 _6392_ (.Y(_2282_),
    .B1(_2235_),
    .B2(_2110_),
    .A2(_2281_),
    .A1(_2111_));
 sg13g2_buf_1 _6393_ (.A(_2282_),
    .X(_2283_));
 sg13g2_or2_1 _6394_ (.X(_2284_),
    .B(_2223_),
    .A(_2216_));
 sg13g2_nor2_1 _6395_ (.A(_2095_),
    .B(net173),
    .Y(_2285_));
 sg13g2_mux2_1 _6396_ (.A0(_2003_),
    .A1(_2096_),
    .S(_2281_),
    .X(_2286_));
 sg13g2_a221oi_1 _6397_ (.B2(_2285_),
    .C1(_2286_),
    .B1(_2235_),
    .A1(_2002_),
    .Y(_2287_),
    .A2(_2284_));
 sg13g2_buf_1 _6398_ (.A(_2287_),
    .X(_2288_));
 sg13g2_or2_1 _6399_ (.X(_2289_),
    .B(_2288_),
    .A(_2283_));
 sg13g2_buf_1 _6400_ (.A(_2289_),
    .X(_2290_));
 sg13g2_nor2_1 _6401_ (.A(_2139_),
    .B(_2290_),
    .Y(_2291_));
 sg13g2_and2_1 _6402_ (.A(_1985_),
    .B(_2144_),
    .X(_2292_));
 sg13g2_nand3_1 _6403_ (.B(_2102_),
    .C(_2106_),
    .A(_2101_),
    .Y(_2293_));
 sg13g2_buf_1 _6404_ (.A(_2293_),
    .X(_2294_));
 sg13g2_nor2_1 _6405_ (.A(net173),
    .B(net96),
    .Y(_2295_));
 sg13g2_nor2_1 _6406_ (.A(_2093_),
    .B(_2295_),
    .Y(_2296_));
 sg13g2_a21oi_1 _6407_ (.A1(_2089_),
    .A2(_2091_),
    .Y(_2297_),
    .B1(_1993_));
 sg13g2_and2_1 _6408_ (.A(_2095_),
    .B(_2297_),
    .X(_2298_));
 sg13g2_a22oi_1 _6409_ (.Y(_2299_),
    .B1(_2298_),
    .B2(_2144_),
    .A2(_2296_),
    .A1(_2292_));
 sg13g2_buf_1 _6410_ (.A(_2299_),
    .X(_2300_));
 sg13g2_or2_1 _6411_ (.X(_2301_),
    .B(_2144_),
    .A(_1985_));
 sg13g2_a21o_1 _6412_ (.A2(_2301_),
    .A1(_2091_),
    .B1(_2292_),
    .X(_2302_));
 sg13g2_nand2_1 _6413_ (.Y(_2303_),
    .A(net96),
    .B(_2302_));
 sg13g2_nand3_1 _6414_ (.B(net96),
    .C(_2302_),
    .A(_2089_),
    .Y(_2304_));
 sg13g2_nand2_1 _6415_ (.Y(_2305_),
    .A(_1985_),
    .B(_2144_));
 sg13g2_a22oi_1 _6416_ (.Y(_2306_),
    .B1(_2304_),
    .B2(_2305_),
    .A2(_2303_),
    .A1(_2297_));
 sg13g2_nor2_1 _6417_ (.A(_2298_),
    .B(_2306_),
    .Y(_2307_));
 sg13g2_nor2_1 _6418_ (.A(_2093_),
    .B(_2108_),
    .Y(_2308_));
 sg13g2_o21ai_1 _6419_ (.B1(_2002_),
    .Y(_2309_),
    .A1(_2144_),
    .A2(_2308_));
 sg13g2_mux2_1 _6420_ (.A0(_2307_),
    .A1(_2309_),
    .S(_1982_),
    .X(_2310_));
 sg13g2_buf_2 _6421_ (.A(_2310_),
    .X(_2311_));
 sg13g2_and2_1 _6422_ (.A(_2300_),
    .B(_2311_),
    .X(_2312_));
 sg13g2_buf_1 _6423_ (.A(_2312_),
    .X(_2313_));
 sg13g2_a21oi_1 _6424_ (.A1(_2148_),
    .A2(_2313_),
    .Y(_2314_),
    .B1(_2142_));
 sg13g2_or2_1 _6425_ (.X(_2315_),
    .B(_2313_),
    .A(_2138_));
 sg13g2_xnor2_1 _6426_ (.Y(_2316_),
    .A(net51),
    .B(net50));
 sg13g2_mux2_1 _6427_ (.A0(_2314_),
    .A1(_2315_),
    .S(_2316_),
    .X(_2317_));
 sg13g2_nor2b_2 _6428_ (.A(_2291_),
    .B_N(_2317_),
    .Y(_2318_));
 sg13g2_nor2_1 _6429_ (.A(net175),
    .B(_2318_),
    .Y(_2319_));
 sg13g2_a21oi_1 _6430_ (.A1(net175),
    .A2(_2235_),
    .Y(_2320_),
    .B1(_2319_));
 sg13g2_nand2_1 _6431_ (.Y(_2321_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29] ),
    .B(net74));
 sg13g2_o21ai_1 _6432_ (.B1(_2321_),
    .Y(_1235_),
    .A1(net75),
    .A2(_2320_));
 sg13g2_buf_1 _6433_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[2] ),
    .X(_2322_));
 sg13g2_nand2_1 _6434_ (.Y(_2323_),
    .A(_2322_),
    .B(net74));
 sg13g2_o21ai_1 _6435_ (.B1(_2323_),
    .Y(_1236_),
    .A1(_1778_),
    .A2(net75));
 sg13g2_buf_1 _6436_ (.A(_2095_),
    .X(_2324_));
 sg13g2_a221oi_1 _6437_ (.B2(_1819_),
    .C1(_1478_),
    .B1(_1825_),
    .A1(_1820_),
    .Y(_2325_),
    .A2(_1823_));
 sg13g2_a21oi_1 _6438_ (.A1(_1821_),
    .A2(_1823_),
    .Y(_2326_),
    .B1(net330));
 sg13g2_nand2_1 _6439_ (.Y(_2327_),
    .A(_1843_),
    .B(_1837_));
 sg13g2_nor3_1 _6440_ (.A(_2325_),
    .B(_2326_),
    .C(_2327_),
    .Y(_2328_));
 sg13g2_nand2_1 _6441_ (.Y(_2329_),
    .A(_1847_),
    .B(_1848_));
 sg13g2_nor2_1 _6442_ (.A(_1751_),
    .B(_1824_),
    .Y(_2330_));
 sg13g2_nor2_1 _6443_ (.A(_1843_),
    .B(_2330_),
    .Y(_2331_));
 sg13g2_nand3_1 _6444_ (.B(_2329_),
    .C(_2331_),
    .A(_1850_),
    .Y(_2332_));
 sg13g2_o21ai_1 _6445_ (.B1(_1700_),
    .Y(_2333_),
    .A1(net305),
    .A2(net174));
 sg13g2_a22oi_1 _6446_ (.Y(_2334_),
    .B1(_2331_),
    .B2(_1756_),
    .A2(_2333_),
    .A1(_1785_));
 sg13g2_nand3b_1 _6447_ (.B(_2332_),
    .C(_2334_),
    .Y(_2335_),
    .A_N(net319));
 sg13g2_or4_1 _6448_ (.A(_1686_),
    .B(_1817_),
    .C(_2328_),
    .D(_2335_),
    .X(_2336_));
 sg13g2_buf_1 _6449_ (.A(_2336_),
    .X(_2337_));
 sg13g2_a21oi_1 _6450_ (.A1(net319),
    .A2(_1701_),
    .Y(_2338_),
    .B1(_1882_));
 sg13g2_o21ai_1 _6451_ (.B1(_2338_),
    .Y(_2339_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .A2(_1878_));
 sg13g2_a22oi_1 _6452_ (.Y(_2340_),
    .B1(_1721_),
    .B2(_1730_),
    .A2(_1715_),
    .A1(net306));
 sg13g2_a21o_1 _6453_ (.A2(_2340_),
    .A1(_1713_),
    .B1(_1368_),
    .X(_2341_));
 sg13g2_nor4_1 _6454_ (.A(_2325_),
    .B(_2326_),
    .C(_2327_),
    .D(_2341_),
    .Y(_2342_));
 sg13g2_a21oi_1 _6455_ (.A1(_2332_),
    .A2(_2334_),
    .Y(_2343_),
    .B1(_2341_));
 sg13g2_nor3_2 _6456_ (.A(_2339_),
    .B(_2342_),
    .C(_2343_),
    .Y(_2344_));
 sg13g2_mux2_1 _6457_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ),
    .S(net264),
    .X(_2345_));
 sg13g2_a22oi_1 _6458_ (.Y(_2346_),
    .B1(_2345_),
    .B2(_1428_),
    .A2(_1950_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ));
 sg13g2_mux2_1 _6459_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ),
    .S(net264),
    .X(_2347_));
 sg13g2_a22oi_1 _6460_ (.Y(_2348_),
    .B1(_2347_),
    .B2(_1428_),
    .A2(_1950_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ));
 sg13g2_or2_1 _6461_ (.X(_2349_),
    .B(_2348_),
    .A(net280));
 sg13g2_o21ai_1 _6462_ (.B1(_2349_),
    .Y(_2350_),
    .A1(net302),
    .A2(_2346_));
 sg13g2_a22oi_1 _6463_ (.Y(_2351_),
    .B1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ),
    .B2(_1439_),
    .A2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ),
    .A1(_1960_));
 sg13g2_nand3_1 _6464_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ),
    .C(_1965_),
    .A(_1960_),
    .Y(_2352_));
 sg13g2_o21ai_1 _6465_ (.B1(_2352_),
    .Y(_2353_),
    .A1(_2184_),
    .A2(_2351_));
 sg13g2_nand3_1 _6466_ (.B(_1965_),
    .C(_2176_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ),
    .Y(_2354_));
 sg13g2_nand2_1 _6467_ (.Y(_2355_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ),
    .B(_1932_));
 sg13g2_a22oi_1 _6468_ (.Y(_2356_),
    .B1(_1929_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ),
    .A2(_1941_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2] ));
 sg13g2_nand2b_1 _6469_ (.Y(_2357_),
    .B(_1900_),
    .A_N(_2356_));
 sg13g2_nand3_1 _6470_ (.B(_2355_),
    .C(_2357_),
    .A(_2354_),
    .Y(_2358_));
 sg13g2_a221oi_1 _6471_ (.B2(_1902_),
    .C1(_2358_),
    .B1(_2353_),
    .A1(_1963_),
    .Y(_2359_),
    .A2(_2350_));
 sg13g2_a22oi_1 _6472_ (.Y(_2360_),
    .B1(_1900_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ),
    .A2(_1955_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ));
 sg13g2_nand3_1 _6473_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ),
    .C(_1894_),
    .A(net284),
    .Y(_2361_));
 sg13g2_o21ai_1 _6474_ (.B1(_2361_),
    .Y(_2362_),
    .A1(net284),
    .A2(_2360_));
 sg13g2_a22oi_1 _6475_ (.Y(_2363_),
    .B1(_1950_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ),
    .A2(_1962_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ));
 sg13g2_nor2_1 _6476_ (.A(net304),
    .B(net280),
    .Y(_2364_));
 sg13g2_nand2b_1 _6477_ (.Y(_2365_),
    .B(_2364_),
    .A_N(_2363_));
 sg13g2_nand3_1 _6478_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ),
    .C(_1954_),
    .A(net282),
    .Y(_2366_));
 sg13g2_nand3_1 _6479_ (.B(_2365_),
    .C(_2366_),
    .A(_1436_),
    .Y(_2367_));
 sg13g2_a221oi_1 _6480_ (.B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ),
    .C1(net284),
    .B1(_1955_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ),
    .Y(_2368_),
    .A2(_1894_));
 sg13g2_a21oi_1 _6481_ (.A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ),
    .A2(_1954_),
    .Y(_2369_),
    .B1(net282));
 sg13g2_o21ai_1 _6482_ (.B1(net261),
    .Y(_2370_),
    .A1(_2368_),
    .A2(_2369_));
 sg13g2_o21ai_1 _6483_ (.B1(_2370_),
    .Y(_2371_),
    .A1(_2362_),
    .A2(_2367_));
 sg13g2_nand2_1 _6484_ (.Y(_2372_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2] ),
    .B(_2176_));
 sg13g2_nand3_1 _6485_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ),
    .C(_1935_),
    .A(_1914_),
    .Y(_2373_));
 sg13g2_o21ai_1 _6486_ (.B1(_2373_),
    .Y(_2374_),
    .A1(net261),
    .A2(_2372_));
 sg13g2_and2_1 _6487_ (.A(_1914_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ),
    .X(_2375_));
 sg13g2_nor2b_1 _6488_ (.A(net261),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ),
    .Y(_2376_));
 sg13g2_a22oi_1 _6489_ (.Y(_2377_),
    .B1(_2376_),
    .B2(_1894_),
    .A2(_2375_),
    .A1(_1954_));
 sg13g2_nor2b_1 _6490_ (.A(net261),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ),
    .Y(_2378_));
 sg13g2_a22oi_1 _6491_ (.Y(_2379_),
    .B1(_2378_),
    .B2(_1944_),
    .A2(_1968_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ));
 sg13g2_and2_1 _6492_ (.A(net281),
    .B(net260),
    .X(_2380_));
 sg13g2_mux2_1 _6493_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ),
    .S(_1424_),
    .X(_2381_));
 sg13g2_a22oi_1 _6494_ (.Y(_2382_),
    .B1(_2380_),
    .B2(_2381_),
    .A2(_1947_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ));
 sg13g2_or2_1 _6495_ (.X(_2383_),
    .B(_2382_),
    .A(net280));
 sg13g2_nand4_1 _6496_ (.B(_2377_),
    .C(_2379_),
    .A(net282),
    .Y(_2384_),
    .D(_2383_));
 sg13g2_o21ai_1 _6497_ (.B1(_2384_),
    .Y(_2385_),
    .A1(_1891_),
    .A2(_2374_));
 sg13g2_nand3_1 _6498_ (.B(_2371_),
    .C(_2385_),
    .A(_2359_),
    .Y(_2386_));
 sg13g2_a22oi_1 _6499_ (.Y(_2387_),
    .B1(_2157_),
    .B2(_2386_),
    .A2(_1997_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ));
 sg13g2_inv_1 _6500_ (.Y(_2388_),
    .A(_2387_));
 sg13g2_a21oi_2 _6501_ (.B1(_2388_),
    .Y(_2389_),
    .A2(_2344_),
    .A1(_2337_));
 sg13g2_buf_1 _6502_ (.A(_2389_),
    .X(_2390_));
 sg13g2_nor2_1 _6503_ (.A(net97),
    .B(net96),
    .Y(_2391_));
 sg13g2_nand3_1 _6504_ (.B(net258),
    .C(_2241_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ),
    .Y(_2392_));
 sg13g2_and3_1 _6505_ (.X(_2393_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ),
    .B(net278),
    .C(net276));
 sg13g2_a21o_1 _6506_ (.A2(_2007_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ),
    .B1(_2393_),
    .X(_2394_));
 sg13g2_mux2_1 _6507_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ),
    .S(net276),
    .X(_2395_));
 sg13g2_and3_1 _6508_ (.X(_2396_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ),
    .B(net278),
    .C(net276));
 sg13g2_a21o_1 _6509_ (.A2(_2395_),
    .A1(_1407_),
    .B1(_2396_),
    .X(_2397_));
 sg13g2_a22oi_1 _6510_ (.Y(_2398_),
    .B1(_2397_),
    .B2(net313),
    .A2(_2394_),
    .A1(_2021_));
 sg13g2_mux2_1 _6511_ (.A0(_2392_),
    .A1(_2398_),
    .S(net259),
    .X(_2399_));
 sg13g2_nand3_1 _6512_ (.B(net259),
    .C(_2035_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ),
    .Y(_2400_));
 sg13g2_nand3_1 _6513_ (.B(net287),
    .C(net242),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ),
    .Y(_2401_));
 sg13g2_nand2_1 _6514_ (.Y(_2402_),
    .A(_2400_),
    .B(_2401_));
 sg13g2_a22oi_1 _6515_ (.Y(_2403_),
    .B1(_2064_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ),
    .A2(_2062_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ));
 sg13g2_inv_1 _6516_ (.Y(_2404_),
    .A(_2403_));
 sg13g2_a221oi_1 _6517_ (.B2(_2032_),
    .C1(net265),
    .B1(_2404_),
    .A1(net258),
    .Y(_2405_),
    .A2(_2402_));
 sg13g2_a21oi_1 _6518_ (.A1(net265),
    .A2(_2399_),
    .Y(_2406_),
    .B1(_2405_));
 sg13g2_mux2_1 _6519_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ),
    .S(net276),
    .X(_2407_));
 sg13g2_nand3_1 _6520_ (.B(net313),
    .C(_2407_),
    .A(_1407_),
    .Y(_2408_));
 sg13g2_nand3_1 _6521_ (.B(net258),
    .C(net242),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ),
    .Y(_2409_));
 sg13g2_nand2_1 _6522_ (.Y(_2410_),
    .A(net287),
    .B(net265));
 sg13g2_a21oi_1 _6523_ (.A1(_2408_),
    .A2(_2409_),
    .Y(_2411_),
    .B1(_2410_));
 sg13g2_nand3_1 _6524_ (.B(net259),
    .C(net258),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ),
    .Y(_2412_));
 sg13g2_mux2_1 _6525_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ),
    .S(net278),
    .X(_2413_));
 sg13g2_a22oi_1 _6526_ (.Y(_2414_),
    .B1(_2413_),
    .B2(net287),
    .A2(_2064_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ));
 sg13g2_mux2_1 _6527_ (.A0(_2412_),
    .A1(_2414_),
    .S(net265),
    .X(_2415_));
 sg13g2_nor2b_1 _6528_ (.A(_2415_),
    .B_N(_2032_),
    .Y(_2416_));
 sg13g2_mux2_1 _6529_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ),
    .S(net276),
    .X(_2417_));
 sg13g2_nand3_1 _6530_ (.B(_2036_),
    .C(_2417_),
    .A(_1419_),
    .Y(_2418_));
 sg13g2_and2_1 _6531_ (.A(_1410_),
    .B(net316),
    .X(_2419_));
 sg13g2_buf_2 _6532_ (.A(_2419_),
    .X(_2420_));
 sg13g2_nand3_1 _6533_ (.B(net242),
    .C(_2420_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ),
    .Y(_2421_));
 sg13g2_a21o_1 _6534_ (.A2(_2421_),
    .A1(_2418_),
    .B1(net287),
    .X(_2422_));
 sg13g2_inv_1 _6535_ (.Y(_2423_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2] ));
 sg13g2_nand3b_1 _6536_ (.B(_1411_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ),
    .Y(_2424_),
    .A_N(net276));
 sg13g2_o21ai_1 _6537_ (.B1(_2424_),
    .Y(_2425_),
    .A1(_2423_),
    .A2(_2086_));
 sg13g2_or2_1 _6538_ (.X(_2426_),
    .B(net278),
    .A(net314));
 sg13g2_nor2_1 _6539_ (.A(net300),
    .B(_2426_),
    .Y(_2427_));
 sg13g2_mux2_1 _6540_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ),
    .S(net279),
    .X(_2428_));
 sg13g2_and2_1 _6541_ (.A(_2035_),
    .B(_2420_),
    .X(_2429_));
 sg13g2_mux2_1 _6542_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ),
    .S(_2078_),
    .X(_2430_));
 sg13g2_and3_1 _6543_ (.X(_2431_),
    .A(net242),
    .B(_2053_),
    .C(_2430_));
 sg13g2_a221oi_1 _6544_ (.B2(_2429_),
    .C1(_2431_),
    .B1(_2428_),
    .A1(_2425_),
    .Y(_2432_),
    .A2(_2427_));
 sg13g2_nand2b_1 _6545_ (.Y(_2433_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ),
    .A_N(net278));
 sg13g2_nand3b_1 _6546_ (.B(_2244_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ),
    .Y(_2434_),
    .A_N(_2004_));
 sg13g2_o21ai_1 _6547_ (.B1(_2434_),
    .Y(_2435_),
    .A1(_2010_),
    .A2(_2433_));
 sg13g2_nand3_1 _6548_ (.B(_2057_),
    .C(_2435_),
    .A(_1397_),
    .Y(_2436_));
 sg13g2_inv_1 _6549_ (.Y(_2437_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2] ));
 sg13g2_nand3_1 _6550_ (.B(net279),
    .C(net278),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ),
    .Y(_2438_));
 sg13g2_o21ai_1 _6551_ (.B1(_2438_),
    .Y(_2439_),
    .A1(_2437_),
    .A2(_2426_));
 sg13g2_nand2b_1 _6552_ (.Y(_2440_),
    .B(net276),
    .A_N(net301));
 sg13g2_nor2_1 _6553_ (.A(net288),
    .B(_2440_),
    .Y(_2441_));
 sg13g2_a22oi_1 _6554_ (.Y(_2442_),
    .B1(_2439_),
    .B2(_2441_),
    .A2(_2059_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ));
 sg13g2_nand4_1 _6555_ (.B(_2432_),
    .C(_2436_),
    .A(_2422_),
    .Y(_2443_),
    .D(_2442_));
 sg13g2_or4_1 _6556_ (.A(_2077_),
    .B(_2411_),
    .C(_2416_),
    .D(_2443_),
    .X(_2444_));
 sg13g2_nand2b_1 _6557_ (.Y(_2445_),
    .B(_2077_),
    .A_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i ));
 sg13g2_o21ai_1 _6558_ (.B1(_2445_),
    .Y(_2446_),
    .A1(_2406_),
    .A2(_2444_));
 sg13g2_buf_1 _6559_ (.A(_2446_),
    .X(_2447_));
 sg13g2_o21ai_1 _6560_ (.B1(net80),
    .Y(_2448_),
    .A1(net52),
    .A2(_2391_));
 sg13g2_or2_1 _6561_ (.X(_2449_),
    .B(net80),
    .A(_2108_));
 sg13g2_buf_1 _6562_ (.A(_2449_),
    .X(_2450_));
 sg13g2_a21o_1 _6563_ (.A2(_2344_),
    .A1(_2337_),
    .B1(_2388_),
    .X(_2451_));
 sg13g2_nand2b_1 _6564_ (.Y(_2452_),
    .B(_2451_),
    .A_N(_2450_));
 sg13g2_buf_2 _6565_ (.A(_2452_),
    .X(_2453_));
 sg13g2_nand2_1 _6566_ (.Y(_2454_),
    .A(_2295_),
    .B(_2390_));
 sg13g2_nand3_1 _6567_ (.B(_2453_),
    .C(_2454_),
    .A(_2448_),
    .Y(_2455_));
 sg13g2_xnor2_1 _6568_ (.Y(_2456_),
    .A(net241),
    .B(_2455_));
 sg13g2_and2_1 _6569_ (.A(net51),
    .B(net50),
    .X(_2457_));
 sg13g2_a21oi_1 _6570_ (.A1(_2290_),
    .A2(_2313_),
    .Y(_2458_),
    .B1(_2457_));
 sg13g2_xnor2_1 _6571_ (.Y(_2459_),
    .A(_2456_),
    .B(_2458_));
 sg13g2_and2_1 _6572_ (.A(net173),
    .B(net80),
    .X(_2460_));
 sg13g2_inv_1 _6573_ (.Y(_2461_),
    .A(_2460_));
 sg13g2_nand2b_1 _6574_ (.Y(_2462_),
    .B(net97),
    .A_N(net80));
 sg13g2_mux2_1 _6575_ (.A0(_2461_),
    .A1(_2462_),
    .S(_2389_),
    .X(_2463_));
 sg13g2_or3_1 _6576_ (.A(net241),
    .B(net52),
    .C(net80),
    .X(_2464_));
 sg13g2_o21ai_1 _6577_ (.B1(_2464_),
    .Y(_2465_),
    .A1(net243),
    .A2(_2463_));
 sg13g2_nor2_1 _6578_ (.A(net86),
    .B(_2118_),
    .Y(_2466_));
 sg13g2_a221oi_1 _6579_ (.B2(_2140_),
    .C1(_2148_),
    .B1(_2456_),
    .A1(_2465_),
    .Y(_2467_),
    .A2(_2466_));
 sg13g2_a21oi_2 _6580_ (.B1(_2467_),
    .Y(_2468_),
    .A2(_2459_),
    .A1(_2148_));
 sg13g2_nand2_1 _6581_ (.Y(_2469_),
    .A(net175),
    .B(_2390_));
 sg13g2_o21ai_1 _6582_ (.B1(_2469_),
    .Y(_2470_),
    .A1(net175),
    .A2(_2468_));
 sg13g2_nand2_1 _6583_ (.Y(_2471_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30] ),
    .B(net74));
 sg13g2_o21ai_1 _6584_ (.B1(_2471_),
    .Y(_1237_),
    .A1(net75),
    .A2(_2470_));
 sg13g2_nand2b_1 _6585_ (.Y(_2472_),
    .B(_1764_),
    .A_N(_1831_));
 sg13g2_nand2_1 _6586_ (.Y(_2473_),
    .A(_1750_),
    .B(_1478_));
 sg13g2_nand2_1 _6587_ (.Y(_2474_),
    .A(_1751_),
    .B(_1477_));
 sg13g2_nor3_1 _6588_ (.A(_1766_),
    .B(_1773_),
    .C(_1783_),
    .Y(_2475_));
 sg13g2_a221oi_1 _6589_ (.B2(_2474_),
    .C1(_2475_),
    .B1(_2473_),
    .A1(_1835_),
    .Y(_2476_),
    .A2(_2472_));
 sg13g2_o21ai_1 _6590_ (.B1(net223),
    .Y(_2477_),
    .A1(_1824_),
    .A2(_1753_));
 sg13g2_a21o_1 _6591_ (.A2(_2330_),
    .A1(_1823_),
    .B1(_2477_),
    .X(_2478_));
 sg13g2_nor2_1 _6592_ (.A(_2476_),
    .B(_2478_),
    .Y(_2479_));
 sg13g2_nor2_1 _6593_ (.A(net260),
    .B(net280),
    .Y(_2480_));
 sg13g2_nor2b_1 _6594_ (.A(_1921_),
    .B_N(_1427_),
    .Y(_2481_));
 sg13g2_and2_1 _6595_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ),
    .B(_2481_),
    .X(_2482_));
 sg13g2_a21o_1 _6596_ (.A2(_2480_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ),
    .B1(_2482_),
    .X(_2483_));
 sg13g2_a22oi_1 _6597_ (.Y(_2484_),
    .B1(_2480_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ),
    .A2(_2481_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ));
 sg13g2_nor3_1 _6598_ (.A(net264),
    .B(_2184_),
    .C(_2484_),
    .Y(_2485_));
 sg13g2_a221oi_1 _6599_ (.B2(_2483_),
    .C1(_2485_),
    .B1(_2187_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ),
    .Y(_2486_),
    .A2(_1932_));
 sg13g2_buf_1 _6600_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[3] ),
    .X(_2487_));
 sg13g2_a22oi_1 _6601_ (.Y(_2488_),
    .B1(_1929_),
    .B2(_2487_),
    .A2(_1941_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ));
 sg13g2_nand2b_1 _6602_ (.Y(_2489_),
    .B(_1935_),
    .A_N(_2488_));
 sg13g2_nand2_1 _6603_ (.Y(_2490_),
    .A(net286),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ));
 sg13g2_nand3b_1 _6604_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ),
    .C(net310),
    .Y(_2491_),
    .A_N(_1423_));
 sg13g2_o21ai_1 _6605_ (.B1(_2491_),
    .Y(_2492_),
    .A1(_1913_),
    .A2(_2490_));
 sg13g2_nand3_1 _6606_ (.B(_2364_),
    .C(_2492_),
    .A(_1915_),
    .Y(_2493_));
 sg13g2_mux2_1 _6607_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ),
    .S(net260),
    .X(_2494_));
 sg13g2_nand3_1 _6608_ (.B(_2195_),
    .C(_2494_),
    .A(_1929_),
    .Y(_2495_));
 sg13g2_buf_1 _6609_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[3] ),
    .X(_2496_));
 sg13g2_a22oi_1 _6610_ (.Y(_2497_),
    .B1(_1929_),
    .B2(_2496_),
    .A2(_1941_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ));
 sg13g2_nand2b_1 _6611_ (.Y(_2498_),
    .B(_2176_),
    .A_N(_2497_));
 sg13g2_and4_1 _6612_ (.A(_2489_),
    .B(_2493_),
    .C(_2495_),
    .D(_2498_),
    .X(_2499_));
 sg13g2_nand2_1 _6613_ (.Y(_2500_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ),
    .B(_2161_));
 sg13g2_nand3_1 _6614_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ),
    .C(_2195_),
    .A(net260),
    .Y(_2501_));
 sg13g2_o21ai_1 _6615_ (.B1(_2501_),
    .Y(_2502_),
    .A1(_1915_),
    .A2(_2500_));
 sg13g2_a22oi_1 _6616_ (.Y(_2503_),
    .B1(_1950_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ),
    .A2(_1962_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ));
 sg13g2_nor2_1 _6617_ (.A(_1924_),
    .B(_2503_),
    .Y(_2504_));
 sg13g2_o21ai_1 _6618_ (.B1(_1965_),
    .Y(_2505_),
    .A1(_2502_),
    .A2(_2504_));
 sg13g2_and3_1 _6619_ (.X(_2506_),
    .A(_2486_),
    .B(_2499_),
    .C(_2505_));
 sg13g2_nor2_1 _6620_ (.A(_1428_),
    .B(net280),
    .Y(_2507_));
 sg13g2_nor2_1 _6621_ (.A(net260),
    .B(net302),
    .Y(_2508_));
 sg13g2_a22oi_1 _6622_ (.Y(_2509_),
    .B1(_2508_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ),
    .A2(_2507_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ));
 sg13g2_mux2_1 _6623_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ),
    .S(net260),
    .X(_2510_));
 sg13g2_nor2b_1 _6624_ (.A(net302),
    .B_N(net264),
    .Y(_2511_));
 sg13g2_a21oi_1 _6625_ (.A1(_2510_),
    .A2(_2511_),
    .Y(_2512_),
    .B1(net281));
 sg13g2_o21ai_1 _6626_ (.B1(_2512_),
    .Y(_2513_),
    .A1(net264),
    .A2(_2509_));
 sg13g2_inv_1 _6627_ (.Y(_2514_),
    .A(_0028_));
 sg13g2_nand2_1 _6628_ (.Y(_2515_),
    .A(_2514_),
    .B(_1944_));
 sg13g2_a21oi_1 _6629_ (.A1(net261),
    .A2(_2515_),
    .Y(_2516_),
    .B1(_1432_));
 sg13g2_mux2_1 _6630_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ),
    .S(net260),
    .X(_2517_));
 sg13g2_a22oi_1 _6631_ (.Y(_2518_),
    .B1(_2195_),
    .B2(_2517_),
    .A2(_1900_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ));
 sg13g2_and3_1 _6632_ (.X(_2519_),
    .A(net285),
    .B(_1423_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ));
 sg13g2_a21o_1 _6633_ (.A2(_1962_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ),
    .B1(_2519_),
    .X(_2520_));
 sg13g2_nand2b_1 _6634_ (.Y(_2521_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ),
    .A_N(net302));
 sg13g2_nand3b_1 _6635_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ),
    .C(net304),
    .Y(_2522_),
    .A_N(_1924_));
 sg13g2_o21ai_1 _6636_ (.B1(_2522_),
    .Y(_2523_),
    .A1(net304),
    .A2(_2521_));
 sg13g2_mux2_1 _6637_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ),
    .S(_1890_),
    .X(_2524_));
 sg13g2_and3_1 _6638_ (.X(_2525_),
    .A(_1439_),
    .B(_1950_),
    .C(_2524_));
 sg13g2_a221oi_1 _6639_ (.B2(_1942_),
    .C1(_2525_),
    .B1(_2523_),
    .A1(_2364_),
    .Y(_2526_),
    .A2(_2520_));
 sg13g2_o21ai_1 _6640_ (.B1(_2526_),
    .Y(_2527_),
    .A1(net282),
    .A2(_2518_));
 sg13g2_a22oi_1 _6641_ (.Y(_2528_),
    .B1(_2527_),
    .B2(net261),
    .A2(_2516_),
    .A1(_2513_));
 sg13g2_a21oi_1 _6642_ (.A1(_2506_),
    .A2(_2528_),
    .Y(_2529_),
    .B1(_1979_));
 sg13g2_a221oi_1 _6643_ (.B2(_1851_),
    .C1(_1853_),
    .B1(_1850_),
    .A1(_1785_),
    .Y(_2530_),
    .A2(_1840_));
 sg13g2_nand2b_1 _6644_ (.Y(_2531_),
    .B(_1878_),
    .A_N(_1367_));
 sg13g2_or3_1 _6645_ (.A(_2529_),
    .B(_2530_),
    .C(_2531_),
    .X(_2532_));
 sg13g2_or4_1 _6646_ (.A(_1686_),
    .B(_1817_),
    .C(_2479_),
    .D(_2532_),
    .X(_2533_));
 sg13g2_a21o_1 _6647_ (.A2(_2528_),
    .A1(_2506_),
    .B1(_1979_),
    .X(_2534_));
 sg13g2_a21oi_1 _6648_ (.A1(net319),
    .A2(_1739_),
    .Y(_2535_),
    .B1(_1882_));
 sg13g2_nor2_1 _6649_ (.A(_1997_),
    .B(_2535_),
    .Y(_2536_));
 sg13g2_nor2_1 _6650_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .B(_1878_),
    .Y(_2537_));
 sg13g2_a21o_1 _6651_ (.A2(_2536_),
    .A1(_2534_),
    .B1(_2537_),
    .X(_2538_));
 sg13g2_nand2_1 _6652_ (.Y(_2539_),
    .A(_1795_),
    .B(_1800_));
 sg13g2_a21oi_1 _6653_ (.A1(net277),
    .A2(_2225_),
    .Y(_2540_),
    .B1(_0004_));
 sg13g2_or3_1 _6654_ (.A(_2539_),
    .B(_2540_),
    .C(_2531_),
    .X(_2541_));
 sg13g2_nor4_1 _6655_ (.A(_2529_),
    .B(_2476_),
    .C(_2478_),
    .D(_2541_),
    .Y(_2542_));
 sg13g2_nor3_1 _6656_ (.A(_2539_),
    .B(_2540_),
    .C(_2531_),
    .Y(_2543_));
 sg13g2_and3_1 _6657_ (.X(_2544_),
    .A(_2534_),
    .B(_2530_),
    .C(_2543_));
 sg13g2_nor3_1 _6658_ (.A(_2538_),
    .B(_2542_),
    .C(_2544_),
    .Y(_2545_));
 sg13g2_nand2_1 _6659_ (.Y(_2546_),
    .A(_2533_),
    .B(_2545_));
 sg13g2_nand2b_1 _6660_ (.Y(_2547_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ),
    .A_N(net314));
 sg13g2_nand3b_1 _6661_ (.B(_1415_),
    .C(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ),
    .Y(_2548_),
    .A_N(net300));
 sg13g2_o21ai_1 _6662_ (.B1(_2548_),
    .Y(_2549_),
    .A1(net301),
    .A2(_2547_));
 sg13g2_nor2b_1 _6663_ (.A(_2010_),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ),
    .Y(_2550_));
 sg13g2_a22oi_1 _6664_ (.Y(_2551_),
    .B1(_2550_),
    .B2(_2057_),
    .A2(_2549_),
    .A1(net288));
 sg13g2_nand3_1 _6665_ (.B(net242),
    .C(_2057_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ),
    .Y(_2552_));
 sg13g2_o21ai_1 _6666_ (.B1(_2552_),
    .Y(_2553_),
    .A1(_1397_),
    .A2(_2551_));
 sg13g2_and2_1 _6667_ (.A(_1407_),
    .B(_2553_),
    .X(_2554_));
 sg13g2_a22oi_1 _6668_ (.Y(_2555_),
    .B1(_1419_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ),
    .A2(_2021_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ));
 sg13g2_nand3_1 _6669_ (.B(_1411_),
    .C(_2039_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ),
    .Y(_2556_));
 sg13g2_o21ai_1 _6670_ (.B1(_2556_),
    .Y(_2557_),
    .A1(_2086_),
    .A2(_2555_));
 sg13g2_and2_1 _6671_ (.A(_2032_),
    .B(_2041_),
    .X(_2558_));
 sg13g2_a22oi_1 _6672_ (.Y(_2559_),
    .B1(_2558_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ),
    .A2(_2557_),
    .A1(net258));
 sg13g2_a22oi_1 _6673_ (.Y(_2560_),
    .B1(_2420_),
    .B2(_2487_),
    .A2(_2036_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ));
 sg13g2_nor2b_1 _6674_ (.A(_2560_),
    .B_N(net242),
    .Y(_2561_));
 sg13g2_a22oi_1 _6675_ (.Y(_2562_),
    .B1(_2420_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ),
    .A2(_2036_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ));
 sg13g2_nor2b_1 _6676_ (.A(_2562_),
    .B_N(_2035_),
    .Y(_2563_));
 sg13g2_o21ai_1 _6677_ (.B1(_2019_),
    .Y(_2564_),
    .A1(_2561_),
    .A2(_2563_));
 sg13g2_o21ai_1 _6678_ (.B1(_2564_),
    .Y(_2565_),
    .A1(_2019_),
    .A2(_2559_));
 sg13g2_nand2_1 _6679_ (.Y(_2566_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ),
    .B(_2420_));
 sg13g2_nand3_1 _6680_ (.B(net279),
    .C(_2036_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ),
    .Y(_2567_));
 sg13g2_o21ai_1 _6681_ (.B1(_2567_),
    .Y(_2568_),
    .A1(net259),
    .A2(_2566_));
 sg13g2_nand3_1 _6682_ (.B(_2018_),
    .C(_2030_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ),
    .Y(_2569_));
 sg13g2_nand3_1 _6683_ (.B(_1416_),
    .C(_2041_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ),
    .Y(_2570_));
 sg13g2_nand2_1 _6684_ (.Y(_2571_),
    .A(_2569_),
    .B(_2570_));
 sg13g2_a22oi_1 _6685_ (.Y(_2572_),
    .B1(_2571_),
    .B2(_2035_),
    .A2(_2568_),
    .A1(_2032_));
 sg13g2_a22oi_1 _6686_ (.Y(_2573_),
    .B1(_2007_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ),
    .A2(_2006_),
    .A1(_2514_));
 sg13g2_nor3_1 _6687_ (.A(net287),
    .B(net300),
    .C(_2573_),
    .Y(_2574_));
 sg13g2_a22oi_1 _6688_ (.Y(_2575_),
    .B1(_2064_),
    .B2(_2496_),
    .A2(_2062_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ));
 sg13g2_nor2_1 _6689_ (.A(_2440_),
    .B(_2575_),
    .Y(_2576_));
 sg13g2_o21ai_1 _6690_ (.B1(_1413_),
    .Y(_2577_),
    .A1(_2574_),
    .A2(_2576_));
 sg13g2_a22oi_1 _6691_ (.Y(_2578_),
    .B1(_2041_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ),
    .A2(_2030_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ));
 sg13g2_nand3_1 _6692_ (.B(_2018_),
    .C(_2030_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ),
    .Y(_2579_));
 sg13g2_o21ai_1 _6693_ (.B1(_2579_),
    .Y(_2580_),
    .A1(net259),
    .A2(_2578_));
 sg13g2_nand3_1 _6694_ (.B(_2026_),
    .C(_2051_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ),
    .Y(_2581_));
 sg13g2_nand4_1 _6695_ (.B(net279),
    .C(_2021_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ),
    .Y(_2582_),
    .D(_2006_));
 sg13g2_a21oi_1 _6696_ (.A1(_2581_),
    .A2(_2582_),
    .Y(_2583_),
    .B1(_1412_));
 sg13g2_a21oi_1 _6697_ (.A1(_2067_),
    .A2(_2580_),
    .Y(_2584_),
    .B1(_2583_));
 sg13g2_nand3_1 _6698_ (.B(_2577_),
    .C(_2584_),
    .A(_2572_),
    .Y(_2585_));
 sg13g2_mux2_1 _6699_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ),
    .S(net258),
    .X(_2586_));
 sg13g2_nand3_1 _6700_ (.B(_2053_),
    .C(_2586_),
    .A(_2270_),
    .Y(_2587_));
 sg13g2_nand3_1 _6701_ (.B(net279),
    .C(_2270_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ),
    .Y(_2588_));
 sg13g2_nand3_1 _6702_ (.B(net287),
    .C(_1397_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ),
    .Y(_2589_));
 sg13g2_nand2_1 _6703_ (.Y(_2590_),
    .A(_2588_),
    .B(_2589_));
 sg13g2_nand3_1 _6704_ (.B(net279),
    .C(_2041_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ),
    .Y(_2591_));
 sg13g2_nand3_1 _6705_ (.B(_1416_),
    .C(_2030_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ),
    .Y(_2592_));
 sg13g2_nand2_1 _6706_ (.Y(_2593_),
    .A(_2591_),
    .B(_2592_));
 sg13g2_a22oi_1 _6707_ (.Y(_2594_),
    .B1(_2593_),
    .B2(_1397_),
    .A2(_2590_),
    .A1(_2420_));
 sg13g2_a21oi_1 _6708_ (.A1(_2587_),
    .A2(_2594_),
    .Y(_2595_),
    .B1(_2004_));
 sg13g2_nor4_1 _6709_ (.A(_2554_),
    .B(_2565_),
    .C(_2585_),
    .D(_2595_),
    .Y(_2596_));
 sg13g2_inv_1 _6710_ (.Y(_2597_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i ));
 sg13g2_mux2_1 _6711_ (.A0(_2596_),
    .A1(_2597_),
    .S(_2077_),
    .X(_2598_));
 sg13g2_buf_2 _6712_ (.A(_2598_),
    .X(_2599_));
 sg13g2_or2_1 _6713_ (.X(_2600_),
    .B(_2599_),
    .A(_1993_));
 sg13g2_and2_1 _6714_ (.A(net86),
    .B(_2600_),
    .X(_2601_));
 sg13g2_nand3_1 _6715_ (.B(_2533_),
    .C(_2545_),
    .A(_1993_),
    .Y(_2602_));
 sg13g2_nor3_1 _6716_ (.A(net86),
    .B(_2538_),
    .C(_2599_),
    .Y(_2603_));
 sg13g2_a221oi_1 _6717_ (.B2(_2602_),
    .C1(_2603_),
    .B1(_2601_),
    .A1(_2546_),
    .Y(_2604_),
    .A2(_2599_));
 sg13g2_buf_1 _6718_ (.A(_2604_),
    .X(_2605_));
 sg13g2_xnor2_1 _6719_ (.Y(_2606_),
    .A(_2324_),
    .B(_2605_));
 sg13g2_and2_1 _6720_ (.A(_2148_),
    .B(_2606_),
    .X(_2607_));
 sg13g2_inv_1 _6721_ (.Y(_2608_),
    .A(_2607_));
 sg13g2_nor2_1 _6722_ (.A(net241),
    .B(_2453_),
    .Y(_2609_));
 sg13g2_o21ai_1 _6723_ (.B1(_2462_),
    .Y(_2610_),
    .A1(net97),
    .A2(net52));
 sg13g2_nand2_1 _6724_ (.Y(_2611_),
    .A(net96),
    .B(_2610_));
 sg13g2_a21oi_1 _6725_ (.A1(net97),
    .A2(net52),
    .Y(_2612_),
    .B1(_2460_));
 sg13g2_nand2_1 _6726_ (.Y(_2613_),
    .A(net243),
    .B(_2612_));
 sg13g2_a221oi_1 _6727_ (.B2(_2613_),
    .C1(_2457_),
    .B1(_2611_),
    .A1(_2290_),
    .Y(_2614_),
    .A2(_2313_));
 sg13g2_or4_1 _6728_ (.A(_2138_),
    .B(_2606_),
    .C(_2609_),
    .D(_2614_),
    .X(_2615_));
 sg13g2_nand4_1 _6729_ (.B(_2300_),
    .C(_2311_),
    .A(net50),
    .Y(_2616_),
    .D(_2450_));
 sg13g2_nand4_1 _6730_ (.B(_2300_),
    .C(_2311_),
    .A(net51),
    .Y(_2617_),
    .D(_2450_));
 sg13g2_nand3_1 _6731_ (.B(net50),
    .C(_2450_),
    .A(net51),
    .Y(_2618_));
 sg13g2_and4_1 _6732_ (.A(net52),
    .B(_2616_),
    .C(_2617_),
    .D(_2618_),
    .X(_2619_));
 sg13g2_nand4_1 _6733_ (.B(_2300_),
    .C(_2311_),
    .A(net50),
    .Y(_2620_),
    .D(net52));
 sg13g2_nand4_1 _6734_ (.B(_2300_),
    .C(_2311_),
    .A(net51),
    .Y(_2621_),
    .D(net52));
 sg13g2_nand3_1 _6735_ (.B(net50),
    .C(net52),
    .A(net51),
    .Y(_2622_));
 sg13g2_and4_1 _6736_ (.A(_2447_),
    .B(_2620_),
    .C(_2621_),
    .D(_2622_),
    .X(_2623_));
 sg13g2_a22oi_1 _6737_ (.Y(_2624_),
    .B1(_2623_),
    .B2(_2003_),
    .A2(_2619_),
    .A1(_2002_));
 sg13g2_mux2_1 _6738_ (.A0(_2608_),
    .A1(_2615_),
    .S(_2624_),
    .X(_2625_));
 sg13g2_inv_1 _6739_ (.Y(_2626_),
    .A(_2606_));
 sg13g2_nor4_1 _6740_ (.A(_2138_),
    .B(net241),
    .C(_2453_),
    .D(_2605_),
    .Y(_2627_));
 sg13g2_a221oi_1 _6741_ (.B2(_2607_),
    .C1(_2627_),
    .B1(_2614_),
    .A1(_2142_),
    .Y(_2628_),
    .A2(_2626_));
 sg13g2_nand2_1 _6742_ (.Y(_2629_),
    .A(_2625_),
    .B(_2628_));
 sg13g2_buf_1 _6743_ (.A(_2599_),
    .X(_2630_));
 sg13g2_and2_1 _6744_ (.A(net173),
    .B(net71),
    .X(_2631_));
 sg13g2_nor2_1 _6745_ (.A(net173),
    .B(_2630_),
    .Y(_2632_));
 sg13g2_buf_8 _6746_ (.A(_2546_),
    .X(_2633_));
 sg13g2_mux2_1 _6747_ (.A0(_2631_),
    .A1(_2632_),
    .S(net56),
    .X(_2634_));
 sg13g2_nor3_1 _6748_ (.A(_2324_),
    .B(net56),
    .C(_2630_),
    .Y(_2635_));
 sg13g2_a21oi_1 _6749_ (.A1(net241),
    .A2(_2634_),
    .Y(_2636_),
    .B1(_2635_));
 sg13g2_nor3_1 _6750_ (.A(net86),
    .B(_2139_),
    .C(_2636_),
    .Y(_2637_));
 sg13g2_or2_1 _6751_ (.X(_2638_),
    .B(_2637_),
    .A(_1461_));
 sg13g2_a21oi_1 _6752_ (.A1(net175),
    .A2(_2633_),
    .Y(_2639_),
    .B1(_1492_));
 sg13g2_o21ai_1 _6753_ (.B1(_2639_),
    .Y(_2640_),
    .A1(_2629_),
    .A2(_2638_));
 sg13g2_nand2_1 _6754_ (.Y(_2641_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31] ),
    .B(net74));
 sg13g2_nand2_1 _6755_ (.Y(_1238_),
    .A(_2640_),
    .B(_2641_));
 sg13g2_buf_2 _6756_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[3] ),
    .X(_2642_));
 sg13g2_nand2_1 _6757_ (.Y(_2643_),
    .A(_2642_),
    .B(_1496_));
 sg13g2_o21ai_1 _6758_ (.B1(_2643_),
    .Y(_1239_),
    .A1(_1770_),
    .A2(_1493_));
 sg13g2_nand2_1 _6759_ (.Y(_2644_),
    .A(net305),
    .B(_1496_));
 sg13g2_o21ai_1 _6760_ (.B1(_2644_),
    .Y(_1240_),
    .A1(_1751_),
    .A2(_1493_));
 sg13g2_mux2_1 _6761_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9] ),
    .A1(_1498_),
    .S(_1685_),
    .X(_1241_));
 sg13g2_mux2_1 _6762_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10] ),
    .A1(_1370_),
    .S(net72),
    .X(_1242_));
 sg13g2_mux2_1 _6763_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11] ),
    .A1(net323),
    .S(net72),
    .X(_1243_));
 sg13g2_mux2_1 _6764_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12] ),
    .A1(_1750_),
    .S(_1685_),
    .X(_1244_));
 sg13g2_mux2_1 _6765_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9] ),
    .S(net74),
    .X(_1245_));
 sg13g2_nand4_1 _6766_ (.B(net336),
    .C(_1744_),
    .A(_2116_),
    .Y(_2645_),
    .D(_1859_));
 sg13g2_buf_2 _6767_ (.A(_2645_),
    .X(_2646_));
 sg13g2_nand3_1 _6768_ (.B(net322),
    .C(_2128_),
    .A(_1494_),
    .Y(_2647_));
 sg13g2_o21ai_1 _6769_ (.B1(_2647_),
    .Y(_2648_),
    .A1(_1494_),
    .A2(net322));
 sg13g2_nor2_1 _6770_ (.A(net322),
    .B(_2128_),
    .Y(_2649_));
 sg13g2_a21oi_1 _6771_ (.A1(_1500_),
    .A2(_2648_),
    .Y(_2650_),
    .B1(_2649_));
 sg13g2_inv_1 _6772_ (.Y(_2651_),
    .A(_1824_));
 sg13g2_nor2_1 _6773_ (.A(net327),
    .B(_2651_),
    .Y(_2652_));
 sg13g2_xnor2_1 _6774_ (.Y(_2653_),
    .A(net307),
    .B(net322));
 sg13g2_nand3_1 _6775_ (.B(_2652_),
    .C(_2653_),
    .A(_2128_),
    .Y(_2654_));
 sg13g2_o21ai_1 _6776_ (.B1(_2654_),
    .Y(_2655_),
    .A1(_1824_),
    .A2(_2650_));
 sg13g2_and2_1 _6777_ (.A(_1474_),
    .B(_2655_),
    .X(_2656_));
 sg13g2_inv_1 _6778_ (.Y(_2657_),
    .A(_0042_));
 sg13g2_a21oi_1 _6779_ (.A1(net327),
    .A2(_2657_),
    .Y(_2658_),
    .B1(_2128_));
 sg13g2_nand3_1 _6780_ (.B(_1475_),
    .C(_2128_),
    .A(net307),
    .Y(_2659_));
 sg13g2_o21ai_1 _6781_ (.B1(net330),
    .Y(_2660_),
    .A1(_1824_),
    .A2(_2659_));
 sg13g2_nand4_1 _6782_ (.B(_1475_),
    .C(_2128_),
    .A(net307),
    .Y(_2661_),
    .D(_2652_));
 sg13g2_o21ai_1 _6783_ (.B1(_2661_),
    .Y(_2662_),
    .A1(net330),
    .A2(_2128_));
 sg13g2_a21oi_1 _6784_ (.A1(net327),
    .A2(_2660_),
    .Y(_2663_),
    .B1(_2662_));
 sg13g2_nor4_1 _6785_ (.A(_2646_),
    .B(_2656_),
    .C(_2658_),
    .D(_2663_),
    .Y(_2664_));
 sg13g2_buf_1 _6786_ (.A(_2664_),
    .X(_2665_));
 sg13g2_buf_1 _6787_ (.A(_2665_),
    .X(_2666_));
 sg13g2_and2_1 _6788_ (.A(net230),
    .B(_1470_),
    .X(_2667_));
 sg13g2_buf_2 _6789_ (.A(_2667_),
    .X(_2668_));
 sg13g2_a21oi_1 _6790_ (.A1(net318),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ),
    .Y(_2669_),
    .B1(_1463_));
 sg13g2_buf_2 _6791_ (.A(_2669_),
    .X(_2670_));
 sg13g2_buf_1 _6792_ (.A(_2670_),
    .X(_2671_));
 sg13g2_buf_1 _6793_ (.A(_1467_),
    .X(_2672_));
 sg13g2_buf_1 _6794_ (.A(net257),
    .X(_2673_));
 sg13g2_nand2b_1 _6795_ (.Y(_2674_),
    .B(net239),
    .A_N(\i_exotiny.i_wb_spi.dat_rx_r[4] ));
 sg13g2_o21ai_1 _6796_ (.B1(_2674_),
    .Y(_2675_),
    .A1(_1512_),
    .A2(net239));
 sg13g2_nor2b_1 _6797_ (.A(net305),
    .B_N(_2322_),
    .Y(_2676_));
 sg13g2_nor2b_1 _6798_ (.A(_2642_),
    .B_N(_2676_),
    .Y(_2677_));
 sg13g2_buf_1 _6799_ (.A(_2677_),
    .X(_2678_));
 sg13g2_or2_1 _6800_ (.X(_2679_),
    .B(net305),
    .A(_2322_));
 sg13g2_buf_1 _6801_ (.A(_2679_),
    .X(_2680_));
 sg13g2_and2_1 _6802_ (.A(_2322_),
    .B(_1797_),
    .X(_2681_));
 sg13g2_a21oi_1 _6803_ (.A1(_2642_),
    .A2(_2680_),
    .Y(_2682_),
    .B1(_2681_));
 sg13g2_o21ai_1 _6804_ (.B1(_2682_),
    .Y(_2683_),
    .A1(_2642_),
    .A2(_2680_));
 sg13g2_buf_1 _6805_ (.A(_2683_),
    .X(_2684_));
 sg13g2_a221oi_1 _6806_ (.B2(net31),
    .C1(_2670_),
    .B1(_2684_),
    .A1(net5),
    .Y(_2685_),
    .A2(_2678_));
 sg13g2_a21oi_1 _6807_ (.A1(net240),
    .A2(_2675_),
    .Y(_2686_),
    .B1(_2685_));
 sg13g2_nand2_1 _6808_ (.Y(_2687_),
    .A(net230),
    .B(_1470_));
 sg13g2_buf_1 _6809_ (.A(_2687_),
    .X(_2688_));
 sg13g2_nand2_1 _6810_ (.Y(_2689_),
    .A(net306),
    .B(_0021_));
 sg13g2_buf_1 _6811_ (.A(_0032_),
    .X(_2690_));
 sg13g2_nor2b_1 _6812_ (.A(_1469_),
    .B_N(_2690_),
    .Y(_2691_));
 sg13g2_o21ai_1 _6813_ (.B1(_2691_),
    .Y(_2692_),
    .A1(net329),
    .A2(_2689_));
 sg13g2_and2_1 _6814_ (.A(_2688_),
    .B(_2692_),
    .X(_2693_));
 sg13g2_buf_1 _6815_ (.A(_2693_),
    .X(_2694_));
 sg13g2_buf_1 _6816_ (.A(_2694_),
    .X(_2695_));
 sg13g2_buf_1 _6817_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[4] ),
    .X(_2696_));
 sg13g2_a22oi_1 _6818_ (.Y(_2697_),
    .B1(_2695_),
    .B2(_2696_),
    .A2(_2686_),
    .A1(_2668_));
 sg13g2_inv_1 _6819_ (.Y(_2698_),
    .A(_2665_));
 sg13g2_o21ai_1 _6820_ (.B1(_2698_),
    .Y(_2699_),
    .A1(_2668_),
    .A2(_2692_));
 sg13g2_buf_1 _6821_ (.A(_2699_),
    .X(_2700_));
 sg13g2_buf_1 _6822_ (.A(_2700_),
    .X(_2701_));
 sg13g2_buf_1 _6823_ (.A(net58),
    .X(_2702_));
 sg13g2_nand2_1 _6824_ (.Y(_2703_),
    .A(_1727_),
    .B(_2702_));
 sg13g2_o21ai_1 _6825_ (.B1(_2703_),
    .Y(_1246_),
    .A1(_2666_),
    .A2(_2697_));
 sg13g2_nor2_1 _6826_ (.A(_1465_),
    .B(_2688_),
    .Y(_2704_));
 sg13g2_buf_1 _6827_ (.A(_2704_),
    .X(_2705_));
 sg13g2_buf_1 _6828_ (.A(net85),
    .X(_2706_));
 sg13g2_buf_1 _6829_ (.A(net239),
    .X(_2707_));
 sg13g2_mux2_1 _6830_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[14] ),
    .S(net221),
    .X(_2708_));
 sg13g2_a22oi_1 _6831_ (.Y(_2709_),
    .B1(_2706_),
    .B2(_2708_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ));
 sg13g2_buf_1 _6832_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[10] ),
    .X(_2710_));
 sg13g2_nand2_1 _6833_ (.Y(_2711_),
    .A(_2710_),
    .B(net55));
 sg13g2_o21ai_1 _6834_ (.B1(_2711_),
    .Y(_1247_),
    .A1(net70),
    .A2(_2709_));
 sg13g2_mux2_1 _6835_ (.A0(_1402_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[15] ),
    .S(_2707_),
    .X(_2712_));
 sg13g2_a22oi_1 _6836_ (.Y(_2713_),
    .B1(_2706_),
    .B2(_2712_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ));
 sg13g2_nand2_1 _6837_ (.Y(_2714_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ),
    .B(net55));
 sg13g2_o21ai_1 _6838_ (.B1(_2714_),
    .Y(_1248_),
    .A1(net70),
    .A2(_2713_));
 sg13g2_buf_1 _6839_ (.A(net58),
    .X(_2715_));
 sg13g2_buf_1 _6840_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[16] ),
    .X(_2716_));
 sg13g2_buf_1 _6841_ (.A(_2688_),
    .X(_2717_));
 sg13g2_inv_1 _6842_ (.Y(_2718_),
    .A(_0003_));
 sg13g2_nand3b_1 _6843_ (.B(_1442_),
    .C(_2642_),
    .Y(_2719_),
    .A_N(_2322_));
 sg13g2_buf_1 _6844_ (.A(_2719_),
    .X(_2720_));
 sg13g2_nor2_1 _6845_ (.A(_2670_),
    .B(_2720_),
    .Y(_2721_));
 sg13g2_mux2_1 _6846_ (.A0(_1408_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[16] ),
    .S(net239),
    .X(_2722_));
 sg13g2_a22oi_1 _6847_ (.Y(_2723_),
    .B1(_2722_),
    .B2(net240),
    .A2(_2721_),
    .A1(_2718_));
 sg13g2_nor2_1 _6848_ (.A(net95),
    .B(_2723_),
    .Y(_2724_));
 sg13g2_a21oi_1 _6849_ (.A1(_2716_),
    .A2(net95),
    .Y(_2725_),
    .B1(_2724_));
 sg13g2_nand2_1 _6850_ (.Y(_2726_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ),
    .B(net55));
 sg13g2_o21ai_1 _6851_ (.B1(_2726_),
    .Y(_1249_),
    .A1(net54),
    .A2(_2725_));
 sg13g2_buf_1 _6852_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[17] ),
    .X(_2727_));
 sg13g2_buf_1 _6853_ (.A(_2688_),
    .X(_2728_));
 sg13g2_buf_1 _6854_ (.A(\i_exotiny.i_wb_regs.spi_size_o[1] ),
    .X(_2729_));
 sg13g2_mux2_1 _6855_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[17] ),
    .S(net257),
    .X(_2730_));
 sg13g2_a22oi_1 _6856_ (.Y(_2731_),
    .B1(_2730_),
    .B2(net240),
    .A2(_2721_),
    .A1(_2729_));
 sg13g2_nor2_1 _6857_ (.A(net94),
    .B(_2731_),
    .Y(_2732_));
 sg13g2_a21oi_1 _6858_ (.A1(_2727_),
    .A2(net95),
    .Y(_2733_),
    .B1(_2732_));
 sg13g2_nand2_1 _6859_ (.Y(_2734_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ),
    .B(net55));
 sg13g2_o21ai_1 _6860_ (.B1(_2734_),
    .Y(_1250_),
    .A1(net54),
    .A2(_2733_));
 sg13g2_mux2_1 _6861_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[18] ),
    .S(net221),
    .X(_2735_));
 sg13g2_a22oi_1 _6862_ (.Y(_2736_),
    .B1(net78),
    .B2(_2735_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ));
 sg13g2_nand2_1 _6863_ (.Y(_2737_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ),
    .B(net55));
 sg13g2_o21ai_1 _6864_ (.B1(_2737_),
    .Y(_1251_),
    .A1(net70),
    .A2(_2736_));
 sg13g2_mux2_1 _6865_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .S(net221),
    .X(_2738_));
 sg13g2_a22oi_1 _6866_ (.Y(_2739_),
    .B1(net78),
    .B2(_2738_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ));
 sg13g2_nand2_1 _6867_ (.Y(_2740_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ),
    .B(net55));
 sg13g2_o21ai_1 _6868_ (.B1(_2740_),
    .Y(_1252_),
    .A1(net70),
    .A2(_2739_));
 sg13g2_mux2_1 _6869_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[20] ),
    .S(net221),
    .X(_2741_));
 sg13g2_a22oi_1 _6870_ (.Y(_2742_),
    .B1(net78),
    .B2(_2741_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ));
 sg13g2_buf_1 _6871_ (.A(net58),
    .X(_2743_));
 sg13g2_nand2_1 _6872_ (.Y(_2744_),
    .A(_2716_),
    .B(_2743_));
 sg13g2_o21ai_1 _6873_ (.B1(_2744_),
    .Y(_1253_),
    .A1(net70),
    .A2(_2742_));
 sg13g2_mux2_1 _6874_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[21] ),
    .S(net221),
    .X(_2745_));
 sg13g2_a22oi_1 _6875_ (.Y(_2746_),
    .B1(net78),
    .B2(_2745_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ));
 sg13g2_nand2_1 _6876_ (.Y(_2747_),
    .A(_2727_),
    .B(net53));
 sg13g2_o21ai_1 _6877_ (.B1(_2747_),
    .Y(_1254_),
    .A1(net70),
    .A2(_2746_));
 sg13g2_mux2_1 _6878_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .S(net221),
    .X(_2748_));
 sg13g2_a22oi_1 _6879_ (.Y(_2749_),
    .B1(net78),
    .B2(_2748_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ));
 sg13g2_nand2_1 _6880_ (.Y(_2750_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ),
    .B(net53));
 sg13g2_o21ai_1 _6881_ (.B1(_2750_),
    .Y(_1255_),
    .A1(net70),
    .A2(_2749_));
 sg13g2_mux2_1 _6882_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .S(net221),
    .X(_2751_));
 sg13g2_a22oi_1 _6883_ (.Y(_2752_),
    .B1(net78),
    .B2(_2751_),
    .A2(net79),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ));
 sg13g2_nand2_1 _6884_ (.Y(_2753_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ),
    .B(net53));
 sg13g2_o21ai_1 _6885_ (.B1(_2753_),
    .Y(_1256_),
    .A1(net70),
    .A2(_2752_));
 sg13g2_buf_1 _6886_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[5] ),
    .X(_2754_));
 sg13g2_buf_1 _6887_ (.A(net257),
    .X(_2755_));
 sg13g2_nor2_1 _6888_ (.A(_1528_),
    .B(net239),
    .Y(_2756_));
 sg13g2_a21oi_1 _6889_ (.A1(\i_exotiny.i_wb_spi.dat_rx_r[5] ),
    .A2(net238),
    .Y(_2757_),
    .B1(_2756_));
 sg13g2_a221oi_1 _6890_ (.B2(net32),
    .C1(_2670_),
    .B1(_2684_),
    .A1(net6),
    .Y(_2758_),
    .A2(_2678_));
 sg13g2_a21oi_1 _6891_ (.A1(net240),
    .A2(_2757_),
    .Y(_2759_),
    .B1(_2758_));
 sg13g2_a22oi_1 _6892_ (.Y(_2760_),
    .B1(_2759_),
    .B2(_2668_),
    .A2(_2695_),
    .A1(_2754_));
 sg13g2_nand2_1 _6893_ (.Y(_2761_),
    .A(_1724_),
    .B(_2743_));
 sg13g2_o21ai_1 _6894_ (.B1(_2761_),
    .Y(_1257_),
    .A1(_2666_),
    .A2(_2760_));
 sg13g2_buf_1 _6895_ (.A(_2665_),
    .X(_2762_));
 sg13g2_buf_1 _6896_ (.A(_2694_),
    .X(_2763_));
 sg13g2_mux2_1 _6897_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .S(_2707_),
    .X(_2764_));
 sg13g2_a22oi_1 _6898_ (.Y(_2765_),
    .B1(net78),
    .B2(_2764_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ));
 sg13g2_nand2_1 _6899_ (.Y(_2766_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ),
    .B(net53));
 sg13g2_o21ai_1 _6900_ (.B1(_2766_),
    .Y(_1258_),
    .A1(net69),
    .A2(_2765_));
 sg13g2_mux2_1 _6901_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .S(net221),
    .X(_2767_));
 sg13g2_a22oi_1 _6902_ (.Y(_2768_),
    .B1(net78),
    .B2(_2767_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ));
 sg13g2_nand2_1 _6903_ (.Y(_2769_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ),
    .B(net53));
 sg13g2_o21ai_1 _6904_ (.B1(_2769_),
    .Y(_1259_),
    .A1(net69),
    .A2(_2768_));
 sg13g2_mux2_1 _6905_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .S(net238),
    .X(_2770_));
 sg13g2_a22oi_1 _6906_ (.Y(_2771_),
    .B1(net85),
    .B2(_2770_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ));
 sg13g2_nand2_1 _6907_ (.Y(_2772_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ),
    .B(net53));
 sg13g2_o21ai_1 _6908_ (.B1(_2772_),
    .Y(_1260_),
    .A1(net69),
    .A2(_2771_));
 sg13g2_mux2_1 _6909_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[27] ),
    .S(net238),
    .X(_2773_));
 sg13g2_a22oi_1 _6910_ (.Y(_2774_),
    .B1(net85),
    .B2(_2773_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ));
 sg13g2_nand2_1 _6911_ (.Y(_2775_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ),
    .B(net53));
 sg13g2_o21ai_1 _6912_ (.B1(_2775_),
    .Y(_1261_),
    .A1(net69),
    .A2(_2774_));
 sg13g2_mux2_1 _6913_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[28] ),
    .S(net238),
    .X(_2776_));
 sg13g2_a22oi_1 _6914_ (.Y(_2777_),
    .B1(net85),
    .B2(_2776_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ));
 sg13g2_nand2_1 _6915_ (.Y(_2778_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ),
    .B(net53));
 sg13g2_o21ai_1 _6916_ (.B1(_2778_),
    .Y(_1262_),
    .A1(net69),
    .A2(_2777_));
 sg13g2_mux2_1 _6917_ (.A0(_1502_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .S(net238),
    .X(_2779_));
 sg13g2_a22oi_1 _6918_ (.Y(_2780_),
    .B1(net85),
    .B2(_2779_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ));
 sg13g2_buf_1 _6919_ (.A(_2700_),
    .X(_2781_));
 sg13g2_nand2_1 _6920_ (.Y(_2782_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ),
    .B(net57));
 sg13g2_o21ai_1 _6921_ (.B1(_2782_),
    .Y(_1263_),
    .A1(net69),
    .A2(_2780_));
 sg13g2_mux2_1 _6922_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .S(net238),
    .X(_2783_));
 sg13g2_a22oi_1 _6923_ (.Y(_2784_),
    .B1(net85),
    .B2(_2783_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ));
 sg13g2_nand2_1 _6924_ (.Y(_2785_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ),
    .B(net57));
 sg13g2_o21ai_1 _6925_ (.B1(_2785_),
    .Y(_1264_),
    .A1(net69),
    .A2(_2784_));
 sg13g2_mux2_1 _6926_ (.A0(_1585_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[31] ),
    .S(net238),
    .X(_2786_));
 sg13g2_a22oi_1 _6927_ (.Y(_2787_),
    .B1(net85),
    .B2(_2786_),
    .A2(net77),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ));
 sg13g2_nand2_1 _6928_ (.Y(_2788_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ),
    .B(net57));
 sg13g2_o21ai_1 _6929_ (.B1(_2788_),
    .Y(_1265_),
    .A1(net69),
    .A2(_2787_));
 sg13g2_nand3_1 _6930_ (.B(_2688_),
    .C(_2692_),
    .A(_2698_),
    .Y(_2789_));
 sg13g2_buf_1 _6931_ (.A(_2789_),
    .X(_2790_));
 sg13g2_nor2b_1 _6932_ (.A(_2790_),
    .B_N(_2153_),
    .Y(_2791_));
 sg13g2_a21o_1 _6933_ (.A2(net54),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ),
    .B1(_2791_),
    .X(_1266_));
 sg13g2_nand2_1 _6934_ (.Y(_2792_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ),
    .B(net57));
 sg13g2_o21ai_1 _6935_ (.B1(_2792_),
    .Y(_1267_),
    .A1(_2318_),
    .A2(_2790_));
 sg13g2_nand3_1 _6936_ (.B(_1465_),
    .C(_2678_),
    .A(net7),
    .Y(_2793_));
 sg13g2_mux2_1 _6937_ (.A0(_1515_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[6] ),
    .S(_2672_),
    .X(_2794_));
 sg13g2_nand2_1 _6938_ (.Y(_2795_),
    .A(net240),
    .B(_2794_));
 sg13g2_a21oi_1 _6939_ (.A1(_2793_),
    .A2(_2795_),
    .Y(_2796_),
    .B1(_2728_));
 sg13g2_a21oi_1 _6940_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ),
    .A2(net95),
    .Y(_2797_),
    .B1(_2796_));
 sg13g2_nand2_1 _6941_ (.Y(_2798_),
    .A(_1709_),
    .B(net57));
 sg13g2_o21ai_1 _6942_ (.B1(_2798_),
    .Y(_1268_),
    .A1(net54),
    .A2(_2797_));
 sg13g2_nor2b_1 _6943_ (.A(_2790_),
    .B_N(_2468_),
    .Y(_2799_));
 sg13g2_a21o_1 _6944_ (.A2(net55),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ),
    .B1(_2799_),
    .X(_1269_));
 sg13g2_nor2_1 _6945_ (.A(_2629_),
    .B(_2637_),
    .Y(_2800_));
 sg13g2_nand2_1 _6946_ (.Y(_2801_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ),
    .B(_2781_));
 sg13g2_o21ai_1 _6947_ (.B1(_2801_),
    .Y(_1270_),
    .A1(_2800_),
    .A2(_2790_));
 sg13g2_mux2_1 _6948_ (.A0(_1386_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[7] ),
    .S(_2755_),
    .X(_2802_));
 sg13g2_a22oi_1 _6949_ (.Y(_2803_),
    .B1(net85),
    .B2(_2802_),
    .A2(_2763_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ));
 sg13g2_buf_2 _6950_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[3] ),
    .X(_2804_));
 sg13g2_nand2_1 _6951_ (.Y(_2805_),
    .A(_2804_),
    .B(net57));
 sg13g2_o21ai_1 _6952_ (.B1(_2805_),
    .Y(_1271_),
    .A1(_2762_),
    .A2(_2803_));
 sg13g2_mux2_1 _6953_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[8] ),
    .S(_2755_),
    .X(_2806_));
 sg13g2_a22oi_1 _6954_ (.Y(_2807_),
    .B1(_2705_),
    .B2(_2806_),
    .A2(_2763_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ));
 sg13g2_nand2_1 _6955_ (.Y(_2808_),
    .A(_2696_),
    .B(_2781_));
 sg13g2_o21ai_1 _6956_ (.B1(_2808_),
    .Y(_1272_),
    .A1(_2762_),
    .A2(_2807_));
 sg13g2_buf_1 _6957_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[9] ),
    .X(_2809_));
 sg13g2_mux2_1 _6958_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[9] ),
    .S(net257),
    .X(_2810_));
 sg13g2_a22oi_1 _6959_ (.Y(_2811_),
    .B1(_2810_),
    .B2(_2671_),
    .A2(_2721_),
    .A1(\i_exotiny.i_wb_regs.spi_cpol_o ));
 sg13g2_nor2_1 _6960_ (.A(net94),
    .B(_2811_),
    .Y(_2812_));
 sg13g2_a21oi_1 _6961_ (.A1(_2809_),
    .A2(net95),
    .Y(_2813_),
    .B1(_2812_));
 sg13g2_nand2_1 _6962_ (.Y(_2814_),
    .A(_2754_),
    .B(net57));
 sg13g2_o21ai_1 _6963_ (.B1(_2814_),
    .Y(_1273_),
    .A1(net54),
    .A2(_2813_));
 sg13g2_mux2_1 _6964_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[10] ),
    .S(net257),
    .X(_2815_));
 sg13g2_a22oi_1 _6965_ (.Y(_2816_),
    .B1(_2815_),
    .B2(net240),
    .A2(_2721_),
    .A1(\i_exotiny.i_wb_regs.spi_auto_cs_o ));
 sg13g2_nor2_1 _6966_ (.A(net94),
    .B(_2816_),
    .Y(_2817_));
 sg13g2_a21oi_1 _6967_ (.A1(_2710_),
    .A2(net95),
    .Y(_2818_),
    .B1(_2817_));
 sg13g2_nand2_1 _6968_ (.Y(_2819_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ),
    .B(net57));
 sg13g2_o21ai_1 _6969_ (.B1(_2819_),
    .Y(_1274_),
    .A1(net54),
    .A2(_2818_));
 sg13g2_mux2_1 _6970_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[11] ),
    .S(net238),
    .X(_2820_));
 sg13g2_a22oi_1 _6971_ (.Y(_2821_),
    .B1(_2705_),
    .B2(_2820_),
    .A2(_2694_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ));
 sg13g2_nand2_1 _6972_ (.Y(_2822_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ),
    .B(net58));
 sg13g2_o21ai_1 _6973_ (.B1(_2822_),
    .Y(_1275_),
    .A1(_2665_),
    .A2(_2821_));
 sg13g2_nand2_1 _6974_ (.Y(_2823_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ),
    .B(net94));
 sg13g2_mux2_1 _6975_ (.A0(_1582_),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[12] ),
    .S(net239),
    .X(_2824_));
 sg13g2_nand3_1 _6976_ (.B(_2668_),
    .C(_2824_),
    .A(net240),
    .Y(_2825_));
 sg13g2_a21oi_1 _6977_ (.A1(_2823_),
    .A2(_2825_),
    .Y(_2826_),
    .B1(net58));
 sg13g2_a21o_1 _6978_ (.A2(net55),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ),
    .B1(_2826_),
    .X(_1276_));
 sg13g2_nand2_1 _6979_ (.Y(_2827_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ),
    .B(net94));
 sg13g2_mux2_1 _6980_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[13] ),
    .S(net239),
    .X(_2828_));
 sg13g2_nand3_1 _6981_ (.B(_2668_),
    .C(_2828_),
    .A(net240),
    .Y(_2829_));
 sg13g2_a21oi_1 _6982_ (.A1(_2827_),
    .A2(_2829_),
    .Y(_2830_),
    .B1(net58));
 sg13g2_a21o_1 _6983_ (.A2(_2702_),
    .A1(_2809_),
    .B1(_2830_),
    .X(_1277_));
 sg13g2_mux2_1 _6984_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[0] ),
    .S(net257),
    .X(_2831_));
 sg13g2_nand2b_1 _6985_ (.Y(_2832_),
    .B(net27),
    .A_N(_2682_));
 sg13g2_buf_2 _6986_ (.A(\i_exotiny.i_wb_regs.spi_rdy_i ),
    .X(_2833_));
 sg13g2_and2_1 _6987_ (.A(_2833_),
    .B(_1797_),
    .X(_2834_));
 sg13g2_a21oi_1 _6988_ (.A1(_1442_),
    .A2(net27),
    .Y(_2835_),
    .B1(_2834_));
 sg13g2_nand2_1 _6989_ (.Y(_2836_),
    .A(net1),
    .B(_2676_));
 sg13g2_o21ai_1 _6990_ (.B1(_2836_),
    .Y(_2837_),
    .A1(_2322_),
    .A2(_2835_));
 sg13g2_o21ai_1 _6991_ (.B1(_2642_),
    .Y(_2838_),
    .A1(_0095_),
    .A2(_2680_));
 sg13g2_o21ai_1 _6992_ (.B1(_2838_),
    .Y(_2839_),
    .A1(_2642_),
    .A2(_2837_));
 sg13g2_nand3_1 _6993_ (.B(_2832_),
    .C(_2839_),
    .A(_1465_),
    .Y(_2840_));
 sg13g2_o21ai_1 _6994_ (.B1(_2840_),
    .Y(_2841_),
    .A1(_1465_),
    .A2(_2831_));
 sg13g2_nor2_1 _6995_ (.A(net94),
    .B(_2841_),
    .Y(_2842_));
 sg13g2_a21oi_1 _6996_ (.A1(_1727_),
    .A2(net95),
    .Y(_2843_),
    .B1(_2842_));
 sg13g2_nand2_1 _6997_ (.Y(_2844_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0] ),
    .B(net58));
 sg13g2_o21ai_1 _6998_ (.B1(_2844_),
    .Y(_1278_),
    .A1(net54),
    .A2(_2843_));
 sg13g2_mux2_1 _6999_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[1] ),
    .S(net257),
    .X(_2845_));
 sg13g2_nor2_1 _7000_ (.A(_1465_),
    .B(_2845_),
    .Y(_2846_));
 sg13g2_a21oi_1 _7001_ (.A1(net2),
    .A2(_2678_),
    .Y(_2847_),
    .B1(_2670_));
 sg13g2_o21ai_1 _7002_ (.B1(_2847_),
    .Y(_2848_),
    .A1(_0094_),
    .A2(_2720_));
 sg13g2_a21oi_1 _7003_ (.A1(net28),
    .A2(_2684_),
    .Y(_2849_),
    .B1(_2848_));
 sg13g2_nor3_1 _7004_ (.A(net94),
    .B(_2846_),
    .C(_2849_),
    .Y(_2850_));
 sg13g2_a21oi_1 _7005_ (.A1(_1724_),
    .A2(net95),
    .Y(_2851_),
    .B1(_2850_));
 sg13g2_nand2_1 _7006_ (.Y(_2852_),
    .A(_1732_),
    .B(net58));
 sg13g2_o21ai_1 _7007_ (.B1(_2852_),
    .Y(_1279_),
    .A1(net54),
    .A2(_2851_));
 sg13g2_nand2_1 _7008_ (.Y(_2853_),
    .A(\i_exotiny.i_wb_spi.dat_rx_r[2] ),
    .B(net257));
 sg13g2_o21ai_1 _7009_ (.B1(_2853_),
    .Y(_2854_),
    .A1(_1544_),
    .A2(net239));
 sg13g2_nor2_1 _7010_ (.A(_1465_),
    .B(_2854_),
    .Y(_2855_));
 sg13g2_a21oi_1 _7011_ (.A1(net3),
    .A2(_2678_),
    .Y(_2856_),
    .B1(_2670_));
 sg13g2_o21ai_1 _7012_ (.B1(_2856_),
    .Y(_2857_),
    .A1(_0093_),
    .A2(_2720_));
 sg13g2_a21oi_1 _7013_ (.A1(net29),
    .A2(_2684_),
    .Y(_2858_),
    .B1(_2857_));
 sg13g2_nor3_1 _7014_ (.A(net94),
    .B(_2855_),
    .C(_2858_),
    .Y(_2859_));
 sg13g2_a21oi_1 _7015_ (.A1(_1709_),
    .A2(_2717_),
    .Y(_2860_),
    .B1(_2859_));
 sg13g2_nand2_1 _7016_ (.Y(_2861_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2] ),
    .B(_2701_));
 sg13g2_o21ai_1 _7017_ (.B1(_2861_),
    .Y(_1280_),
    .A1(_2715_),
    .A2(_2860_));
 sg13g2_nor2_1 _7018_ (.A(_1531_),
    .B(_2673_),
    .Y(_2862_));
 sg13g2_a21oi_1 _7019_ (.A1(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .A2(_2673_),
    .Y(_2863_),
    .B1(_2862_));
 sg13g2_inv_1 _7020_ (.Y(_2864_),
    .A(_2720_));
 sg13g2_a221oi_1 _7021_ (.B2(\i_exotiny.i_wb_regs.spi_presc_o[3] ),
    .C1(_2670_),
    .B1(_2864_),
    .A1(net4),
    .Y(_2865_),
    .A2(_2678_));
 sg13g2_nand2_1 _7022_ (.Y(_2866_),
    .A(net30),
    .B(_2684_));
 sg13g2_a221oi_1 _7023_ (.B2(_2866_),
    .C1(_2728_),
    .B1(_2865_),
    .A1(_2671_),
    .Y(_2867_),
    .A2(_2863_));
 sg13g2_a21oi_1 _7024_ (.A1(_2804_),
    .A2(_2717_),
    .Y(_2868_),
    .B1(_2867_));
 sg13g2_nand2_1 _7025_ (.Y(_2869_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3] ),
    .B(_2701_));
 sg13g2_o21ai_1 _7026_ (.B1(_2869_),
    .Y(_1281_),
    .A1(_2715_),
    .A2(_2868_));
 sg13g2_nor2_1 _7027_ (.A(net331),
    .B(net307),
    .Y(_2870_));
 sg13g2_o21ai_1 _7028_ (.B1(_0115_),
    .Y(_2871_),
    .A1(net327),
    .A2(_2870_));
 sg13g2_nor4_2 _7029_ (.A(_1469_),
    .B(_2670_),
    .C(_2646_),
    .Y(_2872_),
    .D(_2720_));
 sg13g2_nand3_1 _7030_ (.B(_2871_),
    .C(_2872_),
    .A(net326),
    .Y(_2873_));
 sg13g2_mux2_1 _7031_ (.A0(_2710_),
    .A1(\i_exotiny.i_wb_regs.spi_auto_cs_o ),
    .S(_2873_),
    .X(_1287_));
 sg13g2_inv_1 _7032_ (.Y(_2874_),
    .A(net327));
 sg13g2_o21ai_1 _7033_ (.B1(_0115_),
    .Y(_2875_),
    .A1(_2874_),
    .A2(_1495_));
 sg13g2_nand3_1 _7034_ (.B(_2872_),
    .C(_2875_),
    .A(net326),
    .Y(_2876_));
 sg13g2_mux2_1 _7035_ (.A0(_2716_),
    .A1(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .S(_2876_),
    .X(_1293_));
 sg13g2_mux2_1 _7036_ (.A0(_2727_),
    .A1(_2729_),
    .S(_2876_),
    .X(_1294_));
 sg13g2_buf_1 _7037_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[0] ),
    .X(_2877_));
 sg13g2_buf_1 _7038_ (.A(\i_exotiny.i_wb_spi.state_r_reg[1] ),
    .X(_2878_));
 sg13g2_inv_1 _7039_ (.Y(_2879_),
    .A(net321));
 sg13g2_buf_1 _7040_ (.A(_2879_),
    .X(_2880_));
 sg13g2_buf_1 _7041_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[0] ),
    .X(_2881_));
 sg13g2_nor3_1 _7042_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[2] ),
    .B(\i_exotiny.i_wb_spi.cnt_presc_r[1] ),
    .C(_2881_),
    .Y(_2882_));
 sg13g2_nor2b_1 _7043_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[3] ),
    .B_N(_2882_),
    .Y(_2883_));
 sg13g2_nor2b_1 _7044_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[4] ),
    .B_N(_2883_),
    .Y(_2884_));
 sg13g2_nor2b_1 _7045_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[5] ),
    .B_N(_2884_),
    .Y(_2885_));
 sg13g2_nor2b_1 _7046_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[6] ),
    .B_N(_2885_),
    .Y(_2886_));
 sg13g2_buf_2 _7047_ (.A(_2886_),
    .X(_2887_));
 sg13g2_nor2_1 _7048_ (.A(_1469_),
    .B(_2646_),
    .Y(_2888_));
 sg13g2_nand3_1 _7049_ (.B(_1467_),
    .C(_2888_),
    .A(_2833_),
    .Y(_2889_));
 sg13g2_buf_2 _7050_ (.A(_2889_),
    .X(_2890_));
 sg13g2_nand2b_1 _7051_ (.Y(_2891_),
    .B(net321),
    .A_N(_2833_));
 sg13g2_and2_1 _7052_ (.A(_2890_),
    .B(_2891_),
    .X(_2892_));
 sg13g2_inv_1 _7053_ (.Y(_2893_),
    .A(_2892_));
 sg13g2_o21ai_1 _7054_ (.B1(_2893_),
    .Y(_2894_),
    .A1(net275),
    .A2(_2887_));
 sg13g2_nand2_1 _7055_ (.Y(_2895_),
    .A(net321),
    .B(_2887_));
 sg13g2_nand2_1 _7056_ (.Y(_2896_),
    .A(_2672_),
    .B(_2888_));
 sg13g2_nand2_1 _7057_ (.Y(_2897_),
    .A(_2833_),
    .B(_2896_));
 sg13g2_nor2b_2 _7058_ (.A(_2895_),
    .B_N(_2897_),
    .Y(_2898_));
 sg13g2_a22oi_1 _7059_ (.Y(_2899_),
    .B1(_2898_),
    .B2(\i_exotiny._2358_[0] ),
    .A2(_2894_),
    .A1(_2877_));
 sg13g2_inv_1 _7060_ (.Y(_1295_),
    .A(_2899_));
 sg13g2_a21o_1 _7061_ (.A2(_2898_),
    .A1(_2877_),
    .B1(_2894_),
    .X(_2900_));
 sg13g2_nor2_1 _7062_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .B(_2877_),
    .Y(_2901_));
 sg13g2_a22oi_1 _7063_ (.Y(_2902_),
    .B1(_2901_),
    .B2(_2898_),
    .A2(_2900_),
    .A1(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ));
 sg13g2_inv_1 _7064_ (.Y(_1296_),
    .A(_2902_));
 sg13g2_xnor2_1 _7065_ (.Y(_2903_),
    .A(_0050_),
    .B(_2901_));
 sg13g2_and2_1 _7066_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ),
    .B(_2894_),
    .X(_2904_));
 sg13g2_a21o_1 _7067_ (.A2(_2903_),
    .A1(_2898_),
    .B1(_2904_),
    .X(_1297_));
 sg13g2_buf_1 _7068_ (.A(net321),
    .X(_2905_));
 sg13g2_nor2_1 _7069_ (.A(net299),
    .B(_2890_),
    .Y(_2906_));
 sg13g2_nand2b_1 _7070_ (.Y(_2907_),
    .B(_2885_),
    .A_N(\i_exotiny.i_wb_spi.cnt_presc_r[6] ));
 sg13g2_a21oi_1 _7071_ (.A1(net321),
    .A2(_2907_),
    .Y(_2908_),
    .B1(_2892_));
 sg13g2_buf_1 _7072_ (.A(_2908_),
    .X(_2909_));
 sg13g2_buf_1 _7073_ (.A(_2909_),
    .X(_2910_));
 sg13g2_nand3_1 _7074_ (.B(net68),
    .C(_2901_),
    .A(_0050_),
    .Y(_2911_));
 sg13g2_xor2_1 _7075_ (.B(_2911_),
    .A(\i_exotiny.i_wb_spi.cnt_hbit_r[3] ),
    .X(_2912_));
 sg13g2_nor2_1 _7076_ (.A(_2906_),
    .B(_2912_),
    .Y(_1298_));
 sg13g2_buf_1 _7077_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[4] ),
    .X(_2913_));
 sg13g2_nor4_2 _7078_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[3] ),
    .B(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ),
    .C(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .Y(_2914_),
    .D(_2877_));
 sg13g2_nand3_1 _7079_ (.B(_2909_),
    .C(_2914_),
    .A(_2913_),
    .Y(_2915_));
 sg13g2_o21ai_1 _7080_ (.B1(_2915_),
    .Y(_2916_),
    .A1(_2913_),
    .A2(_2914_));
 sg13g2_nor2_1 _7081_ (.A(_2913_),
    .B(net68),
    .Y(_2917_));
 sg13g2_a221oi_1 _7082_ (.B2(net299),
    .C1(_2917_),
    .B1(_2916_),
    .A1(_2718_),
    .Y(_1299_),
    .A2(_2906_));
 sg13g2_xnor2_1 _7083_ (.Y(_2918_),
    .A(_2729_),
    .B(\i_exotiny.i_wb_regs.spi_size_o[0] ));
 sg13g2_buf_1 _7084_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ),
    .X(_2919_));
 sg13g2_nor2b_1 _7085_ (.A(_2913_),
    .B_N(_2914_),
    .Y(_2920_));
 sg13g2_nand3_1 _7086_ (.B(_2909_),
    .C(_2920_),
    .A(_2919_),
    .Y(_2921_));
 sg13g2_o21ai_1 _7087_ (.B1(_2921_),
    .Y(_2922_),
    .A1(_2919_),
    .A2(_2920_));
 sg13g2_nor2_1 _7088_ (.A(_2919_),
    .B(net68),
    .Y(_2923_));
 sg13g2_a221oi_1 _7089_ (.B2(net299),
    .C1(_2923_),
    .B1(_2922_),
    .A1(_2906_),
    .Y(_1300_),
    .A2(_2918_));
 sg13g2_nand2_1 _7090_ (.Y(_2924_),
    .A(_2729_),
    .B(\i_exotiny.i_wb_regs.spi_size_o[0] ));
 sg13g2_buf_1 _7091_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[6] ),
    .X(_2925_));
 sg13g2_nor2b_1 _7092_ (.A(_2919_),
    .B_N(_2920_),
    .Y(_2926_));
 sg13g2_nand3_1 _7093_ (.B(_2909_),
    .C(_2926_),
    .A(_2925_),
    .Y(_2927_));
 sg13g2_o21ai_1 _7094_ (.B1(_2927_),
    .Y(_2928_),
    .A1(_2925_),
    .A2(_2926_));
 sg13g2_nor2_1 _7095_ (.A(_2925_),
    .B(net68),
    .Y(_2929_));
 sg13g2_a221oi_1 _7096_ (.B2(net299),
    .C1(_2929_),
    .B1(_2928_),
    .A1(_2906_),
    .Y(_1301_),
    .A2(_2924_));
 sg13g2_nand3_1 _7097_ (.B(_2877_),
    .C(_2887_),
    .A(_2878_),
    .Y(_2930_));
 sg13g2_buf_1 _7098_ (.A(_2930_),
    .X(_2931_));
 sg13g2_buf_1 _7099_ (.A(_2931_),
    .X(_2932_));
 sg13g2_mux2_1 _7100_ (.A0(net8),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[0] ),
    .S(_2932_),
    .X(_1302_));
 sg13g2_mux2_1 _7101_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[9] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[10] ),
    .S(_2932_),
    .X(_1303_));
 sg13g2_mux2_1 _7102_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[10] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[11] ),
    .S(net84),
    .X(_1304_));
 sg13g2_mux2_1 _7103_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[11] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[12] ),
    .S(net84),
    .X(_1305_));
 sg13g2_mux2_1 _7104_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[12] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[13] ),
    .S(net84),
    .X(_1306_));
 sg13g2_mux2_1 _7105_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[13] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[14] ),
    .S(net84),
    .X(_1307_));
 sg13g2_mux2_1 _7106_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[14] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[15] ),
    .S(net84),
    .X(_1308_));
 sg13g2_mux2_1 _7107_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[15] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[16] ),
    .S(net84),
    .X(_1309_));
 sg13g2_mux2_1 _7108_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[16] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[17] ),
    .S(net84),
    .X(_1310_));
 sg13g2_mux2_1 _7109_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[17] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[18] ),
    .S(net84),
    .X(_1311_));
 sg13g2_buf_1 _7110_ (.A(_2931_),
    .X(_2933_));
 sg13g2_mux2_1 _7111_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[18] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .S(net83),
    .X(_1312_));
 sg13g2_mux2_1 _7112_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[0] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[1] ),
    .S(_2933_),
    .X(_1313_));
 sg13g2_mux2_1 _7113_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[20] ),
    .S(net83),
    .X(_1314_));
 sg13g2_mux2_1 _7114_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[20] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[21] ),
    .S(net83),
    .X(_1315_));
 sg13g2_mux2_1 _7115_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[21] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .S(net83),
    .X(_1316_));
 sg13g2_mux2_1 _7116_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .S(net83),
    .X(_1317_));
 sg13g2_mux2_1 _7117_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .S(net83),
    .X(_1318_));
 sg13g2_mux2_1 _7118_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .S(net83),
    .X(_1319_));
 sg13g2_mux2_1 _7119_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .S(net83),
    .X(_1320_));
 sg13g2_mux2_1 _7120_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[27] ),
    .S(_2933_),
    .X(_1321_));
 sg13g2_buf_1 _7121_ (.A(_2931_),
    .X(_2934_));
 sg13g2_mux2_1 _7122_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[27] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[28] ),
    .S(net82),
    .X(_1322_));
 sg13g2_mux2_1 _7123_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[28] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .S(net82),
    .X(_1323_));
 sg13g2_mux2_1 _7124_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[1] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[2] ),
    .S(net82),
    .X(_1324_));
 sg13g2_mux2_1 _7125_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .S(net82),
    .X(_1325_));
 sg13g2_mux2_1 _7126_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[31] ),
    .S(net82),
    .X(_1326_));
 sg13g2_mux2_1 _7127_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[2] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .S(net82),
    .X(_1327_));
 sg13g2_mux2_1 _7128_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[4] ),
    .S(net82),
    .X(_1328_));
 sg13g2_mux2_1 _7129_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[4] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[5] ),
    .S(net82),
    .X(_1329_));
 sg13g2_mux2_1 _7130_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[5] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[6] ),
    .S(_2934_),
    .X(_1330_));
 sg13g2_mux2_1 _7131_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[6] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[7] ),
    .S(_2934_),
    .X(_1331_));
 sg13g2_mux2_1 _7132_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[7] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[8] ),
    .S(_2931_),
    .X(_1332_));
 sg13g2_mux2_1 _7133_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[8] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[9] ),
    .S(_2931_),
    .X(_1333_));
 sg13g2_o21ai_1 _7134_ (.B1(_2909_),
    .Y(_2935_),
    .A1(_2877_),
    .A2(_2895_));
 sg13g2_buf_1 _7135_ (.A(_2935_),
    .X(_2936_));
 sg13g2_buf_1 _7136_ (.A(net66),
    .X(_2937_));
 sg13g2_nor3_1 _7137_ (.A(net299),
    .B(_1728_),
    .C(_2890_),
    .Y(_2938_));
 sg13g2_a21o_1 _7138_ (.A2(_2937_),
    .A1(\i_exotiny.i_wb_spi.dat_tx_r_reg[0] ),
    .B1(_2938_),
    .X(_1334_));
 sg13g2_buf_1 _7139_ (.A(net66),
    .X(_2939_));
 sg13g2_buf_1 _7140_ (.A(net275),
    .X(_2940_));
 sg13g2_and2_1 _7141_ (.A(net299),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[9] ),
    .X(_2941_));
 sg13g2_a21oi_1 _7142_ (.A1(net256),
    .A2(_2710_),
    .Y(_2942_),
    .B1(_2941_));
 sg13g2_nand2_1 _7143_ (.Y(_2943_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[10] ),
    .B(net65));
 sg13g2_o21ai_1 _7144_ (.B1(_2943_),
    .Y(_1335_),
    .A1(net64),
    .A2(_2942_));
 sg13g2_and2_1 _7145_ (.A(net299),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[10] ),
    .X(_2944_));
 sg13g2_a21oi_1 _7146_ (.A1(net256),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ),
    .Y(_2945_),
    .B1(_2944_));
 sg13g2_nand2_1 _7147_ (.Y(_2946_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[11] ),
    .B(net65));
 sg13g2_o21ai_1 _7148_ (.B1(_2946_),
    .Y(_1336_),
    .A1(net64),
    .A2(_2945_));
 sg13g2_buf_1 _7149_ (.A(net321),
    .X(_2947_));
 sg13g2_and2_1 _7150_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[11] ),
    .X(_2948_));
 sg13g2_a21oi_1 _7151_ (.A1(_2940_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ),
    .Y(_2949_),
    .B1(_2948_));
 sg13g2_nand2_1 _7152_ (.Y(_2950_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[12] ),
    .B(net65));
 sg13g2_o21ai_1 _7153_ (.B1(_2950_),
    .Y(_1337_),
    .A1(_2939_),
    .A2(_2949_));
 sg13g2_and2_1 _7154_ (.A(_2947_),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[12] ),
    .X(_2951_));
 sg13g2_a21oi_1 _7155_ (.A1(_2940_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ),
    .Y(_2952_),
    .B1(_2951_));
 sg13g2_nand2_1 _7156_ (.Y(_2953_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[13] ),
    .B(net65));
 sg13g2_o21ai_1 _7157_ (.B1(_2953_),
    .Y(_1338_),
    .A1(_2939_),
    .A2(_2952_));
 sg13g2_and2_1 _7158_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[13] ),
    .X(_2954_));
 sg13g2_a21oi_1 _7159_ (.A1(net256),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ),
    .Y(_2955_),
    .B1(_2954_));
 sg13g2_nand2_1 _7160_ (.Y(_2956_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[14] ),
    .B(net65));
 sg13g2_o21ai_1 _7161_ (.B1(_2956_),
    .Y(_1339_),
    .A1(net64),
    .A2(_2955_));
 sg13g2_and2_1 _7162_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[14] ),
    .X(_2957_));
 sg13g2_a21oi_1 _7163_ (.A1(net256),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ),
    .Y(_2958_),
    .B1(_2957_));
 sg13g2_nand2_1 _7164_ (.Y(_2959_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[15] ),
    .B(net65));
 sg13g2_o21ai_1 _7165_ (.B1(_2959_),
    .Y(_1340_),
    .A1(net64),
    .A2(_2958_));
 sg13g2_and2_1 _7166_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[15] ),
    .X(_2960_));
 sg13g2_a21oi_1 _7167_ (.A1(net256),
    .A2(_2716_),
    .Y(_2961_),
    .B1(_2960_));
 sg13g2_nand2_1 _7168_ (.Y(_2962_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[16] ),
    .B(net65));
 sg13g2_o21ai_1 _7169_ (.B1(_2962_),
    .Y(_1341_),
    .A1(net64),
    .A2(_2961_));
 sg13g2_and2_1 _7170_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[16] ),
    .X(_2963_));
 sg13g2_a21oi_1 _7171_ (.A1(net256),
    .A2(_2727_),
    .Y(_2964_),
    .B1(_2963_));
 sg13g2_nand2_1 _7172_ (.Y(_2965_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[17] ),
    .B(net65));
 sg13g2_o21ai_1 _7173_ (.B1(_2965_),
    .Y(_1342_),
    .A1(net64),
    .A2(_2964_));
 sg13g2_and2_1 _7174_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[17] ),
    .X(_2966_));
 sg13g2_a21oi_1 _7175_ (.A1(net256),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ),
    .Y(_2967_),
    .B1(_2966_));
 sg13g2_buf_1 _7176_ (.A(net66),
    .X(_2968_));
 sg13g2_nand2_1 _7177_ (.Y(_2969_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[18] ),
    .B(_2968_));
 sg13g2_o21ai_1 _7178_ (.B1(_2969_),
    .Y(_1343_),
    .A1(net64),
    .A2(_2967_));
 sg13g2_and2_1 _7179_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[18] ),
    .X(_2970_));
 sg13g2_a21oi_1 _7180_ (.A1(net256),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ),
    .Y(_2971_),
    .B1(_2970_));
 sg13g2_nand2_1 _7181_ (.Y(_2972_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[19] ),
    .B(net63));
 sg13g2_o21ai_1 _7182_ (.B1(_2972_),
    .Y(_1344_),
    .A1(net64),
    .A2(_2971_));
 sg13g2_buf_1 _7183_ (.A(net66),
    .X(_2973_));
 sg13g2_buf_1 _7184_ (.A(net275),
    .X(_2974_));
 sg13g2_and2_1 _7185_ (.A(_2947_),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[0] ),
    .X(_2975_));
 sg13g2_a21oi_1 _7186_ (.A1(net255),
    .A2(_1724_),
    .Y(_2976_),
    .B1(_2975_));
 sg13g2_nand2_1 _7187_ (.Y(_2977_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[1] ),
    .B(net63));
 sg13g2_o21ai_1 _7188_ (.B1(_2977_),
    .Y(_1345_),
    .A1(net62),
    .A2(_2976_));
 sg13g2_and2_1 _7189_ (.A(net298),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[19] ),
    .X(_2978_));
 sg13g2_a21oi_1 _7190_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ),
    .Y(_2979_),
    .B1(_2978_));
 sg13g2_nand2_1 _7191_ (.Y(_2980_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[20] ),
    .B(net63));
 sg13g2_o21ai_1 _7192_ (.B1(_2980_),
    .Y(_1346_),
    .A1(net62),
    .A2(_2979_));
 sg13g2_buf_1 _7193_ (.A(net321),
    .X(_2981_));
 sg13g2_and2_1 _7194_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[20] ),
    .X(_2982_));
 sg13g2_a21oi_1 _7195_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ),
    .Y(_2983_),
    .B1(_2982_));
 sg13g2_nand2_1 _7196_ (.Y(_2984_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[21] ),
    .B(net63));
 sg13g2_o21ai_1 _7197_ (.B1(_2984_),
    .Y(_1347_),
    .A1(net62),
    .A2(_2983_));
 sg13g2_and2_1 _7198_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[21] ),
    .X(_2985_));
 sg13g2_a21oi_1 _7199_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ),
    .Y(_2986_),
    .B1(_2985_));
 sg13g2_nand2_1 _7200_ (.Y(_2987_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[22] ),
    .B(net63));
 sg13g2_o21ai_1 _7201_ (.B1(_2987_),
    .Y(_1348_),
    .A1(net62),
    .A2(_2986_));
 sg13g2_and2_1 _7202_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[22] ),
    .X(_2988_));
 sg13g2_a21oi_1 _7203_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ),
    .Y(_2989_),
    .B1(_2988_));
 sg13g2_nand2_1 _7204_ (.Y(_2990_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[23] ),
    .B(net63));
 sg13g2_o21ai_1 _7205_ (.B1(_2990_),
    .Y(_1349_),
    .A1(net62),
    .A2(_2989_));
 sg13g2_and2_1 _7206_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[23] ),
    .X(_2991_));
 sg13g2_a21oi_1 _7207_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ),
    .Y(_2992_),
    .B1(_2991_));
 sg13g2_nand2_1 _7208_ (.Y(_2993_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[24] ),
    .B(net63));
 sg13g2_o21ai_1 _7209_ (.B1(_2993_),
    .Y(_1350_),
    .A1(net62),
    .A2(_2992_));
 sg13g2_and2_1 _7210_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[24] ),
    .X(_2994_));
 sg13g2_a21oi_1 _7211_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ),
    .Y(_2995_),
    .B1(_2994_));
 sg13g2_nand2_1 _7212_ (.Y(_2996_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[25] ),
    .B(net63));
 sg13g2_o21ai_1 _7213_ (.B1(_2996_),
    .Y(_1351_),
    .A1(net62),
    .A2(_2995_));
 sg13g2_and2_1 _7214_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[25] ),
    .X(_2997_));
 sg13g2_a21oi_1 _7215_ (.A1(_2974_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ),
    .Y(_2998_),
    .B1(_2997_));
 sg13g2_nand2_1 _7216_ (.Y(_2999_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[26] ),
    .B(_2968_));
 sg13g2_o21ai_1 _7217_ (.B1(_2999_),
    .Y(_1352_),
    .A1(_2973_),
    .A2(_2998_));
 sg13g2_and2_1 _7218_ (.A(_2981_),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[26] ),
    .X(_3000_));
 sg13g2_a21oi_1 _7219_ (.A1(_2974_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ),
    .Y(_3001_),
    .B1(_3000_));
 sg13g2_buf_1 _7220_ (.A(net66),
    .X(_3002_));
 sg13g2_nand2_1 _7221_ (.Y(_3003_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[27] ),
    .B(net61));
 sg13g2_o21ai_1 _7222_ (.B1(_3003_),
    .Y(_1353_),
    .A1(net62),
    .A2(_3001_));
 sg13g2_and2_1 _7223_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[27] ),
    .X(_3004_));
 sg13g2_a21oi_1 _7224_ (.A1(net255),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ),
    .Y(_3005_),
    .B1(_3004_));
 sg13g2_nand2_1 _7225_ (.Y(_3006_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[28] ),
    .B(net61));
 sg13g2_o21ai_1 _7226_ (.B1(_3006_),
    .Y(_1354_),
    .A1(_2973_),
    .A2(_3005_));
 sg13g2_buf_1 _7227_ (.A(net66),
    .X(_3007_));
 sg13g2_buf_1 _7228_ (.A(net275),
    .X(_3008_));
 sg13g2_and2_1 _7229_ (.A(net297),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[28] ),
    .X(_3009_));
 sg13g2_a21oi_1 _7230_ (.A1(net254),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ),
    .Y(_3010_),
    .B1(_3009_));
 sg13g2_nand2_1 _7231_ (.Y(_3011_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[29] ),
    .B(net61));
 sg13g2_o21ai_1 _7232_ (.B1(_3011_),
    .Y(_1355_),
    .A1(net60),
    .A2(_3010_));
 sg13g2_and2_1 _7233_ (.A(_2981_),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[1] ),
    .X(_3012_));
 sg13g2_a21oi_1 _7234_ (.A1(net254),
    .A2(_1709_),
    .Y(_3013_),
    .B1(_3012_));
 sg13g2_nand2_1 _7235_ (.Y(_3014_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[2] ),
    .B(net61));
 sg13g2_o21ai_1 _7236_ (.B1(_3014_),
    .Y(_1356_),
    .A1(net60),
    .A2(_3013_));
 sg13g2_buf_1 _7237_ (.A(net321),
    .X(_3015_));
 sg13g2_and2_1 _7238_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[29] ),
    .X(_3016_));
 sg13g2_a21oi_1 _7239_ (.A1(net254),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ),
    .Y(_3017_),
    .B1(_3016_));
 sg13g2_nand2_1 _7240_ (.Y(_3018_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[30] ),
    .B(net61));
 sg13g2_o21ai_1 _7241_ (.B1(_3018_),
    .Y(_1357_),
    .A1(net60),
    .A2(_3017_));
 sg13g2_and2_1 _7242_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[2] ),
    .X(_3019_));
 sg13g2_a21oi_1 _7243_ (.A1(net254),
    .A2(_2804_),
    .Y(_3020_),
    .B1(_3019_));
 sg13g2_nand2_1 _7244_ (.Y(_3021_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[3] ),
    .B(net61));
 sg13g2_o21ai_1 _7245_ (.B1(_3021_),
    .Y(_1358_),
    .A1(net60),
    .A2(_3020_));
 sg13g2_and2_1 _7246_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[3] ),
    .X(_3022_));
 sg13g2_a21oi_1 _7247_ (.A1(net254),
    .A2(_2696_),
    .Y(_3023_),
    .B1(_3022_));
 sg13g2_nand2_1 _7248_ (.Y(_3024_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[4] ),
    .B(net61));
 sg13g2_o21ai_1 _7249_ (.B1(_3024_),
    .Y(_1359_),
    .A1(net60),
    .A2(_3023_));
 sg13g2_and2_1 _7250_ (.A(_3015_),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[4] ),
    .X(_3025_));
 sg13g2_a21oi_1 _7251_ (.A1(net254),
    .A2(_2754_),
    .Y(_3026_),
    .B1(_3025_));
 sg13g2_nand2_1 _7252_ (.Y(_3027_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[5] ),
    .B(net61));
 sg13g2_o21ai_1 _7253_ (.B1(_3027_),
    .Y(_1360_),
    .A1(net60),
    .A2(_3026_));
 sg13g2_and2_1 _7254_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[5] ),
    .X(_3028_));
 sg13g2_a21oi_1 _7255_ (.A1(_3008_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ),
    .Y(_3029_),
    .B1(_3028_));
 sg13g2_nand2_1 _7256_ (.Y(_3030_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[6] ),
    .B(_3002_));
 sg13g2_o21ai_1 _7257_ (.B1(_3030_),
    .Y(_1361_),
    .A1(_3007_),
    .A2(_3029_));
 sg13g2_and2_1 _7258_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[6] ),
    .X(_3031_));
 sg13g2_a21oi_1 _7259_ (.A1(net254),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ),
    .Y(_3032_),
    .B1(_3031_));
 sg13g2_nand2_1 _7260_ (.Y(_3033_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[7] ),
    .B(_3002_));
 sg13g2_o21ai_1 _7261_ (.B1(_3033_),
    .Y(_1362_),
    .A1(net60),
    .A2(_3032_));
 sg13g2_and2_1 _7262_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[7] ),
    .X(_3034_));
 sg13g2_a21oi_1 _7263_ (.A1(net254),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ),
    .Y(_3035_),
    .B1(_3034_));
 sg13g2_nand2_1 _7264_ (.Y(_3036_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[8] ),
    .B(net66));
 sg13g2_o21ai_1 _7265_ (.B1(_3036_),
    .Y(_1363_),
    .A1(net60),
    .A2(_3035_));
 sg13g2_and2_1 _7266_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[8] ),
    .X(_3037_));
 sg13g2_a21oi_1 _7267_ (.A1(_3008_),
    .A2(_2809_),
    .Y(_3038_),
    .B1(_3037_));
 sg13g2_nand2_1 _7268_ (.Y(_3039_),
    .A(\i_exotiny.i_wb_spi.dat_tx_r_reg[9] ),
    .B(_2936_));
 sg13g2_o21ai_1 _7269_ (.B1(_3039_),
    .Y(_1364_),
    .A1(_3007_),
    .A2(_3038_));
 sg13g2_inv_1 _7270_ (.Y(_3040_),
    .A(_1503_));
 sg13g2_buf_2 _7271_ (.A(_3040_),
    .X(_3041_));
 sg13g2_nor2_1 _7272_ (.A(_2833_),
    .B(_3041_),
    .Y(_3042_));
 sg13g2_nor2b_1 _7273_ (.A(_2925_),
    .B_N(_2926_),
    .Y(_3043_));
 sg13g2_o21ai_1 _7274_ (.B1(_3015_),
    .Y(_3044_),
    .A1(_0092_),
    .A2(_3043_));
 sg13g2_nand3b_1 _7275_ (.B(_2887_),
    .C(_3044_),
    .Y(_3045_),
    .A_N(_0002_));
 sg13g2_o21ai_1 _7276_ (.B1(_3045_),
    .Y(_3046_),
    .A1(\i_exotiny.spi_sck_o ),
    .A2(_2887_));
 sg13g2_o21ai_1 _7277_ (.B1(_3042_),
    .Y(_3047_),
    .A1(_2907_),
    .A2(_3044_));
 sg13g2_inv_1 _7278_ (.Y(_3048_),
    .A(\i_exotiny.i_wb_regs.spi_cpol_o ));
 sg13g2_a22oi_1 _7279_ (.Y(_1365_),
    .B1(_3047_),
    .B2(_3048_),
    .A2(_3046_),
    .A1(_3042_));
 sg13g2_and2_1 _7280_ (.A(net296),
    .B(\i_exotiny.i_wb_spi.dat_tx_r_reg[30] ),
    .X(_3049_));
 sg13g2_a21oi_1 _7281_ (.A1(net275),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ),
    .Y(_3050_),
    .B1(_3049_));
 sg13g2_nand2_1 _7282_ (.Y(_3051_),
    .A(\i_exotiny.spi_sdo_o ),
    .B(net66));
 sg13g2_o21ai_1 _7283_ (.B1(_3051_),
    .Y(_1366_),
    .A1(_2937_),
    .A2(_3050_));
 sg13g2_inv_1 _7284_ (.Y(_3052_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0] ));
 sg13g2_buf_1 _7285_ (.A(_1487_),
    .X(_3053_));
 sg13g2_buf_1 _7286_ (.A(net237),
    .X(_3054_));
 sg13g2_buf_1 _7287_ (.A(net220),
    .X(_3055_));
 sg13g2_buf_1 _7288_ (.A(net237),
    .X(_3056_));
 sg13g2_nand2_1 _7289_ (.Y(_3057_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4] ),
    .B(net219));
 sg13g2_o21ai_1 _7290_ (.B1(_3057_),
    .Y(_0122_),
    .A1(_3052_),
    .A2(net172));
 sg13g2_buf_1 _7291_ (.A(net220),
    .X(_3058_));
 sg13g2_mux2_1 _7292_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5] ),
    .S(net171),
    .X(_0123_));
 sg13g2_mux2_1 _7293_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6] ),
    .S(net171),
    .X(_0124_));
 sg13g2_mux2_1 _7294_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7] ),
    .S(net171),
    .X(_0125_));
 sg13g2_buf_1 _7295_ (.A(_3054_),
    .X(_3059_));
 sg13g2_mux2_1 _7296_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4] ),
    .S(net170),
    .X(_0126_));
 sg13g2_mux2_1 _7297_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5] ),
    .S(_3059_),
    .X(_0127_));
 sg13g2_mux2_1 _7298_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6] ),
    .S(net170),
    .X(_0128_));
 sg13g2_mux2_1 _7299_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7] ),
    .S(_3059_),
    .X(_0129_));
 sg13g2_inv_1 _7300_ (.Y(_3060_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0] ));
 sg13g2_nand2_1 _7301_ (.Y(_3061_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4] ),
    .B(net219));
 sg13g2_o21ai_1 _7302_ (.B1(_3061_),
    .Y(_0130_),
    .A1(_3060_),
    .A2(net172));
 sg13g2_mux2_1 _7303_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5] ),
    .S(net170),
    .X(_0131_));
 sg13g2_mux2_1 _7304_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6] ),
    .S(net170),
    .X(_0132_));
 sg13g2_mux2_1 _7305_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7] ),
    .S(net170),
    .X(_0133_));
 sg13g2_mux2_1 _7306_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4] ),
    .S(net170),
    .X(_0134_));
 sg13g2_mux2_1 _7307_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5] ),
    .S(net170),
    .X(_0135_));
 sg13g2_mux2_1 _7308_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6] ),
    .S(net170),
    .X(_0136_));
 sg13g2_buf_2 _7309_ (.A(_1487_),
    .X(_3062_));
 sg13g2_buf_2 _7310_ (.A(_3062_),
    .X(_3063_));
 sg13g2_buf_1 _7311_ (.A(_3063_),
    .X(_3064_));
 sg13g2_mux2_1 _7312_ (.A0(_2496_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7] ),
    .S(net169),
    .X(_0137_));
 sg13g2_inv_1 _7313_ (.Y(_3065_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0] ));
 sg13g2_nand2_1 _7314_ (.Y(_3066_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4] ),
    .B(net219));
 sg13g2_o21ai_1 _7315_ (.B1(_3066_),
    .Y(_0138_),
    .A1(_3065_),
    .A2(net172));
 sg13g2_mux2_1 _7316_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5] ),
    .S(_3064_),
    .X(_0139_));
 sg13g2_mux2_1 _7317_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6] ),
    .S(net169),
    .X(_0140_));
 sg13g2_mux2_1 _7318_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7] ),
    .S(net169),
    .X(_0141_));
 sg13g2_buf_1 _7319_ (.A(_1487_),
    .X(_3067_));
 sg13g2_buf_1 _7320_ (.A(_3067_),
    .X(_3068_));
 sg13g2_nand2_1 _7321_ (.Y(_3069_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7322_ (.B1(_3069_),
    .Y(_0142_),
    .A1(_1922_),
    .A2(net172));
 sg13g2_mux2_1 _7323_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5] ),
    .S(net169),
    .X(_0143_));
 sg13g2_mux2_1 _7324_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6] ),
    .S(net169),
    .X(_0144_));
 sg13g2_mux2_1 _7325_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7] ),
    .S(net169),
    .X(_0145_));
 sg13g2_nand2_1 _7326_ (.Y(_3070_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7327_ (.B1(_3070_),
    .Y(_0146_),
    .A1(_2015_),
    .A2(net172));
 sg13g2_mux2_1 _7328_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5] ),
    .S(_3064_),
    .X(_0147_));
 sg13g2_mux2_1 _7329_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6] ),
    .S(net169),
    .X(_0148_));
 sg13g2_mux2_1 _7330_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7] ),
    .S(net169),
    .X(_0149_));
 sg13g2_buf_1 _7331_ (.A(_3063_),
    .X(_3071_));
 sg13g2_mux2_1 _7332_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4] ),
    .S(net168),
    .X(_0150_));
 sg13g2_mux2_1 _7333_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5] ),
    .S(net168),
    .X(_0151_));
 sg13g2_nand2_1 _7334_ (.Y(_3072_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6] ),
    .B(net218));
 sg13g2_o21ai_1 _7335_ (.B1(_3072_),
    .Y(_0152_),
    .A1(_2423_),
    .A2(net172));
 sg13g2_mux2_1 _7336_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7] ),
    .S(_3071_),
    .X(_0153_));
 sg13g2_nand2_1 _7337_ (.Y(_3073_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7338_ (.B1(_3073_),
    .Y(_0154_),
    .A1(_2068_),
    .A2(net172));
 sg13g2_mux2_1 _7339_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5] ),
    .S(net168),
    .X(_0155_));
 sg13g2_mux2_1 _7340_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6] ),
    .S(net168),
    .X(_0156_));
 sg13g2_mux2_1 _7341_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7] ),
    .S(_3071_),
    .X(_0157_));
 sg13g2_inv_1 _7342_ (.Y(_3074_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0] ));
 sg13g2_nand2_1 _7343_ (.Y(_3075_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7344_ (.B1(_3075_),
    .Y(_0158_),
    .A1(_3074_),
    .A2(_3055_));
 sg13g2_mux2_1 _7345_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5] ),
    .S(net168),
    .X(_0159_));
 sg13g2_mux2_1 _7346_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6] ),
    .S(net168),
    .X(_0160_));
 sg13g2_mux2_1 _7347_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7] ),
    .S(net168),
    .X(_0161_));
 sg13g2_mux2_1 _7348_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4] ),
    .S(net168),
    .X(_0162_));
 sg13g2_buf_1 _7349_ (.A(_3063_),
    .X(_3076_));
 sg13g2_mux2_1 _7350_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5] ),
    .S(net167),
    .X(_0163_));
 sg13g2_nand2_1 _7351_ (.Y(_3077_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6] ),
    .B(_3068_));
 sg13g2_o21ai_1 _7352_ (.B1(_3077_),
    .Y(_0164_),
    .A1(_2437_),
    .A2(_3055_));
 sg13g2_mux2_1 _7353_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7] ),
    .S(net167),
    .X(_0165_));
 sg13g2_inv_1 _7354_ (.Y(_3078_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0] ));
 sg13g2_nand2_1 _7355_ (.Y(_3079_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7356_ (.B1(_3079_),
    .Y(_0166_),
    .A1(_3078_),
    .A2(net172));
 sg13g2_mux2_1 _7357_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5] ),
    .S(net167),
    .X(_0167_));
 sg13g2_mux2_1 _7358_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6] ),
    .S(net167),
    .X(_0168_));
 sg13g2_mux2_1 _7359_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7] ),
    .S(net167),
    .X(_0169_));
 sg13g2_buf_1 _7360_ (.A(_3054_),
    .X(_3080_));
 sg13g2_nand2_1 _7361_ (.Y(_3081_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7362_ (.B1(_3081_),
    .Y(_0170_),
    .A1(_1925_),
    .A2(net166));
 sg13g2_mux2_1 _7363_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5] ),
    .S(net167),
    .X(_0171_));
 sg13g2_mux2_1 _7364_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6] ),
    .S(net167),
    .X(_0172_));
 sg13g2_mux2_1 _7365_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7] ),
    .S(_3076_),
    .X(_0173_));
 sg13g2_inv_1 _7366_ (.Y(_3082_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0] ));
 sg13g2_nand2_1 _7367_ (.Y(_3083_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4] ),
    .B(_3068_));
 sg13g2_o21ai_1 _7368_ (.B1(_3083_),
    .Y(_0174_),
    .A1(_3082_),
    .A2(net166));
 sg13g2_mux2_1 _7369_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5] ),
    .S(net167),
    .X(_0175_));
 sg13g2_mux2_1 _7370_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6] ),
    .S(_3076_),
    .X(_0176_));
 sg13g2_buf_1 _7371_ (.A(_3063_),
    .X(_3084_));
 sg13g2_mux2_1 _7372_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7] ),
    .S(net165),
    .X(_0177_));
 sg13g2_mux2_1 _7373_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4] ),
    .S(net165),
    .X(_0178_));
 sg13g2_mux2_1 _7374_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5] ),
    .S(net165),
    .X(_0179_));
 sg13g2_mux2_1 _7375_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6] ),
    .S(net165),
    .X(_0180_));
 sg13g2_mux2_1 _7376_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7] ),
    .S(_3084_),
    .X(_0181_));
 sg13g2_inv_1 _7377_ (.Y(_3085_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0] ));
 sg13g2_nand2_1 _7378_ (.Y(_3086_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4] ),
    .B(net218));
 sg13g2_o21ai_1 _7379_ (.B1(_3086_),
    .Y(_0182_),
    .A1(_3085_),
    .A2(net166));
 sg13g2_mux2_1 _7380_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5] ),
    .S(net165),
    .X(_0183_));
 sg13g2_mux2_1 _7381_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6] ),
    .S(net165),
    .X(_0184_));
 sg13g2_mux2_1 _7382_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7] ),
    .S(net165),
    .X(_0185_));
 sg13g2_mux2_1 _7383_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4] ),
    .S(_3084_),
    .X(_0186_));
 sg13g2_mux2_1 _7384_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5] ),
    .S(net165),
    .X(_0187_));
 sg13g2_buf_1 _7385_ (.A(_3063_),
    .X(_3087_));
 sg13g2_mux2_1 _7386_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6] ),
    .S(net164),
    .X(_0188_));
 sg13g2_mux2_1 _7387_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7] ),
    .S(net164),
    .X(_0189_));
 sg13g2_inv_1 _7388_ (.Y(_3088_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0] ));
 sg13g2_buf_1 _7389_ (.A(_3067_),
    .X(_3089_));
 sg13g2_nand2_1 _7390_ (.Y(_3090_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4] ),
    .B(_3089_));
 sg13g2_o21ai_1 _7391_ (.B1(_3090_),
    .Y(_0190_),
    .A1(_3088_),
    .A2(_3080_));
 sg13g2_mux2_1 _7392_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5] ),
    .S(net164),
    .X(_0191_));
 sg13g2_mux2_1 _7393_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6] ),
    .S(_3087_),
    .X(_0192_));
 sg13g2_mux2_1 _7394_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7] ),
    .S(net164),
    .X(_0193_));
 sg13g2_inv_1 _7395_ (.Y(_3091_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0] ));
 sg13g2_nand2_1 _7396_ (.Y(_3092_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7397_ (.B1(_3092_),
    .Y(_0194_),
    .A1(_3091_),
    .A2(_3080_));
 sg13g2_mux2_1 _7398_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5] ),
    .S(_3087_),
    .X(_0195_));
 sg13g2_mux2_1 _7399_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6] ),
    .S(net164),
    .X(_0196_));
 sg13g2_mux2_1 _7400_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7] ),
    .S(net164),
    .X(_0197_));
 sg13g2_inv_1 _7401_ (.Y(_3093_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0] ));
 sg13g2_nand2_1 _7402_ (.Y(_3094_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4] ),
    .B(_3089_));
 sg13g2_o21ai_1 _7403_ (.B1(_3094_),
    .Y(_0198_),
    .A1(_3093_),
    .A2(net166));
 sg13g2_mux2_1 _7404_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5] ),
    .S(net164),
    .X(_0199_));
 sg13g2_mux2_1 _7405_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6] ),
    .S(net164),
    .X(_0200_));
 sg13g2_buf_1 _7406_ (.A(_3063_),
    .X(_3095_));
 sg13g2_mux2_1 _7407_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7] ),
    .S(net163),
    .X(_0201_));
 sg13g2_mux2_1 _7408_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4] ),
    .S(net163),
    .X(_0202_));
 sg13g2_mux2_1 _7409_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5] ),
    .S(net163),
    .X(_0203_));
 sg13g2_mux2_1 _7410_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6] ),
    .S(_3095_),
    .X(_0204_));
 sg13g2_mux2_1 _7411_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7] ),
    .S(_3095_),
    .X(_0205_));
 sg13g2_inv_1 _7412_ (.Y(_3096_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0] ));
 sg13g2_nand2_1 _7413_ (.Y(_3097_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7414_ (.B1(_3097_),
    .Y(_0206_),
    .A1(_3096_),
    .A2(net166));
 sg13g2_nand2_1 _7415_ (.Y(_3098_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5] ),
    .B(net217));
 sg13g2_o21ai_1 _7416_ (.B1(_3098_),
    .Y(_0207_),
    .A1(_2182_),
    .A2(net166));
 sg13g2_mux2_1 _7417_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6] ),
    .S(net163),
    .X(_0208_));
 sg13g2_mux2_1 _7418_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7] ),
    .S(net163),
    .X(_0209_));
 sg13g2_inv_1 _7419_ (.Y(_3099_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0] ));
 sg13g2_nand2_1 _7420_ (.Y(_3100_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7421_ (.B1(_3100_),
    .Y(_0210_),
    .A1(_3099_),
    .A2(net166));
 sg13g2_mux2_1 _7422_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5] ),
    .S(net163),
    .X(_0211_));
 sg13g2_mux2_1 _7423_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6] ),
    .S(net163),
    .X(_0212_));
 sg13g2_mux2_1 _7424_ (.A0(_2487_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7] ),
    .S(net163),
    .X(_0213_));
 sg13g2_inv_1 _7425_ (.Y(_3101_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0] ));
 sg13g2_nand2_1 _7426_ (.Y(_3102_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7427_ (.B1(_3102_),
    .Y(_0214_),
    .A1(_3101_),
    .A2(net166));
 sg13g2_buf_1 _7428_ (.A(_1483_),
    .X(_3103_));
 sg13g2_buf_1 _7429_ (.A(net236),
    .X(_3104_));
 sg13g2_buf_1 _7430_ (.A(net216),
    .X(_3105_));
 sg13g2_mux2_1 _7431_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1] ),
    .S(net162),
    .X(_0215_));
 sg13g2_buf_1 _7432_ (.A(_3063_),
    .X(_3106_));
 sg13g2_mux2_1 _7433_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6] ),
    .S(_3106_),
    .X(_0216_));
 sg13g2_mux2_1 _7434_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3] ),
    .S(net162),
    .X(_0217_));
 sg13g2_inv_1 _7435_ (.Y(_3107_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0] ));
 sg13g2_nand2_1 _7436_ (.Y(_3108_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7437_ (.B1(_3108_),
    .Y(_0218_),
    .A1(_3107_),
    .A2(net171));
 sg13g2_mux2_1 _7438_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5] ),
    .S(net161),
    .X(_0219_));
 sg13g2_mux2_1 _7439_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6] ),
    .S(net161),
    .X(_0220_));
 sg13g2_mux2_1 _7440_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7] ),
    .S(_3106_),
    .X(_0221_));
 sg13g2_nand2_1 _7441_ (.Y(_3109_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7442_ (.B1(_3109_),
    .Y(_0222_),
    .A1(_1903_),
    .A2(net171));
 sg13g2_mux2_1 _7443_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5] ),
    .S(net161),
    .X(_0223_));
 sg13g2_mux2_1 _7444_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6] ),
    .S(net161),
    .X(_0224_));
 sg13g2_mux2_1 _7445_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7] ),
    .S(net161),
    .X(_0225_));
 sg13g2_inv_1 _7446_ (.Y(_3110_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0] ));
 sg13g2_nand2_1 _7447_ (.Y(_3111_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4] ),
    .B(net217));
 sg13g2_o21ai_1 _7448_ (.B1(_3111_),
    .Y(_0226_),
    .A1(_3110_),
    .A2(net171));
 sg13g2_mux2_1 _7449_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5] ),
    .S(net161),
    .X(_0227_));
 sg13g2_mux2_1 _7450_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6] ),
    .S(net161),
    .X(_0228_));
 sg13g2_mux2_1 _7451_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7] ),
    .S(net161),
    .X(_0229_));
 sg13g2_inv_1 _7452_ (.Y(_3112_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0] ));
 sg13g2_buf_1 _7453_ (.A(net237),
    .X(_3113_));
 sg13g2_nand2_1 _7454_ (.Y(_3114_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4] ),
    .B(net215));
 sg13g2_o21ai_1 _7455_ (.B1(_3114_),
    .Y(_0230_),
    .A1(_3112_),
    .A2(net171));
 sg13g2_buf_1 _7456_ (.A(_3062_),
    .X(_3115_));
 sg13g2_buf_1 _7457_ (.A(_3115_),
    .X(_3116_));
 sg13g2_mux2_1 _7458_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5] ),
    .S(net160),
    .X(_0231_));
 sg13g2_mux2_1 _7459_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6] ),
    .S(net160),
    .X(_0232_));
 sg13g2_mux2_1 _7460_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7] ),
    .S(net160),
    .X(_0233_));
 sg13g2_inv_1 _7461_ (.Y(_3117_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0] ));
 sg13g2_nand2_1 _7462_ (.Y(_3118_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4] ),
    .B(net215));
 sg13g2_o21ai_1 _7463_ (.B1(_3118_),
    .Y(_0234_),
    .A1(_3117_),
    .A2(net171));
 sg13g2_mux2_1 _7464_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5] ),
    .S(net160),
    .X(_0235_));
 sg13g2_mux2_1 _7465_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6] ),
    .S(net160),
    .X(_0236_));
 sg13g2_mux2_1 _7466_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7] ),
    .S(_3116_),
    .X(_0237_));
 sg13g2_inv_1 _7467_ (.Y(_3119_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0] ));
 sg13g2_nand2_1 _7468_ (.Y(_3120_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4] ),
    .B(net215));
 sg13g2_o21ai_1 _7469_ (.B1(_3120_),
    .Y(_0238_),
    .A1(_3119_),
    .A2(_3058_));
 sg13g2_mux2_1 _7470_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5] ),
    .S(net160),
    .X(_0239_));
 sg13g2_mux2_1 _7471_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6] ),
    .S(net160),
    .X(_0240_));
 sg13g2_mux2_1 _7472_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7] ),
    .S(_3116_),
    .X(_0241_));
 sg13g2_inv_1 _7473_ (.Y(_3121_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0] ));
 sg13g2_nand2_1 _7474_ (.Y(_3122_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4] ),
    .B(net215));
 sg13g2_o21ai_1 _7475_ (.B1(_3122_),
    .Y(_0242_),
    .A1(_3121_),
    .A2(_3058_));
 sg13g2_mux2_1 _7476_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5] ),
    .S(net160),
    .X(_0243_));
 sg13g2_buf_1 _7477_ (.A(_3115_),
    .X(_3123_));
 sg13g2_mux2_1 _7478_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6] ),
    .S(_3123_),
    .X(_0244_));
 sg13g2_mux2_1 _7479_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7] ),
    .S(_3123_),
    .X(_0245_));
 sg13g2_mux2_1 _7480_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10] ),
    .S(net162),
    .X(_0246_));
 sg13g2_mux2_1 _7481_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11] ),
    .S(net162),
    .X(_0247_));
 sg13g2_mux2_1 _7482_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12] ),
    .S(net162),
    .X(_0248_));
 sg13g2_mux2_1 _7483_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13] ),
    .S(net162),
    .X(_0249_));
 sg13g2_mux2_1 _7484_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18] ),
    .S(net159),
    .X(_0250_));
 sg13g2_mux2_1 _7485_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19] ),
    .S(net159),
    .X(_0251_));
 sg13g2_mux2_1 _7486_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20] ),
    .S(net159),
    .X(_0252_));
 sg13g2_mux2_1 _7487_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21] ),
    .S(net159),
    .X(_0253_));
 sg13g2_mux2_1 _7488_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22] ),
    .S(net159),
    .X(_0254_));
 sg13g2_mux2_1 _7489_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23] ),
    .S(net159),
    .X(_0255_));
 sg13g2_mux2_1 _7490_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24] ),
    .S(net159),
    .X(_0256_));
 sg13g2_mux2_1 _7491_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25] ),
    .S(net159),
    .X(_0257_));
 sg13g2_buf_1 _7492_ (.A(_3115_),
    .X(_3124_));
 sg13g2_mux2_1 _7493_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26] ),
    .S(net158),
    .X(_0258_));
 sg13g2_mux2_1 _7494_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27] ),
    .S(net158),
    .X(_0259_));
 sg13g2_mux2_1 _7495_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28] ),
    .S(net158),
    .X(_0260_));
 sg13g2_mux2_1 _7496_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29] ),
    .S(net158),
    .X(_0261_));
 sg13g2_mux2_1 _7497_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30] ),
    .S(net158),
    .X(_0262_));
 sg13g2_mux2_1 _7498_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31] ),
    .S(net158),
    .X(_0263_));
 sg13g2_nor2_1 _7499_ (.A(_0047_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .Y(_3125_));
 sg13g2_buf_2 _7500_ (.A(_3125_),
    .X(_3126_));
 sg13g2_buf_1 _7501_ (.A(_3126_),
    .X(_3127_));
 sg13g2_nand3_1 _7502_ (.B(_1991_),
    .C(_2106_),
    .A(_2132_),
    .Y(_3128_));
 sg13g2_nand2b_1 _7503_ (.Y(_3129_),
    .B(_3128_),
    .A_N(_0049_));
 sg13g2_buf_2 _7504_ (.A(_3129_),
    .X(_3130_));
 sg13g2_nor3_1 _7505_ (.A(_1387_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .C(_3130_),
    .Y(_3131_));
 sg13g2_buf_2 _7506_ (.A(_3131_),
    .X(_3132_));
 sg13g2_buf_1 _7507_ (.A(_1483_),
    .X(_3133_));
 sg13g2_a21oi_1 _7508_ (.A1(net274),
    .A2(_3132_),
    .Y(_3134_),
    .B1(net235));
 sg13g2_nor2b_1 _7509_ (.A(net56),
    .B_N(net71),
    .Y(_3135_));
 sg13g2_a21oi_1 _7510_ (.A1(_2534_),
    .A2(_2536_),
    .Y(_3136_),
    .B1(_2537_));
 sg13g2_o21ai_1 _7511_ (.B1(net96),
    .Y(_3137_),
    .A1(_3136_),
    .A2(net71));
 sg13g2_inv_1 _7512_ (.Y(_3138_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_msb ));
 sg13g2_nor4_1 _7513_ (.A(_1451_),
    .B(_1453_),
    .C(_1457_),
    .D(_1518_),
    .Y(_3139_));
 sg13g2_a21oi_1 _7514_ (.A1(_1682_),
    .A2(_2105_),
    .Y(_3140_),
    .B1(_3139_));
 sg13g2_nor2_1 _7515_ (.A(_3138_),
    .B(_3140_),
    .Y(_3141_));
 sg13g2_and2_1 _7516_ (.A(_2599_),
    .B(_3141_),
    .X(_3142_));
 sg13g2_nor2_1 _7517_ (.A(net71),
    .B(_3141_),
    .Y(_3143_));
 sg13g2_nor3_1 _7518_ (.A(net243),
    .B(_3142_),
    .C(_3143_),
    .Y(_3144_));
 sg13g2_nor4_1 _7519_ (.A(_2463_),
    .B(_3135_),
    .C(_3137_),
    .D(_3144_),
    .Y(_3145_));
 sg13g2_nand2_1 _7520_ (.Y(_3146_),
    .A(_2294_),
    .B(_3136_));
 sg13g2_inv_1 _7521_ (.Y(_3147_),
    .A(_3146_));
 sg13g2_or2_1 _7522_ (.X(_3148_),
    .B(_3140_),
    .A(_3138_));
 sg13g2_buf_1 _7523_ (.A(_3148_),
    .X(_3149_));
 sg13g2_or4_1 _7524_ (.A(_1994_),
    .B(net71),
    .C(_3147_),
    .D(_3149_),
    .X(_3150_));
 sg13g2_nor2_1 _7525_ (.A(_2109_),
    .B(_2599_),
    .Y(_3151_));
 sg13g2_or4_1 _7526_ (.A(net173),
    .B(_2546_),
    .C(_3151_),
    .D(_3149_),
    .X(_3152_));
 sg13g2_nor2_1 _7527_ (.A(_2109_),
    .B(_3141_),
    .Y(_3153_));
 sg13g2_nand3_1 _7528_ (.B(net71),
    .C(_3153_),
    .A(_2001_),
    .Y(_3154_));
 sg13g2_nand3b_1 _7529_ (.B(_3153_),
    .C(net97),
    .Y(_3155_),
    .A_N(net71));
 sg13g2_mux2_1 _7530_ (.A0(_3154_),
    .A1(_3155_),
    .S(net56),
    .X(_3156_));
 sg13g2_nand4_1 _7531_ (.B(_3150_),
    .C(_3152_),
    .A(net243),
    .Y(_3157_),
    .D(_3156_));
 sg13g2_xnor2_1 _7532_ (.Y(_3158_),
    .A(_2633_),
    .B(net71));
 sg13g2_a221oi_1 _7533_ (.B2(net56),
    .C1(_1986_),
    .B1(_3142_),
    .A1(_2603_),
    .Y(_3159_),
    .A2(_3149_));
 sg13g2_o21ai_1 _7534_ (.B1(_3159_),
    .Y(_3160_),
    .A1(_2453_),
    .A2(_3158_));
 sg13g2_o21ai_1 _7535_ (.B1(_3160_),
    .Y(_3161_),
    .A1(_3145_),
    .A2(_3157_));
 sg13g2_nand2_1 _7536_ (.Y(_3162_),
    .A(_2389_),
    .B(net80));
 sg13g2_nand4_1 _7537_ (.B(_2453_),
    .C(_2605_),
    .A(net241),
    .Y(_3163_),
    .D(_3162_));
 sg13g2_nor2_1 _7538_ (.A(_2095_),
    .B(_2450_),
    .Y(_3164_));
 sg13g2_or2_1 _7539_ (.X(_3165_),
    .B(net80),
    .A(_1993_));
 sg13g2_nand3_1 _7540_ (.B(_2387_),
    .C(_3165_),
    .A(net86),
    .Y(_3166_));
 sg13g2_a21oi_1 _7541_ (.A1(_2337_),
    .A2(_2344_),
    .Y(_3167_),
    .B1(_3166_));
 sg13g2_a221oi_1 _7542_ (.B2(_2391_),
    .C1(_3167_),
    .B1(_3165_),
    .A1(_2451_),
    .Y(_3168_),
    .A2(_3164_));
 sg13g2_nand3_1 _7543_ (.B(_2389_),
    .C(net80),
    .A(net243),
    .Y(_3169_));
 sg13g2_a21o_1 _7544_ (.A2(_3169_),
    .A1(_3168_),
    .B1(_2605_),
    .X(_3170_));
 sg13g2_nand2_1 _7545_ (.Y(_3171_),
    .A(_3163_),
    .B(_3170_));
 sg13g2_nor2b_1 _7546_ (.A(_2114_),
    .B_N(_2099_),
    .Y(_3172_));
 sg13g2_nor2b_1 _7547_ (.A(net50),
    .B_N(net51),
    .Y(_3173_));
 sg13g2_nand2b_1 _7548_ (.Y(_3174_),
    .B(net50),
    .A_N(net51));
 sg13g2_o21ai_1 _7549_ (.B1(_3174_),
    .Y(_3175_),
    .A1(_3172_),
    .A2(_3173_));
 sg13g2_inv_1 _7550_ (.Y(_3176_),
    .A(_0043_));
 sg13g2_nand3_1 _7551_ (.B(_2690_),
    .C(_1866_),
    .A(net324),
    .Y(_3177_));
 sg13g2_o21ai_1 _7552_ (.B1(_3177_),
    .Y(_3178_),
    .A1(_2690_),
    .A2(_3176_));
 sg13g2_a21oi_1 _7553_ (.A1(_3171_),
    .A2(_3175_),
    .Y(_3179_),
    .B1(_3178_));
 sg13g2_a22oi_1 _7554_ (.Y(_3180_),
    .B1(_2308_),
    .B2(_1981_),
    .A2(net86),
    .A1(_2297_));
 sg13g2_o21ai_1 _7555_ (.B1(_3180_),
    .Y(_3181_),
    .A1(_2100_),
    .A2(_2296_));
 sg13g2_nor2_1 _7556_ (.A(_2095_),
    .B(_2281_),
    .Y(_3182_));
 sg13g2_and3_1 _7557_ (.X(_3183_),
    .A(net243),
    .B(net96),
    .C(_2281_));
 sg13g2_mux2_1 _7558_ (.A0(_3182_),
    .A1(_3183_),
    .S(_2235_),
    .X(_3184_));
 sg13g2_a221oi_1 _7559_ (.B2(_2295_),
    .C1(_2100_),
    .B1(_2235_),
    .A1(_2093_),
    .Y(_3185_),
    .A2(net96));
 sg13g2_and2_1 _7560_ (.A(_2095_),
    .B(_2281_),
    .X(_3186_));
 sg13g2_o21ai_1 _7561_ (.B1(_3186_),
    .Y(_3187_),
    .A1(_2216_),
    .A2(_2223_));
 sg13g2_or4_1 _7562_ (.A(net243),
    .B(_2281_),
    .C(_2216_),
    .D(_2223_),
    .X(_3188_));
 sg13g2_nor2b_1 _7563_ (.A(_2281_),
    .B_N(_2093_),
    .Y(_3189_));
 sg13g2_o21ai_1 _7564_ (.B1(net86),
    .Y(_3190_),
    .A1(net97),
    .A2(_3189_));
 sg13g2_nand3_1 _7565_ (.B(_3188_),
    .C(_3190_),
    .A(_3187_),
    .Y(_3191_));
 sg13g2_a22oi_1 _7566_ (.Y(_3192_),
    .B1(_3185_),
    .B2(_3191_),
    .A2(_3184_),
    .A1(_3181_));
 sg13g2_nor2_1 _7567_ (.A(_1982_),
    .B(_2308_),
    .Y(_3193_));
 sg13g2_nand3_1 _7568_ (.B(_3187_),
    .C(_3188_),
    .A(net97),
    .Y(_3194_));
 sg13g2_nand3_1 _7569_ (.B(_3191_),
    .C(_3194_),
    .A(_3193_),
    .Y(_3195_));
 sg13g2_a21oi_1 _7570_ (.A1(net324),
    .A2(_1866_),
    .Y(_3196_),
    .B1(net277));
 sg13g2_nand3_1 _7571_ (.B(_3195_),
    .C(_3196_),
    .A(_3192_),
    .Y(_3197_));
 sg13g2_and3_1 _7572_ (.X(_3198_),
    .A(_3171_),
    .B(_3175_),
    .C(_3197_));
 sg13g2_and2_1 _7573_ (.A(_3192_),
    .B(_3195_),
    .X(_3199_));
 sg13g2_nor2_1 _7574_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb ),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ),
    .Y(_3200_));
 sg13g2_and3_1 _7575_ (.X(_3201_),
    .A(net324),
    .B(_2690_),
    .C(_1866_));
 sg13g2_o21ai_1 _7576_ (.B1(_3201_),
    .Y(_3202_),
    .A1(_3199_),
    .A2(_3200_));
 sg13g2_nor3_1 _7577_ (.A(_3161_),
    .B(_3201_),
    .C(_3196_),
    .Y(_3203_));
 sg13g2_a221oi_1 _7578_ (.B2(_3202_),
    .C1(_3203_),
    .B1(_3198_),
    .A1(_3161_),
    .Y(_3204_),
    .A2(_3179_));
 sg13g2_buf_1 _7579_ (.A(_3204_),
    .X(_3205_));
 sg13g2_or2_1 _7580_ (.X(_3206_),
    .B(_3157_),
    .A(_3145_));
 sg13g2_a221oi_1 _7581_ (.B2(_3175_),
    .C1(_3178_),
    .B1(_3171_),
    .A1(_3160_),
    .Y(_3207_),
    .A2(_3206_));
 sg13g2_buf_1 _7582_ (.A(_3207_),
    .X(_3208_));
 sg13g2_nand2b_1 _7583_ (.Y(_3209_),
    .B(_2690_),
    .A_N(_0040_));
 sg13g2_a221oi_1 _7584_ (.B2(_3195_),
    .C1(_3209_),
    .B1(_3192_),
    .A1(_3163_),
    .Y(_3210_),
    .A2(_3170_));
 sg13g2_o21ai_1 _7585_ (.B1(_3177_),
    .Y(_3211_),
    .A1(_0043_),
    .A2(_3210_));
 sg13g2_nor2_2 _7586_ (.A(_3208_),
    .B(_3211_),
    .Y(_3212_));
 sg13g2_nor4_1 _7587_ (.A(_1680_),
    .B(_1682_),
    .C(_1510_),
    .D(_0026_),
    .Y(_3213_));
 sg13g2_a21o_1 _7588_ (.A2(_1866_),
    .A1(_2657_),
    .B1(_3213_),
    .X(_3214_));
 sg13g2_nand2_1 _7589_ (.Y(_3215_),
    .A(net324),
    .B(_3214_));
 sg13g2_nor3_1 _7590_ (.A(_3205_),
    .B(_3212_),
    .C(_3215_),
    .Y(_3216_));
 sg13g2_o21ai_1 _7591_ (.B1(_3215_),
    .Y(_3217_),
    .A1(_3205_),
    .A2(_3212_));
 sg13g2_a21oi_1 _7592_ (.A1(_1444_),
    .A2(_1453_),
    .Y(_3218_),
    .B1(_1758_));
 sg13g2_nor2b_1 _7593_ (.A(_2104_),
    .B_N(_3218_),
    .Y(_3219_));
 sg13g2_and2_1 _7594_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb ),
    .B(_3219_),
    .X(_3220_));
 sg13g2_nand3b_1 _7595_ (.B(_3217_),
    .C(_3220_),
    .Y(_3221_),
    .A_N(_3216_));
 sg13g2_buf_2 _7596_ (.A(_3221_),
    .X(_3222_));
 sg13g2_buf_8 _7597_ (.A(_3222_),
    .X(_3223_));
 sg13g2_buf_1 _7598_ (.A(net236),
    .X(_3224_));
 sg13g2_nand2_2 _7599_ (.Y(_3225_),
    .A(_3126_),
    .B(_3132_));
 sg13g2_nand2b_1 _7600_ (.Y(_3226_),
    .B(_3218_),
    .A_N(_2104_));
 sg13g2_and2_1 _7601_ (.A(_2153_),
    .B(_3226_),
    .X(_3227_));
 sg13g2_buf_1 _7602_ (.A(_3227_),
    .X(_3228_));
 sg13g2_buf_1 _7603_ (.A(_3228_),
    .X(_3229_));
 sg13g2_nor3_1 _7604_ (.A(net214),
    .B(_3225_),
    .C(net49),
    .Y(_3230_));
 sg13g2_nor2_1 _7605_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28] ),
    .B(net215),
    .Y(_3231_));
 sg13g2_a221oi_1 _7606_ (.B2(_3230_),
    .C1(_3231_),
    .B1(net40),
    .A1(_3052_),
    .Y(_0264_),
    .A2(_3134_));
 sg13g2_nor2_1 _7607_ (.A(_2318_),
    .B(_3219_),
    .Y(_3232_));
 sg13g2_buf_1 _7608_ (.A(_3232_),
    .X(_3233_));
 sg13g2_buf_1 _7609_ (.A(_3233_),
    .X(_3234_));
 sg13g2_mux2_1 _7610_ (.A0(net46),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ),
    .S(_3225_),
    .X(_3235_));
 sg13g2_mux2_1 _7611_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29] ),
    .A1(_3235_),
    .S(net158),
    .X(_0265_));
 sg13g2_nand2_1 _7612_ (.Y(_3236_),
    .A(_2468_),
    .B(_3226_));
 sg13g2_buf_1 _7613_ (.A(_3236_),
    .X(_3237_));
 sg13g2_buf_1 _7614_ (.A(_3237_),
    .X(_3238_));
 sg13g2_nand2_1 _7615_ (.Y(_3239_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ),
    .B(_3225_));
 sg13g2_o21ai_1 _7616_ (.B1(_3239_),
    .Y(_3240_),
    .A1(_3225_),
    .A2(net43));
 sg13g2_mux2_1 _7617_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30] ),
    .A1(_3240_),
    .S(net158),
    .X(_0266_));
 sg13g2_nor2_1 _7618_ (.A(_1483_),
    .B(_3219_),
    .Y(_3241_));
 sg13g2_o21ai_1 _7619_ (.B1(_3241_),
    .Y(_3242_),
    .A1(_2629_),
    .A2(_2637_));
 sg13g2_buf_2 _7620_ (.A(_3242_),
    .X(_3243_));
 sg13g2_buf_8 _7621_ (.A(_3243_),
    .X(_3244_));
 sg13g2_buf_1 _7622_ (.A(net235),
    .X(_3245_));
 sg13g2_a22oi_1 _7623_ (.Y(_3246_),
    .B1(_3134_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ),
    .A2(net213),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7624_ (.B1(_3246_),
    .Y(_0267_),
    .A1(_3225_),
    .A2(net39));
 sg13g2_mux2_1 _7625_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8] ),
    .S(_3124_),
    .X(_0268_));
 sg13g2_mux2_1 _7626_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9] ),
    .S(_3124_),
    .X(_0269_));
 sg13g2_buf_1 _7627_ (.A(_3115_),
    .X(_3247_));
 sg13g2_mux2_1 _7628_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10] ),
    .S(net157),
    .X(_0270_));
 sg13g2_mux2_1 _7629_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11] ),
    .S(net157),
    .X(_0271_));
 sg13g2_mux2_1 _7630_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8] ),
    .S(net162),
    .X(_0272_));
 sg13g2_mux2_1 _7631_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9] ),
    .S(net162),
    .X(_0273_));
 sg13g2_buf_1 _7632_ (.A(net236),
    .X(_3248_));
 sg13g2_buf_1 _7633_ (.A(net212),
    .X(_3249_));
 sg13g2_mux2_1 _7634_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10] ),
    .S(net156),
    .X(_0274_));
 sg13g2_mux2_1 _7635_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11] ),
    .S(net156),
    .X(_0275_));
 sg13g2_mux2_1 _7636_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12] ),
    .S(net156),
    .X(_0276_));
 sg13g2_mux2_1 _7637_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13] ),
    .S(net156),
    .X(_0277_));
 sg13g2_mux2_1 _7638_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18] ),
    .S(net157),
    .X(_0278_));
 sg13g2_mux2_1 _7639_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19] ),
    .S(net157),
    .X(_0279_));
 sg13g2_mux2_1 _7640_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20] ),
    .S(net157),
    .X(_0280_));
 sg13g2_mux2_1 _7641_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21] ),
    .S(net157),
    .X(_0281_));
 sg13g2_mux2_1 _7642_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22] ),
    .S(net157),
    .X(_0282_));
 sg13g2_mux2_1 _7643_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23] ),
    .S(net157),
    .X(_0283_));
 sg13g2_mux2_1 _7644_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24] ),
    .S(_3247_),
    .X(_0284_));
 sg13g2_mux2_1 _7645_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25] ),
    .S(_3247_),
    .X(_0285_));
 sg13g2_buf_1 _7646_ (.A(_3115_),
    .X(_3250_));
 sg13g2_mux2_1 _7647_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26] ),
    .S(net155),
    .X(_0286_));
 sg13g2_mux2_1 _7648_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27] ),
    .S(net155),
    .X(_0287_));
 sg13g2_inv_1 _7649_ (.Y(_3251_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[28] ));
 sg13g2_buf_1 _7650_ (.A(net236),
    .X(_3252_));
 sg13g2_buf_1 _7651_ (.A(net211),
    .X(_3253_));
 sg13g2_buf_1 _7652_ (.A(_1483_),
    .X(_3254_));
 sg13g2_buf_1 _7653_ (.A(_3254_),
    .X(_3255_));
 sg13g2_nand2_1 _7654_ (.Y(_3256_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24] ),
    .B(net210));
 sg13g2_o21ai_1 _7655_ (.B1(_3256_),
    .Y(_0288_),
    .A1(_3251_),
    .A2(net154));
 sg13g2_mux2_1 _7656_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29] ),
    .S(net155),
    .X(_0289_));
 sg13g2_mux2_1 _7657_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30] ),
    .S(net155),
    .X(_0290_));
 sg13g2_mux2_1 _7658_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31] ),
    .S(net155),
    .X(_0291_));
 sg13g2_buf_1 _7659_ (.A(net216),
    .X(_3257_));
 sg13g2_buf_1 _7660_ (.A(_3228_),
    .X(_3258_));
 sg13g2_nand2b_1 _7661_ (.Y(_3259_),
    .B(_1387_),
    .A_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ));
 sg13g2_buf_1 _7662_ (.A(_3259_),
    .X(_3260_));
 sg13g2_nor2_1 _7663_ (.A(_3130_),
    .B(_3260_),
    .Y(_3261_));
 sg13g2_buf_2 _7664_ (.A(_3261_),
    .X(_3262_));
 sg13g2_nand2_1 _7665_ (.Y(_3263_),
    .A(net274),
    .B(_3262_));
 sg13g2_nor3_1 _7666_ (.A(net214),
    .B(net48),
    .C(_3263_),
    .Y(_3264_));
 sg13g2_buf_1 _7667_ (.A(net236),
    .X(_3265_));
 sg13g2_or2_1 _7668_ (.X(_3266_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .A(_0047_));
 sg13g2_nor3_2 _7669_ (.A(_3266_),
    .B(_3130_),
    .C(_3260_),
    .Y(_3267_));
 sg13g2_nor3_1 _7670_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ),
    .B(net209),
    .C(_3267_),
    .Y(_3268_));
 sg13g2_a221oi_1 _7671_ (.B2(_3264_),
    .C1(_3268_),
    .B1(net40),
    .A1(_3251_),
    .Y(_0292_),
    .A2(net153));
 sg13g2_nor2b_1 _7672_ (.A(_3267_),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ),
    .Y(_3269_));
 sg13g2_a21oi_1 _7673_ (.A1(net46),
    .A2(_3267_),
    .Y(_3270_),
    .B1(_3269_));
 sg13g2_nand2_1 _7674_ (.Y(_3271_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29] ),
    .B(net210));
 sg13g2_o21ai_1 _7675_ (.B1(_3271_),
    .Y(_0293_),
    .A1(net154),
    .A2(_3270_));
 sg13g2_nand2_1 _7676_ (.Y(_3272_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ),
    .B(_3263_));
 sg13g2_o21ai_1 _7677_ (.B1(_3272_),
    .Y(_3273_),
    .A1(net43),
    .A2(_3263_));
 sg13g2_mux2_1 _7678_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30] ),
    .A1(_3273_),
    .S(net155),
    .X(_0294_));
 sg13g2_nor2_1 _7679_ (.A(net216),
    .B(_3267_),
    .Y(_3274_));
 sg13g2_a22oi_1 _7680_ (.Y(_3275_),
    .B1(_3274_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ),
    .A2(net213),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7681_ (.B1(_3275_),
    .Y(_0295_),
    .A1(net39),
    .A2(_3263_));
 sg13g2_mux2_1 _7682_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8] ),
    .S(net155),
    .X(_0296_));
 sg13g2_mux2_1 _7683_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9] ),
    .S(_3250_),
    .X(_0297_));
 sg13g2_mux2_1 _7684_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10] ),
    .S(_3250_),
    .X(_0298_));
 sg13g2_mux2_1 _7685_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11] ),
    .S(net155),
    .X(_0299_));
 sg13g2_mux2_1 _7686_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8] ),
    .S(_3249_),
    .X(_0300_));
 sg13g2_mux2_1 _7687_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9] ),
    .S(_3249_),
    .X(_0301_));
 sg13g2_mux2_1 _7688_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10] ),
    .S(net156),
    .X(_0302_));
 sg13g2_mux2_1 _7689_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11] ),
    .S(net156),
    .X(_0303_));
 sg13g2_mux2_1 _7690_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12] ),
    .S(net156),
    .X(_0304_));
 sg13g2_mux2_1 _7691_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13] ),
    .S(net156),
    .X(_0305_));
 sg13g2_buf_1 _7692_ (.A(_3115_),
    .X(_3276_));
 sg13g2_mux2_1 _7693_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18] ),
    .S(net152),
    .X(_0306_));
 sg13g2_mux2_1 _7694_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19] ),
    .S(_3276_),
    .X(_0307_));
 sg13g2_mux2_1 _7695_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20] ),
    .S(net152),
    .X(_0308_));
 sg13g2_mux2_1 _7696_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21] ),
    .S(net152),
    .X(_0309_));
 sg13g2_mux2_1 _7697_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22] ),
    .S(net152),
    .X(_0310_));
 sg13g2_mux2_1 _7698_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23] ),
    .S(_3276_),
    .X(_0311_));
 sg13g2_mux2_1 _7699_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24] ),
    .S(net152),
    .X(_0312_));
 sg13g2_mux2_1 _7700_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25] ),
    .S(net152),
    .X(_0313_));
 sg13g2_mux2_1 _7701_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26] ),
    .S(net152),
    .X(_0314_));
 sg13g2_mux2_1 _7702_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27] ),
    .S(net152),
    .X(_0315_));
 sg13g2_buf_1 _7703_ (.A(_3115_),
    .X(_3277_));
 sg13g2_mux2_1 _7704_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28] ),
    .S(net151),
    .X(_0316_));
 sg13g2_mux2_1 _7705_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29] ),
    .S(net151),
    .X(_0317_));
 sg13g2_mux2_1 _7706_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30] ),
    .S(net151),
    .X(_0318_));
 sg13g2_mux2_1 _7707_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31] ),
    .S(net151),
    .X(_0319_));
 sg13g2_buf_8 _7708_ (.A(_3222_),
    .X(_3278_));
 sg13g2_buf_1 _7709_ (.A(net236),
    .X(_3279_));
 sg13g2_nand2b_1 _7710_ (.Y(_3280_),
    .B(_3128_),
    .A_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ));
 sg13g2_buf_1 _7711_ (.A(_3280_),
    .X(_3281_));
 sg13g2_nor3_1 _7712_ (.A(_1387_),
    .B(_0048_),
    .C(_3281_),
    .Y(_3282_));
 sg13g2_buf_2 _7713_ (.A(_3282_),
    .X(_3283_));
 sg13g2_nand2_2 _7714_ (.Y(_3284_),
    .A(net274),
    .B(_3283_));
 sg13g2_nor3_1 _7715_ (.A(net208),
    .B(net48),
    .C(_3284_),
    .Y(_3285_));
 sg13g2_buf_1 _7716_ (.A(_1483_),
    .X(_3286_));
 sg13g2_a21oi_1 _7717_ (.A1(net274),
    .A2(_3283_),
    .Y(_3287_),
    .B1(net234));
 sg13g2_nor2_1 _7718_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28] ),
    .B(net215),
    .Y(_3288_));
 sg13g2_a221oi_1 _7719_ (.B2(_3060_),
    .C1(_3288_),
    .B1(_3287_),
    .A1(net38),
    .Y(_0320_),
    .A2(_3285_));
 sg13g2_mux2_1 _7720_ (.A0(net46),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ),
    .S(_3284_),
    .X(_3289_));
 sg13g2_mux2_1 _7721_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29] ),
    .A1(_3289_),
    .S(net151),
    .X(_0321_));
 sg13g2_nand2_1 _7722_ (.Y(_3290_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ),
    .B(_3284_));
 sg13g2_o21ai_1 _7723_ (.B1(_3290_),
    .Y(_3291_),
    .A1(net43),
    .A2(_3284_));
 sg13g2_mux2_1 _7724_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30] ),
    .A1(_3291_),
    .S(net151),
    .X(_0322_));
 sg13g2_a22oi_1 _7725_ (.Y(_3292_),
    .B1(_3287_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ),
    .A2(net213),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7726_ (.B1(_3292_),
    .Y(_0323_),
    .A1(net39),
    .A2(_3284_));
 sg13g2_mux2_1 _7727_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8] ),
    .S(net151),
    .X(_0324_));
 sg13g2_mux2_1 _7728_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9] ),
    .S(_3277_),
    .X(_0325_));
 sg13g2_mux2_1 _7729_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10] ),
    .S(_3277_),
    .X(_0326_));
 sg13g2_mux2_1 _7730_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11] ),
    .S(net151),
    .X(_0327_));
 sg13g2_buf_1 _7731_ (.A(net212),
    .X(_3293_));
 sg13g2_mux2_1 _7732_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8] ),
    .S(net150),
    .X(_0328_));
 sg13g2_mux2_1 _7733_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9] ),
    .S(net150),
    .X(_0329_));
 sg13g2_mux2_1 _7734_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10] ),
    .S(net150),
    .X(_0330_));
 sg13g2_mux2_1 _7735_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11] ),
    .S(net150),
    .X(_0331_));
 sg13g2_mux2_1 _7736_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12] ),
    .S(net150),
    .X(_0332_));
 sg13g2_mux2_1 _7737_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13] ),
    .S(net150),
    .X(_0333_));
 sg13g2_buf_1 _7738_ (.A(_3062_),
    .X(_3294_));
 sg13g2_buf_1 _7739_ (.A(_3294_),
    .X(_3295_));
 sg13g2_mux2_1 _7740_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18] ),
    .S(net149),
    .X(_0334_));
 sg13g2_mux2_1 _7741_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19] ),
    .S(net149),
    .X(_0335_));
 sg13g2_mux2_1 _7742_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20] ),
    .S(net149),
    .X(_0336_));
 sg13g2_mux2_1 _7743_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21] ),
    .S(net149),
    .X(_0337_));
 sg13g2_mux2_1 _7744_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22] ),
    .S(net149),
    .X(_0338_));
 sg13g2_mux2_1 _7745_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23] ),
    .S(_3295_),
    .X(_0339_));
 sg13g2_mux2_1 _7746_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24] ),
    .S(net149),
    .X(_0340_));
 sg13g2_mux2_1 _7747_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25] ),
    .S(net149),
    .X(_0341_));
 sg13g2_mux2_1 _7748_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26] ),
    .S(net149),
    .X(_0342_));
 sg13g2_mux2_1 _7749_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27] ),
    .S(_3295_),
    .X(_0343_));
 sg13g2_inv_1 _7750_ (.Y(_3296_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _7751_ (.Y(_3297_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24] ),
    .B(net210));
 sg13g2_o21ai_1 _7752_ (.B1(_3297_),
    .Y(_0344_),
    .A1(_3296_),
    .A2(net154));
 sg13g2_buf_1 _7753_ (.A(_3294_),
    .X(_3298_));
 sg13g2_mux2_1 _7754_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29] ),
    .S(net148),
    .X(_0345_));
 sg13g2_mux2_1 _7755_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30] ),
    .S(net148),
    .X(_0346_));
 sg13g2_mux2_1 _7756_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31] ),
    .S(net148),
    .X(_0347_));
 sg13g2_nand2b_1 _7757_ (.Y(_3299_),
    .B(_1387_),
    .A_N(_0048_));
 sg13g2_buf_1 _7758_ (.A(_3299_),
    .X(_3300_));
 sg13g2_nor2_1 _7759_ (.A(_3281_),
    .B(_3300_),
    .Y(_3301_));
 sg13g2_buf_2 _7760_ (.A(_3301_),
    .X(_3302_));
 sg13g2_nand2_2 _7761_ (.Y(_3303_),
    .A(_3126_),
    .B(_3302_));
 sg13g2_nor3_1 _7762_ (.A(net214),
    .B(net48),
    .C(_3303_),
    .Y(_3304_));
 sg13g2_or2_1 _7763_ (.X(_3305_),
    .B(_3300_),
    .A(_3281_));
 sg13g2_buf_1 _7764_ (.A(_3305_),
    .X(_3306_));
 sg13g2_nor2_1 _7765_ (.A(_3266_),
    .B(_3306_),
    .Y(_3307_));
 sg13g2_nor3_1 _7766_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ),
    .B(net209),
    .C(_3307_),
    .Y(_3308_));
 sg13g2_a221oi_1 _7767_ (.B2(_3304_),
    .C1(_3308_),
    .B1(net40),
    .A1(_3296_),
    .Y(_0348_),
    .A2(net153));
 sg13g2_and2_1 _7768_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ),
    .B(_3303_),
    .X(_3309_));
 sg13g2_a21oi_1 _7769_ (.A1(net46),
    .A2(_3307_),
    .Y(_3310_),
    .B1(_3309_));
 sg13g2_nand2_1 _7770_ (.Y(_3311_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29] ),
    .B(net210));
 sg13g2_o21ai_1 _7771_ (.B1(_3311_),
    .Y(_0349_),
    .A1(net154),
    .A2(_3310_));
 sg13g2_nand2_1 _7772_ (.Y(_3312_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ),
    .B(_3303_));
 sg13g2_o21ai_1 _7773_ (.B1(_3312_),
    .Y(_3313_),
    .A1(net43),
    .A2(_3303_));
 sg13g2_mux2_1 _7774_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30] ),
    .A1(_3313_),
    .S(net148),
    .X(_0350_));
 sg13g2_nor2_1 _7775_ (.A(net216),
    .B(_3307_),
    .Y(_3314_));
 sg13g2_a22oi_1 _7776_ (.Y(_3315_),
    .B1(_3314_),
    .B2(_2496_),
    .A2(net213),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7777_ (.B1(_3315_),
    .Y(_0351_),
    .A1(net39),
    .A2(_3303_));
 sg13g2_mux2_1 _7778_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8] ),
    .S(net148),
    .X(_0352_));
 sg13g2_mux2_1 _7779_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9] ),
    .S(net148),
    .X(_0353_));
 sg13g2_mux2_1 _7780_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10] ),
    .S(net148),
    .X(_0354_));
 sg13g2_mux2_1 _7781_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11] ),
    .S(_3298_),
    .X(_0355_));
 sg13g2_mux2_1 _7782_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8] ),
    .S(net150),
    .X(_0356_));
 sg13g2_mux2_1 _7783_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9] ),
    .S(net150),
    .X(_0357_));
 sg13g2_mux2_1 _7784_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10] ),
    .S(_3293_),
    .X(_0358_));
 sg13g2_mux2_1 _7785_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11] ),
    .S(_3293_),
    .X(_0359_));
 sg13g2_buf_1 _7786_ (.A(net212),
    .X(_3316_));
 sg13g2_mux2_1 _7787_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12] ),
    .S(net147),
    .X(_0360_));
 sg13g2_mux2_1 _7788_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13] ),
    .S(net147),
    .X(_0361_));
 sg13g2_mux2_1 _7789_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18] ),
    .S(net148),
    .X(_0362_));
 sg13g2_mux2_1 _7790_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19] ),
    .S(_3298_),
    .X(_0363_));
 sg13g2_buf_1 _7791_ (.A(_3294_),
    .X(_3317_));
 sg13g2_mux2_1 _7792_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20] ),
    .S(net146),
    .X(_0364_));
 sg13g2_mux2_1 _7793_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21] ),
    .S(net146),
    .X(_0365_));
 sg13g2_mux2_1 _7794_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22] ),
    .S(net146),
    .X(_0366_));
 sg13g2_mux2_1 _7795_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23] ),
    .S(net146),
    .X(_0367_));
 sg13g2_mux2_1 _7796_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24] ),
    .S(_3317_),
    .X(_0368_));
 sg13g2_mux2_1 _7797_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25] ),
    .S(_3317_),
    .X(_0369_));
 sg13g2_mux2_1 _7798_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26] ),
    .S(net146),
    .X(_0370_));
 sg13g2_mux2_1 _7799_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27] ),
    .S(net146),
    .X(_0371_));
 sg13g2_mux2_1 _7800_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28] ),
    .S(net146),
    .X(_0372_));
 sg13g2_mux2_1 _7801_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29] ),
    .S(net146),
    .X(_0373_));
 sg13g2_buf_1 _7802_ (.A(_3294_),
    .X(_3318_));
 sg13g2_mux2_1 _7803_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30] ),
    .S(net145),
    .X(_0374_));
 sg13g2_mux2_1 _7804_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31] ),
    .S(net145),
    .X(_0375_));
 sg13g2_nor3_1 _7805_ (.A(_1387_),
    .B(_0048_),
    .C(_3130_),
    .Y(_3319_));
 sg13g2_buf_2 _7806_ (.A(_3319_),
    .X(_3320_));
 sg13g2_buf_1 _7807_ (.A(_1483_),
    .X(_3321_));
 sg13g2_a21oi_1 _7808_ (.A1(net274),
    .A2(_3320_),
    .Y(_3322_),
    .B1(net233));
 sg13g2_nand2_2 _7809_ (.Y(_3323_),
    .A(net274),
    .B(_3320_));
 sg13g2_nor3_1 _7810_ (.A(net211),
    .B(net49),
    .C(_3323_),
    .Y(_3324_));
 sg13g2_nor2_1 _7811_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28] ),
    .B(net215),
    .Y(_3325_));
 sg13g2_a221oi_1 _7812_ (.B2(net40),
    .C1(_3325_),
    .B1(_3324_),
    .A1(_3065_),
    .Y(_0376_),
    .A2(_3322_));
 sg13g2_buf_1 _7813_ (.A(_3233_),
    .X(_3326_));
 sg13g2_mux2_1 _7814_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ),
    .S(_3323_),
    .X(_3327_));
 sg13g2_mux2_1 _7815_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29] ),
    .A1(_3327_),
    .S(net145),
    .X(_0377_));
 sg13g2_nand2_1 _7816_ (.Y(_3328_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ),
    .B(_3323_));
 sg13g2_o21ai_1 _7817_ (.B1(_3328_),
    .Y(_3329_),
    .A1(_3238_),
    .A2(_3323_));
 sg13g2_mux2_1 _7818_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30] ),
    .A1(_3329_),
    .S(net145),
    .X(_0378_));
 sg13g2_a22oi_1 _7819_ (.Y(_3330_),
    .B1(_3322_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ),
    .A2(net213),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7820_ (.B1(_3330_),
    .Y(_0379_),
    .A1(net39),
    .A2(_3323_));
 sg13g2_mux2_1 _7821_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8] ),
    .S(_3318_),
    .X(_0380_));
 sg13g2_mux2_1 _7822_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9] ),
    .S(net145),
    .X(_0381_));
 sg13g2_mux2_1 _7823_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10] ),
    .S(net145),
    .X(_0382_));
 sg13g2_mux2_1 _7824_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11] ),
    .S(net145),
    .X(_0383_));
 sg13g2_mux2_1 _7825_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8] ),
    .S(net147),
    .X(_0384_));
 sg13g2_mux2_1 _7826_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9] ),
    .S(net147),
    .X(_0385_));
 sg13g2_mux2_1 _7827_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10] ),
    .S(net147),
    .X(_0386_));
 sg13g2_mux2_1 _7828_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11] ),
    .S(net147),
    .X(_0387_));
 sg13g2_mux2_1 _7829_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12] ),
    .S(net147),
    .X(_0388_));
 sg13g2_mux2_1 _7830_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13] ),
    .S(net147),
    .X(_0389_));
 sg13g2_mux2_1 _7831_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18] ),
    .S(net145),
    .X(_0390_));
 sg13g2_mux2_1 _7832_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19] ),
    .S(_3318_),
    .X(_0391_));
 sg13g2_buf_1 _7833_ (.A(_3294_),
    .X(_3331_));
 sg13g2_mux2_1 _7834_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20] ),
    .S(net144),
    .X(_0392_));
 sg13g2_mux2_1 _7835_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21] ),
    .S(net144),
    .X(_0393_));
 sg13g2_mux2_1 _7836_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22] ),
    .S(net144),
    .X(_0394_));
 sg13g2_mux2_1 _7837_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23] ),
    .S(net144),
    .X(_0395_));
 sg13g2_mux2_1 _7838_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24] ),
    .S(_3331_),
    .X(_0396_));
 sg13g2_mux2_1 _7839_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25] ),
    .S(_3331_),
    .X(_0397_));
 sg13g2_mux2_1 _7840_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26] ),
    .S(net144),
    .X(_0398_));
 sg13g2_mux2_1 _7841_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27] ),
    .S(net144),
    .X(_0399_));
 sg13g2_mux2_1 _7842_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28] ),
    .S(net144),
    .X(_0400_));
 sg13g2_mux2_1 _7843_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29] ),
    .S(net144),
    .X(_0401_));
 sg13g2_buf_1 _7844_ (.A(_3294_),
    .X(_3332_));
 sg13g2_mux2_1 _7845_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30] ),
    .S(net143),
    .X(_0402_));
 sg13g2_mux2_1 _7846_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31] ),
    .S(net143),
    .X(_0403_));
 sg13g2_nor2_1 _7847_ (.A(_3130_),
    .B(_3300_),
    .Y(_3333_));
 sg13g2_buf_2 _7848_ (.A(_3333_),
    .X(_3334_));
 sg13g2_a21oi_1 _7849_ (.A1(net274),
    .A2(_3334_),
    .Y(_3335_),
    .B1(net233));
 sg13g2_nand2_2 _7850_ (.Y(_3336_),
    .A(net274),
    .B(_3334_));
 sg13g2_nor3_1 _7851_ (.A(net211),
    .B(net49),
    .C(_3336_),
    .Y(_3337_));
 sg13g2_nor2_1 _7852_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28] ),
    .B(net215),
    .Y(_3338_));
 sg13g2_a221oi_1 _7853_ (.B2(net40),
    .C1(_3338_),
    .B1(_3337_),
    .A1(_1922_),
    .Y(_0404_),
    .A2(_3335_));
 sg13g2_mux2_1 _7854_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ),
    .S(_3336_),
    .X(_3339_));
 sg13g2_mux2_1 _7855_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29] ),
    .A1(_3339_),
    .S(net143),
    .X(_0405_));
 sg13g2_nand2_1 _7856_ (.Y(_3340_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ),
    .B(_3336_));
 sg13g2_o21ai_1 _7857_ (.B1(_3340_),
    .Y(_3341_),
    .A1(net43),
    .A2(_3336_));
 sg13g2_mux2_1 _7858_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30] ),
    .A1(_3341_),
    .S(net143),
    .X(_0406_));
 sg13g2_a22oi_1 _7859_ (.Y(_3342_),
    .B1(_3335_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ),
    .A2(_3245_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7860_ (.B1(_3342_),
    .Y(_0407_),
    .A1(net39),
    .A2(_3336_));
 sg13g2_mux2_1 _7861_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8] ),
    .S(net143),
    .X(_0408_));
 sg13g2_mux2_1 _7862_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9] ),
    .S(net143),
    .X(_0409_));
 sg13g2_mux2_1 _7863_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10] ),
    .S(net143),
    .X(_0410_));
 sg13g2_mux2_1 _7864_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11] ),
    .S(net143),
    .X(_0411_));
 sg13g2_mux2_1 _7865_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8] ),
    .S(_3316_),
    .X(_0412_));
 sg13g2_mux2_1 _7866_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9] ),
    .S(_3316_),
    .X(_0413_));
 sg13g2_buf_1 _7867_ (.A(net212),
    .X(_3343_));
 sg13g2_mux2_1 _7868_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10] ),
    .S(net142),
    .X(_0414_));
 sg13g2_mux2_1 _7869_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11] ),
    .S(_3343_),
    .X(_0415_));
 sg13g2_mux2_1 _7870_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12] ),
    .S(net142),
    .X(_0416_));
 sg13g2_mux2_1 _7871_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13] ),
    .S(net142),
    .X(_0417_));
 sg13g2_mux2_1 _7872_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18] ),
    .S(_3332_),
    .X(_0418_));
 sg13g2_mux2_1 _7873_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19] ),
    .S(_3332_),
    .X(_0419_));
 sg13g2_buf_1 _7874_ (.A(_3294_),
    .X(_3344_));
 sg13g2_mux2_1 _7875_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20] ),
    .S(net141),
    .X(_0420_));
 sg13g2_mux2_1 _7876_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21] ),
    .S(net141),
    .X(_0421_));
 sg13g2_mux2_1 _7877_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22] ),
    .S(net141),
    .X(_0422_));
 sg13g2_mux2_1 _7878_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23] ),
    .S(_3344_),
    .X(_0423_));
 sg13g2_mux2_1 _7879_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24] ),
    .S(net141),
    .X(_0424_));
 sg13g2_mux2_1 _7880_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25] ),
    .S(net141),
    .X(_0425_));
 sg13g2_mux2_1 _7881_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26] ),
    .S(net141),
    .X(_0426_));
 sg13g2_mux2_1 _7882_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27] ),
    .S(net141),
    .X(_0427_));
 sg13g2_mux2_1 _7883_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28] ),
    .S(net141),
    .X(_0428_));
 sg13g2_mux2_1 _7884_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29] ),
    .S(_3344_),
    .X(_0429_));
 sg13g2_buf_1 _7885_ (.A(_3062_),
    .X(_3345_));
 sg13g2_buf_1 _7886_ (.A(_3345_),
    .X(_3346_));
 sg13g2_mux2_1 _7887_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30] ),
    .S(_3346_),
    .X(_0430_));
 sg13g2_mux2_1 _7888_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31] ),
    .S(net140),
    .X(_0431_));
 sg13g2_buf_8 _7889_ (.A(_3222_),
    .X(_3347_));
 sg13g2_buf_1 _7890_ (.A(_3228_),
    .X(_3348_));
 sg13g2_nor2_1 _7891_ (.A(_0046_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .Y(_3349_));
 sg13g2_buf_1 _7892_ (.A(_3349_),
    .X(_3350_));
 sg13g2_buf_1 _7893_ (.A(_3350_),
    .X(_3351_));
 sg13g2_nor3_1 _7894_ (.A(_1387_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .C(_3281_),
    .Y(_3352_));
 sg13g2_buf_2 _7895_ (.A(_3352_),
    .X(_3353_));
 sg13g2_nand2_2 _7896_ (.Y(_3354_),
    .A(net273),
    .B(_3353_));
 sg13g2_nor3_1 _7897_ (.A(net208),
    .B(net47),
    .C(_3354_),
    .Y(_3355_));
 sg13g2_a21oi_1 _7898_ (.A1(net273),
    .A2(_3353_),
    .Y(_3356_),
    .B1(net234));
 sg13g2_nor2_1 _7899_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28] ),
    .B(_3113_),
    .Y(_3357_));
 sg13g2_a221oi_1 _7900_ (.B2(_2015_),
    .C1(_3357_),
    .B1(_3356_),
    .A1(net37),
    .Y(_0432_),
    .A2(_3355_));
 sg13g2_mux2_1 _7901_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ),
    .S(_3354_),
    .X(_3358_));
 sg13g2_mux2_1 _7902_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29] ),
    .A1(_3358_),
    .S(net140),
    .X(_0433_));
 sg13g2_nand2_1 _7903_ (.Y(_3359_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ),
    .B(_3354_));
 sg13g2_o21ai_1 _7904_ (.B1(_3359_),
    .Y(_3360_),
    .A1(net43),
    .A2(_3354_));
 sg13g2_mux2_1 _7905_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30] ),
    .A1(_3360_),
    .S(net140),
    .X(_0434_));
 sg13g2_a22oi_1 _7906_ (.Y(_3361_),
    .B1(_3356_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ),
    .A2(_3245_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7907_ (.B1(_3361_),
    .Y(_0435_),
    .A1(net39),
    .A2(_3354_));
 sg13g2_mux2_1 _7908_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8] ),
    .S(net140),
    .X(_0436_));
 sg13g2_mux2_1 _7909_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9] ),
    .S(net140),
    .X(_0437_));
 sg13g2_mux2_1 _7910_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10] ),
    .S(net140),
    .X(_0438_));
 sg13g2_mux2_1 _7911_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11] ),
    .S(_3346_),
    .X(_0439_));
 sg13g2_mux2_1 _7912_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8] ),
    .S(net142),
    .X(_0440_));
 sg13g2_mux2_1 _7913_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9] ),
    .S(_3343_),
    .X(_0441_));
 sg13g2_mux2_1 _7914_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10] ),
    .S(net142),
    .X(_0442_));
 sg13g2_mux2_1 _7915_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11] ),
    .S(net142),
    .X(_0443_));
 sg13g2_mux2_1 _7916_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12] ),
    .S(net142),
    .X(_0444_));
 sg13g2_mux2_1 _7917_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13] ),
    .S(net142),
    .X(_0445_));
 sg13g2_mux2_1 _7918_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18] ),
    .S(net140),
    .X(_0446_));
 sg13g2_mux2_1 _7919_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19] ),
    .S(net140),
    .X(_0447_));
 sg13g2_buf_1 _7920_ (.A(_3345_),
    .X(_3362_));
 sg13g2_mux2_1 _7921_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20] ),
    .S(net139),
    .X(_0448_));
 sg13g2_mux2_1 _7922_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21] ),
    .S(net139),
    .X(_0449_));
 sg13g2_mux2_1 _7923_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22] ),
    .S(net139),
    .X(_0450_));
 sg13g2_mux2_1 _7924_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23] ),
    .S(net139),
    .X(_0451_));
 sg13g2_mux2_1 _7925_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24] ),
    .S(net139),
    .X(_0452_));
 sg13g2_mux2_1 _7926_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25] ),
    .S(net139),
    .X(_0453_));
 sg13g2_mux2_1 _7927_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26] ),
    .S(net139),
    .X(_0454_));
 sg13g2_mux2_1 _7928_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27] ),
    .S(net139),
    .X(_0455_));
 sg13g2_inv_1 _7929_ (.Y(_3363_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _7930_ (.Y(_3364_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24] ),
    .B(net210));
 sg13g2_o21ai_1 _7931_ (.B1(_3364_),
    .Y(_0456_),
    .A1(_3363_),
    .A2(net154));
 sg13g2_mux2_1 _7932_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29] ),
    .S(_3362_),
    .X(_0457_));
 sg13g2_mux2_1 _7933_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30] ),
    .S(_3362_),
    .X(_0458_));
 sg13g2_buf_1 _7934_ (.A(_3345_),
    .X(_3365_));
 sg13g2_mux2_1 _7935_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31] ),
    .S(net138),
    .X(_0459_));
 sg13g2_nor2_1 _7936_ (.A(_3260_),
    .B(_3281_),
    .Y(_3366_));
 sg13g2_buf_2 _7937_ (.A(_3366_),
    .X(_3367_));
 sg13g2_nand2_2 _7938_ (.Y(_3368_),
    .A(_3350_),
    .B(_3367_));
 sg13g2_nor3_1 _7939_ (.A(net214),
    .B(net48),
    .C(_3368_),
    .Y(_3369_));
 sg13g2_or2_1 _7940_ (.X(_3370_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .A(_0046_));
 sg13g2_buf_1 _7941_ (.A(_3370_),
    .X(_3371_));
 sg13g2_or2_1 _7942_ (.X(_3372_),
    .B(_3281_),
    .A(_3260_));
 sg13g2_nor2_1 _7943_ (.A(_3371_),
    .B(_3372_),
    .Y(_3373_));
 sg13g2_nor3_1 _7944_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ),
    .B(net209),
    .C(_3373_),
    .Y(_3374_));
 sg13g2_a221oi_1 _7945_ (.B2(_3369_),
    .C1(_3374_),
    .B1(net40),
    .A1(_3363_),
    .Y(_0460_),
    .A2(net153));
 sg13g2_and2_1 _7946_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ),
    .B(_3368_),
    .X(_3375_));
 sg13g2_a21oi_1 _7947_ (.A1(net46),
    .A2(_3373_),
    .Y(_3376_),
    .B1(_3375_));
 sg13g2_nand2_1 _7948_ (.Y(_3377_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29] ),
    .B(net210));
 sg13g2_o21ai_1 _7949_ (.B1(_3377_),
    .Y(_0461_),
    .A1(net154),
    .A2(_3376_));
 sg13g2_nand2_1 _7950_ (.Y(_3378_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2] ),
    .B(_3368_));
 sg13g2_o21ai_1 _7951_ (.B1(_3378_),
    .Y(_3379_),
    .A1(net43),
    .A2(_3368_));
 sg13g2_mux2_1 _7952_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30] ),
    .A1(_3379_),
    .S(net138),
    .X(_0462_));
 sg13g2_buf_1 _7953_ (.A(net235),
    .X(_3380_));
 sg13g2_nor2_1 _7954_ (.A(net216),
    .B(_3373_),
    .Y(_3381_));
 sg13g2_a22oi_1 _7955_ (.Y(_3382_),
    .B1(_3381_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7956_ (.B1(_3382_),
    .Y(_0463_),
    .A1(net39),
    .A2(_3368_));
 sg13g2_mux2_1 _7957_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8] ),
    .S(net138),
    .X(_0464_));
 sg13g2_mux2_1 _7958_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9] ),
    .S(net138),
    .X(_0465_));
 sg13g2_mux2_1 _7959_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10] ),
    .S(_3365_),
    .X(_0466_));
 sg13g2_mux2_1 _7960_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11] ),
    .S(net138),
    .X(_0467_));
 sg13g2_buf_1 _7961_ (.A(net212),
    .X(_3383_));
 sg13g2_mux2_1 _7962_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8] ),
    .S(net137),
    .X(_0468_));
 sg13g2_mux2_1 _7963_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9] ),
    .S(_3383_),
    .X(_0469_));
 sg13g2_mux2_1 _7964_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10] ),
    .S(net137),
    .X(_0470_));
 sg13g2_mux2_1 _7965_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11] ),
    .S(net137),
    .X(_0471_));
 sg13g2_mux2_1 _7966_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12] ),
    .S(net137),
    .X(_0472_));
 sg13g2_mux2_1 _7967_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13] ),
    .S(net137),
    .X(_0473_));
 sg13g2_mux2_1 _7968_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18] ),
    .S(net138),
    .X(_0474_));
 sg13g2_mux2_1 _7969_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19] ),
    .S(net138),
    .X(_0475_));
 sg13g2_mux2_1 _7970_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20] ),
    .S(net138),
    .X(_0476_));
 sg13g2_mux2_1 _7971_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21] ),
    .S(_3365_),
    .X(_0477_));
 sg13g2_buf_1 _7972_ (.A(_3345_),
    .X(_3384_));
 sg13g2_mux2_1 _7973_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22] ),
    .S(net136),
    .X(_0478_));
 sg13g2_mux2_1 _7974_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23] ),
    .S(net136),
    .X(_0479_));
 sg13g2_mux2_1 _7975_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24] ),
    .S(net136),
    .X(_0480_));
 sg13g2_mux2_1 _7976_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25] ),
    .S(net136),
    .X(_0481_));
 sg13g2_mux2_1 _7977_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26] ),
    .S(net136),
    .X(_0482_));
 sg13g2_mux2_1 _7978_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27] ),
    .S(net136),
    .X(_0483_));
 sg13g2_mux2_1 _7979_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28] ),
    .S(net136),
    .X(_0484_));
 sg13g2_mux2_1 _7980_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29] ),
    .S(_3384_),
    .X(_0485_));
 sg13g2_mux2_1 _7981_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30] ),
    .S(_3384_),
    .X(_0486_));
 sg13g2_mux2_1 _7982_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31] ),
    .S(net136),
    .X(_0487_));
 sg13g2_nand2_2 _7983_ (.Y(_3385_),
    .A(_3132_),
    .B(net273));
 sg13g2_nor3_1 _7984_ (.A(net208),
    .B(net47),
    .C(_3385_),
    .Y(_3386_));
 sg13g2_a21oi_1 _7985_ (.A1(_3132_),
    .A2(net273),
    .Y(_3387_),
    .B1(net234));
 sg13g2_nor2_1 _7986_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28] ),
    .B(_3113_),
    .Y(_3388_));
 sg13g2_a221oi_1 _7987_ (.B2(_2068_),
    .C1(_3388_),
    .B1(_3387_),
    .A1(net37),
    .Y(_0488_),
    .A2(_3386_));
 sg13g2_mux2_1 _7988_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ),
    .S(_3385_),
    .X(_3389_));
 sg13g2_buf_1 _7989_ (.A(_3345_),
    .X(_3390_));
 sg13g2_mux2_1 _7990_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29] ),
    .A1(_3389_),
    .S(net135),
    .X(_0489_));
 sg13g2_nand2_1 _7991_ (.Y(_3391_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ),
    .B(_3385_));
 sg13g2_o21ai_1 _7992_ (.B1(_3391_),
    .Y(_3392_),
    .A1(net43),
    .A2(_3385_));
 sg13g2_mux2_1 _7993_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30] ),
    .A1(_3392_),
    .S(net135),
    .X(_0490_));
 sg13g2_a22oi_1 _7994_ (.Y(_3393_),
    .B1(_3387_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _7995_ (.B1(_3393_),
    .Y(_0491_),
    .A1(_3244_),
    .A2(_3385_));
 sg13g2_mux2_1 _7996_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8] ),
    .S(net135),
    .X(_0492_));
 sg13g2_mux2_1 _7997_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9] ),
    .S(_3390_),
    .X(_0493_));
 sg13g2_mux2_1 _7998_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10] ),
    .S(_3390_),
    .X(_0494_));
 sg13g2_mux2_1 _7999_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11] ),
    .S(net135),
    .X(_0495_));
 sg13g2_mux2_1 _8000_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8] ),
    .S(net137),
    .X(_0496_));
 sg13g2_mux2_1 _8001_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9] ),
    .S(net137),
    .X(_0497_));
 sg13g2_mux2_1 _8002_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10] ),
    .S(_3383_),
    .X(_0498_));
 sg13g2_mux2_1 _8003_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11] ),
    .S(net137),
    .X(_0499_));
 sg13g2_buf_1 _8004_ (.A(net212),
    .X(_3394_));
 sg13g2_mux2_1 _8005_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12] ),
    .S(net134),
    .X(_0500_));
 sg13g2_mux2_1 _8006_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13] ),
    .S(net134),
    .X(_0501_));
 sg13g2_mux2_1 _8007_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18] ),
    .S(net135),
    .X(_0502_));
 sg13g2_mux2_1 _8008_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19] ),
    .S(net135),
    .X(_0503_));
 sg13g2_mux2_1 _8009_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20] ),
    .S(net135),
    .X(_0504_));
 sg13g2_mux2_1 _8010_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21] ),
    .S(net135),
    .X(_0505_));
 sg13g2_buf_1 _8011_ (.A(_3345_),
    .X(_3395_));
 sg13g2_mux2_1 _8012_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22] ),
    .S(net133),
    .X(_0506_));
 sg13g2_mux2_1 _8013_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23] ),
    .S(net133),
    .X(_0507_));
 sg13g2_mux2_1 _8014_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24] ),
    .S(net133),
    .X(_0508_));
 sg13g2_mux2_1 _8015_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25] ),
    .S(net133),
    .X(_0509_));
 sg13g2_mux2_1 _8016_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26] ),
    .S(net133),
    .X(_0510_));
 sg13g2_mux2_1 _8017_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27] ),
    .S(net133),
    .X(_0511_));
 sg13g2_mux2_1 _8018_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28] ),
    .S(net133),
    .X(_0512_));
 sg13g2_mux2_1 _8019_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29] ),
    .S(_3395_),
    .X(_0513_));
 sg13g2_mux2_1 _8020_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30] ),
    .S(_3395_),
    .X(_0514_));
 sg13g2_mux2_1 _8021_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31] ),
    .S(net133),
    .X(_0515_));
 sg13g2_a21oi_1 _8022_ (.A1(_3262_),
    .A2(net273),
    .Y(_3396_),
    .B1(_3321_));
 sg13g2_nand2_2 _8023_ (.Y(_3397_),
    .A(_3262_),
    .B(net273));
 sg13g2_nor3_1 _8024_ (.A(net211),
    .B(_3229_),
    .C(_3397_),
    .Y(_3398_));
 sg13g2_buf_1 _8025_ (.A(_3053_),
    .X(_3399_));
 sg13g2_nor2_1 _8026_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28] ),
    .B(_3399_),
    .Y(_3400_));
 sg13g2_a221oi_1 _8027_ (.B2(net38),
    .C1(_3400_),
    .B1(_3398_),
    .A1(_3074_),
    .Y(_0516_),
    .A2(_3396_));
 sg13g2_mux2_1 _8028_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ),
    .S(_3397_),
    .X(_3401_));
 sg13g2_buf_1 _8029_ (.A(_3345_),
    .X(_3402_));
 sg13g2_mux2_1 _8030_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29] ),
    .A1(_3401_),
    .S(net132),
    .X(_0517_));
 sg13g2_nand2_1 _8031_ (.Y(_3403_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ),
    .B(_3397_));
 sg13g2_o21ai_1 _8032_ (.B1(_3403_),
    .Y(_3404_),
    .A1(_3238_),
    .A2(_3397_));
 sg13g2_mux2_1 _8033_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30] ),
    .A1(_3404_),
    .S(net132),
    .X(_0518_));
 sg13g2_a22oi_1 _8034_ (.Y(_3405_),
    .B1(_3396_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8035_ (.B1(_3405_),
    .Y(_0519_),
    .A1(_3244_),
    .A2(_3397_));
 sg13g2_mux2_1 _8036_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8] ),
    .S(net132),
    .X(_0520_));
 sg13g2_mux2_1 _8037_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9] ),
    .S(net132),
    .X(_0521_));
 sg13g2_mux2_1 _8038_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10] ),
    .S(net132),
    .X(_0522_));
 sg13g2_mux2_1 _8039_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11] ),
    .S(net132),
    .X(_0523_));
 sg13g2_mux2_1 _8040_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8] ),
    .S(net134),
    .X(_0524_));
 sg13g2_mux2_1 _8041_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9] ),
    .S(net134),
    .X(_0525_));
 sg13g2_mux2_1 _8042_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10] ),
    .S(net134),
    .X(_0526_));
 sg13g2_mux2_1 _8043_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11] ),
    .S(net134),
    .X(_0527_));
 sg13g2_mux2_1 _8044_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12] ),
    .S(net134),
    .X(_0528_));
 sg13g2_mux2_1 _8045_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13] ),
    .S(net134),
    .X(_0529_));
 sg13g2_mux2_1 _8046_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18] ),
    .S(net132),
    .X(_0530_));
 sg13g2_mux2_1 _8047_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19] ),
    .S(net132),
    .X(_0531_));
 sg13g2_mux2_1 _8048_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20] ),
    .S(_3402_),
    .X(_0532_));
 sg13g2_mux2_1 _8049_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21] ),
    .S(_3402_),
    .X(_0533_));
 sg13g2_buf_1 _8050_ (.A(_3062_),
    .X(_3406_));
 sg13g2_buf_1 _8051_ (.A(_3406_),
    .X(_3407_));
 sg13g2_mux2_1 _8052_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22] ),
    .S(net131),
    .X(_0534_));
 sg13g2_mux2_1 _8053_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23] ),
    .S(net131),
    .X(_0535_));
 sg13g2_mux2_1 _8054_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24] ),
    .S(net131),
    .X(_0536_));
 sg13g2_mux2_1 _8055_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25] ),
    .S(net131),
    .X(_0537_));
 sg13g2_mux2_1 _8056_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26] ),
    .S(_3407_),
    .X(_0538_));
 sg13g2_mux2_1 _8057_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27] ),
    .S(_3407_),
    .X(_0539_));
 sg13g2_inv_1 _8058_ (.Y(_3408_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _8059_ (.Y(_3409_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24] ),
    .B(net210));
 sg13g2_o21ai_1 _8060_ (.B1(_3409_),
    .Y(_0540_),
    .A1(_3408_),
    .A2(net154));
 sg13g2_mux2_1 _8061_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29] ),
    .S(net131),
    .X(_0541_));
 sg13g2_mux2_1 _8062_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30] ),
    .S(net131),
    .X(_0542_));
 sg13g2_mux2_1 _8063_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31] ),
    .S(net131),
    .X(_0543_));
 sg13g2_nor2_1 _8064_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .Y(_3410_));
 sg13g2_buf_2 _8065_ (.A(_3410_),
    .X(_3411_));
 sg13g2_nand2_2 _8066_ (.Y(_3412_),
    .A(_3367_),
    .B(_3411_));
 sg13g2_nor3_1 _8067_ (.A(net214),
    .B(net48),
    .C(_3412_),
    .Y(_3413_));
 sg13g2_and2_1 _8068_ (.A(_3367_),
    .B(_3411_),
    .X(_3414_));
 sg13g2_buf_1 _8069_ (.A(_3414_),
    .X(_3415_));
 sg13g2_nor3_1 _8070_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ),
    .B(net209),
    .C(_3415_),
    .Y(_3416_));
 sg13g2_a221oi_1 _8071_ (.B2(_3413_),
    .C1(_3416_),
    .B1(net40),
    .A1(_3408_),
    .Y(_0544_),
    .A2(net153));
 sg13g2_and2_1 _8072_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ),
    .B(_3412_),
    .X(_3417_));
 sg13g2_a21oi_1 _8073_ (.A1(net46),
    .A2(_3415_),
    .Y(_3418_),
    .B1(_3417_));
 sg13g2_nand2_1 _8074_ (.Y(_3419_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29] ),
    .B(net210));
 sg13g2_o21ai_1 _8075_ (.B1(_3419_),
    .Y(_0545_),
    .A1(net153),
    .A2(_3418_));
 sg13g2_buf_1 _8076_ (.A(_3237_),
    .X(_3420_));
 sg13g2_nand2_1 _8077_ (.Y(_3421_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2] ),
    .B(_3412_));
 sg13g2_o21ai_1 _8078_ (.B1(_3421_),
    .Y(_3422_),
    .A1(net42),
    .A2(_3412_));
 sg13g2_mux2_1 _8079_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30] ),
    .A1(_3422_),
    .S(net131),
    .X(_0546_));
 sg13g2_buf_8 _8080_ (.A(_3243_),
    .X(_3423_));
 sg13g2_nor2_1 _8081_ (.A(_3104_),
    .B(_3415_),
    .Y(_3424_));
 sg13g2_a22oi_1 _8082_ (.Y(_3425_),
    .B1(_3424_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8083_ (.B1(_3425_),
    .Y(_0547_),
    .A1(net36),
    .A2(_3412_));
 sg13g2_buf_1 _8084_ (.A(_3406_),
    .X(_3426_));
 sg13g2_mux2_1 _8085_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8] ),
    .S(net130),
    .X(_0548_));
 sg13g2_mux2_1 _8086_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9] ),
    .S(net130),
    .X(_0549_));
 sg13g2_mux2_1 _8087_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10] ),
    .S(net130),
    .X(_0550_));
 sg13g2_mux2_1 _8088_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11] ),
    .S(net130),
    .X(_0551_));
 sg13g2_mux2_1 _8089_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8] ),
    .S(_3394_),
    .X(_0552_));
 sg13g2_mux2_1 _8090_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9] ),
    .S(_3394_),
    .X(_0553_));
 sg13g2_buf_1 _8091_ (.A(net212),
    .X(_3427_));
 sg13g2_mux2_1 _8092_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10] ),
    .S(_3427_),
    .X(_0554_));
 sg13g2_mux2_1 _8093_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11] ),
    .S(net129),
    .X(_0555_));
 sg13g2_mux2_1 _8094_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12] ),
    .S(net129),
    .X(_0556_));
 sg13g2_mux2_1 _8095_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13] ),
    .S(net129),
    .X(_0557_));
 sg13g2_mux2_1 _8096_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18] ),
    .S(net130),
    .X(_0558_));
 sg13g2_mux2_1 _8097_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19] ),
    .S(_3426_),
    .X(_0559_));
 sg13g2_mux2_1 _8098_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20] ),
    .S(net130),
    .X(_0560_));
 sg13g2_mux2_1 _8099_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21] ),
    .S(net130),
    .X(_0561_));
 sg13g2_mux2_1 _8100_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22] ),
    .S(net130),
    .X(_0562_));
 sg13g2_mux2_1 _8101_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23] ),
    .S(_3426_),
    .X(_0563_));
 sg13g2_buf_1 _8102_ (.A(_3406_),
    .X(_3428_));
 sg13g2_mux2_1 _8103_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24] ),
    .S(net128),
    .X(_0564_));
 sg13g2_mux2_1 _8104_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25] ),
    .S(net128),
    .X(_0565_));
 sg13g2_mux2_1 _8105_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26] ),
    .S(_3428_),
    .X(_0566_));
 sg13g2_mux2_1 _8106_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27] ),
    .S(net128),
    .X(_0567_));
 sg13g2_mux2_1 _8107_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28] ),
    .S(net128),
    .X(_0568_));
 sg13g2_mux2_1 _8108_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29] ),
    .S(_3428_),
    .X(_0569_));
 sg13g2_mux2_1 _8109_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30] ),
    .S(net128),
    .X(_0570_));
 sg13g2_mux2_1 _8110_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31] ),
    .S(net128),
    .X(_0571_));
 sg13g2_nand2_2 _8111_ (.Y(_3429_),
    .A(_3283_),
    .B(net273));
 sg13g2_nor3_1 _8112_ (.A(net208),
    .B(net47),
    .C(_3429_),
    .Y(_3430_));
 sg13g2_a21oi_1 _8113_ (.A1(_3283_),
    .A2(net273),
    .Y(_3431_),
    .B1(net234));
 sg13g2_nor2_1 _8114_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3432_));
 sg13g2_a221oi_1 _8115_ (.B2(_3078_),
    .C1(_3432_),
    .B1(_3431_),
    .A1(net37),
    .Y(_0572_),
    .A2(_3430_));
 sg13g2_mux2_1 _8116_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ),
    .S(_3429_),
    .X(_3433_));
 sg13g2_mux2_1 _8117_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29] ),
    .A1(_3433_),
    .S(net128),
    .X(_0573_));
 sg13g2_nand2_1 _8118_ (.Y(_3434_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ),
    .B(_3429_));
 sg13g2_o21ai_1 _8119_ (.B1(_3434_),
    .Y(_3435_),
    .A1(net42),
    .A2(_3429_));
 sg13g2_mux2_1 _8120_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30] ),
    .A1(_3435_),
    .S(net128),
    .X(_0574_));
 sg13g2_a22oi_1 _8121_ (.Y(_3436_),
    .B1(_3431_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ),
    .A2(_3380_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8122_ (.B1(_3436_),
    .Y(_0575_),
    .A1(net36),
    .A2(_3429_));
 sg13g2_buf_1 _8123_ (.A(_3406_),
    .X(_3437_));
 sg13g2_mux2_1 _8124_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8] ),
    .S(net127),
    .X(_0576_));
 sg13g2_mux2_1 _8125_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9] ),
    .S(net127),
    .X(_0577_));
 sg13g2_mux2_1 _8126_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10] ),
    .S(net127),
    .X(_0578_));
 sg13g2_mux2_1 _8127_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11] ),
    .S(net127),
    .X(_0579_));
 sg13g2_mux2_1 _8128_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8] ),
    .S(_3427_),
    .X(_0580_));
 sg13g2_mux2_1 _8129_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9] ),
    .S(net129),
    .X(_0581_));
 sg13g2_mux2_1 _8130_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10] ),
    .S(net129),
    .X(_0582_));
 sg13g2_mux2_1 _8131_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11] ),
    .S(net129),
    .X(_0583_));
 sg13g2_mux2_1 _8132_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12] ),
    .S(net129),
    .X(_0584_));
 sg13g2_mux2_1 _8133_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13] ),
    .S(net129),
    .X(_0585_));
 sg13g2_mux2_1 _8134_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18] ),
    .S(net127),
    .X(_0586_));
 sg13g2_mux2_1 _8135_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19] ),
    .S(_3437_),
    .X(_0587_));
 sg13g2_mux2_1 _8136_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20] ),
    .S(net127),
    .X(_0588_));
 sg13g2_mux2_1 _8137_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21] ),
    .S(net127),
    .X(_0589_));
 sg13g2_mux2_1 _8138_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22] ),
    .S(net127),
    .X(_0590_));
 sg13g2_mux2_1 _8139_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23] ),
    .S(_3437_),
    .X(_0591_));
 sg13g2_buf_1 _8140_ (.A(_3406_),
    .X(_3438_));
 sg13g2_mux2_1 _8141_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24] ),
    .S(net126),
    .X(_0592_));
 sg13g2_mux2_1 _8142_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25] ),
    .S(net126),
    .X(_0593_));
 sg13g2_mux2_1 _8143_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26] ),
    .S(net126),
    .X(_0594_));
 sg13g2_mux2_1 _8144_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27] ),
    .S(_3438_),
    .X(_0595_));
 sg13g2_mux2_1 _8145_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28] ),
    .S(net126),
    .X(_0596_));
 sg13g2_mux2_1 _8146_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29] ),
    .S(net126),
    .X(_0597_));
 sg13g2_mux2_1 _8147_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30] ),
    .S(net126),
    .X(_0598_));
 sg13g2_mux2_1 _8148_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31] ),
    .S(_3438_),
    .X(_0599_));
 sg13g2_nand2_2 _8149_ (.Y(_3439_),
    .A(_3302_),
    .B(_3350_));
 sg13g2_nor3_1 _8150_ (.A(_3279_),
    .B(net47),
    .C(_3439_),
    .Y(_3440_));
 sg13g2_nor2_1 _8151_ (.A(_3306_),
    .B(_3371_),
    .Y(_3441_));
 sg13g2_nor2_1 _8152_ (.A(_3286_),
    .B(_3441_),
    .Y(_3442_));
 sg13g2_nor2_1 _8153_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3443_));
 sg13g2_a221oi_1 _8154_ (.B2(_1925_),
    .C1(_3443_),
    .B1(_3442_),
    .A1(_3347_),
    .Y(_0600_),
    .A2(_3440_));
 sg13g2_and2_1 _8155_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ),
    .B(_3439_),
    .X(_3444_));
 sg13g2_a21oi_1 _8156_ (.A1(net46),
    .A2(_3441_),
    .Y(_3445_),
    .B1(_3444_));
 sg13g2_nand2_1 _8157_ (.Y(_3446_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29] ),
    .B(_3255_));
 sg13g2_o21ai_1 _8158_ (.B1(_3446_),
    .Y(_0601_),
    .A1(net153),
    .A2(_3445_));
 sg13g2_nand2_1 _8159_ (.Y(_3447_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ),
    .B(_3439_));
 sg13g2_o21ai_1 _8160_ (.B1(_3447_),
    .Y(_3448_),
    .A1(net42),
    .A2(_3439_));
 sg13g2_mux2_1 _8161_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30] ),
    .A1(_3448_),
    .S(net126),
    .X(_0602_));
 sg13g2_a22oi_1 _8162_ (.Y(_3449_),
    .B1(_3442_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8163_ (.B1(_3449_),
    .Y(_0603_),
    .A1(net36),
    .A2(_3439_));
 sg13g2_mux2_1 _8164_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8] ),
    .S(net126),
    .X(_0604_));
 sg13g2_buf_1 _8165_ (.A(_3406_),
    .X(_3450_));
 sg13g2_mux2_1 _8166_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9] ),
    .S(net125),
    .X(_0605_));
 sg13g2_mux2_1 _8167_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10] ),
    .S(net125),
    .X(_0606_));
 sg13g2_mux2_1 _8168_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11] ),
    .S(net125),
    .X(_0607_));
 sg13g2_buf_2 _8169_ (.A(net236),
    .X(_3451_));
 sg13g2_buf_1 _8170_ (.A(_3451_),
    .X(_3452_));
 sg13g2_mux2_1 _8171_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8] ),
    .S(net124),
    .X(_0608_));
 sg13g2_mux2_1 _8172_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9] ),
    .S(net124),
    .X(_0609_));
 sg13g2_mux2_1 _8173_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10] ),
    .S(net124),
    .X(_0610_));
 sg13g2_mux2_1 _8174_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11] ),
    .S(_3452_),
    .X(_0611_));
 sg13g2_mux2_1 _8175_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12] ),
    .S(net124),
    .X(_0612_));
 sg13g2_mux2_1 _8176_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13] ),
    .S(net124),
    .X(_0613_));
 sg13g2_mux2_1 _8177_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18] ),
    .S(net125),
    .X(_0614_));
 sg13g2_mux2_1 _8178_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19] ),
    .S(net125),
    .X(_0615_));
 sg13g2_mux2_1 _8179_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20] ),
    .S(net125),
    .X(_0616_));
 sg13g2_mux2_1 _8180_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21] ),
    .S(net125),
    .X(_0617_));
 sg13g2_mux2_1 _8181_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22] ),
    .S(_3450_),
    .X(_0618_));
 sg13g2_mux2_1 _8182_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23] ),
    .S(_3450_),
    .X(_0619_));
 sg13g2_mux2_1 _8183_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24] ),
    .S(net125),
    .X(_0620_));
 sg13g2_buf_1 _8184_ (.A(_3406_),
    .X(_3453_));
 sg13g2_mux2_1 _8185_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25] ),
    .S(_3453_),
    .X(_0621_));
 sg13g2_mux2_1 _8186_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26] ),
    .S(net123),
    .X(_0622_));
 sg13g2_mux2_1 _8187_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27] ),
    .S(net123),
    .X(_0623_));
 sg13g2_mux2_1 _8188_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28] ),
    .S(net123),
    .X(_0624_));
 sg13g2_mux2_1 _8189_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29] ),
    .S(_3453_),
    .X(_0625_));
 sg13g2_mux2_1 _8190_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30] ),
    .S(net123),
    .X(_0626_));
 sg13g2_mux2_1 _8191_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31] ),
    .S(net123),
    .X(_0627_));
 sg13g2_nand2_2 _8192_ (.Y(_3454_),
    .A(_3320_),
    .B(_3350_));
 sg13g2_nor3_1 _8193_ (.A(_3279_),
    .B(net47),
    .C(_3454_),
    .Y(_3455_));
 sg13g2_a21oi_1 _8194_ (.A1(_3320_),
    .A2(_3351_),
    .Y(_3456_),
    .B1(_3286_));
 sg13g2_nor2_1 _8195_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28] ),
    .B(_3399_),
    .Y(_3457_));
 sg13g2_a221oi_1 _8196_ (.B2(_3082_),
    .C1(_3457_),
    .B1(_3456_),
    .A1(_3347_),
    .Y(_0628_),
    .A2(_3455_));
 sg13g2_mux2_1 _8197_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ),
    .S(_3454_),
    .X(_3458_));
 sg13g2_mux2_1 _8198_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29] ),
    .A1(_3458_),
    .S(net123),
    .X(_0629_));
 sg13g2_nand2_1 _8199_ (.Y(_3459_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ),
    .B(_3454_));
 sg13g2_o21ai_1 _8200_ (.B1(_3459_),
    .Y(_3460_),
    .A1(net42),
    .A2(_3454_));
 sg13g2_mux2_1 _8201_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30] ),
    .A1(_3460_),
    .S(net123),
    .X(_0630_));
 sg13g2_a22oi_1 _8202_ (.Y(_3461_),
    .B1(_3456_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ),
    .A2(_3380_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8203_ (.B1(_3461_),
    .Y(_0631_),
    .A1(net36),
    .A2(_3454_));
 sg13g2_mux2_1 _8204_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8] ),
    .S(net123),
    .X(_0632_));
 sg13g2_buf_1 _8205_ (.A(_3062_),
    .X(_3462_));
 sg13g2_buf_1 _8206_ (.A(_3462_),
    .X(_3463_));
 sg13g2_mux2_1 _8207_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9] ),
    .S(net122),
    .X(_0633_));
 sg13g2_mux2_1 _8208_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10] ),
    .S(net122),
    .X(_0634_));
 sg13g2_mux2_1 _8209_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11] ),
    .S(net122),
    .X(_0635_));
 sg13g2_mux2_1 _8210_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8] ),
    .S(net124),
    .X(_0636_));
 sg13g2_mux2_1 _8211_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9] ),
    .S(net124),
    .X(_0637_));
 sg13g2_mux2_1 _8212_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10] ),
    .S(net124),
    .X(_0638_));
 sg13g2_mux2_1 _8213_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11] ),
    .S(_3452_),
    .X(_0639_));
 sg13g2_buf_1 _8214_ (.A(_3451_),
    .X(_3464_));
 sg13g2_mux2_1 _8215_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12] ),
    .S(net121),
    .X(_0640_));
 sg13g2_mux2_1 _8216_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13] ),
    .S(net121),
    .X(_0641_));
 sg13g2_mux2_1 _8217_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18] ),
    .S(net122),
    .X(_0642_));
 sg13g2_mux2_1 _8218_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19] ),
    .S(net122),
    .X(_0643_));
 sg13g2_mux2_1 _8219_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20] ),
    .S(net122),
    .X(_0644_));
 sg13g2_mux2_1 _8220_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21] ),
    .S(net122),
    .X(_0645_));
 sg13g2_mux2_1 _8221_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22] ),
    .S(_3463_),
    .X(_0646_));
 sg13g2_mux2_1 _8222_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23] ),
    .S(net122),
    .X(_0647_));
 sg13g2_mux2_1 _8223_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24] ),
    .S(_3463_),
    .X(_0648_));
 sg13g2_buf_1 _8224_ (.A(_3462_),
    .X(_3465_));
 sg13g2_mux2_1 _8225_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25] ),
    .S(net120),
    .X(_0649_));
 sg13g2_mux2_1 _8226_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26] ),
    .S(net120),
    .X(_0650_));
 sg13g2_mux2_1 _8227_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27] ),
    .S(net120),
    .X(_0651_));
 sg13g2_inv_1 _8228_ (.Y(_3466_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _8229_ (.Y(_3467_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24] ),
    .B(_3255_));
 sg13g2_o21ai_1 _8230_ (.B1(_3467_),
    .Y(_0652_),
    .A1(_3466_),
    .A2(_3253_));
 sg13g2_mux2_1 _8231_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29] ),
    .S(net120),
    .X(_0653_));
 sg13g2_mux2_1 _8232_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30] ),
    .S(_3465_),
    .X(_0654_));
 sg13g2_mux2_1 _8233_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31] ),
    .S(net120),
    .X(_0655_));
 sg13g2_nand2_1 _8234_ (.Y(_3468_),
    .A(_3334_),
    .B(_3351_));
 sg13g2_nor3_1 _8235_ (.A(net214),
    .B(_3258_),
    .C(_3468_),
    .Y(_3469_));
 sg13g2_nor3_2 _8236_ (.A(_3130_),
    .B(_3300_),
    .C(_3371_),
    .Y(_3470_));
 sg13g2_nor3_1 _8237_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ),
    .B(_3265_),
    .C(_3470_),
    .Y(_3471_));
 sg13g2_a221oi_1 _8238_ (.B2(_3469_),
    .C1(_3471_),
    .B1(_3223_),
    .A1(_3466_),
    .Y(_0656_),
    .A2(net153));
 sg13g2_nor2b_1 _8239_ (.A(_3470_),
    .B_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ),
    .Y(_3472_));
 sg13g2_a21oi_1 _8240_ (.A1(_3234_),
    .A2(_3470_),
    .Y(_3473_),
    .B1(_3472_));
 sg13g2_buf_1 _8241_ (.A(_3254_),
    .X(_3474_));
 sg13g2_nand2_1 _8242_ (.Y(_3475_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29] ),
    .B(net205));
 sg13g2_o21ai_1 _8243_ (.B1(_3475_),
    .Y(_0657_),
    .A1(net153),
    .A2(_3473_));
 sg13g2_nand2_1 _8244_ (.Y(_3476_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ),
    .B(_3468_));
 sg13g2_o21ai_1 _8245_ (.B1(_3476_),
    .Y(_3477_),
    .A1(net42),
    .A2(_3468_));
 sg13g2_mux2_1 _8246_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30] ),
    .A1(_3477_),
    .S(net120),
    .X(_0658_));
 sg13g2_nor2_1 _8247_ (.A(net216),
    .B(_3470_),
    .Y(_3478_));
 sg13g2_a22oi_1 _8248_ (.Y(_3479_),
    .B1(_3478_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8249_ (.B1(_3479_),
    .Y(_0659_),
    .A1(net36),
    .A2(_3468_));
 sg13g2_mux2_1 _8250_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8] ),
    .S(net120),
    .X(_0660_));
 sg13g2_mux2_1 _8251_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9] ),
    .S(net120),
    .X(_0661_));
 sg13g2_mux2_1 _8252_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10] ),
    .S(_3465_),
    .X(_0662_));
 sg13g2_buf_1 _8253_ (.A(_3462_),
    .X(_3480_));
 sg13g2_mux2_1 _8254_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11] ),
    .S(net119),
    .X(_0663_));
 sg13g2_mux2_1 _8255_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8] ),
    .S(net121),
    .X(_0664_));
 sg13g2_mux2_1 _8256_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9] ),
    .S(net121),
    .X(_0665_));
 sg13g2_mux2_1 _8257_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10] ),
    .S(net121),
    .X(_0666_));
 sg13g2_mux2_1 _8258_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11] ),
    .S(net121),
    .X(_0667_));
 sg13g2_mux2_1 _8259_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12] ),
    .S(_3464_),
    .X(_0668_));
 sg13g2_mux2_1 _8260_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13] ),
    .S(net121),
    .X(_0669_));
 sg13g2_mux2_1 _8261_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18] ),
    .S(net119),
    .X(_0670_));
 sg13g2_mux2_1 _8262_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19] ),
    .S(net119),
    .X(_0671_));
 sg13g2_mux2_1 _8263_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20] ),
    .S(net119),
    .X(_0672_));
 sg13g2_mux2_1 _8264_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21] ),
    .S(net119),
    .X(_0673_));
 sg13g2_mux2_1 _8265_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22] ),
    .S(net119),
    .X(_0674_));
 sg13g2_mux2_1 _8266_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23] ),
    .S(net119),
    .X(_0675_));
 sg13g2_mux2_1 _8267_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24] ),
    .S(net119),
    .X(_0676_));
 sg13g2_mux2_1 _8268_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25] ),
    .S(_3480_),
    .X(_0677_));
 sg13g2_mux2_1 _8269_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26] ),
    .S(_3480_),
    .X(_0678_));
 sg13g2_buf_1 _8270_ (.A(_3462_),
    .X(_3481_));
 sg13g2_mux2_1 _8271_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27] ),
    .S(net118),
    .X(_0679_));
 sg13g2_mux2_1 _8272_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28] ),
    .S(net118),
    .X(_0680_));
 sg13g2_mux2_1 _8273_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29] ),
    .S(net118),
    .X(_0681_));
 sg13g2_mux2_1 _8274_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30] ),
    .S(net118),
    .X(_0682_));
 sg13g2_mux2_1 _8275_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31] ),
    .S(net118),
    .X(_0683_));
 sg13g2_nor2_1 _8276_ (.A(_0047_),
    .B(_0046_),
    .Y(_3482_));
 sg13g2_buf_2 _8277_ (.A(_3482_),
    .X(_3483_));
 sg13g2_buf_1 _8278_ (.A(_3483_),
    .X(_3484_));
 sg13g2_nand2_2 _8279_ (.Y(_3485_),
    .A(_3353_),
    .B(net272));
 sg13g2_nor3_1 _8280_ (.A(net208),
    .B(_3348_),
    .C(_3485_),
    .Y(_3486_));
 sg13g2_a21oi_1 _8281_ (.A1(_3353_),
    .A2(net272),
    .Y(_3487_),
    .B1(net235));
 sg13g2_nor2_1 _8282_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3488_));
 sg13g2_a221oi_1 _8283_ (.B2(_3085_),
    .C1(_3488_),
    .B1(_3487_),
    .A1(net37),
    .Y(_0684_),
    .A2(_3486_));
 sg13g2_mux2_1 _8284_ (.A0(net45),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ),
    .S(_3485_),
    .X(_3489_));
 sg13g2_mux2_1 _8285_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29] ),
    .A1(_3489_),
    .S(_3481_),
    .X(_0685_));
 sg13g2_nand2_1 _8286_ (.Y(_3490_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ),
    .B(_3485_));
 sg13g2_o21ai_1 _8287_ (.B1(_3490_),
    .Y(_3491_),
    .A1(net42),
    .A2(_3485_));
 sg13g2_mux2_1 _8288_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30] ),
    .A1(_3491_),
    .S(net118),
    .X(_0686_));
 sg13g2_a22oi_1 _8289_ (.Y(_3492_),
    .B1(_3487_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8290_ (.B1(_3492_),
    .Y(_0687_),
    .A1(net36),
    .A2(_3485_));
 sg13g2_mux2_1 _8291_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8] ),
    .S(_3481_),
    .X(_0688_));
 sg13g2_mux2_1 _8292_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9] ),
    .S(net118),
    .X(_0689_));
 sg13g2_mux2_1 _8293_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10] ),
    .S(net118),
    .X(_0690_));
 sg13g2_buf_1 _8294_ (.A(_3462_),
    .X(_3493_));
 sg13g2_mux2_1 _8295_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11] ),
    .S(_3493_),
    .X(_0691_));
 sg13g2_mux2_1 _8296_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8] ),
    .S(_3464_),
    .X(_0692_));
 sg13g2_mux2_1 _8297_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9] ),
    .S(net121),
    .X(_0693_));
 sg13g2_buf_1 _8298_ (.A(_3451_),
    .X(_3494_));
 sg13g2_mux2_1 _8299_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10] ),
    .S(net116),
    .X(_0694_));
 sg13g2_mux2_1 _8300_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11] ),
    .S(_3494_),
    .X(_0695_));
 sg13g2_mux2_1 _8301_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12] ),
    .S(net116),
    .X(_0696_));
 sg13g2_mux2_1 _8302_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13] ),
    .S(net116),
    .X(_0697_));
 sg13g2_mux2_1 _8303_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18] ),
    .S(net117),
    .X(_0698_));
 sg13g2_mux2_1 _8304_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19] ),
    .S(net117),
    .X(_0699_));
 sg13g2_mux2_1 _8305_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20] ),
    .S(net117),
    .X(_0700_));
 sg13g2_mux2_1 _8306_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21] ),
    .S(net117),
    .X(_0701_));
 sg13g2_mux2_1 _8307_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22] ),
    .S(net117),
    .X(_0702_));
 sg13g2_mux2_1 _8308_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23] ),
    .S(net117),
    .X(_0703_));
 sg13g2_mux2_1 _8309_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24] ),
    .S(net117),
    .X(_0704_));
 sg13g2_mux2_1 _8310_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25] ),
    .S(net117),
    .X(_0705_));
 sg13g2_mux2_1 _8311_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26] ),
    .S(_3493_),
    .X(_0706_));
 sg13g2_buf_1 _8312_ (.A(_3462_),
    .X(_3495_));
 sg13g2_mux2_1 _8313_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27] ),
    .S(net115),
    .X(_0707_));
 sg13g2_inv_1 _8314_ (.Y(_3496_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _8315_ (.Y(_3497_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24] ),
    .B(net205));
 sg13g2_o21ai_1 _8316_ (.B1(_3497_),
    .Y(_0708_),
    .A1(_3496_),
    .A2(_3253_));
 sg13g2_mux2_1 _8317_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29] ),
    .S(net115),
    .X(_0709_));
 sg13g2_mux2_1 _8318_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30] ),
    .S(net115),
    .X(_0710_));
 sg13g2_mux2_1 _8319_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31] ),
    .S(net115),
    .X(_0711_));
 sg13g2_nand2_2 _8320_ (.Y(_3498_),
    .A(_3367_),
    .B(_3483_));
 sg13g2_nor3_1 _8321_ (.A(net214),
    .B(_3258_),
    .C(_3498_),
    .Y(_3499_));
 sg13g2_or2_1 _8322_ (.X(_3500_),
    .B(_0046_),
    .A(_0047_));
 sg13g2_nor2_1 _8323_ (.A(_3372_),
    .B(_3500_),
    .Y(_3501_));
 sg13g2_nor3_1 _8324_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ),
    .B(_3265_),
    .C(_3501_),
    .Y(_3502_));
 sg13g2_a221oi_1 _8325_ (.B2(_3499_),
    .C1(_3502_),
    .B1(_3223_),
    .A1(_3496_),
    .Y(_0712_),
    .A2(_3105_));
 sg13g2_and2_1 _8326_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ),
    .B(_3498_),
    .X(_3503_));
 sg13g2_a21oi_1 _8327_ (.A1(_3234_),
    .A2(_3501_),
    .Y(_3504_),
    .B1(_3503_));
 sg13g2_nand2_1 _8328_ (.Y(_3505_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29] ),
    .B(net205));
 sg13g2_o21ai_1 _8329_ (.B1(_3505_),
    .Y(_0713_),
    .A1(_3257_),
    .A2(_3504_));
 sg13g2_nand2_1 _8330_ (.Y(_3506_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ),
    .B(_3498_));
 sg13g2_o21ai_1 _8331_ (.B1(_3506_),
    .Y(_3507_),
    .A1(net42),
    .A2(_3498_));
 sg13g2_mux2_1 _8332_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30] ),
    .A1(_3507_),
    .S(net115),
    .X(_0714_));
 sg13g2_nor2_1 _8333_ (.A(net212),
    .B(_3501_),
    .Y(_3508_));
 sg13g2_a22oi_1 _8334_ (.Y(_3509_),
    .B1(_3508_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ),
    .A2(net207),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8335_ (.B1(_3509_),
    .Y(_0715_),
    .A1(net36),
    .A2(_3498_));
 sg13g2_mux2_1 _8336_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8] ),
    .S(_3495_),
    .X(_0716_));
 sg13g2_mux2_1 _8337_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9] ),
    .S(net115),
    .X(_0717_));
 sg13g2_mux2_1 _8338_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10] ),
    .S(_3495_),
    .X(_0718_));
 sg13g2_mux2_1 _8339_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11] ),
    .S(net115),
    .X(_0719_));
 sg13g2_mux2_1 _8340_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8] ),
    .S(_3494_),
    .X(_0720_));
 sg13g2_mux2_1 _8341_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9] ),
    .S(net116),
    .X(_0721_));
 sg13g2_mux2_1 _8342_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10] ),
    .S(net116),
    .X(_0722_));
 sg13g2_mux2_1 _8343_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11] ),
    .S(net116),
    .X(_0723_));
 sg13g2_mux2_1 _8344_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12] ),
    .S(net116),
    .X(_0724_));
 sg13g2_mux2_1 _8345_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13] ),
    .S(net116),
    .X(_0725_));
 sg13g2_mux2_1 _8346_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18] ),
    .S(net115),
    .X(_0726_));
 sg13g2_buf_1 _8347_ (.A(_3462_),
    .X(_3510_));
 sg13g2_mux2_1 _8348_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19] ),
    .S(_3510_),
    .X(_0727_));
 sg13g2_mux2_1 _8349_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20] ),
    .S(net114),
    .X(_0728_));
 sg13g2_mux2_1 _8350_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21] ),
    .S(net114),
    .X(_0729_));
 sg13g2_mux2_1 _8351_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22] ),
    .S(net114),
    .X(_0730_));
 sg13g2_mux2_1 _8352_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23] ),
    .S(_3510_),
    .X(_0731_));
 sg13g2_mux2_1 _8353_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24] ),
    .S(net114),
    .X(_0732_));
 sg13g2_mux2_1 _8354_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25] ),
    .S(net114),
    .X(_0733_));
 sg13g2_mux2_1 _8355_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26] ),
    .S(net114),
    .X(_0734_));
 sg13g2_mux2_1 _8356_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27] ),
    .S(net114),
    .X(_0735_));
 sg13g2_mux2_1 _8357_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28] ),
    .S(net114),
    .X(_0736_));
 sg13g2_buf_1 _8358_ (.A(_3062_),
    .X(_3511_));
 sg13g2_buf_1 _8359_ (.A(_3511_),
    .X(_3512_));
 sg13g2_mux2_1 _8360_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29] ),
    .S(net113),
    .X(_0737_));
 sg13g2_mux2_1 _8361_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30] ),
    .S(net113),
    .X(_0738_));
 sg13g2_mux2_1 _8362_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31] ),
    .S(net113),
    .X(_0739_));
 sg13g2_a21oi_1 _8363_ (.A1(_3132_),
    .A2(net272),
    .Y(_3513_),
    .B1(_3321_));
 sg13g2_nand2_2 _8364_ (.Y(_3514_),
    .A(_3132_),
    .B(net272));
 sg13g2_nor3_1 _8365_ (.A(net211),
    .B(_3229_),
    .C(_3514_),
    .Y(_3515_));
 sg13g2_nor2_1 _8366_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3516_));
 sg13g2_a221oi_1 _8367_ (.B2(_3278_),
    .C1(_3516_),
    .B1(_3515_),
    .A1(_3088_),
    .Y(_0740_),
    .A2(_3513_));
 sg13g2_mux2_1 _8368_ (.A0(_3326_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ),
    .S(_3514_),
    .X(_3517_));
 sg13g2_mux2_1 _8369_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29] ),
    .A1(_3517_),
    .S(net113),
    .X(_0741_));
 sg13g2_nand2_1 _8370_ (.Y(_3518_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ),
    .B(_3514_));
 sg13g2_o21ai_1 _8371_ (.B1(_3518_),
    .Y(_3519_),
    .A1(net42),
    .A2(_3514_));
 sg13g2_mux2_1 _8372_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30] ),
    .A1(_3519_),
    .S(net113),
    .X(_0742_));
 sg13g2_buf_1 _8373_ (.A(net235),
    .X(_3520_));
 sg13g2_a22oi_1 _8374_ (.Y(_3521_),
    .B1(_3513_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8375_ (.B1(_3521_),
    .Y(_0743_),
    .A1(net36),
    .A2(_3514_));
 sg13g2_mux2_1 _8376_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8] ),
    .S(net113),
    .X(_0744_));
 sg13g2_mux2_1 _8377_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9] ),
    .S(_3512_),
    .X(_0745_));
 sg13g2_mux2_1 _8378_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10] ),
    .S(_3512_),
    .X(_0746_));
 sg13g2_mux2_1 _8379_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11] ),
    .S(net113),
    .X(_0747_));
 sg13g2_buf_1 _8380_ (.A(_3451_),
    .X(_3522_));
 sg13g2_mux2_1 _8381_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8] ),
    .S(net112),
    .X(_0748_));
 sg13g2_mux2_1 _8382_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9] ),
    .S(_3522_),
    .X(_0749_));
 sg13g2_mux2_1 _8383_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10] ),
    .S(net112),
    .X(_0750_));
 sg13g2_mux2_1 _8384_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11] ),
    .S(net112),
    .X(_0751_));
 sg13g2_mux2_1 _8385_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12] ),
    .S(net112),
    .X(_0752_));
 sg13g2_mux2_1 _8386_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13] ),
    .S(net112),
    .X(_0753_));
 sg13g2_mux2_1 _8387_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18] ),
    .S(net113),
    .X(_0754_));
 sg13g2_buf_1 _8388_ (.A(_3511_),
    .X(_3523_));
 sg13g2_mux2_1 _8389_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19] ),
    .S(net111),
    .X(_0755_));
 sg13g2_mux2_1 _8390_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20] ),
    .S(net111),
    .X(_0756_));
 sg13g2_mux2_1 _8391_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21] ),
    .S(net111),
    .X(_0757_));
 sg13g2_mux2_1 _8392_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22] ),
    .S(net111),
    .X(_0758_));
 sg13g2_mux2_1 _8393_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23] ),
    .S(net111),
    .X(_0759_));
 sg13g2_mux2_1 _8394_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24] ),
    .S(_3523_),
    .X(_0760_));
 sg13g2_mux2_1 _8395_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25] ),
    .S(_3523_),
    .X(_0761_));
 sg13g2_mux2_1 _8396_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26] ),
    .S(net111),
    .X(_0762_));
 sg13g2_mux2_1 _8397_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27] ),
    .S(net111),
    .X(_0763_));
 sg13g2_mux2_1 _8398_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28] ),
    .S(net111),
    .X(_0764_));
 sg13g2_buf_1 _8399_ (.A(_3511_),
    .X(_3524_));
 sg13g2_mux2_1 _8400_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29] ),
    .S(net110),
    .X(_0765_));
 sg13g2_mux2_1 _8401_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30] ),
    .S(net110),
    .X(_0766_));
 sg13g2_mux2_1 _8402_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31] ),
    .S(net110),
    .X(_0767_));
 sg13g2_a21oi_1 _8403_ (.A1(_3262_),
    .A2(net272),
    .Y(_3525_),
    .B1(net233));
 sg13g2_nand2_2 _8404_ (.Y(_3526_),
    .A(_3262_),
    .B(net272));
 sg13g2_nor3_1 _8405_ (.A(_3252_),
    .B(net49),
    .C(_3526_),
    .Y(_3527_));
 sg13g2_nor2_1 _8406_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3528_));
 sg13g2_a221oi_1 _8407_ (.B2(_3278_),
    .C1(_3528_),
    .B1(_3527_),
    .A1(_3091_),
    .Y(_0768_),
    .A2(_3525_));
 sg13g2_mux2_1 _8408_ (.A0(_3326_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ),
    .S(_3526_),
    .X(_3529_));
 sg13g2_mux2_1 _8409_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29] ),
    .A1(_3529_),
    .S(net110),
    .X(_0769_));
 sg13g2_nand2_1 _8410_ (.Y(_3530_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ),
    .B(_3526_));
 sg13g2_o21ai_1 _8411_ (.B1(_3530_),
    .Y(_3531_),
    .A1(_3420_),
    .A2(_3526_));
 sg13g2_mux2_1 _8412_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30] ),
    .A1(_3531_),
    .S(net110),
    .X(_0770_));
 sg13g2_a22oi_1 _8413_ (.Y(_3532_),
    .B1(_3525_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8414_ (.B1(_3532_),
    .Y(_0771_),
    .A1(_3423_),
    .A2(_3526_));
 sg13g2_mux2_1 _8415_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8] ),
    .S(net110),
    .X(_0772_));
 sg13g2_mux2_1 _8416_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9] ),
    .S(net110),
    .X(_0773_));
 sg13g2_mux2_1 _8417_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10] ),
    .S(net110),
    .X(_0774_));
 sg13g2_mux2_1 _8418_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11] ),
    .S(_3524_),
    .X(_0775_));
 sg13g2_mux2_1 _8419_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8] ),
    .S(net112),
    .X(_0776_));
 sg13g2_mux2_1 _8420_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9] ),
    .S(net112),
    .X(_0777_));
 sg13g2_mux2_1 _8421_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10] ),
    .S(_3522_),
    .X(_0778_));
 sg13g2_mux2_1 _8422_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11] ),
    .S(net112),
    .X(_0779_));
 sg13g2_buf_1 _8423_ (.A(_3451_),
    .X(_3533_));
 sg13g2_mux2_1 _8424_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12] ),
    .S(net109),
    .X(_0780_));
 sg13g2_mux2_1 _8425_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13] ),
    .S(net109),
    .X(_0781_));
 sg13g2_mux2_1 _8426_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18] ),
    .S(_3524_),
    .X(_0782_));
 sg13g2_buf_1 _8427_ (.A(_3511_),
    .X(_3534_));
 sg13g2_mux2_1 _8428_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19] ),
    .S(net108),
    .X(_0783_));
 sg13g2_mux2_1 _8429_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20] ),
    .S(net108),
    .X(_0784_));
 sg13g2_mux2_1 _8430_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21] ),
    .S(net108),
    .X(_0785_));
 sg13g2_mux2_1 _8431_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22] ),
    .S(net108),
    .X(_0786_));
 sg13g2_mux2_1 _8432_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23] ),
    .S(net108),
    .X(_0787_));
 sg13g2_mux2_1 _8433_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24] ),
    .S(net108),
    .X(_0788_));
 sg13g2_mux2_1 _8434_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25] ),
    .S(_3534_),
    .X(_0789_));
 sg13g2_mux2_1 _8435_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26] ),
    .S(net108),
    .X(_0790_));
 sg13g2_mux2_1 _8436_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27] ),
    .S(_3534_),
    .X(_0791_));
 sg13g2_mux2_1 _8437_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28] ),
    .S(net108),
    .X(_0792_));
 sg13g2_buf_1 _8438_ (.A(_3511_),
    .X(_3535_));
 sg13g2_mux2_1 _8439_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29] ),
    .S(net107),
    .X(_0793_));
 sg13g2_mux2_1 _8440_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30] ),
    .S(net107),
    .X(_0794_));
 sg13g2_mux2_1 _8441_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31] ),
    .S(net107),
    .X(_0795_));
 sg13g2_nand2_2 _8442_ (.Y(_3536_),
    .A(_3283_),
    .B(_3484_));
 sg13g2_nor3_1 _8443_ (.A(net208),
    .B(net47),
    .C(_3536_),
    .Y(_3537_));
 sg13g2_a21oi_1 _8444_ (.A1(_3283_),
    .A2(_3484_),
    .Y(_3538_),
    .B1(net235));
 sg13g2_nor2_1 _8445_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3539_));
 sg13g2_a221oi_1 _8446_ (.B2(_3093_),
    .C1(_3539_),
    .B1(_3538_),
    .A1(net37),
    .Y(_0796_),
    .A2(_3537_));
 sg13g2_buf_1 _8447_ (.A(_3233_),
    .X(_3540_));
 sg13g2_mux2_1 _8448_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ),
    .S(_3536_),
    .X(_3541_));
 sg13g2_mux2_1 _8449_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29] ),
    .A1(_3541_),
    .S(net107),
    .X(_0797_));
 sg13g2_nand2_1 _8450_ (.Y(_3542_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ),
    .B(_3536_));
 sg13g2_o21ai_1 _8451_ (.B1(_3542_),
    .Y(_3543_),
    .A1(_3420_),
    .A2(_3536_));
 sg13g2_mux2_1 _8452_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30] ),
    .A1(_3543_),
    .S(_3535_),
    .X(_0798_));
 sg13g2_a22oi_1 _8453_ (.Y(_3544_),
    .B1(_3538_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ),
    .A2(_3520_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8454_ (.B1(_3544_),
    .Y(_0799_),
    .A1(_3423_),
    .A2(_3536_));
 sg13g2_mux2_1 _8455_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8] ),
    .S(net107),
    .X(_0800_));
 sg13g2_mux2_1 _8456_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9] ),
    .S(net107),
    .X(_0801_));
 sg13g2_mux2_1 _8457_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10] ),
    .S(net107),
    .X(_0802_));
 sg13g2_mux2_1 _8458_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11] ),
    .S(net107),
    .X(_0803_));
 sg13g2_mux2_1 _8459_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8] ),
    .S(_3533_),
    .X(_0804_));
 sg13g2_mux2_1 _8460_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9] ),
    .S(_3533_),
    .X(_0805_));
 sg13g2_mux2_1 _8461_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10] ),
    .S(net109),
    .X(_0806_));
 sg13g2_mux2_1 _8462_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11] ),
    .S(net109),
    .X(_0807_));
 sg13g2_mux2_1 _8463_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12] ),
    .S(net109),
    .X(_0808_));
 sg13g2_mux2_1 _8464_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13] ),
    .S(net109),
    .X(_0809_));
 sg13g2_mux2_1 _8465_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18] ),
    .S(_3535_),
    .X(_0810_));
 sg13g2_buf_1 _8466_ (.A(_3511_),
    .X(_3545_));
 sg13g2_mux2_1 _8467_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19] ),
    .S(net106),
    .X(_0811_));
 sg13g2_mux2_1 _8468_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20] ),
    .S(net106),
    .X(_0812_));
 sg13g2_mux2_1 _8469_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21] ),
    .S(_3545_),
    .X(_0813_));
 sg13g2_mux2_1 _8470_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22] ),
    .S(net106),
    .X(_0814_));
 sg13g2_mux2_1 _8471_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23] ),
    .S(net106),
    .X(_0815_));
 sg13g2_mux2_1 _8472_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24] ),
    .S(net106),
    .X(_0816_));
 sg13g2_mux2_1 _8473_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25] ),
    .S(net106),
    .X(_0817_));
 sg13g2_mux2_1 _8474_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26] ),
    .S(_3545_),
    .X(_0818_));
 sg13g2_mux2_1 _8475_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27] ),
    .S(net106),
    .X(_0819_));
 sg13g2_inv_1 _8476_ (.Y(_3546_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[28] ));
 sg13g2_nand2_1 _8477_ (.Y(_3547_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24] ),
    .B(_3474_));
 sg13g2_o21ai_1 _8478_ (.B1(_3547_),
    .Y(_0820_),
    .A1(_3546_),
    .A2(net154));
 sg13g2_mux2_1 _8479_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29] ),
    .S(net106),
    .X(_0821_));
 sg13g2_buf_1 _8480_ (.A(_3511_),
    .X(_3548_));
 sg13g2_mux2_1 _8481_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30] ),
    .S(net105),
    .X(_0822_));
 sg13g2_mux2_1 _8482_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31] ),
    .S(net105),
    .X(_0823_));
 sg13g2_nand2_2 _8483_ (.Y(_3549_),
    .A(_3302_),
    .B(_3483_));
 sg13g2_nor3_1 _8484_ (.A(net208),
    .B(net48),
    .C(_3549_),
    .Y(_3550_));
 sg13g2_nor2_1 _8485_ (.A(_3306_),
    .B(_3500_),
    .Y(_3551_));
 sg13g2_nor3_1 _8486_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ),
    .B(_3252_),
    .C(_3551_),
    .Y(_3552_));
 sg13g2_a221oi_1 _8487_ (.B2(_3550_),
    .C1(_3552_),
    .B1(net40),
    .A1(_3546_),
    .Y(_0824_),
    .A2(_3105_));
 sg13g2_and2_1 _8488_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ),
    .B(_3549_),
    .X(_3553_));
 sg13g2_a21oi_1 _8489_ (.A1(net46),
    .A2(_3551_),
    .Y(_3554_),
    .B1(_3553_));
 sg13g2_nand2_1 _8490_ (.Y(_3555_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29] ),
    .B(_3474_));
 sg13g2_o21ai_1 _8491_ (.B1(_3555_),
    .Y(_0825_),
    .A1(_3257_),
    .A2(_3554_));
 sg13g2_buf_1 _8492_ (.A(_3237_),
    .X(_3556_));
 sg13g2_nand2_1 _8493_ (.Y(_3557_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ),
    .B(_3549_));
 sg13g2_o21ai_1 _8494_ (.B1(_3557_),
    .Y(_3558_),
    .A1(_3556_),
    .A2(_3549_));
 sg13g2_mux2_1 _8495_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30] ),
    .A1(_3558_),
    .S(net105),
    .X(_0826_));
 sg13g2_buf_8 _8496_ (.A(_3243_),
    .X(_3559_));
 sg13g2_nor2_1 _8497_ (.A(_3248_),
    .B(_3551_),
    .Y(_3560_));
 sg13g2_a22oi_1 _8498_ (.Y(_3561_),
    .B1(_3560_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ),
    .A2(_3520_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8499_ (.B1(_3561_),
    .Y(_0827_),
    .A1(_3559_),
    .A2(_3549_));
 sg13g2_mux2_1 _8500_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8] ),
    .S(net105),
    .X(_0828_));
 sg13g2_mux2_1 _8501_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9] ),
    .S(net105),
    .X(_0829_));
 sg13g2_mux2_1 _8502_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10] ),
    .S(_3548_),
    .X(_0830_));
 sg13g2_mux2_1 _8503_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11] ),
    .S(_3548_),
    .X(_0831_));
 sg13g2_mux2_1 _8504_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8] ),
    .S(net109),
    .X(_0832_));
 sg13g2_mux2_1 _8505_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9] ),
    .S(net109),
    .X(_0833_));
 sg13g2_buf_1 _8506_ (.A(_3451_),
    .X(_3562_));
 sg13g2_mux2_1 _8507_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10] ),
    .S(net104),
    .X(_0834_));
 sg13g2_mux2_1 _8508_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11] ),
    .S(net104),
    .X(_0835_));
 sg13g2_mux2_1 _8509_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12] ),
    .S(_3562_),
    .X(_0836_));
 sg13g2_mux2_1 _8510_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13] ),
    .S(net104),
    .X(_0837_));
 sg13g2_mux2_1 _8511_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18] ),
    .S(net105),
    .X(_0838_));
 sg13g2_mux2_1 _8512_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19] ),
    .S(net105),
    .X(_0839_));
 sg13g2_mux2_1 _8513_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20] ),
    .S(net105),
    .X(_0840_));
 sg13g2_buf_2 _8514_ (.A(_1487_),
    .X(_3563_));
 sg13g2_buf_1 _8515_ (.A(_3563_),
    .X(_3564_));
 sg13g2_mux2_1 _8516_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21] ),
    .S(net203),
    .X(_0841_));
 sg13g2_mux2_1 _8517_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22] ),
    .S(net203),
    .X(_0842_));
 sg13g2_mux2_1 _8518_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23] ),
    .S(_3564_),
    .X(_0843_));
 sg13g2_mux2_1 _8519_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24] ),
    .S(_3564_),
    .X(_0844_));
 sg13g2_mux2_1 _8520_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25] ),
    .S(net203),
    .X(_0845_));
 sg13g2_mux2_1 _8521_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26] ),
    .S(net203),
    .X(_0846_));
 sg13g2_mux2_1 _8522_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27] ),
    .S(net203),
    .X(_0847_));
 sg13g2_mux2_1 _8523_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28] ),
    .S(net203),
    .X(_0848_));
 sg13g2_mux2_1 _8524_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29] ),
    .S(net203),
    .X(_0849_));
 sg13g2_mux2_1 _8525_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30] ),
    .S(net203),
    .X(_0850_));
 sg13g2_buf_1 _8526_ (.A(_3563_),
    .X(_3565_));
 sg13g2_mux2_1 _8527_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31] ),
    .S(net202),
    .X(_0851_));
 sg13g2_buf_1 _8528_ (.A(_3411_),
    .X(_3566_));
 sg13g2_nand2_2 _8529_ (.Y(_3567_),
    .A(_3132_),
    .B(_3566_));
 sg13g2_nor3_1 _8530_ (.A(net208),
    .B(net47),
    .C(_3567_),
    .Y(_3568_));
 sg13g2_a21oi_1 _8531_ (.A1(_3132_),
    .A2(_3566_),
    .Y(_3569_),
    .B1(_3133_));
 sg13g2_nor2_1 _8532_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3570_));
 sg13g2_a221oi_1 _8533_ (.B2(_3096_),
    .C1(_3570_),
    .B1(_3569_),
    .A1(net37),
    .Y(_0852_),
    .A2(_3568_));
 sg13g2_mux2_1 _8534_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1] ),
    .S(_3567_),
    .X(_3571_));
 sg13g2_mux2_1 _8535_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29] ),
    .A1(_3571_),
    .S(net202),
    .X(_0853_));
 sg13g2_nand2_1 _8536_ (.Y(_3572_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ),
    .B(_3567_));
 sg13g2_o21ai_1 _8537_ (.B1(_3572_),
    .Y(_3573_),
    .A1(net41),
    .A2(_3567_));
 sg13g2_mux2_1 _8538_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30] ),
    .A1(_3573_),
    .S(net202),
    .X(_0854_));
 sg13g2_a22oi_1 _8539_ (.Y(_3574_),
    .B1(_3569_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8540_ (.B1(_3574_),
    .Y(_0855_),
    .A1(net35),
    .A2(_3567_));
 sg13g2_mux2_1 _8541_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8] ),
    .S(net202),
    .X(_0856_));
 sg13g2_mux2_1 _8542_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9] ),
    .S(net202),
    .X(_0857_));
 sg13g2_mux2_1 _8543_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10] ),
    .S(_3565_),
    .X(_0858_));
 sg13g2_mux2_1 _8544_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11] ),
    .S(_3565_),
    .X(_0859_));
 sg13g2_mux2_1 _8545_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8] ),
    .S(_3562_),
    .X(_0860_));
 sg13g2_mux2_1 _8546_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9] ),
    .S(net104),
    .X(_0861_));
 sg13g2_mux2_1 _8547_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10] ),
    .S(net104),
    .X(_0862_));
 sg13g2_mux2_1 _8548_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11] ),
    .S(net104),
    .X(_0863_));
 sg13g2_mux2_1 _8549_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12] ),
    .S(net104),
    .X(_0864_));
 sg13g2_mux2_1 _8550_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13] ),
    .S(net104),
    .X(_0865_));
 sg13g2_mux2_1 _8551_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18] ),
    .S(net202),
    .X(_0866_));
 sg13g2_mux2_1 _8552_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19] ),
    .S(net202),
    .X(_0867_));
 sg13g2_mux2_1 _8553_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20] ),
    .S(net202),
    .X(_0868_));
 sg13g2_buf_1 _8554_ (.A(_3563_),
    .X(_3575_));
 sg13g2_mux2_1 _8555_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21] ),
    .S(net201),
    .X(_0869_));
 sg13g2_mux2_1 _8556_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22] ),
    .S(net201),
    .X(_0870_));
 sg13g2_mux2_1 _8557_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23] ),
    .S(net201),
    .X(_0871_));
 sg13g2_mux2_1 _8558_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24] ),
    .S(_3575_),
    .X(_0872_));
 sg13g2_mux2_1 _8559_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25] ),
    .S(net201),
    .X(_0873_));
 sg13g2_mux2_1 _8560_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26] ),
    .S(net201),
    .X(_0874_));
 sg13g2_mux2_1 _8561_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27] ),
    .S(_3575_),
    .X(_0875_));
 sg13g2_mux2_1 _8562_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28] ),
    .S(net201),
    .X(_0876_));
 sg13g2_mux2_1 _8563_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29] ),
    .S(net201),
    .X(_0877_));
 sg13g2_mux2_1 _8564_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30] ),
    .S(net201),
    .X(_0878_));
 sg13g2_buf_1 _8565_ (.A(_3563_),
    .X(_3576_));
 sg13g2_mux2_1 _8566_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31] ),
    .S(net200),
    .X(_0879_));
 sg13g2_nand2_2 _8567_ (.Y(_3577_),
    .A(_3320_),
    .B(_3483_));
 sg13g2_nor3_1 _8568_ (.A(net216),
    .B(_3348_),
    .C(_3577_),
    .Y(_3578_));
 sg13g2_a21oi_1 _8569_ (.A1(_3320_),
    .A2(net272),
    .Y(_3579_),
    .B1(_3133_));
 sg13g2_nor2_1 _8570_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28] ),
    .B(net206),
    .Y(_3580_));
 sg13g2_a221oi_1 _8571_ (.B2(_3099_),
    .C1(_3580_),
    .B1(_3579_),
    .A1(net37),
    .Y(_0880_),
    .A2(_3578_));
 sg13g2_mux2_1 _8572_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ),
    .S(_3577_),
    .X(_3581_));
 sg13g2_mux2_1 _8573_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29] ),
    .A1(_3581_),
    .S(net200),
    .X(_0881_));
 sg13g2_nand2_1 _8574_ (.Y(_3582_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ),
    .B(_3577_));
 sg13g2_o21ai_1 _8575_ (.B1(_3582_),
    .Y(_3583_),
    .A1(net41),
    .A2(_3577_));
 sg13g2_mux2_1 _8576_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30] ),
    .A1(_3583_),
    .S(net200),
    .X(_0882_));
 sg13g2_a22oi_1 _8577_ (.Y(_3584_),
    .B1(_3579_),
    .B2(_2487_),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8578_ (.B1(_3584_),
    .Y(_0883_),
    .A1(net35),
    .A2(_3577_));
 sg13g2_mux2_1 _8579_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8] ),
    .S(net200),
    .X(_0884_));
 sg13g2_mux2_1 _8580_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9] ),
    .S(net200),
    .X(_0885_));
 sg13g2_mux2_1 _8581_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10] ),
    .S(_3576_),
    .X(_0886_));
 sg13g2_mux2_1 _8582_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11] ),
    .S(_3576_),
    .X(_0887_));
 sg13g2_buf_1 _8583_ (.A(_3451_),
    .X(_3585_));
 sg13g2_mux2_1 _8584_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8] ),
    .S(_3585_),
    .X(_0888_));
 sg13g2_mux2_1 _8585_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9] ),
    .S(_3585_),
    .X(_0889_));
 sg13g2_mux2_1 _8586_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10] ),
    .S(net103),
    .X(_0890_));
 sg13g2_mux2_1 _8587_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11] ),
    .S(net103),
    .X(_0891_));
 sg13g2_mux2_1 _8588_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12] ),
    .S(net103),
    .X(_0892_));
 sg13g2_mux2_1 _8589_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13] ),
    .S(net103),
    .X(_0893_));
 sg13g2_mux2_1 _8590_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18] ),
    .S(net200),
    .X(_0894_));
 sg13g2_mux2_1 _8591_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19] ),
    .S(net200),
    .X(_0895_));
 sg13g2_mux2_1 _8592_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20] ),
    .S(net200),
    .X(_0896_));
 sg13g2_buf_1 _8593_ (.A(_3563_),
    .X(_3586_));
 sg13g2_mux2_1 _8594_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21] ),
    .S(net199),
    .X(_0897_));
 sg13g2_mux2_1 _8595_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22] ),
    .S(net199),
    .X(_0898_));
 sg13g2_mux2_1 _8596_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23] ),
    .S(net199),
    .X(_0899_));
 sg13g2_mux2_1 _8597_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24] ),
    .S(net199),
    .X(_0900_));
 sg13g2_mux2_1 _8598_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25] ),
    .S(net199),
    .X(_0901_));
 sg13g2_mux2_1 _8599_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26] ),
    .S(net199),
    .X(_0902_));
 sg13g2_mux2_1 _8600_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27] ),
    .S(_3586_),
    .X(_0903_));
 sg13g2_mux2_1 _8601_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28] ),
    .S(_3586_),
    .X(_0904_));
 sg13g2_mux2_1 _8602_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29] ),
    .S(net199),
    .X(_0905_));
 sg13g2_mux2_1 _8603_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30] ),
    .S(net199),
    .X(_0906_));
 sg13g2_buf_1 _8604_ (.A(_3563_),
    .X(_3587_));
 sg13g2_mux2_1 _8605_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31] ),
    .S(net198),
    .X(_0907_));
 sg13g2_a21oi_1 _8606_ (.A1(_3334_),
    .A2(net272),
    .Y(_3588_),
    .B1(net233));
 sg13g2_nand2_2 _8607_ (.Y(_3589_),
    .A(_3334_),
    .B(_3483_));
 sg13g2_nor3_1 _8608_ (.A(net211),
    .B(net49),
    .C(_3589_),
    .Y(_3590_));
 sg13g2_buf_1 _8609_ (.A(net237),
    .X(_3591_));
 sg13g2_nor2_1 _8610_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3592_));
 sg13g2_a221oi_1 _8611_ (.B2(net38),
    .C1(_3592_),
    .B1(_3590_),
    .A1(_3101_),
    .Y(_0908_),
    .A2(_3588_));
 sg13g2_mux2_1 _8612_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1] ),
    .S(_3589_),
    .X(_3593_));
 sg13g2_mux2_1 _8613_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29] ),
    .A1(_3593_),
    .S(net198),
    .X(_0909_));
 sg13g2_nand2_1 _8614_ (.Y(_3594_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ),
    .B(_3589_));
 sg13g2_o21ai_1 _8615_ (.B1(_3594_),
    .Y(_3595_),
    .A1(net41),
    .A2(_3589_));
 sg13g2_mux2_1 _8616_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30] ),
    .A1(_3595_),
    .S(_3587_),
    .X(_0910_));
 sg13g2_a22oi_1 _8617_ (.Y(_3596_),
    .B1(_3588_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8618_ (.B1(_3596_),
    .Y(_0911_),
    .A1(net35),
    .A2(_3589_));
 sg13g2_mux2_1 _8619_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8] ),
    .S(net198),
    .X(_0912_));
 sg13g2_mux2_1 _8620_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9] ),
    .S(net198),
    .X(_0913_));
 sg13g2_mux2_1 _8621_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10] ),
    .S(net198),
    .X(_0914_));
 sg13g2_mux2_1 _8622_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11] ),
    .S(_3587_),
    .X(_0915_));
 sg13g2_mux2_1 _8623_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8] ),
    .S(net103),
    .X(_0916_));
 sg13g2_mux2_1 _8624_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9] ),
    .S(net103),
    .X(_0917_));
 sg13g2_mux2_1 _8625_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10] ),
    .S(net103),
    .X(_0918_));
 sg13g2_mux2_1 _8626_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11] ),
    .S(net103),
    .X(_0919_));
 sg13g2_buf_1 _8627_ (.A(_3254_),
    .X(_3597_));
 sg13g2_mux2_1 _8628_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12] ),
    .S(net196),
    .X(_0920_));
 sg13g2_mux2_1 _8629_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13] ),
    .S(net196),
    .X(_0921_));
 sg13g2_mux2_1 _8630_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18] ),
    .S(net198),
    .X(_0922_));
 sg13g2_mux2_1 _8631_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19] ),
    .S(net198),
    .X(_0923_));
 sg13g2_mux2_1 _8632_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20] ),
    .S(net198),
    .X(_0924_));
 sg13g2_buf_1 _8633_ (.A(_3563_),
    .X(_3598_));
 sg13g2_mux2_1 _8634_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21] ),
    .S(net195),
    .X(_0925_));
 sg13g2_mux2_1 _8635_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22] ),
    .S(net195),
    .X(_0926_));
 sg13g2_mux2_1 _8636_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23] ),
    .S(net195),
    .X(_0927_));
 sg13g2_mux2_1 _8637_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24] ),
    .S(_3598_),
    .X(_0928_));
 sg13g2_mux2_1 _8638_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25] ),
    .S(net195),
    .X(_0929_));
 sg13g2_mux2_1 _8639_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26] ),
    .S(net195),
    .X(_0930_));
 sg13g2_mux2_1 _8640_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27] ),
    .S(net195),
    .X(_0931_));
 sg13g2_mux2_1 _8641_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28] ),
    .S(_3598_),
    .X(_0932_));
 sg13g2_mux2_1 _8642_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29] ),
    .S(net195),
    .X(_0933_));
 sg13g2_mux2_1 _8643_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30] ),
    .S(net195),
    .X(_0934_));
 sg13g2_buf_1 _8644_ (.A(_1487_),
    .X(_3599_));
 sg13g2_buf_1 _8645_ (.A(_3599_),
    .X(_3600_));
 sg13g2_mux2_1 _8646_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31] ),
    .S(net194),
    .X(_0935_));
 sg13g2_a21oi_1 _8647_ (.A1(_3262_),
    .A2(net271),
    .Y(_3601_),
    .B1(net233));
 sg13g2_nand2_2 _8648_ (.Y(_3602_),
    .A(_3262_),
    .B(net271));
 sg13g2_nor3_1 _8649_ (.A(net211),
    .B(net49),
    .C(_3602_),
    .Y(_3603_));
 sg13g2_nor2_1 _8650_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3604_));
 sg13g2_a221oi_1 _8651_ (.B2(net38),
    .C1(_3604_),
    .B1(_3603_),
    .A1(_3107_),
    .Y(_0936_),
    .A2(_3601_));
 sg13g2_mux2_1 _8652_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ),
    .S(_3602_),
    .X(_3605_));
 sg13g2_mux2_1 _8653_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29] ),
    .A1(_3605_),
    .S(net194),
    .X(_0937_));
 sg13g2_nand2_1 _8654_ (.Y(_3606_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ),
    .B(_3602_));
 sg13g2_o21ai_1 _8655_ (.B1(_3606_),
    .Y(_3607_),
    .A1(net41),
    .A2(_3602_));
 sg13g2_mux2_1 _8656_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30] ),
    .A1(_3607_),
    .S(net194),
    .X(_0938_));
 sg13g2_a22oi_1 _8657_ (.Y(_3608_),
    .B1(_3601_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8658_ (.B1(_3608_),
    .Y(_0939_),
    .A1(net35),
    .A2(_3602_));
 sg13g2_mux2_1 _8659_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8] ),
    .S(net194),
    .X(_0940_));
 sg13g2_mux2_1 _8660_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9] ),
    .S(net194),
    .X(_0941_));
 sg13g2_mux2_1 _8661_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10] ),
    .S(_3600_),
    .X(_0942_));
 sg13g2_mux2_1 _8662_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11] ),
    .S(_3600_),
    .X(_0943_));
 sg13g2_mux2_1 _8663_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8] ),
    .S(net196),
    .X(_0944_));
 sg13g2_mux2_1 _8664_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9] ),
    .S(net196),
    .X(_0945_));
 sg13g2_mux2_1 _8665_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10] ),
    .S(net196),
    .X(_0946_));
 sg13g2_mux2_1 _8666_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11] ),
    .S(_3597_),
    .X(_0947_));
 sg13g2_mux2_1 _8667_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12] ),
    .S(_3597_),
    .X(_0948_));
 sg13g2_mux2_1 _8668_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13] ),
    .S(net196),
    .X(_0949_));
 sg13g2_mux2_1 _8669_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18] ),
    .S(net194),
    .X(_0950_));
 sg13g2_mux2_1 _8670_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19] ),
    .S(net194),
    .X(_0951_));
 sg13g2_mux2_1 _8671_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20] ),
    .S(net194),
    .X(_0952_));
 sg13g2_buf_1 _8672_ (.A(_3599_),
    .X(_3609_));
 sg13g2_mux2_1 _8673_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21] ),
    .S(net193),
    .X(_0953_));
 sg13g2_mux2_1 _8674_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22] ),
    .S(net193),
    .X(_0954_));
 sg13g2_mux2_1 _8675_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23] ),
    .S(net193),
    .X(_0955_));
 sg13g2_mux2_1 _8676_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24] ),
    .S(_3609_),
    .X(_0956_));
 sg13g2_mux2_1 _8677_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25] ),
    .S(net193),
    .X(_0957_));
 sg13g2_mux2_1 _8678_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26] ),
    .S(net193),
    .X(_0958_));
 sg13g2_mux2_1 _8679_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27] ),
    .S(_3609_),
    .X(_0959_));
 sg13g2_mux2_1 _8680_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28] ),
    .S(net193),
    .X(_0960_));
 sg13g2_mux2_1 _8681_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29] ),
    .S(net193),
    .X(_0961_));
 sg13g2_mux2_1 _8682_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30] ),
    .S(net193),
    .X(_0962_));
 sg13g2_buf_1 _8683_ (.A(_3599_),
    .X(_3610_));
 sg13g2_mux2_1 _8684_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31] ),
    .S(net192),
    .X(_0963_));
 sg13g2_nand2_2 _8685_ (.Y(_3611_),
    .A(_3283_),
    .B(net271));
 sg13g2_nor3_1 _8686_ (.A(net216),
    .B(net47),
    .C(_3611_),
    .Y(_3612_));
 sg13g2_a21oi_1 _8687_ (.A1(_3283_),
    .A2(net271),
    .Y(_3613_),
    .B1(net235));
 sg13g2_nor2_1 _8688_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3614_));
 sg13g2_a221oi_1 _8689_ (.B2(_1903_),
    .C1(_3614_),
    .B1(_3613_),
    .A1(net37),
    .Y(_0964_),
    .A2(_3612_));
 sg13g2_mux2_1 _8690_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ),
    .S(_3611_),
    .X(_3615_));
 sg13g2_mux2_1 _8691_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29] ),
    .A1(_3615_),
    .S(net192),
    .X(_0965_));
 sg13g2_nand2_1 _8692_ (.Y(_3616_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ),
    .B(_3611_));
 sg13g2_o21ai_1 _8693_ (.B1(_3616_),
    .Y(_3617_),
    .A1(net41),
    .A2(_3611_));
 sg13g2_mux2_1 _8694_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30] ),
    .A1(_3617_),
    .S(net192),
    .X(_0966_));
 sg13g2_a22oi_1 _8695_ (.Y(_3618_),
    .B1(_3613_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8696_ (.B1(_3618_),
    .Y(_0967_),
    .A1(net35),
    .A2(_3611_));
 sg13g2_mux2_1 _8697_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8] ),
    .S(net192),
    .X(_0968_));
 sg13g2_mux2_1 _8698_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9] ),
    .S(net192),
    .X(_0969_));
 sg13g2_mux2_1 _8699_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10] ),
    .S(_3610_),
    .X(_0970_));
 sg13g2_mux2_1 _8700_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11] ),
    .S(net192),
    .X(_0971_));
 sg13g2_mux2_1 _8701_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8] ),
    .S(net196),
    .X(_0972_));
 sg13g2_mux2_1 _8702_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9] ),
    .S(net196),
    .X(_0973_));
 sg13g2_buf_1 _8703_ (.A(_3254_),
    .X(_3619_));
 sg13g2_mux2_1 _8704_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10] ),
    .S(net191),
    .X(_0974_));
 sg13g2_mux2_1 _8705_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11] ),
    .S(net191),
    .X(_0975_));
 sg13g2_mux2_1 _8706_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12] ),
    .S(net191),
    .X(_0976_));
 sg13g2_mux2_1 _8707_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13] ),
    .S(net191),
    .X(_0977_));
 sg13g2_mux2_1 _8708_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18] ),
    .S(_3610_),
    .X(_0978_));
 sg13g2_mux2_1 _8709_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19] ),
    .S(net192),
    .X(_0979_));
 sg13g2_mux2_1 _8710_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20] ),
    .S(net192),
    .X(_0980_));
 sg13g2_buf_1 _8711_ (.A(_3599_),
    .X(_3620_));
 sg13g2_mux2_1 _8712_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21] ),
    .S(net190),
    .X(_0981_));
 sg13g2_mux2_1 _8713_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22] ),
    .S(net190),
    .X(_0982_));
 sg13g2_mux2_1 _8714_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23] ),
    .S(net190),
    .X(_0983_));
 sg13g2_mux2_1 _8715_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24] ),
    .S(_3620_),
    .X(_0984_));
 sg13g2_mux2_1 _8716_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25] ),
    .S(net190),
    .X(_0985_));
 sg13g2_mux2_1 _8717_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26] ),
    .S(net190),
    .X(_0986_));
 sg13g2_mux2_1 _8718_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27] ),
    .S(net190),
    .X(_0987_));
 sg13g2_mux2_1 _8719_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28] ),
    .S(_3620_),
    .X(_0988_));
 sg13g2_mux2_1 _8720_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29] ),
    .S(net190),
    .X(_0989_));
 sg13g2_mux2_1 _8721_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30] ),
    .S(net190),
    .X(_0990_));
 sg13g2_buf_1 _8722_ (.A(_3599_),
    .X(_3621_));
 sg13g2_mux2_1 _8723_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31] ),
    .S(net189),
    .X(_0991_));
 sg13g2_a21oi_1 _8724_ (.A1(_3302_),
    .A2(net271),
    .Y(_3622_),
    .B1(net233));
 sg13g2_nand2_2 _8725_ (.Y(_3623_),
    .A(_3302_),
    .B(net271));
 sg13g2_nor3_1 _8726_ (.A(net211),
    .B(net49),
    .C(_3623_),
    .Y(_3624_));
 sg13g2_nor2_1 _8727_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3625_));
 sg13g2_a221oi_1 _8728_ (.B2(net38),
    .C1(_3625_),
    .B1(_3624_),
    .A1(_3110_),
    .Y(_0992_),
    .A2(_3622_));
 sg13g2_mux2_1 _8729_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ),
    .S(_3623_),
    .X(_3626_));
 sg13g2_mux2_1 _8730_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29] ),
    .A1(_3626_),
    .S(net189),
    .X(_0993_));
 sg13g2_nand2_1 _8731_ (.Y(_3627_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ),
    .B(_3623_));
 sg13g2_o21ai_1 _8732_ (.B1(_3627_),
    .Y(_3628_),
    .A1(net41),
    .A2(_3623_));
 sg13g2_mux2_1 _8733_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30] ),
    .A1(_3628_),
    .S(net189),
    .X(_0994_));
 sg13g2_a22oi_1 _8734_ (.Y(_3629_),
    .B1(_3622_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ),
    .A2(net204),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8735_ (.B1(_3629_),
    .Y(_0995_),
    .A1(net35),
    .A2(_3623_));
 sg13g2_mux2_1 _8736_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8] ),
    .S(net189),
    .X(_0996_));
 sg13g2_mux2_1 _8737_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9] ),
    .S(net189),
    .X(_0997_));
 sg13g2_mux2_1 _8738_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10] ),
    .S(net189),
    .X(_0998_));
 sg13g2_mux2_1 _8739_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11] ),
    .S(net189),
    .X(_0999_));
 sg13g2_mux2_1 _8740_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8] ),
    .S(net191),
    .X(_1000_));
 sg13g2_mux2_1 _8741_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9] ),
    .S(net191),
    .X(_1001_));
 sg13g2_mux2_1 _8742_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10] ),
    .S(net191),
    .X(_1002_));
 sg13g2_mux2_1 _8743_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11] ),
    .S(net191),
    .X(_1003_));
 sg13g2_mux2_1 _8744_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12] ),
    .S(_3619_),
    .X(_1004_));
 sg13g2_mux2_1 _8745_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13] ),
    .S(_3619_),
    .X(_1005_));
 sg13g2_mux2_1 _8746_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18] ),
    .S(net189),
    .X(_1006_));
 sg13g2_mux2_1 _8747_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19] ),
    .S(_3621_),
    .X(_1007_));
 sg13g2_mux2_1 _8748_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20] ),
    .S(_3621_),
    .X(_1008_));
 sg13g2_buf_1 _8749_ (.A(_3599_),
    .X(_3630_));
 sg13g2_mux2_1 _8750_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21] ),
    .S(net188),
    .X(_1009_));
 sg13g2_mux2_1 _8751_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22] ),
    .S(net188),
    .X(_1010_));
 sg13g2_mux2_1 _8752_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23] ),
    .S(net188),
    .X(_1011_));
 sg13g2_mux2_1 _8753_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24] ),
    .S(_3630_),
    .X(_1012_));
 sg13g2_mux2_1 _8754_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25] ),
    .S(net188),
    .X(_1013_));
 sg13g2_mux2_1 _8755_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26] ),
    .S(net188),
    .X(_1014_));
 sg13g2_mux2_1 _8756_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27] ),
    .S(net188),
    .X(_1015_));
 sg13g2_mux2_1 _8757_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28] ),
    .S(_3630_),
    .X(_1016_));
 sg13g2_mux2_1 _8758_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29] ),
    .S(net188),
    .X(_1017_));
 sg13g2_mux2_1 _8759_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30] ),
    .S(net188),
    .X(_1018_));
 sg13g2_buf_1 _8760_ (.A(_3599_),
    .X(_3631_));
 sg13g2_mux2_1 _8761_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31] ),
    .S(net187),
    .X(_1019_));
 sg13g2_a21oi_1 _8762_ (.A1(_3320_),
    .A2(net271),
    .Y(_3632_),
    .B1(net233));
 sg13g2_nand2_2 _8763_ (.Y(_3633_),
    .A(_3320_),
    .B(_3411_));
 sg13g2_nor3_1 _8764_ (.A(net214),
    .B(net49),
    .C(_3633_),
    .Y(_3634_));
 sg13g2_nor2_1 _8765_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3635_));
 sg13g2_a221oi_1 _8766_ (.B2(net38),
    .C1(_3635_),
    .B1(_3634_),
    .A1(_3112_),
    .Y(_1020_),
    .A2(_3632_));
 sg13g2_mux2_1 _8767_ (.A0(net44),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ),
    .S(_3633_),
    .X(_3636_));
 sg13g2_mux2_1 _8768_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29] ),
    .A1(_3636_),
    .S(net187),
    .X(_1021_));
 sg13g2_nand2_1 _8769_ (.Y(_3637_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ),
    .B(_3633_));
 sg13g2_o21ai_1 _8770_ (.B1(_3637_),
    .Y(_3638_),
    .A1(net41),
    .A2(_3633_));
 sg13g2_mux2_1 _8771_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30] ),
    .A1(_3638_),
    .S(net187),
    .X(_1022_));
 sg13g2_a22oi_1 _8772_ (.Y(_3639_),
    .B1(_3632_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ),
    .A2(net209),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8773_ (.B1(_3639_),
    .Y(_1023_),
    .A1(net35),
    .A2(_3633_));
 sg13g2_mux2_1 _8774_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8] ),
    .S(net187),
    .X(_1024_));
 sg13g2_mux2_1 _8775_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9] ),
    .S(net187),
    .X(_1025_));
 sg13g2_mux2_1 _8776_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10] ),
    .S(net187),
    .X(_1026_));
 sg13g2_mux2_1 _8777_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11] ),
    .S(net187),
    .X(_1027_));
 sg13g2_buf_1 _8778_ (.A(_3254_),
    .X(_3640_));
 sg13g2_mux2_1 _8779_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8] ),
    .S(net186),
    .X(_1028_));
 sg13g2_mux2_1 _8780_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9] ),
    .S(net186),
    .X(_1029_));
 sg13g2_mux2_1 _8781_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10] ),
    .S(net186),
    .X(_1030_));
 sg13g2_mux2_1 _8782_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11] ),
    .S(net186),
    .X(_1031_));
 sg13g2_mux2_1 _8783_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12] ),
    .S(_3640_),
    .X(_1032_));
 sg13g2_mux2_1 _8784_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13] ),
    .S(net186),
    .X(_1033_));
 sg13g2_mux2_1 _8785_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18] ),
    .S(net187),
    .X(_1034_));
 sg13g2_mux2_1 _8786_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19] ),
    .S(_3631_),
    .X(_1035_));
 sg13g2_mux2_1 _8787_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20] ),
    .S(_3631_),
    .X(_1036_));
 sg13g2_buf_1 _8788_ (.A(_3067_),
    .X(_3641_));
 sg13g2_mux2_1 _8789_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21] ),
    .S(net185),
    .X(_1037_));
 sg13g2_mux2_1 _8790_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22] ),
    .S(net185),
    .X(_1038_));
 sg13g2_mux2_1 _8791_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23] ),
    .S(net185),
    .X(_1039_));
 sg13g2_mux2_1 _8792_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24] ),
    .S(net185),
    .X(_1040_));
 sg13g2_mux2_1 _8793_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25] ),
    .S(net185),
    .X(_1041_));
 sg13g2_mux2_1 _8794_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26] ),
    .S(net185),
    .X(_1042_));
 sg13g2_mux2_1 _8795_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27] ),
    .S(net185),
    .X(_1043_));
 sg13g2_mux2_1 _8796_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28] ),
    .S(net185),
    .X(_1044_));
 sg13g2_mux2_1 _8797_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29] ),
    .S(_3641_),
    .X(_1045_));
 sg13g2_mux2_1 _8798_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30] ),
    .S(_3641_),
    .X(_1046_));
 sg13g2_buf_1 _8799_ (.A(_3067_),
    .X(_3642_));
 sg13g2_mux2_1 _8800_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31] ),
    .S(net184),
    .X(_1047_));
 sg13g2_a21oi_1 _8801_ (.A1(_3334_),
    .A2(net271),
    .Y(_3643_),
    .B1(net233));
 sg13g2_nand2_2 _8802_ (.Y(_3644_),
    .A(_3334_),
    .B(_3411_));
 sg13g2_nor3_1 _8803_ (.A(_3224_),
    .B(net48),
    .C(_3644_),
    .Y(_3645_));
 sg13g2_nor2_1 _8804_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28] ),
    .B(_3591_),
    .Y(_3646_));
 sg13g2_a221oi_1 _8805_ (.B2(net38),
    .C1(_3646_),
    .B1(_3645_),
    .A1(_3117_),
    .Y(_1048_),
    .A2(_3643_));
 sg13g2_mux2_1 _8806_ (.A0(_3540_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ),
    .S(_3644_),
    .X(_3647_));
 sg13g2_mux2_1 _8807_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29] ),
    .A1(_3647_),
    .S(net184),
    .X(_1049_));
 sg13g2_nand2_1 _8808_ (.Y(_3648_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ),
    .B(_3644_));
 sg13g2_o21ai_1 _8809_ (.B1(_3648_),
    .Y(_3649_),
    .A1(_3556_),
    .A2(_3644_));
 sg13g2_mux2_1 _8810_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30] ),
    .A1(_3649_),
    .S(net184),
    .X(_1050_));
 sg13g2_a22oi_1 _8811_ (.Y(_3650_),
    .B1(_3643_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ),
    .A2(net209),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8812_ (.B1(_3650_),
    .Y(_1051_),
    .A1(_3559_),
    .A2(_3644_));
 sg13g2_mux2_1 _8813_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8] ),
    .S(net184),
    .X(_1052_));
 sg13g2_mux2_1 _8814_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9] ),
    .S(net184),
    .X(_1053_));
 sg13g2_mux2_1 _8815_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10] ),
    .S(net184),
    .X(_1054_));
 sg13g2_mux2_1 _8816_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11] ),
    .S(net184),
    .X(_1055_));
 sg13g2_mux2_1 _8817_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8] ),
    .S(net186),
    .X(_1056_));
 sg13g2_mux2_1 _8818_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9] ),
    .S(net186),
    .X(_1057_));
 sg13g2_mux2_1 _8819_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10] ),
    .S(_3640_),
    .X(_1058_));
 sg13g2_mux2_1 _8820_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11] ),
    .S(net186),
    .X(_1059_));
 sg13g2_buf_1 _8821_ (.A(_3254_),
    .X(_3651_));
 sg13g2_mux2_1 _8822_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12] ),
    .S(net183),
    .X(_1060_));
 sg13g2_mux2_1 _8823_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13] ),
    .S(net183),
    .X(_1061_));
 sg13g2_mux2_1 _8824_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18] ),
    .S(_3642_),
    .X(_1062_));
 sg13g2_mux2_1 _8825_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19] ),
    .S(net184),
    .X(_1063_));
 sg13g2_mux2_1 _8826_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20] ),
    .S(_3642_),
    .X(_1064_));
 sg13g2_buf_1 _8827_ (.A(_3067_),
    .X(_3652_));
 sg13g2_mux2_1 _8828_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21] ),
    .S(net182),
    .X(_1065_));
 sg13g2_mux2_1 _8829_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22] ),
    .S(_3652_),
    .X(_1066_));
 sg13g2_mux2_1 _8830_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23] ),
    .S(net182),
    .X(_1067_));
 sg13g2_mux2_1 _8831_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24] ),
    .S(net182),
    .X(_1068_));
 sg13g2_mux2_1 _8832_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25] ),
    .S(net182),
    .X(_1069_));
 sg13g2_mux2_1 _8833_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26] ),
    .S(_3652_),
    .X(_1070_));
 sg13g2_mux2_1 _8834_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27] ),
    .S(net182),
    .X(_1071_));
 sg13g2_mux2_1 _8835_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28] ),
    .S(net182),
    .X(_1072_));
 sg13g2_mux2_1 _8836_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29] ),
    .S(net182),
    .X(_1073_));
 sg13g2_mux2_1 _8837_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30] ),
    .S(net182),
    .X(_1074_));
 sg13g2_buf_1 _8838_ (.A(_3067_),
    .X(_3653_));
 sg13g2_mux2_1 _8839_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31] ),
    .S(net181),
    .X(_1075_));
 sg13g2_nand2_2 _8840_ (.Y(_3654_),
    .A(_3126_),
    .B(_3353_));
 sg13g2_nor3_1 _8841_ (.A(_3104_),
    .B(_3228_),
    .C(_3654_),
    .Y(_3655_));
 sg13g2_a21oi_1 _8842_ (.A1(_3127_),
    .A2(_3353_),
    .Y(_3656_),
    .B1(net235));
 sg13g2_nor2_1 _8843_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28] ),
    .B(net197),
    .Y(_3657_));
 sg13g2_a221oi_1 _8844_ (.B2(_3119_),
    .C1(_3657_),
    .B1(_3656_),
    .A1(_3222_),
    .Y(_1076_),
    .A2(_3655_));
 sg13g2_mux2_1 _8845_ (.A0(_3540_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ),
    .S(_3654_),
    .X(_3658_));
 sg13g2_mux2_1 _8846_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29] ),
    .A1(_3658_),
    .S(_3653_),
    .X(_1077_));
 sg13g2_nand2_1 _8847_ (.Y(_3659_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ),
    .B(_3654_));
 sg13g2_o21ai_1 _8848_ (.B1(_3659_),
    .Y(_3660_),
    .A1(net41),
    .A2(_3654_));
 sg13g2_mux2_1 _8849_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30] ),
    .A1(_3660_),
    .S(net181),
    .X(_1078_));
 sg13g2_a22oi_1 _8850_ (.Y(_3661_),
    .B1(_3656_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ),
    .A2(net209),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8851_ (.B1(_3661_),
    .Y(_1079_),
    .A1(net35),
    .A2(_3654_));
 sg13g2_mux2_1 _8852_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8] ),
    .S(net181),
    .X(_1080_));
 sg13g2_mux2_1 _8853_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9] ),
    .S(_3653_),
    .X(_1081_));
 sg13g2_mux2_1 _8854_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10] ),
    .S(net181),
    .X(_1082_));
 sg13g2_mux2_1 _8855_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11] ),
    .S(net181),
    .X(_1083_));
 sg13g2_mux2_1 _8856_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8] ),
    .S(_3651_),
    .X(_1084_));
 sg13g2_mux2_1 _8857_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9] ),
    .S(_3651_),
    .X(_1085_));
 sg13g2_mux2_1 _8858_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10] ),
    .S(net183),
    .X(_1086_));
 sg13g2_mux2_1 _8859_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11] ),
    .S(net183),
    .X(_1087_));
 sg13g2_mux2_1 _8860_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12] ),
    .S(net183),
    .X(_1088_));
 sg13g2_mux2_1 _8861_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13] ),
    .S(net183),
    .X(_1089_));
 sg13g2_mux2_1 _8862_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18] ),
    .S(net181),
    .X(_1090_));
 sg13g2_mux2_1 _8863_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19] ),
    .S(net181),
    .X(_1091_));
 sg13g2_mux2_1 _8864_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20] ),
    .S(net181),
    .X(_1092_));
 sg13g2_buf_1 _8865_ (.A(_3067_),
    .X(_3662_));
 sg13g2_mux2_1 _8866_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21] ),
    .S(net180),
    .X(_1093_));
 sg13g2_mux2_1 _8867_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22] ),
    .S(net180),
    .X(_1094_));
 sg13g2_mux2_1 _8868_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23] ),
    .S(_3662_),
    .X(_1095_));
 sg13g2_mux2_1 _8869_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24] ),
    .S(net180),
    .X(_1096_));
 sg13g2_mux2_1 _8870_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25] ),
    .S(net180),
    .X(_1097_));
 sg13g2_mux2_1 _8871_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26] ),
    .S(net180),
    .X(_1098_));
 sg13g2_mux2_1 _8872_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27] ),
    .S(_3662_),
    .X(_1099_));
 sg13g2_mux2_1 _8873_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28] ),
    .S(net180),
    .X(_1100_));
 sg13g2_mux2_1 _8874_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29] ),
    .S(net180),
    .X(_1101_));
 sg13g2_mux2_1 _8875_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30] ),
    .S(net180),
    .X(_1102_));
 sg13g2_mux2_1 _8876_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31] ),
    .S(net219),
    .X(_1103_));
 sg13g2_a21oi_1 _8877_ (.A1(_3127_),
    .A2(_3367_),
    .Y(_3663_),
    .B1(_3103_));
 sg13g2_nand2_2 _8878_ (.Y(_3664_),
    .A(_3126_),
    .B(_3367_));
 sg13g2_nor3_1 _8879_ (.A(_3224_),
    .B(net48),
    .C(_3664_),
    .Y(_3665_));
 sg13g2_nor2_1 _8880_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28] ),
    .B(_3591_),
    .Y(_3666_));
 sg13g2_a221oi_1 _8881_ (.B2(net38),
    .C1(_3666_),
    .B1(_3665_),
    .A1(_3121_),
    .Y(_1104_),
    .A2(_3663_));
 sg13g2_mux2_1 _8882_ (.A0(_3233_),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ),
    .S(_3664_),
    .X(_3667_));
 sg13g2_mux2_1 _8883_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29] ),
    .A1(_3667_),
    .S(net219),
    .X(_1105_));
 sg13g2_nand2_1 _8884_ (.Y(_3668_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ),
    .B(_3664_));
 sg13g2_o21ai_1 _8885_ (.B1(_3668_),
    .Y(_3669_),
    .A1(_3237_),
    .A2(_3664_));
 sg13g2_mux2_1 _8886_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30] ),
    .A1(_3669_),
    .S(net219),
    .X(_1106_));
 sg13g2_a22oi_1 _8887_ (.Y(_3670_),
    .B1(_3663_),
    .B2(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ),
    .A2(net209),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31] ));
 sg13g2_o21ai_1 _8888_ (.B1(_3670_),
    .Y(_1107_),
    .A1(_3243_),
    .A2(_3664_));
 sg13g2_mux2_1 _8889_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8] ),
    .S(net219),
    .X(_1108_));
 sg13g2_mux2_1 _8890_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9] ),
    .S(net219),
    .X(_1109_));
 sg13g2_mux2_1 _8891_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10] ),
    .S(_3056_),
    .X(_1110_));
 sg13g2_mux2_1 _8892_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11] ),
    .S(_3056_),
    .X(_1111_));
 sg13g2_mux2_1 _8893_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8] ),
    .S(net183),
    .X(_1112_));
 sg13g2_mux2_1 _8894_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13] ),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9] ),
    .S(net183),
    .X(_1113_));
 sg13g2_buf_1 _8895_ (.A(net289),
    .X(_3671_));
 sg13g2_buf_1 _8896_ (.A(net253),
    .X(_3672_));
 sg13g2_nor4_1 _8897_ (.A(_3672_),
    .B(_1485_),
    .C(net290),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3] ),
    .Y(_3673_));
 sg13g2_nand2_1 _8898_ (.Y(_3674_),
    .A(_1504_),
    .B(_3673_));
 sg13g2_nor2_1 _8899_ (.A(_1776_),
    .B(_3674_),
    .Y(_1129_));
 sg13g2_xnor2_1 _8900_ (.Y(_3675_),
    .A(_1474_),
    .B(_1475_));
 sg13g2_nor2_1 _8901_ (.A(_3674_),
    .B(_3675_),
    .Y(_1130_));
 sg13g2_xnor2_1 _8902_ (.Y(_3676_),
    .A(_2651_),
    .B(_1476_));
 sg13g2_nor2_1 _8903_ (.A(_3674_),
    .B(_3676_),
    .Y(_1131_));
 sg13g2_inv_1 _8904_ (.Y(_3677_),
    .A(net307));
 sg13g2_nand2_2 _8905_ (.Y(_3678_),
    .A(_2874_),
    .B(_3677_));
 sg13g2_nor3_1 _8906_ (.A(_2642_),
    .B(_2322_),
    .C(_3678_),
    .Y(_3679_));
 sg13g2_and4_1 _8907_ (.A(_0112_),
    .B(_1465_),
    .C(_2888_),
    .D(_3679_),
    .X(_3680_));
 sg13g2_buf_1 _8908_ (.A(_3680_),
    .X(_3681_));
 sg13g2_buf_1 _8909_ (.A(_3681_),
    .X(_3682_));
 sg13g2_nand2_1 _8910_ (.Y(_3683_),
    .A(_1727_),
    .B(net93));
 sg13g2_nand2b_1 _8911_ (.Y(_3684_),
    .B(net27),
    .A_N(net93));
 sg13g2_buf_1 _8912_ (.A(_3041_),
    .X(_3685_));
 sg13g2_a21oi_1 _8913_ (.A1(_3683_),
    .A2(_3684_),
    .Y(_0116_),
    .B1(net270));
 sg13g2_nand2_1 _8914_ (.Y(_3686_),
    .A(_1724_),
    .B(_3682_));
 sg13g2_nand2b_1 _8915_ (.Y(_3687_),
    .B(net28),
    .A_N(net93));
 sg13g2_a21oi_1 _8916_ (.A1(_3686_),
    .A2(_3687_),
    .Y(_0117_),
    .B1(net270));
 sg13g2_nand2_1 _8917_ (.Y(_3688_),
    .A(_1709_),
    .B(_3682_));
 sg13g2_nand2b_1 _8918_ (.Y(_3689_),
    .B(net29),
    .A_N(net93));
 sg13g2_a21oi_1 _8919_ (.A1(_3688_),
    .A2(_3689_),
    .Y(_0118_),
    .B1(net270));
 sg13g2_nand2_1 _8920_ (.Y(_3690_),
    .A(_2804_),
    .B(net93));
 sg13g2_nand2b_1 _8921_ (.Y(_3691_),
    .B(net30),
    .A_N(net93));
 sg13g2_a21oi_1 _8922_ (.A1(_3690_),
    .A2(_3691_),
    .Y(_0119_),
    .B1(net270));
 sg13g2_nand2_1 _8923_ (.Y(_3692_),
    .A(_2696_),
    .B(net93));
 sg13g2_nand2b_1 _8924_ (.Y(_3693_),
    .B(net31),
    .A_N(_3681_));
 sg13g2_a21oi_1 _8925_ (.A1(_3692_),
    .A2(_3693_),
    .Y(_0120_),
    .B1(_3685_));
 sg13g2_nand2_1 _8926_ (.Y(_3694_),
    .A(_2754_),
    .B(net93));
 sg13g2_nand2b_1 _8927_ (.Y(_3695_),
    .B(net32),
    .A_N(_3681_));
 sg13g2_a21oi_1 _8928_ (.A1(_3694_),
    .A2(_3695_),
    .Y(_0121_),
    .B1(_3685_));
 sg13g2_buf_1 _8929_ (.A(_3041_),
    .X(_3696_));
 sg13g2_buf_1 _8930_ (.A(\i_exotiny.i_wb_qspi_mem.cnt_r[1] ),
    .X(_3697_));
 sg13g2_inv_1 _8931_ (.Y(_3698_),
    .A(_0097_));
 sg13g2_buf_1 _8932_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[28] ),
    .X(_3699_));
 sg13g2_nor2b_1 _8933_ (.A(net318),
    .B_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28] ),
    .Y(_3700_));
 sg13g2_a21o_1 _8934_ (.A2(_3699_),
    .A1(net318),
    .B1(_3700_),
    .X(_3701_));
 sg13g2_buf_2 _8935_ (.A(_3701_),
    .X(_3702_));
 sg13g2_buf_2 _8936_ (.A(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ),
    .X(_3703_));
 sg13g2_nor2_1 _8937_ (.A(_3697_),
    .B(_3703_),
    .Y(_3704_));
 sg13g2_a22oi_1 _8938_ (.Y(_3705_),
    .B1(_3702_),
    .B2(_3704_),
    .A2(_3698_),
    .A1(_3697_));
 sg13g2_buf_2 _8939_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[2] ),
    .X(_3706_));
 sg13g2_buf_1 _8940_ (.A(\i_exotiny.i_wb_qspi_mem.cnt_r[0] ),
    .X(_3707_));
 sg13g2_nand3b_1 _8941_ (.B(_3706_),
    .C(_3707_),
    .Y(_3708_),
    .A_N(_3705_));
 sg13g2_buf_2 _8942_ (.A(_3708_),
    .X(_3709_));
 sg13g2_buf_2 _8943_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[4] ),
    .X(_3710_));
 sg13g2_inv_1 _8944_ (.Y(_3711_),
    .A(_3710_));
 sg13g2_o21ai_1 _8945_ (.B1(_1468_),
    .Y(_3712_),
    .A1(net318),
    .A2(net329));
 sg13g2_buf_1 _8946_ (.A(_3712_),
    .X(_3713_));
 sg13g2_and2_1 _8947_ (.A(net329),
    .B(_2135_),
    .X(_3714_));
 sg13g2_buf_1 _8948_ (.A(_3714_),
    .X(_3715_));
 sg13g2_nor3_1 _8949_ (.A(_3711_),
    .B(_3713_),
    .C(_3715_),
    .Y(_3716_));
 sg13g2_buf_1 _8950_ (.A(_0099_),
    .X(_3717_));
 sg13g2_buf_1 _8951_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[5] ),
    .X(_3718_));
 sg13g2_nor2_1 _8952_ (.A(_3706_),
    .B(net320),
    .Y(_3719_));
 sg13g2_nand2_1 _8953_ (.Y(_3720_),
    .A(_3717_),
    .B(_3719_));
 sg13g2_buf_2 _8954_ (.A(\i_exotiny.i_wb_qspi_mem.crm_r ),
    .X(_3721_));
 sg13g2_inv_1 _8955_ (.Y(_3722_),
    .A(_3721_));
 sg13g2_nor2_1 _8956_ (.A(_3722_),
    .B(_3702_),
    .Y(_3723_));
 sg13g2_nand3_1 _8957_ (.B(_3720_),
    .C(_3723_),
    .A(_3716_),
    .Y(_3724_));
 sg13g2_inv_1 _8958_ (.Y(_3725_),
    .A(_0110_));
 sg13g2_nor2_1 _8959_ (.A(net232),
    .B(_3725_),
    .Y(_3726_));
 sg13g2_a221oi_1 _8960_ (.B2(_3724_),
    .C1(_3726_),
    .B1(_3709_),
    .A1(net232),
    .Y(_3727_),
    .A2(_0109_));
 sg13g2_nand2b_1 _8961_ (.Y(_3728_),
    .B(_3720_),
    .A_N(net320));
 sg13g2_buf_1 _8962_ (.A(_3728_),
    .X(_3729_));
 sg13g2_and2_1 _8963_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ),
    .B(_3729_),
    .X(_3730_));
 sg13g2_and2_1 _8964_ (.A(_3717_),
    .B(_3719_),
    .X(_3731_));
 sg13g2_buf_2 _8965_ (.A(_3731_),
    .X(_3732_));
 sg13g2_nand2b_1 _8966_ (.Y(_3733_),
    .B(_3707_),
    .A_N(_3705_));
 sg13g2_buf_1 _8967_ (.A(_3733_),
    .X(_3734_));
 sg13g2_and2_1 _8968_ (.A(_3706_),
    .B(net99),
    .X(_3735_));
 sg13g2_buf_1 _8969_ (.A(_3735_),
    .X(_3736_));
 sg13g2_and2_1 _8970_ (.A(_3710_),
    .B(net102),
    .X(_3737_));
 sg13g2_buf_1 _8971_ (.A(_3737_),
    .X(_3738_));
 sg13g2_nor2_2 _8972_ (.A(_3736_),
    .B(_3738_),
    .Y(_3739_));
 sg13g2_nor3_1 _8973_ (.A(_0108_),
    .B(_3732_),
    .C(_3739_),
    .Y(_3740_));
 sg13g2_or4_1 _8974_ (.A(net269),
    .B(_3727_),
    .C(_3730_),
    .D(_3740_),
    .X(_1134_));
 sg13g2_buf_1 _8975_ (.A(net326),
    .X(_3741_));
 sg13g2_buf_1 _8976_ (.A(net295),
    .X(_3742_));
 sg13g2_nor3_2 _8977_ (.A(_3702_),
    .B(net102),
    .C(_3715_),
    .Y(_3743_));
 sg13g2_a22oi_1 _8978_ (.Y(_3744_),
    .B1(_3743_),
    .B2(_3722_),
    .A2(net102),
    .A1(_1659_));
 sg13g2_nand2_1 _8979_ (.Y(_3745_),
    .A(_3710_),
    .B(_3720_));
 sg13g2_o21ai_1 _8980_ (.B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ),
    .Y(_3746_),
    .A1(_3729_),
    .A2(_3736_));
 sg13g2_o21ai_1 _8981_ (.B1(_3746_),
    .Y(_3747_),
    .A1(_3744_),
    .A2(_3745_));
 sg13g2_and2_1 _8982_ (.A(net268),
    .B(_3747_),
    .X(_1135_));
 sg13g2_nor2_1 _8983_ (.A(_0111_),
    .B(_3739_),
    .Y(_3748_));
 sg13g2_nand2_1 _8984_ (.Y(_3749_),
    .A(_3710_),
    .B(_3743_));
 sg13g2_nor2b_1 _8985_ (.A(net232),
    .B_N(_0112_),
    .Y(_3750_));
 sg13g2_a221oi_1 _8986_ (.B2(_3749_),
    .C1(_3750_),
    .B1(_3709_),
    .A1(net232),
    .Y(_3751_),
    .A2(_0113_));
 sg13g2_a21oi_1 _8987_ (.A1(_3718_),
    .A2(_1408_),
    .Y(_3752_),
    .B1(_3732_));
 sg13g2_o21ai_1 _8988_ (.B1(_3752_),
    .Y(_3753_),
    .A1(_3721_),
    .A2(_3749_));
 sg13g2_nor3_1 _8989_ (.A(_3748_),
    .B(_3751_),
    .C(_3753_),
    .Y(_3754_));
 sg13g2_buf_1 _8990_ (.A(_3720_),
    .X(_3755_));
 sg13g2_o21ai_1 _8991_ (.B1(net295),
    .Y(_3756_),
    .A1(_1408_),
    .A2(net252));
 sg13g2_nor2_1 _8992_ (.A(_3754_),
    .B(_3756_),
    .Y(_1136_));
 sg13g2_buf_1 _8993_ (.A(net320),
    .X(_3757_));
 sg13g2_a21oi_1 _8994_ (.A1(net294),
    .A2(net9),
    .Y(_3758_),
    .B1(net269));
 sg13g2_nand2b_1 _8995_ (.Y(_3759_),
    .B(_3743_),
    .A_N(_3717_));
 sg13g2_nand3_1 _8996_ (.B(_3758_),
    .C(_3759_),
    .A(_3709_),
    .Y(_1137_));
 sg13g2_nor2b_1 _8997_ (.A(net289),
    .B_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16] ),
    .Y(_3760_));
 sg13g2_a21oi_1 _8998_ (.A1(net289),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16] ),
    .Y(_3761_),
    .B1(_3760_));
 sg13g2_nor3_1 _8999_ (.A(net99),
    .B(_3732_),
    .C(_3761_),
    .Y(_3762_));
 sg13g2_a21oi_1 _9000_ (.A1(_1582_),
    .A2(net99),
    .Y(_3763_),
    .B1(_3762_));
 sg13g2_or2_1 _9001_ (.X(_3764_),
    .B(_3763_),
    .A(_0104_));
 sg13g2_nor2_1 _9002_ (.A(_3713_),
    .B(_3715_),
    .Y(_3765_));
 sg13g2_a21oi_1 _9003_ (.A1(_3723_),
    .A2(_3761_),
    .Y(_3766_),
    .B1(_3732_));
 sg13g2_a22oi_1 _9004_ (.Y(_3767_),
    .B1(_3765_),
    .B2(_3766_),
    .A2(net102),
    .A1(_1582_));
 sg13g2_nor2_1 _9005_ (.A(_3717_),
    .B(_3767_),
    .Y(_3768_));
 sg13g2_a21oi_1 _9006_ (.A1(_1582_),
    .A2(_3729_),
    .Y(_3769_),
    .B1(_3768_));
 sg13g2_a21oi_1 _9007_ (.A1(_3764_),
    .A2(_3769_),
    .Y(_1177_),
    .B1(net270));
 sg13g2_mux2_1 _9008_ (.A0(_0107_),
    .A1(_0106_),
    .S(_3671_),
    .X(_3770_));
 sg13g2_o21ai_1 _9009_ (.B1(_3749_),
    .Y(_3771_),
    .A1(_3709_),
    .A2(_3770_));
 sg13g2_nand2_1 _9010_ (.Y(_3772_),
    .A(_3721_),
    .B(_3770_));
 sg13g2_nor2_1 _9011_ (.A(_0105_),
    .B(_3739_),
    .Y(_3773_));
 sg13g2_a21oi_1 _9012_ (.A1(_3771_),
    .A2(_3772_),
    .Y(_3774_),
    .B1(_3773_));
 sg13g2_a21oi_1 _9013_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1] ),
    .A2(_3729_),
    .Y(_3775_),
    .B1(_3696_));
 sg13g2_o21ai_1 _9014_ (.B1(_3775_),
    .Y(_1178_),
    .A1(_3732_),
    .A2(_3774_));
 sg13g2_inv_1 _9015_ (.Y(_3776_),
    .A(_0115_));
 sg13g2_nand2_1 _9016_ (.Y(_3777_),
    .A(net329),
    .B(_2135_));
 sg13g2_nor3_1 _9017_ (.A(_1389_),
    .B(_3776_),
    .C(_3777_),
    .Y(_3778_));
 sg13g2_nand2_1 _9018_ (.Y(_3779_),
    .A(net307),
    .B(_3778_));
 sg13g2_o21ai_1 _9019_ (.B1(_3709_),
    .Y(_3780_),
    .A1(_3722_),
    .A2(_3749_));
 sg13g2_buf_1 _9020_ (.A(_3780_),
    .X(_3781_));
 sg13g2_nor2b_1 _9021_ (.A(_3779_),
    .B_N(_3781_),
    .Y(_3782_));
 sg13g2_nor2_1 _9022_ (.A(_0114_),
    .B(_3739_),
    .Y(_3783_));
 sg13g2_o21ai_1 _9023_ (.B1(net252),
    .Y(_3784_),
    .A1(_3782_),
    .A2(_3783_));
 sg13g2_a21oi_1 _9024_ (.A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8] ),
    .A2(_3729_),
    .Y(_3785_),
    .B1(net269));
 sg13g2_nand2_1 _9025_ (.Y(_1179_),
    .A(_3784_),
    .B(_3785_));
 sg13g2_buf_1 _9026_ (.A(net269),
    .X(_3786_));
 sg13g2_mux2_1 _9027_ (.A0(_0101_),
    .A1(_0102_),
    .S(net289),
    .X(_3787_));
 sg13g2_a21o_1 _9028_ (.A2(_3787_),
    .A1(_3721_),
    .B1(_3702_),
    .X(_3788_));
 sg13g2_a22oi_1 _9029_ (.Y(_3789_),
    .B1(_3765_),
    .B2(_3788_),
    .A2(net102),
    .A1(_0100_));
 sg13g2_nor2b_1 _9030_ (.A(net99),
    .B_N(_3787_),
    .Y(_3790_));
 sg13g2_a21oi_1 _9031_ (.A1(_0100_),
    .A2(net99),
    .Y(_3791_),
    .B1(_3790_));
 sg13g2_a22oi_1 _9032_ (.Y(_3792_),
    .B1(_3791_),
    .B2(_3706_),
    .A2(_3789_),
    .A1(_3710_));
 sg13g2_inv_1 _9033_ (.Y(_3793_),
    .A(_3792_));
 sg13g2_a22oi_1 _9034_ (.Y(_3794_),
    .B1(_3793_),
    .B2(_3755_),
    .A2(_3729_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0] ));
 sg13g2_nor2_1 _9035_ (.A(net251),
    .B(_3794_),
    .Y(_1180_));
 sg13g2_nand2_1 _9036_ (.Y(_3795_),
    .A(_2090_),
    .B(net205));
 sg13g2_nand2_1 _9037_ (.Y(_3796_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4] ),
    .B(net197));
 sg13g2_a21oi_1 _9038_ (.A1(_3795_),
    .A2(_3796_),
    .Y(_1184_),
    .B1(net270));
 sg13g2_nand2_1 _9039_ (.Y(_3797_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .B(net205));
 sg13g2_nand2_1 _9040_ (.Y(_3798_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5] ),
    .B(net197));
 sg13g2_a21oi_1 _9041_ (.A1(_3797_),
    .A2(_3798_),
    .Y(_1185_),
    .B1(net270));
 sg13g2_nand2_1 _9042_ (.Y(_3799_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i ),
    .B(net205));
 sg13g2_buf_1 _9043_ (.A(net237),
    .X(_3800_));
 sg13g2_nand2_1 _9044_ (.Y(_3801_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6] ),
    .B(_3800_));
 sg13g2_buf_1 _9045_ (.A(_3696_),
    .X(_3802_));
 sg13g2_a21oi_1 _9046_ (.A1(_3799_),
    .A2(_3801_),
    .Y(_1186_),
    .B1(_3802_));
 sg13g2_nand2_1 _9047_ (.Y(_3803_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i ),
    .B(net205));
 sg13g2_nand2_1 _9048_ (.Y(_3804_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7] ),
    .B(net179));
 sg13g2_a21oi_1 _9049_ (.A1(_3803_),
    .A2(_3804_),
    .Y(_1187_),
    .B1(_3802_));
 sg13g2_nand2_1 _9050_ (.Y(_3805_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10] ),
    .B(net205));
 sg13g2_nand2_1 _9051_ (.Y(_3806_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14] ),
    .B(net179));
 sg13g2_a21oi_1 _9052_ (.A1(_3805_),
    .A2(_3806_),
    .Y(_1188_),
    .B1(net250));
 sg13g2_buf_1 _9053_ (.A(_3254_),
    .X(_3807_));
 sg13g2_nand2_1 _9054_ (.Y(_3808_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11] ),
    .B(net178));
 sg13g2_nand2_1 _9055_ (.Y(_3809_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15] ),
    .B(net179));
 sg13g2_a21oi_1 _9056_ (.A1(_3808_),
    .A2(_3809_),
    .Y(_1189_),
    .B1(net250));
 sg13g2_nand2_1 _9057_ (.Y(_3810_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12] ),
    .B(net178));
 sg13g2_nand2_1 _9058_ (.Y(_3811_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16] ),
    .B(net179));
 sg13g2_a21oi_1 _9059_ (.A1(_3810_),
    .A2(_3811_),
    .Y(_1190_),
    .B1(net250));
 sg13g2_nand2_1 _9060_ (.Y(_3812_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13] ),
    .B(net178));
 sg13g2_nand2_1 _9061_ (.Y(_3813_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17] ),
    .B(net179));
 sg13g2_a21oi_1 _9062_ (.A1(_3812_),
    .A2(_3813_),
    .Y(_1191_),
    .B1(net250));
 sg13g2_nand2_1 _9063_ (.Y(_3814_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14] ),
    .B(net178));
 sg13g2_nand2_1 _9064_ (.Y(_3815_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18] ),
    .B(_3800_));
 sg13g2_a21oi_1 _9065_ (.A1(_3814_),
    .A2(_3815_),
    .Y(_1192_),
    .B1(net250));
 sg13g2_nand2_1 _9066_ (.Y(_3816_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15] ),
    .B(net178));
 sg13g2_nand2_1 _9067_ (.Y(_3817_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19] ),
    .B(net179));
 sg13g2_a21oi_1 _9068_ (.A1(_3816_),
    .A2(_3817_),
    .Y(_1193_),
    .B1(net250));
 sg13g2_nand2_1 _9069_ (.Y(_3818_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16] ),
    .B(net178));
 sg13g2_nand2_1 _9070_ (.Y(_3819_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20] ),
    .B(net179));
 sg13g2_a21oi_1 _9071_ (.A1(_3818_),
    .A2(_3819_),
    .Y(_1194_),
    .B1(net250));
 sg13g2_nand2_1 _9072_ (.Y(_3820_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17] ),
    .B(net178));
 sg13g2_nand2_1 _9073_ (.Y(_3821_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21] ),
    .B(net179));
 sg13g2_a21oi_1 _9074_ (.A1(_3820_),
    .A2(_3821_),
    .Y(_1195_),
    .B1(net250));
 sg13g2_nand2_1 _9075_ (.Y(_3822_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18] ),
    .B(_3807_));
 sg13g2_buf_1 _9076_ (.A(net237),
    .X(_3823_));
 sg13g2_nand2_1 _9077_ (.Y(_3824_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22] ),
    .B(net177));
 sg13g2_buf_1 _9078_ (.A(_3041_),
    .X(_3825_));
 sg13g2_a21oi_1 _9079_ (.A1(_3822_),
    .A2(_3824_),
    .Y(_1196_),
    .B1(net267));
 sg13g2_nand2_1 _9080_ (.Y(_3826_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19] ),
    .B(_3807_));
 sg13g2_nand2_1 _9081_ (.Y(_3827_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23] ),
    .B(net177));
 sg13g2_a21oi_1 _9082_ (.A1(_3826_),
    .A2(_3827_),
    .Y(_1197_),
    .B1(net267));
 sg13g2_nand2_1 _9083_ (.Y(_3828_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20] ),
    .B(net178));
 sg13g2_nand2_1 _9084_ (.Y(_3829_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24] ),
    .B(net177));
 sg13g2_a21oi_1 _9085_ (.A1(_3828_),
    .A2(_3829_),
    .Y(_1198_),
    .B1(net267));
 sg13g2_buf_1 _9086_ (.A(net234),
    .X(_3830_));
 sg13g2_nand2_1 _9087_ (.Y(_3831_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21] ),
    .B(net176));
 sg13g2_nand2_1 _9088_ (.Y(_3832_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25] ),
    .B(net177));
 sg13g2_a21oi_1 _9089_ (.A1(_3831_),
    .A2(_3832_),
    .Y(_1199_),
    .B1(_3825_));
 sg13g2_nand2_1 _9090_ (.Y(_3833_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22] ),
    .B(net176));
 sg13g2_nand2_1 _9091_ (.Y(_3834_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26] ),
    .B(net177));
 sg13g2_a21oi_1 _9092_ (.A1(_3833_),
    .A2(_3834_),
    .Y(_1200_),
    .B1(net267));
 sg13g2_nand2_1 _9093_ (.Y(_3835_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23] ),
    .B(net176));
 sg13g2_nand2_1 _9094_ (.Y(_3836_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27] ),
    .B(net177));
 sg13g2_a21oi_1 _9095_ (.A1(_3835_),
    .A2(_3836_),
    .Y(_1201_),
    .B1(net267));
 sg13g2_nand2_1 _9096_ (.Y(_3837_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24] ),
    .B(net176));
 sg13g2_nand2_1 _9097_ (.Y(_3838_),
    .A(_3699_),
    .B(_3823_));
 sg13g2_a21oi_1 _9098_ (.A1(_3837_),
    .A2(_3838_),
    .Y(_1202_),
    .B1(_3825_));
 sg13g2_nand2_1 _9099_ (.Y(_3839_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25] ),
    .B(_3830_));
 sg13g2_nand2_1 _9100_ (.Y(_3840_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ),
    .B(net177));
 sg13g2_a21oi_1 _9101_ (.A1(_3839_),
    .A2(_3840_),
    .Y(_1203_),
    .B1(net267));
 sg13g2_nand2_1 _9102_ (.Y(_3841_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26] ),
    .B(net176));
 sg13g2_nand2_1 _9103_ (.Y(_3842_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30] ),
    .B(net177));
 sg13g2_a21oi_1 _9104_ (.A1(_3841_),
    .A2(_3842_),
    .Y(_1204_),
    .B1(net267));
 sg13g2_nand2_1 _9105_ (.Y(_3843_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27] ),
    .B(net176));
 sg13g2_nand2_1 _9106_ (.Y(_3844_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31] ),
    .B(_3823_));
 sg13g2_a21oi_1 _9107_ (.A1(_3843_),
    .A2(_3844_),
    .Y(_1205_),
    .B1(net267));
 sg13g2_and2_1 _9108_ (.A(_1688_),
    .B(_3214_),
    .X(_3845_));
 sg13g2_nand2_1 _9109_ (.Y(_3846_),
    .A(net277),
    .B(_1521_));
 sg13g2_or4_1 _9110_ (.A(_3205_),
    .B(_3212_),
    .C(_3845_),
    .D(_3846_),
    .X(_3847_));
 sg13g2_buf_1 _9111_ (.A(_3847_),
    .X(_3848_));
 sg13g2_or2_1 _9112_ (.X(_3849_),
    .B(_3846_),
    .A(_3215_));
 sg13g2_inv_1 _9113_ (.Y(_3850_),
    .A(_3849_));
 sg13g2_o21ai_1 _9114_ (.B1(_3850_),
    .Y(_3851_),
    .A1(_3205_),
    .A2(_3212_));
 sg13g2_buf_1 _9115_ (.A(_3851_),
    .X(_3852_));
 sg13g2_a21oi_1 _9116_ (.A1(_3848_),
    .A2(_3852_),
    .Y(_3853_),
    .B1(_2153_));
 sg13g2_nor2_1 _9117_ (.A(_3845_),
    .B(_3846_),
    .Y(_3854_));
 sg13g2_nand2_1 _9118_ (.Y(_3855_),
    .A(_3211_),
    .B(_3854_));
 sg13g2_nand2b_1 _9119_ (.Y(_3856_),
    .B(_3850_),
    .A_N(_3208_));
 sg13g2_a21oi_1 _9120_ (.A1(_3198_),
    .A2(_3202_),
    .Y(_3857_),
    .B1(_3203_));
 sg13g2_mux2_1 _9121_ (.A0(_3855_),
    .A1(_3856_),
    .S(_3857_),
    .X(_3858_));
 sg13g2_xor2_1 _9122_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ),
    .A(_2090_),
    .X(_3859_));
 sg13g2_nor3_1 _9123_ (.A(_3208_),
    .B(_3211_),
    .C(_3849_),
    .Y(_3860_));
 sg13g2_and2_1 _9124_ (.A(_3208_),
    .B(_3854_),
    .X(_3861_));
 sg13g2_nor3_1 _9125_ (.A(_3859_),
    .B(_3860_),
    .C(_3861_),
    .Y(_3862_));
 sg13g2_nand2_1 _9126_ (.Y(_3863_),
    .A(net277),
    .B(_2133_));
 sg13g2_nand4_1 _9127_ (.B(_0040_),
    .C(net237),
    .A(net326),
    .Y(_3864_),
    .D(_3863_));
 sg13g2_a21o_1 _9128_ (.A2(_3862_),
    .A1(_3858_),
    .B1(_3864_),
    .X(_3865_));
 sg13g2_and2_1 _9129_ (.A(net277),
    .B(_2133_),
    .X(_3866_));
 sg13g2_buf_1 _9130_ (.A(_3866_),
    .X(_3867_));
 sg13g2_nor2b_1 _9131_ (.A(_0008_),
    .B_N(_0040_),
    .Y(_3868_));
 sg13g2_a22oi_1 _9132_ (.Y(_3869_),
    .B1(_3867_),
    .B2(_3868_),
    .A2(net234),
    .A1(_3699_));
 sg13g2_nand2b_1 _9133_ (.Y(_3870_),
    .B(net295),
    .A_N(_3869_));
 sg13g2_o21ai_1 _9134_ (.B1(_3870_),
    .Y(_1206_),
    .A1(_3853_),
    .A2(_3865_));
 sg13g2_inv_1 _9135_ (.Y(_3871_),
    .A(_2318_));
 sg13g2_a21oi_1 _9136_ (.A1(_3848_),
    .A2(_3852_),
    .Y(_3872_),
    .B1(_3871_));
 sg13g2_a21o_1 _9137_ (.A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ),
    .A1(_2090_),
    .B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .X(_3873_));
 sg13g2_nand3_1 _9138_ (.B(_2090_),
    .C(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .Y(_3874_));
 sg13g2_a221oi_1 _9139_ (.B2(_3874_),
    .C1(_3860_),
    .B1(_3873_),
    .A1(_3208_),
    .Y(_3875_),
    .A2(_3854_));
 sg13g2_nand3_1 _9140_ (.B(net237),
    .C(_3863_),
    .A(net326),
    .Y(_3876_));
 sg13g2_a21o_1 _9141_ (.A2(_3875_),
    .A1(_3858_),
    .B1(_3876_),
    .X(_3877_));
 sg13g2_a22oi_1 _9142_ (.Y(_3878_),
    .B1(_3867_),
    .B2(_1724_),
    .A2(net234),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ));
 sg13g2_nand2b_1 _9143_ (.Y(_3879_),
    .B(_3741_),
    .A_N(_3878_));
 sg13g2_o21ai_1 _9144_ (.B1(_3879_),
    .Y(_1207_),
    .A1(_3872_),
    .A2(_3877_));
 sg13g2_a21oi_1 _9145_ (.A1(_3848_),
    .A2(_3852_),
    .Y(_3880_),
    .B1(_2468_));
 sg13g2_nand3_1 _9146_ (.B(_2101_),
    .C(_2646_),
    .A(net222),
    .Y(_3881_));
 sg13g2_mux2_1 _9147_ (.A0(_0041_),
    .A1(_2690_),
    .S(_3881_),
    .X(_3882_));
 sg13g2_o21ai_1 _9148_ (.B1(_3874_),
    .Y(_3883_),
    .A1(_0040_),
    .A2(_3882_));
 sg13g2_xnor2_1 _9149_ (.Y(_3884_),
    .A(_0045_),
    .B(_3883_));
 sg13g2_nor3_1 _9150_ (.A(_3860_),
    .B(_3861_),
    .C(_3884_),
    .Y(_3885_));
 sg13g2_a21o_1 _9151_ (.A2(_3885_),
    .A1(_3858_),
    .B1(_3876_),
    .X(_3886_));
 sg13g2_a22oi_1 _9152_ (.Y(_3887_),
    .B1(_3867_),
    .B2(_1709_),
    .A2(net234),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30] ));
 sg13g2_nand2b_1 _9153_ (.Y(_3888_),
    .B(_3741_),
    .A_N(_3887_));
 sg13g2_o21ai_1 _9154_ (.B1(_3888_),
    .Y(_1208_),
    .A1(_3880_),
    .A2(_3886_));
 sg13g2_o21ai_1 _9155_ (.B1(_1503_),
    .Y(_3889_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31] ),
    .A2(_1487_));
 sg13g2_nand2b_1 _9156_ (.Y(_3890_),
    .B(_3863_),
    .A_N(_3889_));
 sg13g2_nand2_1 _9157_ (.Y(_3891_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i ),
    .B(_3883_));
 sg13g2_xnor2_1 _9158_ (.Y(_3892_),
    .A(_2597_),
    .B(_3891_));
 sg13g2_nor2_1 _9159_ (.A(_3890_),
    .B(_3892_),
    .Y(_3893_));
 sg13g2_nand3_1 _9160_ (.B(_3852_),
    .C(_3893_),
    .A(_3848_),
    .Y(_3894_));
 sg13g2_a21o_1 _9161_ (.A2(_2628_),
    .A1(_2625_),
    .B1(_3890_),
    .X(_3895_));
 sg13g2_a21o_1 _9162_ (.A2(_3852_),
    .A1(_3848_),
    .B1(_3895_),
    .X(_3896_));
 sg13g2_a21oi_1 _9163_ (.A1(_2804_),
    .A2(_3867_),
    .Y(_3897_),
    .B1(net236));
 sg13g2_or2_1 _9164_ (.X(_3898_),
    .B(_3897_),
    .A(_3889_));
 sg13g2_nand3_1 _9165_ (.B(_3896_),
    .C(_3898_),
    .A(_3894_),
    .Y(_1209_));
 sg13g2_nand2_1 _9166_ (.Y(_3899_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4] ),
    .B(net176));
 sg13g2_nand2_1 _9167_ (.Y(_3900_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8] ),
    .B(net220));
 sg13g2_buf_1 _9168_ (.A(_3041_),
    .X(_3901_));
 sg13g2_a21oi_1 _9169_ (.A1(_3899_),
    .A2(_3900_),
    .Y(_1210_),
    .B1(net266));
 sg13g2_nand2_1 _9170_ (.Y(_3902_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5] ),
    .B(_3830_));
 sg13g2_nand2_1 _9171_ (.Y(_3903_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9] ),
    .B(net220));
 sg13g2_a21oi_1 _9172_ (.A1(_3902_),
    .A2(_3903_),
    .Y(_1211_),
    .B1(net266));
 sg13g2_nand2_1 _9173_ (.Y(_3904_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6] ),
    .B(net176));
 sg13g2_nand2_1 _9174_ (.Y(_3905_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10] ),
    .B(net220));
 sg13g2_a21oi_1 _9175_ (.A1(_3904_),
    .A2(_3905_),
    .Y(_1212_),
    .B1(net266));
 sg13g2_nand2_1 _9176_ (.Y(_3906_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7] ),
    .B(net213));
 sg13g2_nand2_1 _9177_ (.Y(_3907_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11] ),
    .B(net220));
 sg13g2_a21oi_1 _9178_ (.A1(_3906_),
    .A2(_3907_),
    .Y(_1213_),
    .B1(net266));
 sg13g2_nand2_1 _9179_ (.Y(_3908_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8] ),
    .B(net213));
 sg13g2_nand2_1 _9180_ (.Y(_3909_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12] ),
    .B(net220));
 sg13g2_a21oi_1 _9181_ (.A1(_3908_),
    .A2(_3909_),
    .Y(_1214_),
    .B1(net266));
 sg13g2_nand2_1 _9182_ (.Y(_3910_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9] ),
    .B(net213));
 sg13g2_nand2_1 _9183_ (.Y(_3911_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13] ),
    .B(net220));
 sg13g2_a21oi_1 _9184_ (.A1(_3910_),
    .A2(_3911_),
    .Y(_1215_),
    .B1(net266));
 sg13g2_inv_1 _9185_ (.Y(_3912_),
    .A(_1785_));
 sg13g2_a21oi_1 _9186_ (.A1(_1686_),
    .A2(_3912_),
    .Y(_3913_),
    .B1(_1817_));
 sg13g2_nor2_1 _9187_ (.A(_1714_),
    .B(_3913_),
    .Y(_1282_));
 sg13g2_buf_1 _9188_ (.A(_3707_),
    .X(_3914_));
 sg13g2_buf_1 _9189_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[6] ),
    .X(_3915_));
 sg13g2_buf_1 _9190_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[1] ),
    .X(_3916_));
 sg13g2_nor3_1 _9191_ (.A(_3915_),
    .B(_3916_),
    .C(_3738_),
    .Y(_3917_));
 sg13g2_nor4_1 _9192_ (.A(_3710_),
    .B(_3706_),
    .C(_3915_),
    .D(_3916_),
    .Y(_3918_));
 sg13g2_buf_2 _9193_ (.A(_0098_),
    .X(_3919_));
 sg13g2_o21ai_1 _9194_ (.B1(_3919_),
    .Y(_3920_),
    .A1(_3736_),
    .A2(_3918_));
 sg13g2_o21ai_1 _9195_ (.B1(_3920_),
    .Y(_3921_),
    .A1(net293),
    .A2(_3917_));
 sg13g2_and2_1 _9196_ (.A(net268),
    .B(_3921_),
    .X(_1283_));
 sg13g2_inv_1 _9197_ (.Y(_3922_),
    .A(_3916_));
 sg13g2_nor2b_1 _9198_ (.A(_0097_),
    .B_N(_3707_),
    .Y(_3923_));
 sg13g2_o21ai_1 _9199_ (.B1(_3923_),
    .Y(_3924_),
    .A1(_3697_),
    .A2(_3702_));
 sg13g2_a21oi_1 _9200_ (.A1(_3915_),
    .A2(_3924_),
    .Y(_3925_),
    .B1(_3918_));
 sg13g2_and2_1 _9201_ (.A(_3739_),
    .B(_3925_),
    .X(_3926_));
 sg13g2_or2_1 _9202_ (.X(_3927_),
    .B(net293),
    .A(_3697_));
 sg13g2_nand2_2 _9203_ (.Y(_3928_),
    .A(_3697_),
    .B(net293));
 sg13g2_nand3_1 _9204_ (.B(_3927_),
    .C(_3928_),
    .A(net295),
    .Y(_3929_));
 sg13g2_a21oi_1 _9205_ (.A1(_3922_),
    .A2(_3926_),
    .Y(_1284_),
    .B1(_3929_));
 sg13g2_xor2_1 _9206_ (.B(_3928_),
    .A(_3703_),
    .X(_3930_));
 sg13g2_nand3_1 _9207_ (.B(_3916_),
    .C(_3928_),
    .A(_3698_),
    .Y(_3931_));
 sg13g2_o21ai_1 _9208_ (.B1(_3931_),
    .Y(_3932_),
    .A1(_3926_),
    .A2(_3930_));
 sg13g2_and2_1 _9209_ (.A(net268),
    .B(_3932_),
    .X(_1285_));
 sg13g2_o21ai_1 _9210_ (.B1(_3722_),
    .Y(_3933_),
    .A1(_3702_),
    .A2(_3709_));
 sg13g2_nand2_1 _9211_ (.Y(_3934_),
    .A(net295),
    .B(_3933_));
 sg13g2_inv_1 _9212_ (.Y(_1286_),
    .A(_3934_));
 sg13g2_nand3_1 _9213_ (.B(_2871_),
    .C(_2872_),
    .A(_2809_),
    .Y(_3935_));
 sg13g2_a21o_1 _9214_ (.A2(_2872_),
    .A1(_2871_),
    .B1(_3048_),
    .X(_3936_));
 sg13g2_a21oi_1 _9215_ (.A1(_3935_),
    .A2(_3936_),
    .Y(_1288_),
    .B1(net266));
 sg13g2_nand3_1 _9216_ (.B(_3677_),
    .C(_2872_),
    .A(_2874_),
    .Y(_3937_));
 sg13g2_buf_2 _9217_ (.A(_3937_),
    .X(_3938_));
 sg13g2_nor2_1 _9218_ (.A(_1727_),
    .B(_3938_),
    .Y(_3939_));
 sg13g2_nor2b_1 _9219_ (.A(\i_exotiny.i_wb_regs.spi_presc_o[0] ),
    .B_N(_3938_),
    .Y(_3940_));
 sg13g2_o21ai_1 _9220_ (.B1(net268),
    .Y(_1289_),
    .A1(_3939_),
    .A2(_3940_));
 sg13g2_nor2_1 _9221_ (.A(_1724_),
    .B(_3938_),
    .Y(_3941_));
 sg13g2_nor2b_1 _9222_ (.A(\i_exotiny.i_wb_regs.spi_presc_o[1] ),
    .B_N(_3938_),
    .Y(_3942_));
 sg13g2_o21ai_1 _9223_ (.B1(net268),
    .Y(_1290_),
    .A1(_3941_),
    .A2(_3942_));
 sg13g2_nand2_1 _9224_ (.Y(_3943_),
    .A(\i_exotiny.i_wb_regs.spi_presc_o[2] ),
    .B(_3938_));
 sg13g2_o21ai_1 _9225_ (.B1(_3943_),
    .Y(_3944_),
    .A1(_1715_),
    .A2(_3938_));
 sg13g2_and2_1 _9226_ (.A(net268),
    .B(_3944_),
    .X(_1291_));
 sg13g2_nor2_1 _9227_ (.A(_2804_),
    .B(_3938_),
    .Y(_3945_));
 sg13g2_inv_1 _9228_ (.Y(_3946_),
    .A(\i_exotiny.i_wb_regs.spi_presc_o[3] ));
 sg13g2_and2_1 _9229_ (.A(_3946_),
    .B(_3938_),
    .X(_3947_));
 sg13g2_o21ai_1 _9230_ (.B1(_3742_),
    .Y(_1292_),
    .A1(_3945_),
    .A2(_3947_));
 sg13g2_a21oi_2 _9231_ (.B1(_3700_),
    .Y(_3948_),
    .A2(_3699_),
    .A1(net289));
 sg13g2_inv_1 _9232_ (.Y(_3949_),
    .A(\i_exotiny.i_wb_qspi_mem.state_r_reg[0] ));
 sg13g2_nor3_1 _9233_ (.A(_3949_),
    .B(_1504_),
    .C(_0001_),
    .Y(_3950_));
 sg13g2_a21oi_1 _9234_ (.A1(_0001_),
    .A2(_3948_),
    .Y(_3951_),
    .B1(_3950_));
 sg13g2_nand3_1 _9235_ (.B(_1462_),
    .C(_3951_),
    .A(_3711_),
    .Y(cs_ram_n));
 sg13g2_nand4_1 _9236_ (.B(_3949_),
    .C(_1462_),
    .A(_3711_),
    .Y(cs_rom_n),
    .D(_3948_));
 sg13g2_nor2_1 _9237_ (.A(_3786_),
    .B(net229),
    .Y(\i_exotiny._0000_ ));
 sg13g2_nor2_1 _9238_ (.A(_1477_),
    .B(_1476_),
    .Y(_3952_));
 sg13g2_and2_1 _9239_ (.A(_1443_),
    .B(_3952_),
    .X(_3953_));
 sg13g2_nand3b_1 _9240_ (.B(_2125_),
    .C(_3953_),
    .Y(_3954_),
    .A_N(_2119_));
 sg13g2_nand2_1 _9241_ (.Y(_3955_),
    .A(_2136_),
    .B(_3226_));
 sg13g2_nand3_1 _9242_ (.B(_3952_),
    .C(_2646_),
    .A(_2120_),
    .Y(_3956_));
 sg13g2_a21oi_1 _9243_ (.A1(_3672_),
    .A2(_1462_),
    .Y(_3957_),
    .B1(_3041_));
 sg13g2_nand3_1 _9244_ (.B(net222),
    .C(_1470_),
    .A(net329),
    .Y(_3958_));
 sg13g2_and3_1 _9245_ (.X(_3959_),
    .A(_3956_),
    .B(_3957_),
    .C(_3958_));
 sg13g2_o21ai_1 _9246_ (.B1(_3959_),
    .Y(\i_exotiny._0001_ ),
    .A1(_3954_),
    .A2(_3955_));
 sg13g2_a21oi_1 _9247_ (.A1(_1443_),
    .A2(_1479_),
    .Y(_3960_),
    .B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3] ));
 sg13g2_nor2_1 _9248_ (.A(_3786_),
    .B(_3960_),
    .Y(\i_exotiny._0002_ ));
 sg13g2_a22oi_1 _9249_ (.Y(_3961_),
    .B1(_2135_),
    .B2(net277),
    .A2(net230),
    .A1(_1443_));
 sg13g2_nand2b_1 _9250_ (.Y(_3962_),
    .B(_3952_),
    .A_N(_3961_));
 sg13g2_nand2b_1 _9251_ (.Y(_3963_),
    .B(net329),
    .A_N(_1470_));
 sg13g2_a21oi_1 _9252_ (.A1(_3962_),
    .A2(_3963_),
    .Y(\i_exotiny._0003_ ),
    .B1(_3901_));
 sg13g2_a22oi_1 _9253_ (.Y(_3964_),
    .B1(_3953_),
    .B2(_1461_),
    .A2(_2668_),
    .A1(_1485_));
 sg13g2_nand2b_1 _9254_ (.Y(_3965_),
    .B(net326),
    .A_N(_3964_));
 sg13g2_nor2_1 _9255_ (.A(_1370_),
    .B(net323),
    .Y(_3966_));
 sg13g2_nand4_1 _9256_ (.B(net222),
    .C(_1710_),
    .A(_0110_),
    .Y(_3967_),
    .D(_3966_));
 sg13g2_o21ai_1 _9257_ (.B1(_3967_),
    .Y(_3968_),
    .A1(net222),
    .A2(_3678_));
 sg13g2_nor2_1 _9258_ (.A(net290),
    .B(_3968_),
    .Y(_3969_));
 sg13g2_a21oi_1 _9259_ (.A1(net290),
    .A2(_1472_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[3] ),
    .B1(_3969_));
 sg13g2_nand2_1 _9260_ (.Y(_3970_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[0] ),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[3] ));
 sg13g2_nor2b_1 _9261_ (.A(_3954_),
    .B_N(_3955_),
    .Y(_3971_));
 sg13g2_a21o_1 _9262_ (.A2(_1479_),
    .A1(_2120_),
    .B1(_1473_),
    .X(_3972_));
 sg13g2_o21ai_1 _9263_ (.B1(net295),
    .Y(_3973_),
    .A1(_3971_),
    .A2(_3972_));
 sg13g2_o21ai_1 _9264_ (.B1(_3973_),
    .Y(\i_exotiny._0004_ ),
    .A1(_3965_),
    .A2(_3970_));
 sg13g2_nand2_1 _9265_ (.Y(_3974_),
    .A(net295),
    .B(net290));
 sg13g2_a22oi_1 _9266_ (.Y(\i_exotiny._0005_ ),
    .B1(_3974_),
    .B2(_3965_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[3] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[0] ));
 sg13g2_nor2_1 _9267_ (.A(_0097_),
    .B(_3928_),
    .Y(_3975_));
 sg13g2_o21ai_1 _9268_ (.B1(net268),
    .Y(\i_exotiny._0006_ ),
    .A1(_3949_),
    .A2(_3975_));
 sg13g2_inv_1 _9269_ (.Y(_3976_),
    .A(_3915_));
 sg13g2_nor2_1 _9270_ (.A(_3976_),
    .B(_3924_),
    .Y(_3977_));
 sg13g2_nor2_1 _9271_ (.A(_3703_),
    .B(_3928_),
    .Y(_3978_));
 sg13g2_nor2_1 _9272_ (.A(_3922_),
    .B(_3978_),
    .Y(_3979_));
 sg13g2_a21oi_1 _9273_ (.A1(_3777_),
    .A2(_3977_),
    .Y(_3980_),
    .B1(_3979_));
 sg13g2_nor2_1 _9274_ (.A(net251),
    .B(_3980_),
    .Y(\i_exotiny._0007_ ));
 sg13g2_nand2_1 _9275_ (.Y(_3981_),
    .A(_3706_),
    .B(net99));
 sg13g2_nand2_1 _9276_ (.Y(_3982_),
    .A(_2646_),
    .B(_3723_));
 sg13g2_nand2_1 _9277_ (.Y(_3983_),
    .A(_3721_),
    .B(_3948_));
 sg13g2_a21o_1 _9278_ (.A2(_3983_),
    .A1(net232),
    .B1(net329),
    .X(_3984_));
 sg13g2_nand4_1 _9279_ (.B(_1468_),
    .C(_3982_),
    .A(_3710_),
    .Y(_3985_),
    .D(_3984_));
 sg13g2_a21oi_1 _9280_ (.A1(_3981_),
    .A2(_3985_),
    .Y(\i_exotiny._0008_ ),
    .B1(net266));
 sg13g2_nor2_1 _9281_ (.A(_0115_),
    .B(_3678_),
    .Y(_3986_));
 sg13g2_o21ai_1 _9282_ (.B1(_3703_),
    .Y(_3987_),
    .A1(_1390_),
    .A2(_3986_));
 sg13g2_or3_1 _9283_ (.A(net289),
    .B(_3703_),
    .C(_3986_),
    .X(_3988_));
 sg13g2_nor2_1 _9284_ (.A(net309),
    .B(_2121_),
    .Y(_3989_));
 sg13g2_o21ai_1 _9285_ (.B1(_3989_),
    .Y(_3990_),
    .A1(_2874_),
    .A2(_2870_));
 sg13g2_nand2_1 _9286_ (.Y(_3991_),
    .A(_1500_),
    .B(_1495_));
 sg13g2_nor3_1 _9287_ (.A(_1682_),
    .B(_3776_),
    .C(_3678_),
    .Y(_3992_));
 sg13g2_a21oi_1 _9288_ (.A1(_3776_),
    .A2(_3678_),
    .Y(_3993_),
    .B1(_3992_));
 sg13g2_a21oi_1 _9289_ (.A1(_3991_),
    .A2(_3993_),
    .Y(_3994_),
    .B1(_1389_));
 sg13g2_xnor2_1 _9290_ (.Y(_3995_),
    .A(_0005_),
    .B(_3994_));
 sg13g2_nand2_1 _9291_ (.Y(_3996_),
    .A(_3990_),
    .B(_3995_));
 sg13g2_a21oi_1 _9292_ (.A1(_3987_),
    .A2(_3988_),
    .Y(_3997_),
    .B1(_3996_));
 sg13g2_nor3_1 _9293_ (.A(_3703_),
    .B(_3990_),
    .C(_3995_),
    .Y(_3998_));
 sg13g2_o21ai_1 _9294_ (.B1(net293),
    .Y(_3999_),
    .A1(_3997_),
    .A2(_3998_));
 sg13g2_buf_1 _9295_ (.A(\i_exotiny.i_wb_qspi_mem.state_r_reg[3] ),
    .X(_4000_));
 sg13g2_a22oi_1 _9296_ (.Y(_4001_),
    .B1(_3999_),
    .B2(_4000_),
    .A2(_3977_),
    .A1(_3715_));
 sg13g2_nor2_1 _9297_ (.A(net251),
    .B(_4001_),
    .Y(\i_exotiny._0009_ ));
 sg13g2_a221oi_1 _9298_ (.B2(\i_exotiny.i_wb_qspi_mem.state_r_reg[0] ),
    .C1(_1391_),
    .B1(_3975_),
    .A1(_3710_),
    .Y(_4002_),
    .A2(net102));
 sg13g2_nor2_1 _9299_ (.A(net251),
    .B(_4002_),
    .Y(\i_exotiny._0010_ ));
 sg13g2_inv_1 _9300_ (.Y(_4003_),
    .A(_3975_));
 sg13g2_a22oi_1 _9301_ (.Y(_4004_),
    .B1(_4003_),
    .B2(_3757_),
    .A2(_3978_),
    .A1(_3916_));
 sg13g2_nor2_1 _9302_ (.A(net251),
    .B(_4004_),
    .Y(\i_exotiny._0011_ ));
 sg13g2_buf_1 _9303_ (.A(net76),
    .X(_4005_));
 sg13g2_a21oi_1 _9304_ (.A1(_3915_),
    .A2(_3924_),
    .Y(_4006_),
    .B1(_4005_));
 sg13g2_nor2_1 _9305_ (.A(net251),
    .B(_4006_),
    .Y(\i_exotiny._0012_ ));
 sg13g2_inv_1 _9306_ (.Y(_4007_),
    .A(_3999_));
 sg13g2_a22oi_1 _9307_ (.Y(_4008_),
    .B1(_4007_),
    .B2(_4000_),
    .A2(_3975_),
    .A1(net294));
 sg13g2_nor2_1 _9308_ (.A(net251),
    .B(_4008_),
    .Y(\i_exotiny._0013_ ));
 sg13g2_nand3_1 _9309_ (.B(_2887_),
    .C(_3043_),
    .A(net299),
    .Y(_4009_));
 sg13g2_nand3_1 _9310_ (.B(_2897_),
    .C(_4009_),
    .A(_3742_),
    .Y(\i_exotiny._0014_ ));
 sg13g2_a21o_1 _9311_ (.A2(_3043_),
    .A1(_2887_),
    .B1(net275),
    .X(_4010_));
 sg13g2_a21oi_1 _9312_ (.A1(_2890_),
    .A2(_4010_),
    .Y(\i_exotiny._0015_ ),
    .B1(_3901_));
 sg13g2_nor2_1 _9313_ (.A(_3732_),
    .B(_3738_),
    .Y(_4011_));
 sg13g2_inv_1 _9314_ (.Y(_4012_),
    .A(_4011_));
 sg13g2_o21ai_1 _9315_ (.B1(net326),
    .Y(_4013_),
    .A1(_3736_),
    .A2(_4012_));
 sg13g2_buf_1 _9316_ (.A(_4013_),
    .X(_4014_));
 sg13g2_buf_1 _9317_ (.A(_4014_),
    .X(_4015_));
 sg13g2_buf_1 _9318_ (.A(net289),
    .X(_4016_));
 sg13g2_nand2b_1 _9319_ (.Y(_4017_),
    .B(net249),
    .A_N(_0045_));
 sg13g2_o21ai_1 _9320_ (.B1(_4017_),
    .Y(_4018_),
    .A1(net232),
    .A2(_0088_));
 sg13g2_a22oi_1 _9321_ (.Y(_4019_),
    .B1(net67),
    .B2(_4018_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ),
    .A1(net294));
 sg13g2_nor2_1 _9322_ (.A(_3041_),
    .B(_3732_),
    .Y(_4020_));
 sg13g2_buf_2 _9323_ (.A(_4020_),
    .X(_4021_));
 sg13g2_buf_1 _9324_ (.A(_4021_),
    .X(_4022_));
 sg13g2_nand2b_1 _9325_ (.Y(_4023_),
    .B(net101),
    .A_N(_4019_));
 sg13g2_o21ai_1 _9326_ (.B1(_4023_),
    .Y(\i_exotiny._0062_ ),
    .A1(_0010_),
    .A2(net59));
 sg13g2_nand2b_1 _9327_ (.Y(_4024_),
    .B(net249),
    .A_N(_0051_));
 sg13g2_o21ai_1 _9328_ (.B1(_4024_),
    .Y(_4025_),
    .A1(net232),
    .A2(_0087_));
 sg13g2_a22oi_1 _9329_ (.Y(_4026_),
    .B1(net67),
    .B2(_4025_),
    .A2(_1585_),
    .A1(net294));
 sg13g2_nand2b_1 _9330_ (.Y(_4027_),
    .B(net101),
    .A_N(_4026_));
 sg13g2_o21ai_1 _9331_ (.B1(_4027_),
    .Y(\i_exotiny._0063_ ),
    .A1(_0009_),
    .A2(net59));
 sg13g2_nand2b_1 _9332_ (.Y(_4028_),
    .B(_4016_),
    .A_N(_0085_));
 sg13g2_o21ai_1 _9333_ (.B1(_4028_),
    .Y(_4029_),
    .A1(net232),
    .A2(_0086_));
 sg13g2_a22oi_1 _9334_ (.Y(_4030_),
    .B1(net67),
    .B2(_4029_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ),
    .A1(net294));
 sg13g2_nand2b_1 _9335_ (.Y(_4031_),
    .B(_4022_),
    .A_N(_4030_));
 sg13g2_o21ai_1 _9336_ (.B1(_4031_),
    .Y(\i_exotiny._0064_ ),
    .A1(_0084_),
    .A2(_4015_));
 sg13g2_buf_1 _9337_ (.A(net320),
    .X(_4032_));
 sg13g2_buf_1 _9338_ (.A(net253),
    .X(_4033_));
 sg13g2_nand2b_1 _9339_ (.Y(_4034_),
    .B(net249),
    .A_N(_0083_));
 sg13g2_o21ai_1 _9340_ (.B1(_4034_),
    .Y(_4035_),
    .A1(_4033_),
    .A2(_1775_));
 sg13g2_a22oi_1 _9341_ (.Y(_4036_),
    .B1(net67),
    .B2(_4035_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ),
    .A1(net292));
 sg13g2_nand2b_1 _9342_ (.Y(_4037_),
    .B(net101),
    .A_N(_4036_));
 sg13g2_o21ai_1 _9343_ (.B1(_4037_),
    .Y(\i_exotiny._0065_ ),
    .A1(_0082_),
    .A2(net59));
 sg13g2_nand2b_1 _9344_ (.Y(_4038_),
    .B(net249),
    .A_N(_0081_));
 sg13g2_o21ai_1 _9345_ (.B1(_4038_),
    .Y(_4039_),
    .A1(net231),
    .A2(_0024_));
 sg13g2_a22oi_1 _9346_ (.Y(_4040_),
    .B1(net67),
    .B2(_4039_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ),
    .A1(net292));
 sg13g2_nand2b_1 _9347_ (.Y(_4041_),
    .B(net101),
    .A_N(_4040_));
 sg13g2_o21ai_1 _9348_ (.B1(_4041_),
    .Y(\i_exotiny._0066_ ),
    .A1(_0080_),
    .A2(net59));
 sg13g2_nand2b_1 _9349_ (.Y(_4042_),
    .B(net249),
    .A_N(_0078_));
 sg13g2_o21ai_1 _9350_ (.B1(_4042_),
    .Y(_4043_),
    .A1(net231),
    .A2(_0079_));
 sg13g2_a22oi_1 _9351_ (.Y(_4044_),
    .B1(net67),
    .B2(_4043_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ),
    .A1(_4032_));
 sg13g2_nand2b_1 _9352_ (.Y(_4045_),
    .B(net101),
    .A_N(_4044_));
 sg13g2_o21ai_1 _9353_ (.B1(_4045_),
    .Y(\i_exotiny._0067_ ),
    .A1(_0020_),
    .A2(net59));
 sg13g2_nand2b_1 _9354_ (.Y(_4046_),
    .B(net249),
    .A_N(_0076_));
 sg13g2_o21ai_1 _9355_ (.B1(_4046_),
    .Y(_4047_),
    .A1(_4033_),
    .A2(_0077_));
 sg13g2_a22oi_1 _9356_ (.Y(_4048_),
    .B1(net76),
    .B2(_4047_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ),
    .A1(net292));
 sg13g2_nand2b_1 _9357_ (.Y(_4049_),
    .B(net101),
    .A_N(_4048_));
 sg13g2_o21ai_1 _9358_ (.B1(_4049_),
    .Y(\i_exotiny._0068_ ),
    .A1(_0018_),
    .A2(net59));
 sg13g2_nand2b_1 _9359_ (.Y(_4050_),
    .B(net249),
    .A_N(_0074_));
 sg13g2_o21ai_1 _9360_ (.B1(_4050_),
    .Y(_4051_),
    .A1(net231),
    .A2(_0075_));
 sg13g2_a22oi_1 _9361_ (.Y(_4052_),
    .B1(net76),
    .B2(_4051_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ),
    .A1(net292));
 sg13g2_nand2b_1 _9362_ (.Y(_4053_),
    .B(net101),
    .A_N(_4052_));
 sg13g2_o21ai_1 _9363_ (.B1(_4053_),
    .Y(\i_exotiny._0069_ ),
    .A1(_0016_),
    .A2(net59));
 sg13g2_and3_1 _9364_ (.X(\i_exotiny._0070_ ),
    .A(net294),
    .B(net268),
    .C(net10));
 sg13g2_nand2b_1 _9365_ (.Y(_4054_),
    .B(net253),
    .A_N(_0072_));
 sg13g2_o21ai_1 _9366_ (.B1(_4054_),
    .Y(_4055_),
    .A1(net231),
    .A2(_0073_));
 sg13g2_a22oi_1 _9367_ (.Y(_4056_),
    .B1(net76),
    .B2(_4055_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2] ),
    .A1(_4032_));
 sg13g2_nand2b_1 _9368_ (.Y(_4057_),
    .B(net101),
    .A_N(_4056_));
 sg13g2_o21ai_1 _9369_ (.B1(_4057_),
    .Y(\i_exotiny._0071_ ),
    .A1(_0019_),
    .A2(_4015_));
 sg13g2_nand2b_1 _9370_ (.Y(_4058_),
    .B(net253),
    .A_N(_0070_));
 sg13g2_o21ai_1 _9371_ (.B1(_4058_),
    .Y(_4059_),
    .A1(net231),
    .A2(_0071_));
 sg13g2_a22oi_1 _9372_ (.Y(_4060_),
    .B1(net76),
    .B2(_4059_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3] ),
    .A1(net292));
 sg13g2_nand2b_1 _9373_ (.Y(_4061_),
    .B(_4021_),
    .A_N(_4060_));
 sg13g2_o21ai_1 _9374_ (.B1(_4061_),
    .Y(\i_exotiny._0072_ ),
    .A1(_0017_),
    .A2(net59));
 sg13g2_nand2b_1 _9375_ (.Y(_4062_),
    .B(net253),
    .A_N(_0068_));
 sg13g2_o21ai_1 _9376_ (.B1(_4062_),
    .Y(_4063_),
    .A1(net231),
    .A2(_0069_));
 sg13g2_a22oi_1 _9377_ (.Y(_4064_),
    .B1(net76),
    .B2(_4063_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4] ),
    .A1(net292));
 sg13g2_nand2b_1 _9378_ (.Y(_4065_),
    .B(_4021_),
    .A_N(_4064_));
 sg13g2_o21ai_1 _9379_ (.B1(_4065_),
    .Y(\i_exotiny._0073_ ),
    .A1(_0015_),
    .A2(_4014_));
 sg13g2_nand2_1 _9380_ (.Y(_4066_),
    .A(_3721_),
    .B(_3716_));
 sg13g2_nor2b_1 _9381_ (.A(_3671_),
    .B_N(_0067_),
    .Y(_4067_));
 sg13g2_a221oi_1 _9382_ (.B2(_4066_),
    .C1(_4067_),
    .B1(_3709_),
    .A1(_4016_),
    .Y(_4068_),
    .A2(_0066_));
 sg13g2_a221oi_1 _9383_ (.B2(_3716_),
    .C1(_4068_),
    .B1(_3702_),
    .A1(net320),
    .Y(_4069_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ));
 sg13g2_nand2b_1 _9384_ (.Y(_4070_),
    .B(_4021_),
    .A_N(_4069_));
 sg13g2_o21ai_1 _9385_ (.B1(_4070_),
    .Y(\i_exotiny._0074_ ),
    .A1(_0065_),
    .A2(_4014_));
 sg13g2_nand2b_1 _9386_ (.Y(_4071_),
    .B(net253),
    .A_N(_0063_));
 sg13g2_o21ai_1 _9387_ (.B1(_4071_),
    .Y(_4072_),
    .A1(net231),
    .A2(_0064_));
 sg13g2_a22oi_1 _9388_ (.Y(_4073_),
    .B1(net76),
    .B2(_4072_),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ),
    .A1(net292));
 sg13g2_nand2b_1 _9389_ (.Y(_4074_),
    .B(_4021_),
    .A_N(_4073_));
 sg13g2_o21ai_1 _9390_ (.B1(_4074_),
    .Y(\i_exotiny._0075_ ),
    .A1(_0062_),
    .A2(_4014_));
 sg13g2_mux2_1 _9391_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19] ),
    .S(net318),
    .X(_4075_));
 sg13g2_nor2b_1 _9392_ (.A(net99),
    .B_N(_4075_),
    .Y(_4076_));
 sg13g2_a21oi_1 _9393_ (.A1(_1402_),
    .A2(net99),
    .Y(_4077_),
    .B1(_4076_));
 sg13g2_nand2_1 _9394_ (.Y(_4078_),
    .A(_3721_),
    .B(_4075_));
 sg13g2_a221oi_1 _9395_ (.B2(_4078_),
    .C1(_3711_),
    .B1(_3743_),
    .A1(_0061_),
    .Y(_4079_),
    .A2(net102));
 sg13g2_a21oi_1 _9396_ (.A1(net320),
    .A2(_1402_),
    .Y(_4080_),
    .B1(_4079_));
 sg13g2_o21ai_1 _9397_ (.B1(_4080_),
    .Y(_4081_),
    .A1(_0104_),
    .A2(_4077_));
 sg13g2_nor2_1 _9398_ (.A(_0061_),
    .B(net252),
    .Y(_4082_));
 sg13g2_a21oi_1 _9399_ (.A1(net252),
    .A2(_4081_),
    .Y(_4083_),
    .B1(_4082_));
 sg13g2_nor2_1 _9400_ (.A(net251),
    .B(_4083_),
    .Y(\i_exotiny._0076_ ));
 sg13g2_mux2_1 _9401_ (.A0(_0060_),
    .A1(_0059_),
    .S(net289),
    .X(_4084_));
 sg13g2_or2_1 _9402_ (.X(_4085_),
    .B(_4084_),
    .A(_3983_));
 sg13g2_a221oi_1 _9403_ (.B2(_4085_),
    .C1(_3711_),
    .B1(_3765_),
    .A1(_0058_),
    .Y(_4086_),
    .A2(net102));
 sg13g2_nand2_1 _9404_ (.Y(_4087_),
    .A(_3718_),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1] ));
 sg13g2_o21ai_1 _9405_ (.B1(_4087_),
    .Y(_4088_),
    .A1(_3709_),
    .A2(_4084_));
 sg13g2_o21ai_1 _9406_ (.B1(net252),
    .Y(_4089_),
    .A1(_4086_),
    .A2(_4088_));
 sg13g2_a21o_1 _9407_ (.A2(_3981_),
    .A1(_3755_),
    .B1(_0058_),
    .X(_4090_));
 sg13g2_a21oi_1 _9408_ (.A1(_4089_),
    .A2(_4090_),
    .Y(\i_exotiny._0077_ ),
    .B1(net269));
 sg13g2_a21oi_1 _9409_ (.A1(net294),
    .A2(net11),
    .Y(_4091_),
    .B1(_4005_));
 sg13g2_nor2b_1 _9410_ (.A(_4091_),
    .B_N(_4022_),
    .Y(\i_exotiny._0078_ ));
 sg13g2_nand2b_1 _9411_ (.Y(_4092_),
    .B(net253),
    .A_N(_0056_));
 sg13g2_o21ai_1 _9412_ (.B1(_4092_),
    .Y(_4093_),
    .A1(net231),
    .A2(_0057_));
 sg13g2_a22oi_1 _9413_ (.Y(_4094_),
    .B1(net76),
    .B2(_4093_),
    .A2(_1508_),
    .A1(net292));
 sg13g2_nand2b_1 _9414_ (.Y(_4095_),
    .B(_4021_),
    .A_N(_4094_));
 sg13g2_o21ai_1 _9415_ (.B1(_4095_),
    .Y(\i_exotiny._0079_ ),
    .A1(_0055_),
    .A2(_4014_));
 sg13g2_nand2b_1 _9416_ (.Y(_4096_),
    .B(net253),
    .A_N(_0053_));
 sg13g2_o21ai_1 _9417_ (.B1(_4096_),
    .Y(_4097_),
    .A1(net249),
    .A2(_0054_));
 sg13g2_a22oi_1 _9418_ (.Y(_4098_),
    .B1(_3781_),
    .B2(_4097_),
    .A2(_1509_),
    .A1(net320));
 sg13g2_nand2b_1 _9419_ (.Y(_4099_),
    .B(_4021_),
    .A_N(_4098_));
 sg13g2_o21ai_1 _9420_ (.B1(_4099_),
    .Y(\i_exotiny._0080_ ),
    .A1(_0052_),
    .A2(_4014_));
 sg13g2_and3_1 _9421_ (.X(\i_exotiny._0081_ ),
    .A(_3757_),
    .B(net295),
    .C(net12));
 sg13g2_or2_1 _9422_ (.X(_4100_),
    .B(_4011_),
    .A(_0014_));
 sg13g2_nor2b_1 _9423_ (.A(_3719_),
    .B_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5] ),
    .Y(_4101_));
 sg13g2_o21ai_1 _9424_ (.B1(net252),
    .Y(_4102_),
    .A1(net67),
    .A2(_4101_));
 sg13g2_a21oi_1 _9425_ (.A1(_4100_),
    .A2(_4102_),
    .Y(\i_exotiny._0082_ ),
    .B1(net269));
 sg13g2_or2_1 _9426_ (.X(_4103_),
    .B(_4011_),
    .A(_0013_));
 sg13g2_o21ai_1 _9427_ (.B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6] ),
    .Y(_4104_),
    .A1(net294),
    .A2(_3736_));
 sg13g2_a21oi_1 _9428_ (.A1(_4103_),
    .A2(_4104_),
    .Y(\i_exotiny._0083_ ),
    .B1(net269));
 sg13g2_or2_1 _9429_ (.X(_4105_),
    .B(_4011_),
    .A(_0012_));
 sg13g2_nor2b_1 _9430_ (.A(_3719_),
    .B_N(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7] ),
    .Y(_4106_));
 sg13g2_o21ai_1 _9431_ (.B1(net252),
    .Y(_4107_),
    .A1(net67),
    .A2(_4106_));
 sg13g2_a21oi_1 _9432_ (.A1(_4105_),
    .A2(_4107_),
    .Y(\i_exotiny._0084_ ),
    .B1(net269));
 sg13g2_inv_1 _9433_ (.Y(_4108_),
    .A(_0011_));
 sg13g2_nor2b_1 _9434_ (.A(_3734_),
    .B_N(_3778_),
    .Y(_4109_));
 sg13g2_a22oi_1 _9435_ (.Y(_4110_),
    .B1(_4109_),
    .B2(net327),
    .A2(_3734_),
    .A1(_1502_));
 sg13g2_nand2_1 _9436_ (.Y(_4111_),
    .A(net320),
    .B(_1502_));
 sg13g2_o21ai_1 _9437_ (.B1(_4111_),
    .Y(_4112_),
    .A1(_0104_),
    .A2(_4110_));
 sg13g2_a22oi_1 _9438_ (.Y(_4113_),
    .B1(_4112_),
    .B2(net252),
    .A2(_4012_),
    .A1(_4108_));
 sg13g2_nor2_1 _9439_ (.A(net270),
    .B(_4113_),
    .Y(\i_exotiny._0085_ ));
 sg13g2_nor2_1 _9440_ (.A(_3205_),
    .B(_3212_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.ex_cmp_tmp ));
 sg13g2_nor2_1 _9441_ (.A(_2609_),
    .B(_2614_),
    .Y(_4114_));
 sg13g2_nand2_1 _9442_ (.Y(_4115_),
    .A(_2624_),
    .B(_4114_));
 sg13g2_o21ai_1 _9443_ (.B1(net56),
    .Y(_4116_),
    .A1(_3151_),
    .A2(_4115_));
 sg13g2_o21ai_1 _9444_ (.B1(_2631_),
    .Y(_4117_),
    .A1(_3147_),
    .A2(_4115_));
 sg13g2_o21ai_1 _9445_ (.B1(_4117_),
    .Y(_4118_),
    .A1(_2001_),
    .A2(_4116_));
 sg13g2_nand2_1 _9446_ (.Y(_4119_),
    .A(_1986_),
    .B(_3151_));
 sg13g2_a21oi_1 _9447_ (.A1(_2602_),
    .A2(_2600_),
    .Y(_4120_),
    .B1(net241));
 sg13g2_nor2_1 _9448_ (.A(_1994_),
    .B(net56),
    .Y(_4121_));
 sg13g2_o21ai_1 _9449_ (.B1(_2294_),
    .Y(_4122_),
    .A1(_2632_),
    .A2(_4121_));
 sg13g2_nand2b_1 _9450_ (.Y(_4123_),
    .B(_4122_),
    .A_N(_4120_));
 sg13g2_nand2_1 _9451_ (.Y(_4124_),
    .A(_4115_),
    .B(_4123_));
 sg13g2_o21ai_1 _9452_ (.B1(_4124_),
    .Y(_4125_),
    .A1(net56),
    .A2(_4119_));
 sg13g2_a21o_1 _9453_ (.A2(_4118_),
    .A1(net241),
    .B1(_4125_),
    .X(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.genblk1[3].i_fazyrv_fadd_x.c_o ));
 sg13g2_nor2_1 _9454_ (.A(_0051_),
    .B(_3891_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.c_o ));
 sg13g2_xor2_1 _9455_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ),
    .X(_4126_));
 sg13g2_xor2_1 _9456_ (.B(_1757_),
    .A(_1370_),
    .X(_4127_));
 sg13g2_nand2_1 _9457_ (.Y(_4128_),
    .A(_0024_),
    .B(net174));
 sg13g2_o21ai_1 _9458_ (.B1(_4128_),
    .Y(_4129_),
    .A1(net174),
    .A2(_4127_));
 sg13g2_nor2_1 _9459_ (.A(_0023_),
    .B(net222),
    .Y(_4130_));
 sg13g2_a21oi_1 _9460_ (.A1(_1792_),
    .A2(_4129_),
    .Y(_4131_),
    .B1(_4130_));
 sg13g2_nor2_1 _9461_ (.A(net290),
    .B(_4131_),
    .Y(_4132_));
 sg13g2_a21oi_1 _9462_ (.A1(_1369_),
    .A2(_4126_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[1] ),
    .B1(_4132_));
 sg13g2_o21ai_1 _9463_ (.B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ),
    .Y(_4133_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ));
 sg13g2_nor2b_1 _9464_ (.A(_1471_),
    .B_N(_4133_),
    .Y(_4134_));
 sg13g2_xnor2_1 _9465_ (.Y(_4135_),
    .A(_3725_),
    .B(_3966_));
 sg13g2_nor2_1 _9466_ (.A(net174),
    .B(_4135_),
    .Y(_4136_));
 sg13g2_a221oi_1 _9467_ (.B2(_1751_),
    .C1(_4136_),
    .B1(net174),
    .A1(_1718_),
    .Y(_4137_),
    .A2(_1380_));
 sg13g2_a21oi_1 _9468_ (.A1(_3678_),
    .A2(_3991_),
    .Y(_4138_),
    .B1(_1792_));
 sg13g2_nor3_1 _9469_ (.A(net290),
    .B(_4137_),
    .C(_4138_),
    .Y(_4139_));
 sg13g2_a21oi_1 _9470_ (.A1(_1369_),
    .A2(_4134_),
    .Y(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[2] ),
    .B1(_4139_));
 sg13g2_o21ai_1 _9471_ (.B1(_2881_),
    .Y(_4140_),
    .A1(_2905_),
    .A2(_2833_));
 sg13g2_inv_1 _9472_ (.Y(_4141_),
    .A(_4140_));
 sg13g2_nor3_1 _9473_ (.A(_2905_),
    .B(_2833_),
    .C(_0096_),
    .Y(_4142_));
 sg13g2_nor3_1 _9474_ (.A(net68),
    .B(_4141_),
    .C(_4142_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[0] ));
 sg13g2_xor2_1 _9475_ (.B(_2881_),
    .A(\i_exotiny.i_wb_spi.cnt_presc_r[1] ),
    .X(_4143_));
 sg13g2_nor2_1 _9476_ (.A(_2910_),
    .B(_4143_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[1] ));
 sg13g2_o21ai_1 _9477_ (.B1(\i_exotiny.i_wb_spi.cnt_presc_r[2] ),
    .Y(_4144_),
    .A1(\i_exotiny.i_wb_spi.cnt_presc_r[1] ),
    .A2(_2881_));
 sg13g2_nor2b_1 _9478_ (.A(_2882_),
    .B_N(_4144_),
    .Y(_4145_));
 sg13g2_nor2_1 _9479_ (.A(_2910_),
    .B(_4145_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[2] ));
 sg13g2_nor2b_1 _9480_ (.A(_2882_),
    .B_N(\i_exotiny.i_wb_spi.cnt_presc_r[3] ),
    .Y(_4146_));
 sg13g2_o21ai_1 _9481_ (.B1(net68),
    .Y(_4147_),
    .A1(net275),
    .A2(_0095_));
 sg13g2_o21ai_1 _9482_ (.B1(_4147_),
    .Y(_4148_),
    .A1(_2883_),
    .A2(_4146_));
 sg13g2_o21ai_1 _9483_ (.B1(_4148_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[3] ),
    .A1(_0095_),
    .A2(_2890_));
 sg13g2_nor2b_1 _9484_ (.A(_2883_),
    .B_N(\i_exotiny.i_wb_spi.cnt_presc_r[4] ),
    .Y(_4149_));
 sg13g2_o21ai_1 _9485_ (.B1(net68),
    .Y(_4150_),
    .A1(net275),
    .A2(_0094_));
 sg13g2_o21ai_1 _9486_ (.B1(_4150_),
    .Y(_4151_),
    .A1(_2884_),
    .A2(_4149_));
 sg13g2_o21ai_1 _9487_ (.B1(_4151_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[4] ),
    .A1(_0094_),
    .A2(_2890_));
 sg13g2_nor2b_1 _9488_ (.A(_2884_),
    .B_N(\i_exotiny.i_wb_spi.cnt_presc_r[5] ),
    .Y(_4152_));
 sg13g2_o21ai_1 _9489_ (.B1(net68),
    .Y(_4153_),
    .A1(_2880_),
    .A2(_0093_));
 sg13g2_o21ai_1 _9490_ (.B1(_4153_),
    .Y(_4154_),
    .A1(_2885_),
    .A2(_4152_));
 sg13g2_o21ai_1 _9491_ (.B1(_4154_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[5] ),
    .A1(_0093_),
    .A2(_2890_));
 sg13g2_nor2b_1 _9492_ (.A(_2885_),
    .B_N(\i_exotiny.i_wb_spi.cnt_presc_r[6] ),
    .Y(_4155_));
 sg13g2_nor2_1 _9493_ (.A(\i_exotiny.i_wb_regs.spi_presc_o[3] ),
    .B(_4155_),
    .Y(_4156_));
 sg13g2_o21ai_1 _9494_ (.B1(_2893_),
    .Y(_4157_),
    .A1(_0092_),
    .A2(_4156_));
 sg13g2_o21ai_1 _9495_ (.B1(_4157_),
    .Y(_4158_),
    .A1(_2887_),
    .A2(_4155_));
 sg13g2_o21ai_1 _9496_ (.B1(_4158_),
    .Y(\i_exotiny.i_wb_spi.cnt_presc_n[6] ),
    .A1(_3946_),
    .A2(_2890_));
 sg13g2_buf_4 clkbuf_leaf_0_clk (.X(clknet_leaf_0_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_1 _9498_ (.A(_4000_),
    .X(_4159_));
 sg13g2_nor3_1 _9499_ (.A(_3949_),
    .B(_3041_),
    .C(_0001_),
    .Y(_4160_));
 sg13g2_or4_1 _9500_ (.A(_3706_),
    .B(_3915_),
    .C(net291),
    .D(_4160_),
    .X(net14));
 sg13g2_nor2b_1 _9501_ (.A(_3706_),
    .B_N(_0001_),
    .Y(_4161_));
 sg13g2_nor3_1 _9502_ (.A(_0104_),
    .B(_3948_),
    .C(_4161_),
    .Y(_4162_));
 sg13g2_or3_1 _9503_ (.A(_3915_),
    .B(net291),
    .C(_4162_),
    .X(net18));
 sg13g2_xnor2_1 _9504_ (.Y(_4163_),
    .A(_0005_),
    .B(_3779_));
 sg13g2_nand2_1 _9505_ (.Y(_4164_),
    .A(_3697_),
    .B(net307));
 sg13g2_xnor2_1 _9506_ (.Y(_4165_),
    .A(net327),
    .B(_4164_));
 sg13g2_nand2_1 _9507_ (.Y(_4166_),
    .A(_3778_),
    .B(_4165_));
 sg13g2_xor2_1 _9508_ (.B(_4166_),
    .A(_3703_),
    .X(_4167_));
 sg13g2_buf_1 _9509_ (.A(_4167_),
    .X(_4168_));
 sg13g2_nand2_1 _9510_ (.Y(_4169_),
    .A(_4163_),
    .B(net81));
 sg13g2_xor2_1 _9511_ (.B(_3779_),
    .A(_0005_),
    .X(_4170_));
 sg13g2_buf_4 _9512_ (.X(_4171_),
    .A(_4170_));
 sg13g2_mux2_1 _9513_ (.A0(_2716_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ),
    .S(_4171_),
    .X(_4172_));
 sg13g2_nand2b_1 _9514_ (.Y(_4173_),
    .B(_4172_),
    .A_N(net81));
 sg13g2_o21ai_1 _9515_ (.B1(_4173_),
    .Y(_4174_),
    .A1(_0008_),
    .A2(_4169_));
 sg13g2_and2_1 _9516_ (.A(net293),
    .B(_4168_),
    .X(_4175_));
 sg13g2_mux2_1 _9517_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ),
    .S(net81),
    .X(_4176_));
 sg13g2_a22oi_1 _9518_ (.Y(_4177_),
    .B1(_4176_),
    .B2(_3919_),
    .A2(_4175_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ));
 sg13g2_a21oi_2 _9519_ (.B1(net293),
    .Y(_4178_),
    .A2(_4169_),
    .A1(_3919_));
 sg13g2_nor2_1 _9520_ (.A(_4171_),
    .B(_4167_),
    .Y(_4179_));
 sg13g2_and2_1 _9521_ (.A(_3919_),
    .B(_4179_),
    .X(_4180_));
 sg13g2_a22oi_1 _9522_ (.Y(_4181_),
    .B1(_4180_),
    .B2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ),
    .A2(_4178_),
    .A1(_2696_));
 sg13g2_o21ai_1 _9523_ (.B1(_4181_),
    .Y(_4182_),
    .A1(_4163_),
    .A2(_4177_));
 sg13g2_a21oi_1 _9524_ (.A1(net293),
    .A2(_4174_),
    .Y(_4183_),
    .B1(_4182_));
 sg13g2_nor2_1 _9525_ (.A(_1512_),
    .B(net291),
    .Y(_4184_));
 sg13g2_a21oi_1 _9526_ (.A1(net291),
    .A2(_4183_),
    .Y(net21),
    .B1(_4184_));
 sg13g2_inv_1 _9527_ (.Y(_4185_),
    .A(_0007_));
 sg13g2_mux4_1 _9528_ (.S0(_4171_),
    .A0(_2727_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ),
    .A2(_4185_),
    .A3(_2809_),
    .S1(_4168_),
    .X(_4186_));
 sg13g2_mux2_1 _9529_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ),
    .S(net81),
    .X(_4187_));
 sg13g2_a22oi_1 _9530_ (.Y(_4188_),
    .B1(_4187_),
    .B2(_4171_),
    .A2(_4179_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ));
 sg13g2_nor2b_1 _9531_ (.A(_4188_),
    .B_N(_3919_),
    .Y(_4189_));
 sg13g2_a221oi_1 _9532_ (.B2(net293),
    .C1(_4189_),
    .B1(_4186_),
    .A1(_2754_),
    .Y(_4190_),
    .A2(_4178_));
 sg13g2_nor2_1 _9533_ (.A(_1514_),
    .B(net291),
    .Y(_4191_));
 sg13g2_a21oi_1 _9534_ (.A1(_4159_),
    .A2(_4190_),
    .Y(net22),
    .B1(_4191_));
 sg13g2_mux4_1 _9535_ (.S0(_4171_),
    .A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ),
    .A2(_1796_),
    .A3(_2710_),
    .S1(net81),
    .X(_4192_));
 sg13g2_mux2_1 _9536_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ),
    .S(net81),
    .X(_4193_));
 sg13g2_a22oi_1 _9537_ (.Y(_4194_),
    .B1(_4193_),
    .B2(_4171_),
    .A2(_4179_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ));
 sg13g2_nor2b_1 _9538_ (.A(_4194_),
    .B_N(_3919_),
    .Y(_4195_));
 sg13g2_a221oi_1 _9539_ (.B2(_3914_),
    .C1(_4195_),
    .B1(_4192_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ),
    .Y(_4196_),
    .A2(_4178_));
 sg13g2_nor2_1 _9540_ (.A(net325),
    .B(net291),
    .Y(_4197_));
 sg13g2_a21oi_1 _9541_ (.A1(_4159_),
    .A2(_4196_),
    .Y(net24),
    .B1(_4197_));
 sg13g2_mux2_1 _9542_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ),
    .S(_4171_),
    .X(_4198_));
 sg13g2_nand2b_1 _9543_ (.Y(_4199_),
    .B(_4198_),
    .A_N(net81));
 sg13g2_o21ai_1 _9544_ (.B1(_4199_),
    .Y(_4200_),
    .A1(_0004_),
    .A2(_4169_));
 sg13g2_mux2_1 _9545_ (.A0(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ),
    .S(net81),
    .X(_4201_));
 sg13g2_a22oi_1 _9546_ (.Y(_4202_),
    .B1(_4201_),
    .B2(_3919_),
    .A2(_4175_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ));
 sg13g2_a22oi_1 _9547_ (.Y(_4203_),
    .B1(_4180_),
    .B2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ),
    .A2(_4178_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ));
 sg13g2_o21ai_1 _9548_ (.B1(_4203_),
    .Y(_4204_),
    .A1(_4163_),
    .A2(_4202_));
 sg13g2_a21oi_1 _9549_ (.A1(_3914_),
    .A2(_4200_),
    .Y(_4205_),
    .B1(_4204_));
 sg13g2_nor2_1 _9550_ (.A(_1386_),
    .B(net291),
    .Y(_4206_));
 sg13g2_a21oi_1 _9551_ (.A1(net291),
    .A2(_4205_),
    .Y(net25),
    .B1(_4206_));
 sg13g2_inv_1 _9497__1 (.Y(net1646),
    .A(clknet_leaf_34_clk));
 sg13g2_tiehi \i_exotiny.gpo_o[0]$_SDFFE_PN0P__340  (.L_HI(net340));
 sg13g2_buf_1 _9554_ (.A(ena),
    .X(net13));
 sg13g2_buf_1 _9555_ (.A(net18),
    .X(net15));
 sg13g2_buf_1 _9556_ (.A(ena),
    .X(net16));
 sg13g2_buf_1 _9557_ (.A(net18),
    .X(net17));
 sg13g2_buf_1 _9558_ (.A(ena),
    .X(net19));
 sg13g2_buf_1 _9559_ (.A(net338),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9560_ (.A(cs_rom_n),
    .X(net20));
 sg13g2_buf_1 _9561_ (.A(net1646),
    .X(net23));
 sg13g2_buf_1 _9562_ (.A(cs_ram_n),
    .X(net26));
 sg13g2_buf_1 _9563_ (.A(net339),
    .X(uio_out[7]));
 sg13g2_buf_1 _9564_ (.A(\i_exotiny.spi_sck_o ),
    .X(net33));
 sg13g2_buf_1 _9565_ (.A(\i_exotiny.spi_sdo_o ),
    .X(net34));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net340),
    .D(_0116_),
    .Q_N(_5373_),
    .Q(net27));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net341),
    .D(_0117_),
    .Q_N(_5372_),
    .Q(net28));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net342),
    .D(_0118_),
    .Q_N(_5371_),
    .Q(net29));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net343),
    .D(_0119_),
    .Q_N(_5370_),
    .Q(net30));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net344),
    .D(_0120_),
    .Q_N(_5369_),
    .Q(net31));
 sg13g2_dfrbp_1 \i_exotiny.gpo_o[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net345),
    .D(_0121_),
    .Q_N(_5368_),
    .Q(net32));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net346),
    .D(_0122_),
    .Q_N(_5367_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net347),
    .D(_0123_),
    .Q_N(_5366_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net348),
    .D(_0124_),
    .Q_N(_5365_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net349),
    .D(_0125_),
    .Q_N(_5364_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net350),
    .D(_0126_),
    .Q_N(_5363_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net351),
    .D(_0127_),
    .Q_N(_5362_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net352),
    .D(_0128_),
    .Q_N(_5361_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net353),
    .D(_0129_),
    .Q_N(_5360_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net354),
    .D(_0130_),
    .Q_N(_5359_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net355),
    .D(_0131_),
    .Q_N(_5358_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net356),
    .D(_0132_),
    .Q_N(_5357_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net357),
    .D(_0133_),
    .Q_N(_5356_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net358),
    .D(_0134_),
    .Q_N(_5355_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net359),
    .D(_0135_),
    .Q_N(_5354_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net360),
    .D(_0136_),
    .Q_N(_5353_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net361),
    .D(_0137_),
    .Q_N(_5352_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net362),
    .D(_0138_),
    .Q_N(_5351_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net363),
    .D(_0139_),
    .Q_N(_5350_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net364),
    .D(_0140_),
    .Q_N(_5349_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net365),
    .D(_0141_),
    .Q_N(_5348_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net366),
    .D(_0142_),
    .Q_N(_5347_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net367),
    .D(_0143_),
    .Q_N(_5346_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net368),
    .D(_0144_),
    .Q_N(_5345_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net369),
    .D(_0145_),
    .Q_N(_5344_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net370),
    .D(_0146_),
    .Q_N(_5343_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net371),
    .D(_0147_),
    .Q_N(_5342_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net372),
    .D(_0148_),
    .Q_N(_5341_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net373),
    .D(_0149_),
    .Q_N(_5340_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net374),
    .D(_0150_),
    .Q_N(_5339_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net375),
    .D(_0151_),
    .Q_N(_5338_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net376),
    .D(_0152_),
    .Q_N(_5337_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net377),
    .D(_0153_),
    .Q_N(_5336_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net378),
    .D(_0154_),
    .Q_N(_5335_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net379),
    .D(_0155_),
    .Q_N(_5334_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net380),
    .D(_0156_),
    .Q_N(_5333_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net381),
    .D(_0157_),
    .Q_N(_5332_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net382),
    .D(_0158_),
    .Q_N(_5331_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net383),
    .D(_0159_),
    .Q_N(_5330_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net384),
    .D(_0160_),
    .Q_N(_5329_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net385),
    .D(_0161_),
    .Q_N(_5328_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net386),
    .D(_0162_),
    .Q_N(_5327_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net387),
    .D(_0163_),
    .Q_N(_5326_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net388),
    .D(_0164_),
    .Q_N(_5325_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net389),
    .D(_0165_),
    .Q_N(_5324_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net390),
    .D(_0166_),
    .Q_N(_5323_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net391),
    .D(_0167_),
    .Q_N(_5322_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net392),
    .D(_0168_),
    .Q_N(_5321_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net393),
    .D(_0169_),
    .Q_N(_5320_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net394),
    .D(_0170_),
    .Q_N(_5319_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net395),
    .D(_0171_),
    .Q_N(_5318_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net396),
    .D(_0172_),
    .Q_N(_5317_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net397),
    .D(_0173_),
    .Q_N(_5316_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net398),
    .D(_0174_),
    .Q_N(_5315_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net399),
    .D(_0175_),
    .Q_N(_5314_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net400),
    .D(_0176_),
    .Q_N(_5313_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net401),
    .D(_0177_),
    .Q_N(_5312_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net402),
    .D(_0178_),
    .Q_N(_5311_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net403),
    .D(_0179_),
    .Q_N(_5310_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net404),
    .D(_0180_),
    .Q_N(_5309_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net405),
    .D(_0181_),
    .Q_N(_5308_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net406),
    .D(_0182_),
    .Q_N(_5307_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net407),
    .D(_0183_),
    .Q_N(_5306_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net408),
    .D(_0184_),
    .Q_N(_5305_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net409),
    .D(_0185_),
    .Q_N(_5304_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net410),
    .D(_0186_),
    .Q_N(_5303_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net411),
    .D(_0187_),
    .Q_N(_5302_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net412),
    .D(_0188_),
    .Q_N(_5301_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net413),
    .D(_0189_),
    .Q_N(_5300_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net414),
    .D(_0190_),
    .Q_N(_5299_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net415),
    .D(_0191_),
    .Q_N(_5298_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net416),
    .D(_0192_),
    .Q_N(_5297_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net417),
    .D(_0193_),
    .Q_N(_5296_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net418),
    .D(_0194_),
    .Q_N(_5295_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net419),
    .D(_0195_),
    .Q_N(_5294_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net420),
    .D(_0196_),
    .Q_N(_5293_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net421),
    .D(_0197_),
    .Q_N(_5292_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net422),
    .D(_0198_),
    .Q_N(_5291_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net423),
    .D(_0199_),
    .Q_N(_5290_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net424),
    .D(_0200_),
    .Q_N(_5289_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net425),
    .D(_0201_),
    .Q_N(_5288_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net426),
    .D(_0202_),
    .Q_N(_5287_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net427),
    .D(_0203_),
    .Q_N(_5286_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net428),
    .D(_0204_),
    .Q_N(_5285_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net429),
    .D(_0205_),
    .Q_N(_5284_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net430),
    .D(_0206_),
    .Q_N(_5283_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net431),
    .D(_0207_),
    .Q_N(_5282_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net432),
    .D(_0208_),
    .Q_N(_5281_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net433),
    .D(_0209_),
    .Q_N(_5280_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net434),
    .D(_0210_),
    .Q_N(_5279_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net435),
    .D(_0211_),
    .Q_N(_5278_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net436),
    .D(_0212_),
    .Q_N(_5277_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net437),
    .D(_0213_),
    .Q_N(_5276_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net438),
    .D(_0214_),
    .Q_N(_5275_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net439),
    .D(_0215_),
    .Q_N(_0039_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net440),
    .D(_0216_),
    .Q_N(_5274_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net441),
    .D(_0217_),
    .Q_N(_0028_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net442),
    .D(_0218_),
    .Q_N(_5273_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net443),
    .D(_0219_),
    .Q_N(_5272_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net444),
    .D(_0220_),
    .Q_N(_5271_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net445),
    .D(_0221_),
    .Q_N(_5270_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net446),
    .D(_0222_),
    .Q_N(_5269_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net447),
    .D(_0223_),
    .Q_N(_5268_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net448),
    .D(_0224_),
    .Q_N(_5267_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net449),
    .D(_0225_),
    .Q_N(_5266_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net450),
    .D(_0226_),
    .Q_N(_5265_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net451),
    .D(_0227_),
    .Q_N(_5264_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net452),
    .D(_0228_),
    .Q_N(_5263_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net453),
    .D(_0229_),
    .Q_N(_5262_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net454),
    .D(_0230_),
    .Q_N(_5261_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net455),
    .D(_0231_),
    .Q_N(_5260_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net456),
    .D(_0232_),
    .Q_N(_5259_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net457),
    .D(_0233_),
    .Q_N(_5258_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net458),
    .D(_0234_),
    .Q_N(_5257_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net459),
    .D(_0235_),
    .Q_N(_5256_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net460),
    .D(_0236_),
    .Q_N(_5255_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net461),
    .D(_0237_),
    .Q_N(_5254_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net462),
    .D(_0238_),
    .Q_N(_5253_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net463),
    .D(_0239_),
    .Q_N(_5252_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net464),
    .D(_0240_),
    .Q_N(_5251_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net465),
    .D(_0241_),
    .Q_N(_5250_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net466),
    .D(_0242_),
    .Q_N(_5249_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net467),
    .D(_0243_),
    .Q_N(_5248_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net468),
    .D(_0244_),
    .Q_N(_5247_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net469),
    .D(_0245_),
    .Q_N(_5246_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net470),
    .D(_0246_),
    .Q_N(_5245_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net471),
    .D(_0247_),
    .Q_N(_5244_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net472),
    .D(_0248_),
    .Q_N(_5243_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net473),
    .D(_0249_),
    .Q_N(_5242_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net474),
    .D(_0250_),
    .Q_N(_5241_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net475),
    .D(_0251_),
    .Q_N(_5240_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net476),
    .D(_0252_),
    .Q_N(_5239_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net477),
    .D(_0253_),
    .Q_N(_5238_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net478),
    .D(_0254_),
    .Q_N(_5237_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net479),
    .D(_0255_),
    .Q_N(_5236_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net480),
    .D(_0256_),
    .Q_N(_5235_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net481),
    .D(_0257_),
    .Q_N(_5234_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net482),
    .D(_0258_),
    .Q_N(_5233_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net483),
    .D(_0259_),
    .Q_N(_5232_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net484),
    .D(_0260_),
    .Q_N(_5231_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net485),
    .D(_0261_),
    .Q_N(_5230_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net486),
    .D(_0262_),
    .Q_N(_5229_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net487),
    .D(_0263_),
    .Q_N(_5228_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net488),
    .D(_0264_),
    .Q_N(_5227_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net489),
    .D(_0265_),
    .Q_N(_5226_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net490),
    .D(_0266_),
    .Q_N(_5225_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net491),
    .D(_0267_),
    .Q_N(_5224_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net492),
    .D(_0268_),
    .Q_N(_5223_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net493),
    .D(_0269_),
    .Q_N(_5222_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net494),
    .D(_0270_),
    .Q_N(_5221_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net495),
    .D(_0271_),
    .Q_N(_5220_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net496),
    .D(_0272_),
    .Q_N(_5219_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net497),
    .D(_0273_),
    .Q_N(_5218_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net498),
    .D(_0274_),
    .Q_N(_5217_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net499),
    .D(_0275_),
    .Q_N(_5216_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net500),
    .D(_0276_),
    .Q_N(_5215_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net501),
    .D(_0277_),
    .Q_N(_5214_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net502),
    .D(_0278_),
    .Q_N(_5213_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net503),
    .D(_0279_),
    .Q_N(_5212_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net504),
    .D(_0280_),
    .Q_N(_5211_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net505),
    .D(_0281_),
    .Q_N(_5210_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net506),
    .D(_0282_),
    .Q_N(_5209_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net507),
    .D(_0283_),
    .Q_N(_5208_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net508),
    .D(_0284_),
    .Q_N(_5207_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net509),
    .D(_0285_),
    .Q_N(_5206_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net510),
    .D(_0286_),
    .Q_N(_5205_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net511),
    .D(_0287_),
    .Q_N(_5204_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net512),
    .D(_0288_),
    .Q_N(_5203_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net513),
    .D(_0289_),
    .Q_N(_5202_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net514),
    .D(_0290_),
    .Q_N(_5201_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net515),
    .D(_0291_),
    .Q_N(_5200_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net516),
    .D(_0292_),
    .Q_N(_5199_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net517),
    .D(_0293_),
    .Q_N(_5198_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net518),
    .D(_0294_),
    .Q_N(_5197_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net519),
    .D(_0295_),
    .Q_N(_5196_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net520),
    .D(_0296_),
    .Q_N(_5195_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net521),
    .D(_0297_),
    .Q_N(_5194_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net522),
    .D(_0298_),
    .Q_N(_5193_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net523),
    .D(_0299_),
    .Q_N(_5192_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net524),
    .D(_0300_),
    .Q_N(_5191_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net525),
    .D(_0301_),
    .Q_N(_5190_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net526),
    .D(_0302_),
    .Q_N(_5189_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net527),
    .D(_0303_),
    .Q_N(_5188_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net528),
    .D(_0304_),
    .Q_N(_5187_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net529),
    .D(_0305_),
    .Q_N(_5186_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net530),
    .D(_0306_),
    .Q_N(_5185_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net531),
    .D(_0307_),
    .Q_N(_5184_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net532),
    .D(_0308_),
    .Q_N(_5183_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net533),
    .D(_0309_),
    .Q_N(_5182_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net534),
    .D(_0310_),
    .Q_N(_5181_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net535),
    .D(_0311_),
    .Q_N(_5180_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net536),
    .D(_0312_),
    .Q_N(_5179_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net537),
    .D(_0313_),
    .Q_N(_5178_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net538),
    .D(_0314_),
    .Q_N(_5177_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net539),
    .D(_0315_),
    .Q_N(_5176_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net540),
    .D(_0316_),
    .Q_N(_5175_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net541),
    .D(_0317_),
    .Q_N(_5174_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net542),
    .D(_0318_),
    .Q_N(_5173_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net543),
    .D(_0319_),
    .Q_N(_5172_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net544),
    .D(_0320_),
    .Q_N(_5171_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net545),
    .D(_0321_),
    .Q_N(_5170_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net546),
    .D(_0322_),
    .Q_N(_5169_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net547),
    .D(_0323_),
    .Q_N(_5168_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net548),
    .D(_0324_),
    .Q_N(_5167_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net549),
    .D(_0325_),
    .Q_N(_5166_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net550),
    .D(_0326_),
    .Q_N(_5165_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net551),
    .D(_0327_),
    .Q_N(_5164_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net552),
    .D(_0328_),
    .Q_N(_5163_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net553),
    .D(_0329_),
    .Q_N(_5162_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net554),
    .D(_0330_),
    .Q_N(_5161_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net555),
    .D(_0331_),
    .Q_N(_5160_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net556),
    .D(_0332_),
    .Q_N(_5159_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net557),
    .D(_0333_),
    .Q_N(_5158_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net558),
    .D(_0334_),
    .Q_N(_5157_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net559),
    .D(_0335_),
    .Q_N(_5156_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net560),
    .D(_0336_),
    .Q_N(_5155_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net561),
    .D(_0337_),
    .Q_N(_5154_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net562),
    .D(_0338_),
    .Q_N(_5153_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net563),
    .D(_0339_),
    .Q_N(_5152_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net564),
    .D(_0340_),
    .Q_N(_5151_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net565),
    .D(_0341_),
    .Q_N(_5150_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net566),
    .D(_0342_),
    .Q_N(_5149_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net567),
    .D(_0343_),
    .Q_N(_5148_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net568),
    .D(_0344_),
    .Q_N(_5147_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net569),
    .D(_0345_),
    .Q_N(_5146_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net570),
    .D(_0346_),
    .Q_N(_5145_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net571),
    .D(_0347_),
    .Q_N(_5144_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net572),
    .D(_0348_),
    .Q_N(_5143_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net573),
    .D(_0349_),
    .Q_N(_5142_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net574),
    .D(_0350_),
    .Q_N(_5141_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net575),
    .D(_0351_),
    .Q_N(_5140_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net576),
    .D(_0352_),
    .Q_N(_5139_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net577),
    .D(_0353_),
    .Q_N(_5138_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net578),
    .D(_0354_),
    .Q_N(_5137_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net579),
    .D(_0355_),
    .Q_N(_5136_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net580),
    .D(_0356_),
    .Q_N(_5135_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net581),
    .D(_0357_),
    .Q_N(_5134_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net582),
    .D(_0358_),
    .Q_N(_5133_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net583),
    .D(_0359_),
    .Q_N(_5132_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net584),
    .D(_0360_),
    .Q_N(_5131_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net585),
    .D(_0361_),
    .Q_N(_5130_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net586),
    .D(_0362_),
    .Q_N(_5129_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net587),
    .D(_0363_),
    .Q_N(_5128_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net588),
    .D(_0364_),
    .Q_N(_5127_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net589),
    .D(_0365_),
    .Q_N(_5126_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net590),
    .D(_0366_),
    .Q_N(_5125_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net591),
    .D(_0367_),
    .Q_N(_5124_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net592),
    .D(_0368_),
    .Q_N(_5123_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net593),
    .D(_0369_),
    .Q_N(_5122_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net594),
    .D(_0370_),
    .Q_N(_5121_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net595),
    .D(_0371_),
    .Q_N(_5120_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net596),
    .D(_0372_),
    .Q_N(_5119_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net597),
    .D(_0373_),
    .Q_N(_5118_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net598),
    .D(_0374_),
    .Q_N(_5117_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net599),
    .D(_0375_),
    .Q_N(_5116_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net600),
    .D(_0376_),
    .Q_N(_5115_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net601),
    .D(_0377_),
    .Q_N(_5114_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net602),
    .D(_0378_),
    .Q_N(_5113_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net603),
    .D(_0379_),
    .Q_N(_5112_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net604),
    .D(_0380_),
    .Q_N(_5111_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net605),
    .D(_0381_),
    .Q_N(_5110_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net606),
    .D(_0382_),
    .Q_N(_5109_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net607),
    .D(_0383_),
    .Q_N(_5108_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net608),
    .D(_0384_),
    .Q_N(_5107_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net609),
    .D(_0385_),
    .Q_N(_5106_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net610),
    .D(_0386_),
    .Q_N(_5105_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net611),
    .D(_0387_),
    .Q_N(_5104_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net612),
    .D(_0388_),
    .Q_N(_5103_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net613),
    .D(_0389_),
    .Q_N(_5102_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net614),
    .D(_0390_),
    .Q_N(_5101_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net615),
    .D(_0391_),
    .Q_N(_5100_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net616),
    .D(_0392_),
    .Q_N(_5099_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net617),
    .D(_0393_),
    .Q_N(_5098_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net618),
    .D(_0394_),
    .Q_N(_5097_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net619),
    .D(_0395_),
    .Q_N(_5096_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net620),
    .D(_0396_),
    .Q_N(_5095_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net621),
    .D(_0397_),
    .Q_N(_5094_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net622),
    .D(_0398_),
    .Q_N(_5093_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net623),
    .D(_0399_),
    .Q_N(_5092_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net624),
    .D(_0400_),
    .Q_N(_5091_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net625),
    .D(_0401_),
    .Q_N(_5090_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net626),
    .D(_0402_),
    .Q_N(_5089_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net627),
    .D(_0403_),
    .Q_N(_5088_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net628),
    .D(_0404_),
    .Q_N(_5087_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net629),
    .D(_0405_),
    .Q_N(_5086_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net630),
    .D(_0406_),
    .Q_N(_5085_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net631),
    .D(_0407_),
    .Q_N(_5084_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net632),
    .D(_0408_),
    .Q_N(_5083_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net633),
    .D(_0409_),
    .Q_N(_5082_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net634),
    .D(_0410_),
    .Q_N(_5081_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net635),
    .D(_0411_),
    .Q_N(_5080_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net636),
    .D(_0412_),
    .Q_N(_5079_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net637),
    .D(_0413_),
    .Q_N(_5078_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net638),
    .D(_0414_),
    .Q_N(_5077_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net639),
    .D(_0415_),
    .Q_N(_5076_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net640),
    .D(_0416_),
    .Q_N(_5075_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net641),
    .D(_0417_),
    .Q_N(_5074_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net642),
    .D(_0418_),
    .Q_N(_5073_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net643),
    .D(_0419_),
    .Q_N(_5072_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net644),
    .D(_0420_),
    .Q_N(_5071_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net645),
    .D(_0421_),
    .Q_N(_5070_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net646),
    .D(_0422_),
    .Q_N(_5069_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net647),
    .D(_0423_),
    .Q_N(_5068_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net648),
    .D(_0424_),
    .Q_N(_5067_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net649),
    .D(_0425_),
    .Q_N(_5066_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net650),
    .D(_0426_),
    .Q_N(_5065_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net651),
    .D(_0427_),
    .Q_N(_5064_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net652),
    .D(_0428_),
    .Q_N(_5063_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net653),
    .D(_0429_),
    .Q_N(_5062_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net654),
    .D(_0430_),
    .Q_N(_5061_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net655),
    .D(_0431_),
    .Q_N(_5060_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net656),
    .D(_0432_),
    .Q_N(_5059_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net657),
    .D(_0433_),
    .Q_N(_5058_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net658),
    .D(_0434_),
    .Q_N(_5057_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net659),
    .D(_0435_),
    .Q_N(_5056_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net660),
    .D(_0436_),
    .Q_N(_5055_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net661),
    .D(_0437_),
    .Q_N(_5054_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net662),
    .D(_0438_),
    .Q_N(_5053_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net663),
    .D(_0439_),
    .Q_N(_5052_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net664),
    .D(_0440_),
    .Q_N(_5051_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net665),
    .D(_0441_),
    .Q_N(_5050_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net666),
    .D(_0442_),
    .Q_N(_5049_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net667),
    .D(_0443_),
    .Q_N(_5048_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net668),
    .D(_0444_),
    .Q_N(_5047_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net669),
    .D(_0445_),
    .Q_N(_5046_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net670),
    .D(_0446_),
    .Q_N(_5045_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net671),
    .D(_0447_),
    .Q_N(_5044_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net672),
    .D(_0448_),
    .Q_N(_5043_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net673),
    .D(_0449_),
    .Q_N(_5042_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net674),
    .D(_0450_),
    .Q_N(_5041_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net675),
    .D(_0451_),
    .Q_N(_5040_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net676),
    .D(_0452_),
    .Q_N(_5039_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net677),
    .D(_0453_),
    .Q_N(_5038_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net678),
    .D(_0454_),
    .Q_N(_5037_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net679),
    .D(_0455_),
    .Q_N(_5036_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net680),
    .D(_0456_),
    .Q_N(_5035_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net681),
    .D(_0457_),
    .Q_N(_5034_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net682),
    .D(_0458_),
    .Q_N(_5033_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net683),
    .D(_0459_),
    .Q_N(_5032_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net684),
    .D(_0460_),
    .Q_N(_5031_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net685),
    .D(_0461_),
    .Q_N(_5030_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net686),
    .D(_0462_),
    .Q_N(_5029_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net687),
    .D(_0463_),
    .Q_N(_5028_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net688),
    .D(_0464_),
    .Q_N(_5027_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net689),
    .D(_0465_),
    .Q_N(_5026_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net690),
    .D(_0466_),
    .Q_N(_5025_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net691),
    .D(_0467_),
    .Q_N(_5024_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net692),
    .D(_0468_),
    .Q_N(_5023_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net693),
    .D(_0469_),
    .Q_N(_5022_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net694),
    .D(_0470_),
    .Q_N(_5021_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net695),
    .D(_0471_),
    .Q_N(_5020_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net696),
    .D(_0472_),
    .Q_N(_5019_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net697),
    .D(_0473_),
    .Q_N(_5018_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net698),
    .D(_0474_),
    .Q_N(_5017_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net699),
    .D(_0475_),
    .Q_N(_5016_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net700),
    .D(_0476_),
    .Q_N(_5015_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net701),
    .D(_0477_),
    .Q_N(_5014_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net702),
    .D(_0478_),
    .Q_N(_5013_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net703),
    .D(_0479_),
    .Q_N(_5012_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net704),
    .D(_0480_),
    .Q_N(_5011_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net705),
    .D(_0481_),
    .Q_N(_5010_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net706),
    .D(_0482_),
    .Q_N(_5009_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net707),
    .D(_0483_),
    .Q_N(_5008_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net708),
    .D(_0484_),
    .Q_N(_5007_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net709),
    .D(_0485_),
    .Q_N(_5006_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net710),
    .D(_0486_),
    .Q_N(_5005_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net711),
    .D(_0487_),
    .Q_N(_5004_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net712),
    .D(_0488_),
    .Q_N(_5003_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net713),
    .D(_0489_),
    .Q_N(_5002_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net714),
    .D(_0490_),
    .Q_N(_5001_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net715),
    .D(_0491_),
    .Q_N(_5000_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net716),
    .D(_0492_),
    .Q_N(_4999_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net717),
    .D(_0493_),
    .Q_N(_4998_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net718),
    .D(_0494_),
    .Q_N(_4997_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net719),
    .D(_0495_),
    .Q_N(_4996_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net720),
    .D(_0496_),
    .Q_N(_4995_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net721),
    .D(_0497_),
    .Q_N(_4994_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net722),
    .D(_0498_),
    .Q_N(_4993_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net723),
    .D(_0499_),
    .Q_N(_4992_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net724),
    .D(_0500_),
    .Q_N(_4991_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net725),
    .D(_0501_),
    .Q_N(_4990_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net726),
    .D(_0502_),
    .Q_N(_4989_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net727),
    .D(_0503_),
    .Q_N(_4988_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net728),
    .D(_0504_),
    .Q_N(_4987_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net729),
    .D(_0505_),
    .Q_N(_4986_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net730),
    .D(_0506_),
    .Q_N(_4985_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net731),
    .D(_0507_),
    .Q_N(_4984_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net732),
    .D(_0508_),
    .Q_N(_4983_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net733),
    .D(_0509_),
    .Q_N(_4982_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net734),
    .D(_0510_),
    .Q_N(_4981_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net735),
    .D(_0511_),
    .Q_N(_4980_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net736),
    .D(_0512_),
    .Q_N(_4979_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net737),
    .D(_0513_),
    .Q_N(_4978_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net738),
    .D(_0514_),
    .Q_N(_4977_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net739),
    .D(_0515_),
    .Q_N(_4976_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net740),
    .D(_0516_),
    .Q_N(_4975_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net741),
    .D(_0517_),
    .Q_N(_4974_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net742),
    .D(_0518_),
    .Q_N(_4973_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net743),
    .D(_0519_),
    .Q_N(_4972_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net744),
    .D(_0520_),
    .Q_N(_4971_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net745),
    .D(_0521_),
    .Q_N(_4970_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net746),
    .D(_0522_),
    .Q_N(_4969_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net747),
    .D(_0523_),
    .Q_N(_4968_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net748),
    .D(_0524_),
    .Q_N(_4967_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net749),
    .D(_0525_),
    .Q_N(_4966_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net750),
    .D(_0526_),
    .Q_N(_4965_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net751),
    .D(_0527_),
    .Q_N(_4964_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net752),
    .D(_0528_),
    .Q_N(_4963_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net753),
    .D(_0529_),
    .Q_N(_4962_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net754),
    .D(_0530_),
    .Q_N(_4961_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net755),
    .D(_0531_),
    .Q_N(_4960_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net756),
    .D(_0532_),
    .Q_N(_4959_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net757),
    .D(_0533_),
    .Q_N(_4958_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net758),
    .D(_0534_),
    .Q_N(_4957_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net759),
    .D(_0535_),
    .Q_N(_4956_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net760),
    .D(_0536_),
    .Q_N(_4955_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net761),
    .D(_0537_),
    .Q_N(_4954_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net762),
    .D(_0538_),
    .Q_N(_4953_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net763),
    .D(_0539_),
    .Q_N(_4952_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net764),
    .D(_0540_),
    .Q_N(_4951_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net765),
    .D(_0541_),
    .Q_N(_4950_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net766),
    .D(_0542_),
    .Q_N(_4949_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net767),
    .D(_0543_),
    .Q_N(_4948_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net768),
    .D(_0544_),
    .Q_N(_4947_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net769),
    .D(_0545_),
    .Q_N(_4946_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net770),
    .D(_0546_),
    .Q_N(_4945_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net771),
    .D(_0547_),
    .Q_N(_4944_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net772),
    .D(_0548_),
    .Q_N(_4943_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net773),
    .D(_0549_),
    .Q_N(_4942_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net774),
    .D(_0550_),
    .Q_N(_4941_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net775),
    .D(_0551_),
    .Q_N(_4940_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net776),
    .D(_0552_),
    .Q_N(_4939_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net777),
    .D(_0553_),
    .Q_N(_4938_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net778),
    .D(_0554_),
    .Q_N(_4937_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net779),
    .D(_0555_),
    .Q_N(_4936_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net780),
    .D(_0556_),
    .Q_N(_4935_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net781),
    .D(_0557_),
    .Q_N(_4934_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net782),
    .D(_0558_),
    .Q_N(_4933_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net783),
    .D(_0559_),
    .Q_N(_4932_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net784),
    .D(_0560_),
    .Q_N(_4931_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net785),
    .D(_0561_),
    .Q_N(_4930_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net786),
    .D(_0562_),
    .Q_N(_4929_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net787),
    .D(_0563_),
    .Q_N(_4928_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net788),
    .D(_0564_),
    .Q_N(_4927_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net789),
    .D(_0565_),
    .Q_N(_4926_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net790),
    .D(_0566_),
    .Q_N(_4925_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net791),
    .D(_0567_),
    .Q_N(_4924_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net792),
    .D(_0568_),
    .Q_N(_4923_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net793),
    .D(_0569_),
    .Q_N(_4922_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net794),
    .D(_0570_),
    .Q_N(_4921_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net795),
    .D(_0571_),
    .Q_N(_4920_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net796),
    .D(_0572_),
    .Q_N(_4919_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net797),
    .D(_0573_),
    .Q_N(_4918_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net798),
    .D(_0574_),
    .Q_N(_4917_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net799),
    .D(_0575_),
    .Q_N(_4916_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net800),
    .D(_0576_),
    .Q_N(_4915_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net801),
    .D(_0577_),
    .Q_N(_4914_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net802),
    .D(_0578_),
    .Q_N(_4913_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net803),
    .D(_0579_),
    .Q_N(_4912_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net804),
    .D(_0580_),
    .Q_N(_4911_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net805),
    .D(_0581_),
    .Q_N(_4910_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net806),
    .D(_0582_),
    .Q_N(_4909_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net807),
    .D(_0583_),
    .Q_N(_4908_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net808),
    .D(_0584_),
    .Q_N(_4907_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net809),
    .D(_0585_),
    .Q_N(_4906_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net810),
    .D(_0586_),
    .Q_N(_4905_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net811),
    .D(_0587_),
    .Q_N(_4904_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net812),
    .D(_0588_),
    .Q_N(_4903_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net813),
    .D(_0589_),
    .Q_N(_4902_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net814),
    .D(_0590_),
    .Q_N(_4901_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net815),
    .D(_0591_),
    .Q_N(_4900_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net816),
    .D(_0592_),
    .Q_N(_4899_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net817),
    .D(_0593_),
    .Q_N(_4898_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net818),
    .D(_0594_),
    .Q_N(_4897_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net819),
    .D(_0595_),
    .Q_N(_4896_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net820),
    .D(_0596_),
    .Q_N(_4895_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net821),
    .D(_0597_),
    .Q_N(_4894_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net822),
    .D(_0598_),
    .Q_N(_4893_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net823),
    .D(_0599_),
    .Q_N(_4892_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net824),
    .D(_0600_),
    .Q_N(_4891_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net825),
    .D(_0601_),
    .Q_N(_4890_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net826),
    .D(_0602_),
    .Q_N(_4889_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net827),
    .D(_0603_),
    .Q_N(_4888_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net828),
    .D(_0604_),
    .Q_N(_4887_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net829),
    .D(_0605_),
    .Q_N(_4886_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net830),
    .D(_0606_),
    .Q_N(_4885_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net831),
    .D(_0607_),
    .Q_N(_4884_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net832),
    .D(_0608_),
    .Q_N(_4883_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net833),
    .D(_0609_),
    .Q_N(_4882_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net834),
    .D(_0610_),
    .Q_N(_4881_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net835),
    .D(_0611_),
    .Q_N(_4880_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net836),
    .D(_0612_),
    .Q_N(_4879_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net837),
    .D(_0613_),
    .Q_N(_4878_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net838),
    .D(_0614_),
    .Q_N(_4877_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net839),
    .D(_0615_),
    .Q_N(_4876_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net840),
    .D(_0616_),
    .Q_N(_4875_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net841),
    .D(_0617_),
    .Q_N(_4874_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net842),
    .D(_0618_),
    .Q_N(_4873_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net843),
    .D(_0619_),
    .Q_N(_4872_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net844),
    .D(_0620_),
    .Q_N(_4871_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net845),
    .D(_0621_),
    .Q_N(_4870_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net846),
    .D(_0622_),
    .Q_N(_4869_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net847),
    .D(_0623_),
    .Q_N(_4868_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net848),
    .D(_0624_),
    .Q_N(_4867_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net849),
    .D(_0625_),
    .Q_N(_4866_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net850),
    .D(_0626_),
    .Q_N(_4865_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net851),
    .D(_0627_),
    .Q_N(_4864_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net852),
    .D(_0628_),
    .Q_N(_4863_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net853),
    .D(_0629_),
    .Q_N(_4862_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net854),
    .D(_0630_),
    .Q_N(_4861_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net855),
    .D(_0631_),
    .Q_N(_4860_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net856),
    .D(_0632_),
    .Q_N(_4859_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net857),
    .D(_0633_),
    .Q_N(_4858_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net858),
    .D(_0634_),
    .Q_N(_4857_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net859),
    .D(_0635_),
    .Q_N(_4856_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net860),
    .D(_0636_),
    .Q_N(_4855_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net861),
    .D(_0637_),
    .Q_N(_4854_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net862),
    .D(_0638_),
    .Q_N(_4853_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net863),
    .D(_0639_),
    .Q_N(_4852_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net864),
    .D(_0640_),
    .Q_N(_4851_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net865),
    .D(_0641_),
    .Q_N(_4850_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net866),
    .D(_0642_),
    .Q_N(_4849_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net867),
    .D(_0643_),
    .Q_N(_4848_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net868),
    .D(_0644_),
    .Q_N(_4847_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net869),
    .D(_0645_),
    .Q_N(_4846_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net870),
    .D(_0646_),
    .Q_N(_4845_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net871),
    .D(_0647_),
    .Q_N(_4844_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net872),
    .D(_0648_),
    .Q_N(_4843_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net873),
    .D(_0649_),
    .Q_N(_4842_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net874),
    .D(_0650_),
    .Q_N(_4841_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net875),
    .D(_0651_),
    .Q_N(_4840_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net876),
    .D(_0652_),
    .Q_N(_4839_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net877),
    .D(_0653_),
    .Q_N(_4838_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net878),
    .D(_0654_),
    .Q_N(_4837_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net879),
    .D(_0655_),
    .Q_N(_4836_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net880),
    .D(_0656_),
    .Q_N(_4835_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net881),
    .D(_0657_),
    .Q_N(_4834_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net882),
    .D(_0658_),
    .Q_N(_4833_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net883),
    .D(_0659_),
    .Q_N(_4832_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net884),
    .D(_0660_),
    .Q_N(_4831_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net885),
    .D(_0661_),
    .Q_N(_4830_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net886),
    .D(_0662_),
    .Q_N(_4829_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net887),
    .D(_0663_),
    .Q_N(_4828_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net888),
    .D(_0664_),
    .Q_N(_4827_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net889),
    .D(_0665_),
    .Q_N(_4826_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net890),
    .D(_0666_),
    .Q_N(_4825_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net891),
    .D(_0667_),
    .Q_N(_4824_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net892),
    .D(_0668_),
    .Q_N(_4823_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net893),
    .D(_0669_),
    .Q_N(_4822_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net894),
    .D(_0670_),
    .Q_N(_4821_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net895),
    .D(_0671_),
    .Q_N(_4820_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net896),
    .D(_0672_),
    .Q_N(_4819_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net897),
    .D(_0673_),
    .Q_N(_4818_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net898),
    .D(_0674_),
    .Q_N(_4817_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net899),
    .D(_0675_),
    .Q_N(_4816_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net900),
    .D(_0676_),
    .Q_N(_4815_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net901),
    .D(_0677_),
    .Q_N(_4814_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net902),
    .D(_0678_),
    .Q_N(_4813_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net903),
    .D(_0679_),
    .Q_N(_4812_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net904),
    .D(_0680_),
    .Q_N(_4811_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net905),
    .D(_0681_),
    .Q_N(_4810_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net906),
    .D(_0682_),
    .Q_N(_4809_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net907),
    .D(_0683_),
    .Q_N(_4808_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net908),
    .D(_0684_),
    .Q_N(_4807_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net909),
    .D(_0685_),
    .Q_N(_4806_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net910),
    .D(_0686_),
    .Q_N(_4805_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net911),
    .D(_0687_),
    .Q_N(_4804_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net912),
    .D(_0688_),
    .Q_N(_4803_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net913),
    .D(_0689_),
    .Q_N(_4802_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net914),
    .D(_0690_),
    .Q_N(_4801_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net915),
    .D(_0691_),
    .Q_N(_4800_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net916),
    .D(_0692_),
    .Q_N(_4799_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net917),
    .D(_0693_),
    .Q_N(_4798_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net918),
    .D(_0694_),
    .Q_N(_4797_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net919),
    .D(_0695_),
    .Q_N(_4796_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net920),
    .D(_0696_),
    .Q_N(_4795_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net921),
    .D(_0697_),
    .Q_N(_4794_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net922),
    .D(_0698_),
    .Q_N(_4793_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net923),
    .D(_0699_),
    .Q_N(_4792_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net924),
    .D(_0700_),
    .Q_N(_4791_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net925),
    .D(_0701_),
    .Q_N(_4790_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net926),
    .D(_0702_),
    .Q_N(_4789_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net927),
    .D(_0703_),
    .Q_N(_4788_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net928),
    .D(_0704_),
    .Q_N(_4787_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net929),
    .D(_0705_),
    .Q_N(_4786_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net930),
    .D(_0706_),
    .Q_N(_4785_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net931),
    .D(_0707_),
    .Q_N(_4784_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net932),
    .D(_0708_),
    .Q_N(_4783_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net933),
    .D(_0709_),
    .Q_N(_4782_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net934),
    .D(_0710_),
    .Q_N(_4781_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net935),
    .D(_0711_),
    .Q_N(_4780_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net936),
    .D(_0712_),
    .Q_N(_4779_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net937),
    .D(_0713_),
    .Q_N(_4778_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net938),
    .D(_0714_),
    .Q_N(_4777_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net939),
    .D(_0715_),
    .Q_N(_4776_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net940),
    .D(_0716_),
    .Q_N(_4775_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net941),
    .D(_0717_),
    .Q_N(_4774_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net942),
    .D(_0718_),
    .Q_N(_4773_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net943),
    .D(_0719_),
    .Q_N(_4772_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net944),
    .D(_0720_),
    .Q_N(_4771_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net945),
    .D(_0721_),
    .Q_N(_4770_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net946),
    .D(_0722_),
    .Q_N(_4769_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net947),
    .D(_0723_),
    .Q_N(_4768_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net948),
    .D(_0724_),
    .Q_N(_4767_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net949),
    .D(_0725_),
    .Q_N(_4766_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net950),
    .D(_0726_),
    .Q_N(_4765_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net951),
    .D(_0727_),
    .Q_N(_4764_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net952),
    .D(_0728_),
    .Q_N(_4763_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net953),
    .D(_0729_),
    .Q_N(_4762_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net954),
    .D(_0730_),
    .Q_N(_4761_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net955),
    .D(_0731_),
    .Q_N(_4760_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net956),
    .D(_0732_),
    .Q_N(_4759_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net957),
    .D(_0733_),
    .Q_N(_4758_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net958),
    .D(_0734_),
    .Q_N(_4757_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net959),
    .D(_0735_),
    .Q_N(_4756_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net960),
    .D(_0736_),
    .Q_N(_4755_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net961),
    .D(_0737_),
    .Q_N(_4754_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net962),
    .D(_0738_),
    .Q_N(_4753_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net963),
    .D(_0739_),
    .Q_N(_4752_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net964),
    .D(_0740_),
    .Q_N(_4751_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net965),
    .D(_0741_),
    .Q_N(_4750_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net966),
    .D(_0742_),
    .Q_N(_4749_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net967),
    .D(_0743_),
    .Q_N(_4748_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net968),
    .D(_0744_),
    .Q_N(_4747_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net969),
    .D(_0745_),
    .Q_N(_4746_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net970),
    .D(_0746_),
    .Q_N(_4745_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net971),
    .D(_0747_),
    .Q_N(_4744_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net972),
    .D(_0748_),
    .Q_N(_4743_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net973),
    .D(_0749_),
    .Q_N(_4742_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net974),
    .D(_0750_),
    .Q_N(_4741_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net975),
    .D(_0751_),
    .Q_N(_4740_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net976),
    .D(_0752_),
    .Q_N(_4739_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net977),
    .D(_0753_),
    .Q_N(_4738_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net978),
    .D(_0754_),
    .Q_N(_4737_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net979),
    .D(_0755_),
    .Q_N(_4736_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net980),
    .D(_0756_),
    .Q_N(_4735_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net981),
    .D(_0757_),
    .Q_N(_4734_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net982),
    .D(_0758_),
    .Q_N(_4733_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net983),
    .D(_0759_),
    .Q_N(_4732_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net984),
    .D(_0760_),
    .Q_N(_4731_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net985),
    .D(_0761_),
    .Q_N(_4730_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net986),
    .D(_0762_),
    .Q_N(_4729_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net987),
    .D(_0763_),
    .Q_N(_4728_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net988),
    .D(_0764_),
    .Q_N(_4727_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net989),
    .D(_0765_),
    .Q_N(_4726_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net990),
    .D(_0766_),
    .Q_N(_4725_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net991),
    .D(_0767_),
    .Q_N(_4724_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net992),
    .D(_0768_),
    .Q_N(_4723_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net993),
    .D(_0769_),
    .Q_N(_4722_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net994),
    .D(_0770_),
    .Q_N(_4721_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net995),
    .D(_0771_),
    .Q_N(_4720_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net996),
    .D(_0772_),
    .Q_N(_4719_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net997),
    .D(_0773_),
    .Q_N(_4718_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net998),
    .D(_0774_),
    .Q_N(_4717_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net999),
    .D(_0775_),
    .Q_N(_4716_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1000),
    .D(_0776_),
    .Q_N(_4715_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1001),
    .D(_0777_),
    .Q_N(_4714_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1002),
    .D(_0778_),
    .Q_N(_4713_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1003),
    .D(_0779_),
    .Q_N(_4712_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1004),
    .D(_0780_),
    .Q_N(_4711_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1005),
    .D(_0781_),
    .Q_N(_4710_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1006),
    .D(_0782_),
    .Q_N(_4709_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1007),
    .D(_0783_),
    .Q_N(_4708_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1008),
    .D(_0784_),
    .Q_N(_4707_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1009),
    .D(_0785_),
    .Q_N(_4706_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1010),
    .D(_0786_),
    .Q_N(_4705_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1011),
    .D(_0787_),
    .Q_N(_4704_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1012),
    .D(_0788_),
    .Q_N(_4703_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1013),
    .D(_0789_),
    .Q_N(_4702_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1014),
    .D(_0790_),
    .Q_N(_4701_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1015),
    .D(_0791_),
    .Q_N(_4700_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1016),
    .D(_0792_),
    .Q_N(_4699_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1017),
    .D(_0793_),
    .Q_N(_4698_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1018),
    .D(_0794_),
    .Q_N(_4697_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1019),
    .D(_0795_),
    .Q_N(_4696_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1020),
    .D(_0796_),
    .Q_N(_4695_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1021),
    .D(_0797_),
    .Q_N(_4694_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1022),
    .D(_0798_),
    .Q_N(_4693_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1023),
    .D(_0799_),
    .Q_N(_4692_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1024),
    .D(_0800_),
    .Q_N(_4691_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1025),
    .D(_0801_),
    .Q_N(_4690_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1026),
    .D(_0802_),
    .Q_N(_4689_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1027),
    .D(_0803_),
    .Q_N(_4688_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1028),
    .D(_0804_),
    .Q_N(_4687_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1029),
    .D(_0805_),
    .Q_N(_4686_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1030),
    .D(_0806_),
    .Q_N(_4685_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1031),
    .D(_0807_),
    .Q_N(_4684_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1032),
    .D(_0808_),
    .Q_N(_4683_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1033),
    .D(_0809_),
    .Q_N(_4682_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1034),
    .D(_0810_),
    .Q_N(_4681_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1035),
    .D(_0811_),
    .Q_N(_4680_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1036),
    .D(_0812_),
    .Q_N(_4679_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1037),
    .D(_0813_),
    .Q_N(_4678_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1038),
    .D(_0814_),
    .Q_N(_4677_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1039),
    .D(_0815_),
    .Q_N(_4676_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1040),
    .D(_0816_),
    .Q_N(_4675_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1041),
    .D(_0817_),
    .Q_N(_4674_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1042),
    .D(_0818_),
    .Q_N(_4673_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1043),
    .D(_0819_),
    .Q_N(_4672_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1044),
    .D(_0820_),
    .Q_N(_4671_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1045),
    .D(_0821_),
    .Q_N(_4670_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1046),
    .D(_0822_),
    .Q_N(_4669_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1047),
    .D(_0823_),
    .Q_N(_4668_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1048),
    .D(_0824_),
    .Q_N(_4667_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1049),
    .D(_0825_),
    .Q_N(_4666_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1050),
    .D(_0826_),
    .Q_N(_4665_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1051),
    .D(_0827_),
    .Q_N(_4664_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1052),
    .D(_0828_),
    .Q_N(_4663_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1053),
    .D(_0829_),
    .Q_N(_4662_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1054),
    .D(_0830_),
    .Q_N(_4661_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1055),
    .D(_0831_),
    .Q_N(_4660_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1056),
    .D(_0832_),
    .Q_N(_4659_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1057),
    .D(_0833_),
    .Q_N(_4658_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1058),
    .D(_0834_),
    .Q_N(_4657_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1059),
    .D(_0835_),
    .Q_N(_4656_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1060),
    .D(_0836_),
    .Q_N(_4655_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1061),
    .D(_0837_),
    .Q_N(_4654_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1062),
    .D(_0838_),
    .Q_N(_4653_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1063),
    .D(_0839_),
    .Q_N(_4652_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1064),
    .D(_0840_),
    .Q_N(_4651_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1065),
    .D(_0841_),
    .Q_N(_4650_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1066),
    .D(_0842_),
    .Q_N(_4649_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1067),
    .D(_0843_),
    .Q_N(_4648_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1068),
    .D(_0844_),
    .Q_N(_4647_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1069),
    .D(_0845_),
    .Q_N(_4646_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1070),
    .D(_0846_),
    .Q_N(_4645_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1071),
    .D(_0847_),
    .Q_N(_4644_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1072),
    .D(_0848_),
    .Q_N(_4643_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1073),
    .D(_0849_),
    .Q_N(_4642_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1074),
    .D(_0850_),
    .Q_N(_4641_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1075),
    .D(_0851_),
    .Q_N(_4640_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1076),
    .D(_0852_),
    .Q_N(_4639_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1077),
    .D(_0853_),
    .Q_N(_4638_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1078),
    .D(_0854_),
    .Q_N(_4637_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1079),
    .D(_0855_),
    .Q_N(_4636_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1080),
    .D(_0856_),
    .Q_N(_4635_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1081),
    .D(_0857_),
    .Q_N(_4634_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1082),
    .D(_0858_),
    .Q_N(_4633_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1083),
    .D(_0859_),
    .Q_N(_4632_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1084),
    .D(_0860_),
    .Q_N(_4631_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1085),
    .D(_0861_),
    .Q_N(_4630_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1086),
    .D(_0862_),
    .Q_N(_4629_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1087),
    .D(_0863_),
    .Q_N(_4628_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1088),
    .D(_0864_),
    .Q_N(_4627_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1089),
    .D(_0865_),
    .Q_N(_4626_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1090),
    .D(_0866_),
    .Q_N(_4625_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1091),
    .D(_0867_),
    .Q_N(_4624_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1092),
    .D(_0868_),
    .Q_N(_4623_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1093),
    .D(_0869_),
    .Q_N(_4622_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1094),
    .D(_0870_),
    .Q_N(_4621_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1095),
    .D(_0871_),
    .Q_N(_4620_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1096),
    .D(_0872_),
    .Q_N(_4619_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1097),
    .D(_0873_),
    .Q_N(_4618_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1098),
    .D(_0874_),
    .Q_N(_4617_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1099),
    .D(_0875_),
    .Q_N(_4616_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1100),
    .D(_0876_),
    .Q_N(_4615_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1101),
    .D(_0877_),
    .Q_N(_4614_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1102),
    .D(_0878_),
    .Q_N(_4613_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1103),
    .D(_0879_),
    .Q_N(_4612_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1104),
    .D(_0880_),
    .Q_N(_4611_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1105),
    .D(_0881_),
    .Q_N(_4610_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1106),
    .D(_0882_),
    .Q_N(_4609_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1107),
    .D(_0883_),
    .Q_N(_4608_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1108),
    .D(_0884_),
    .Q_N(_4607_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1109),
    .D(_0885_),
    .Q_N(_4606_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1110),
    .D(_0886_),
    .Q_N(_4605_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1111),
    .D(_0887_),
    .Q_N(_4604_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1112),
    .D(_0888_),
    .Q_N(_4603_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1113),
    .D(_0889_),
    .Q_N(_4602_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1114),
    .D(_0890_),
    .Q_N(_4601_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1115),
    .D(_0891_),
    .Q_N(_4600_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1116),
    .D(_0892_),
    .Q_N(_4599_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1117),
    .D(_0893_),
    .Q_N(_4598_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1118),
    .D(_0894_),
    .Q_N(_4597_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1119),
    .D(_0895_),
    .Q_N(_4596_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1120),
    .D(_0896_),
    .Q_N(_4595_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1121),
    .D(_0897_),
    .Q_N(_4594_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1122),
    .D(_0898_),
    .Q_N(_4593_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1123),
    .D(_0899_),
    .Q_N(_4592_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1124),
    .D(_0900_),
    .Q_N(_4591_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1125),
    .D(_0901_),
    .Q_N(_4590_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1126),
    .D(_0902_),
    .Q_N(_4589_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1127),
    .D(_0903_),
    .Q_N(_4588_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1128),
    .D(_0904_),
    .Q_N(_4587_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1129),
    .D(_0905_),
    .Q_N(_4586_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1130),
    .D(_0906_),
    .Q_N(_4585_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1131),
    .D(_0907_),
    .Q_N(_4584_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1132),
    .D(_0908_),
    .Q_N(_4583_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1133),
    .D(_0909_),
    .Q_N(_4582_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1134),
    .D(_0910_),
    .Q_N(_4581_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1135),
    .D(_0911_),
    .Q_N(_4580_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1136),
    .D(_0912_),
    .Q_N(_4579_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1137),
    .D(_0913_),
    .Q_N(_4578_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1138),
    .D(_0914_),
    .Q_N(_4577_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1139),
    .D(_0915_),
    .Q_N(_4576_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1140),
    .D(_0916_),
    .Q_N(_4575_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1141),
    .D(_0917_),
    .Q_N(_4574_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1142),
    .D(_0918_),
    .Q_N(_4573_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1143),
    .D(_0919_),
    .Q_N(_4572_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1144),
    .D(_0920_),
    .Q_N(_4571_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1145),
    .D(_0921_),
    .Q_N(_4570_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1146),
    .D(_0922_),
    .Q_N(_4569_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1147),
    .D(_0923_),
    .Q_N(_4568_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1148),
    .D(_0924_),
    .Q_N(_4567_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1149),
    .D(_0925_),
    .Q_N(_4566_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1150),
    .D(_0926_),
    .Q_N(_4565_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1151),
    .D(_0927_),
    .Q_N(_4564_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1152),
    .D(_0928_),
    .Q_N(_4563_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1153),
    .D(_0929_),
    .Q_N(_4562_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1154),
    .D(_0930_),
    .Q_N(_4561_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1155),
    .D(_0931_),
    .Q_N(_4560_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1156),
    .D(_0932_),
    .Q_N(_4559_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1157),
    .D(_0933_),
    .Q_N(_4558_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1158),
    .D(_0934_),
    .Q_N(_4557_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1159),
    .D(_0935_),
    .Q_N(_4556_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1160),
    .D(_0936_),
    .Q_N(_4555_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1161),
    .D(_0937_),
    .Q_N(_4554_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1162),
    .D(_0938_),
    .Q_N(_4553_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1163),
    .D(_0939_),
    .Q_N(_4552_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1164),
    .D(_0940_),
    .Q_N(_4551_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1165),
    .D(_0941_),
    .Q_N(_4550_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1166),
    .D(_0942_),
    .Q_N(_4549_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1167),
    .D(_0943_),
    .Q_N(_4548_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1168),
    .D(_0944_),
    .Q_N(_4547_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1169),
    .D(_0945_),
    .Q_N(_4546_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1170),
    .D(_0946_),
    .Q_N(_4545_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1171),
    .D(_0947_),
    .Q_N(_4544_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1172),
    .D(_0948_),
    .Q_N(_4543_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1173),
    .D(_0949_),
    .Q_N(_4542_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1174),
    .D(_0950_),
    .Q_N(_4541_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1175),
    .D(_0951_),
    .Q_N(_4540_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1176),
    .D(_0952_),
    .Q_N(_4539_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1177),
    .D(_0953_),
    .Q_N(_4538_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1178),
    .D(_0954_),
    .Q_N(_4537_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1179),
    .D(_0955_),
    .Q_N(_4536_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1180),
    .D(_0956_),
    .Q_N(_4535_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1181),
    .D(_0957_),
    .Q_N(_4534_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1182),
    .D(_0958_),
    .Q_N(_4533_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1183),
    .D(_0959_),
    .Q_N(_4532_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1184),
    .D(_0960_),
    .Q_N(_4531_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1185),
    .D(_0961_),
    .Q_N(_4530_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1186),
    .D(_0962_),
    .Q_N(_4529_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1187),
    .D(_0963_),
    .Q_N(_4528_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1188),
    .D(_0964_),
    .Q_N(_4527_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1189),
    .D(_0965_),
    .Q_N(_4526_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1190),
    .D(_0966_),
    .Q_N(_4525_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1191),
    .D(_0967_),
    .Q_N(_4524_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1192),
    .D(_0968_),
    .Q_N(_4523_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1193),
    .D(_0969_),
    .Q_N(_4522_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1194),
    .D(_0970_),
    .Q_N(_4521_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1195),
    .D(_0971_),
    .Q_N(_4520_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1196),
    .D(_0972_),
    .Q_N(_4519_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1197),
    .D(_0973_),
    .Q_N(_4518_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1198),
    .D(_0974_),
    .Q_N(_4517_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1199),
    .D(_0975_),
    .Q_N(_4516_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1200),
    .D(_0976_),
    .Q_N(_4515_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1201),
    .D(_0977_),
    .Q_N(_4514_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1202),
    .D(_0978_),
    .Q_N(_4513_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1203),
    .D(_0979_),
    .Q_N(_4512_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1204),
    .D(_0980_),
    .Q_N(_4511_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1205),
    .D(_0981_),
    .Q_N(_4510_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1206),
    .D(_0982_),
    .Q_N(_4509_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1207),
    .D(_0983_),
    .Q_N(_4508_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1208),
    .D(_0984_),
    .Q_N(_4507_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1209),
    .D(_0985_),
    .Q_N(_4506_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1210),
    .D(_0986_),
    .Q_N(_4505_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1211),
    .D(_0987_),
    .Q_N(_4504_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1212),
    .D(_0988_),
    .Q_N(_4503_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1213),
    .D(_0989_),
    .Q_N(_4502_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1214),
    .D(_0990_),
    .Q_N(_4501_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1215),
    .D(_0991_),
    .Q_N(_4500_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1216),
    .D(_0992_),
    .Q_N(_4499_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1217),
    .D(_0993_),
    .Q_N(_4498_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1218),
    .D(_0994_),
    .Q_N(_4497_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1219),
    .D(_0995_),
    .Q_N(_4496_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1220),
    .D(_0996_),
    .Q_N(_4495_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1221),
    .D(_0997_),
    .Q_N(_4494_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1222),
    .D(_0998_),
    .Q_N(_4493_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1223),
    .D(_0999_),
    .Q_N(_4492_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1224),
    .D(_1000_),
    .Q_N(_4491_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1225),
    .D(_1001_),
    .Q_N(_4490_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1226),
    .D(_1002_),
    .Q_N(_4489_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1227),
    .D(_1003_),
    .Q_N(_4488_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1228),
    .D(_1004_),
    .Q_N(_4487_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1229),
    .D(_1005_),
    .Q_N(_4486_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1230),
    .D(_1006_),
    .Q_N(_4485_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1231),
    .D(_1007_),
    .Q_N(_4484_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1232),
    .D(_1008_),
    .Q_N(_4483_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1233),
    .D(_1009_),
    .Q_N(_4482_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1234),
    .D(_1010_),
    .Q_N(_4481_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1235),
    .D(_1011_),
    .Q_N(_4480_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1236),
    .D(_1012_),
    .Q_N(_4479_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1237),
    .D(_1013_),
    .Q_N(_4478_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1238),
    .D(_1014_),
    .Q_N(_4477_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1239),
    .D(_1015_),
    .Q_N(_4476_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1240),
    .D(_1016_),
    .Q_N(_4475_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1241),
    .D(_1017_),
    .Q_N(_4474_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1242),
    .D(_1018_),
    .Q_N(_4473_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1243),
    .D(_1019_),
    .Q_N(_4472_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1244),
    .D(_1020_),
    .Q_N(_4471_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1245),
    .D(_1021_),
    .Q_N(_4470_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1246),
    .D(_1022_),
    .Q_N(_4469_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1247),
    .D(_1023_),
    .Q_N(_4468_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1248),
    .D(_1024_),
    .Q_N(_4467_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1249),
    .D(_1025_),
    .Q_N(_4466_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1250),
    .D(_1026_),
    .Q_N(_4465_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1251),
    .D(_1027_),
    .Q_N(_4464_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1252),
    .D(_1028_),
    .Q_N(_4463_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1253),
    .D(_1029_),
    .Q_N(_4462_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1254),
    .D(_1030_),
    .Q_N(_4461_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1255),
    .D(_1031_),
    .Q_N(_4460_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1256),
    .D(_1032_),
    .Q_N(_4459_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1257),
    .D(_1033_),
    .Q_N(_4458_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1258),
    .D(_1034_),
    .Q_N(_4457_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1259),
    .D(_1035_),
    .Q_N(_4456_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1260),
    .D(_1036_),
    .Q_N(_4455_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1261),
    .D(_1037_),
    .Q_N(_4454_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1262),
    .D(_1038_),
    .Q_N(_4453_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1263),
    .D(_1039_),
    .Q_N(_4452_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1264),
    .D(_1040_),
    .Q_N(_4451_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1265),
    .D(_1041_),
    .Q_N(_4450_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1266),
    .D(_1042_),
    .Q_N(_4449_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1267),
    .D(_1043_),
    .Q_N(_4448_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1268),
    .D(_1044_),
    .Q_N(_4447_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1269),
    .D(_1045_),
    .Q_N(_4446_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1270),
    .D(_1046_),
    .Q_N(_4445_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1271),
    .D(_1047_),
    .Q_N(_4444_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1272),
    .D(_1048_),
    .Q_N(_4443_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1273),
    .D(_1049_),
    .Q_N(_4442_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1274),
    .D(_1050_),
    .Q_N(_4441_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1275),
    .D(_1051_),
    .Q_N(_4440_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1276),
    .D(_1052_),
    .Q_N(_4439_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1277),
    .D(_1053_),
    .Q_N(_4438_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1278),
    .D(_1054_),
    .Q_N(_4437_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1279),
    .D(_1055_),
    .Q_N(_4436_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1280),
    .D(_1056_),
    .Q_N(_4435_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1281),
    .D(_1057_),
    .Q_N(_4434_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1282),
    .D(_1058_),
    .Q_N(_4433_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1283),
    .D(_1059_),
    .Q_N(_4432_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1284),
    .D(_1060_),
    .Q_N(_4431_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1285),
    .D(_1061_),
    .Q_N(_4430_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1286),
    .D(_1062_),
    .Q_N(_4429_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1287),
    .D(_1063_),
    .Q_N(_4428_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1288),
    .D(_1064_),
    .Q_N(_4427_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1289),
    .D(_1065_),
    .Q_N(_4426_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1290),
    .D(_1066_),
    .Q_N(_4425_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1291),
    .D(_1067_),
    .Q_N(_4424_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1292),
    .D(_1068_),
    .Q_N(_4423_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1293),
    .D(_1069_),
    .Q_N(_4422_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1294),
    .D(_1070_),
    .Q_N(_4421_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1295),
    .D(_1071_),
    .Q_N(_4420_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1296),
    .D(_1072_),
    .Q_N(_4419_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1297),
    .D(_1073_),
    .Q_N(_4418_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1298),
    .D(_1074_),
    .Q_N(_4417_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1299),
    .D(_1075_),
    .Q_N(_4416_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1300),
    .D(_1076_),
    .Q_N(_4415_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1301),
    .D(_1077_),
    .Q_N(_4414_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1302),
    .D(_1078_),
    .Q_N(_4413_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1303),
    .D(_1079_),
    .Q_N(_4412_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1304),
    .D(_1080_),
    .Q_N(_4411_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1305),
    .D(_1081_),
    .Q_N(_4410_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1306),
    .D(_1082_),
    .Q_N(_4409_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1307),
    .D(_1083_),
    .Q_N(_4408_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1308),
    .D(_1084_),
    .Q_N(_4407_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1309),
    .D(_1085_),
    .Q_N(_4406_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1310),
    .D(_1086_),
    .Q_N(_4405_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1311),
    .D(_1087_),
    .Q_N(_4404_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1312),
    .D(_1088_),
    .Q_N(_4403_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1313),
    .D(_1089_),
    .Q_N(_4402_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1314),
    .D(_1090_),
    .Q_N(_4401_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1315),
    .D(_1091_),
    .Q_N(_4400_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1316),
    .D(_1092_),
    .Q_N(_4399_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1317),
    .D(_1093_),
    .Q_N(_4398_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1318),
    .D(_1094_),
    .Q_N(_4397_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1319),
    .D(_1095_),
    .Q_N(_4396_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1320),
    .D(_1096_),
    .Q_N(_4395_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1321),
    .D(_1097_),
    .Q_N(_4394_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22]$_DFFE_PN_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1322),
    .D(_1098_),
    .Q_N(_4393_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1323),
    .D(_1099_),
    .Q_N(_4392_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1324),
    .D(_1100_),
    .Q_N(_4391_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1325),
    .D(_1101_),
    .Q_N(_4390_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26]$_DFFE_PN_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1326),
    .D(_1102_),
    .Q_N(_4389_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1327),
    .D(_1103_),
    .Q_N(_4388_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28]$_DFFE_PN_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1328),
    .D(_1104_),
    .Q_N(_4387_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1329),
    .D(_1105_),
    .Q_N(_4386_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1330),
    .D(_1106_),
    .Q_N(_4385_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1331),
    .D(_1107_),
    .Q_N(_4384_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1332),
    .D(_1108_),
    .Q_N(_4383_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1333),
    .D(_1109_),
    .Q_N(_4382_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6]$_DFFE_PN_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1334),
    .D(_1110_),
    .Q_N(_4381_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7]$_DFFE_PN_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1335),
    .D(_1111_),
    .Q_N(_4380_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8]$_DFFE_PN_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1336),
    .D(_1112_),
    .Q_N(_4379_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9]$_DFFE_PN_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1337),
    .D(_1113_),
    .Q_N(_4378_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1338),
    .D(_1114_),
    .Q_N(_4377_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1339),
    .D(_1115_),
    .Q_N(_0049_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1340),
    .D(_1116_),
    .Q_N(_0048_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1341),
    .D(_1117_),
    .Q_N(_0047_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1342),
    .D(_1118_),
    .Q_N(_0046_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1343),
    .D(_1119_),
    .Q_N(_4376_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[1]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1344),
    .D(_1120_),
    .Q_N(_4375_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1345),
    .D(_1121_),
    .Q_N(_4374_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[3]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1346),
    .D(_1122_),
    .Q_N(_4373_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[4]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1347),
    .D(_1123_),
    .Q_N(_0038_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1348),
    .D(_1124_),
    .Q_N(_4372_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1349),
    .D(_1125_),
    .Q_N(_4371_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1350),
    .D(_1126_),
    .Q_N(_4370_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[3]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1351),
    .D(_1127_),
    .Q_N(_4369_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1352),
    .D(_1128_),
    .Q_N(_0027_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_ack$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1353),
    .D(\i_exotiny._0003_ ),
    .Q_N(_0089_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_ack ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_shft$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1354),
    .D(\i_exotiny._0005_ ),
    .Q_N(_0021_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_shft ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_two$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1355),
    .D(\i_exotiny._0004_ ),
    .Q_N(_0032_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_two ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1356),
    .D(_1129_),
    .Q_N(\i_exotiny._2356_[0] ),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1]$_SDFF_PP0_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1357),
    .D(_1130_),
    .Q_N(_0030_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2]$_SDFF_PP0_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1358),
    .D(_1131_),
    .Q_N(_0029_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1359),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_msb ),
    .Q_N(_0040_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[0]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1360),
    .D(_1132_),
    .Q_N(_0023_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[1]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1361),
    .D(_1133_),
    .Q_N(_5374_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1362),
    .D(\i_exotiny._0083_ ),
    .Q_N(_0010_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[11]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1363),
    .D(\i_exotiny._0080_ ),
    .Q_N(_4368_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1364),
    .D(_1134_),
    .Q_N(_0105_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1365),
    .D(\i_exotiny._0067_ ),
    .Q_N(_0019_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[31]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1366),
    .D(\i_exotiny._0084_ ),
    .Q_N(_0009_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1367),
    .D(\i_exotiny._0068_ ),
    .Q_N(_0017_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1368),
    .D(\i_exotiny._0069_ ),
    .Q_N(_0015_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1369),
    .D(\i_exotiny._0070_ ),
    .Q_N(_0014_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1370),
    .D(\i_exotiny._0078_ ),
    .Q_N(_0013_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1371),
    .D(\i_exotiny._0081_ ),
    .Q_N(_0012_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1372),
    .D(_1135_),
    .Q_N(_0114_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[9]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1373),
    .D(\i_exotiny._0082_ ),
    .Q_N(_0011_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0]$_SDFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1374),
    .D(_1136_),
    .Q_N(_0108_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1375),
    .D(\i_exotiny._0064_ ),
    .Q_N(_0020_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1376),
    .D(\i_exotiny._0065_ ),
    .Q_N(_0018_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1377),
    .D(\i_exotiny._0066_ ),
    .Q_N(_0016_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1378),
    .D(_1137_),
    .Q_N(_0000_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1379),
    .D(_1138_),
    .Q_N(_4367_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1380),
    .D(_1139_),
    .Q_N(_0025_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1381),
    .D(_1140_),
    .Q_N(_0037_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1382),
    .D(_1141_),
    .Q_N(_0022_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1383),
    .D(_1142_),
    .Q_N(_0090_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[5]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1384),
    .D(_1143_),
    .Q_N(_0091_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[6]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1385),
    .D(_1144_),
    .Q_N(_0026_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1386),
    .D(_1145_),
    .Q_N(_4366_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1387),
    .D(_1146_),
    .Q_N(_4365_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1388),
    .D(_1147_),
    .Q_N(_4364_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1389),
    .D(_1148_),
    .Q_N(_4363_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1390),
    .D(_1149_),
    .Q_N(_4362_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1391),
    .D(_1150_),
    .Q_N(_4361_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1392),
    .D(_1151_),
    .Q_N(_4360_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1393),
    .D(_1152_),
    .Q_N(_4359_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1394),
    .D(_1153_),
    .Q_N(_4358_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1395),
    .D(_1154_),
    .Q_N(_4357_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1396),
    .D(_1155_),
    .Q_N(_4356_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1397),
    .D(_1156_),
    .Q_N(_4355_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1398),
    .D(_1157_),
    .Q_N(_4354_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1399),
    .D(_1158_),
    .Q_N(_4353_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1400),
    .D(_1159_),
    .Q_N(_4352_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1401),
    .D(_1160_),
    .Q_N(_4351_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1402),
    .D(_1161_),
    .Q_N(_4350_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1403),
    .D(_1162_),
    .Q_N(_4349_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1404),
    .D(_1163_),
    .Q_N(_4348_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1405),
    .D(_1164_),
    .Q_N(_4347_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1406),
    .D(_1165_),
    .Q_N(_4346_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1407),
    .D(_1166_),
    .Q_N(_4345_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1408),
    .D(_1167_),
    .Q_N(_4344_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1409),
    .D(_1168_),
    .Q_N(_4343_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1410),
    .D(_1169_),
    .Q_N(_4342_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1411),
    .D(_1170_),
    .Q_N(_4341_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1412),
    .D(_1171_),
    .Q_N(_4340_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1413),
    .D(_1172_),
    .Q_N(_4339_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1414),
    .D(_1173_),
    .Q_N(_4338_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1415),
    .D(_1174_),
    .Q_N(_4337_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1416),
    .D(_1175_),
    .Q_N(_4336_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1417),
    .D(_1176_),
    .Q_N(_4335_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0]$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1418),
    .D(_1177_),
    .Q_N(_0100_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[12]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1419),
    .D(_1178_),
    .Q_N(_5375_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1420),
    .D(\i_exotiny._0071_ ),
    .Q_N(_0065_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1421),
    .D(\i_exotiny._0072_ ),
    .Q_N(_0062_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[15]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1422),
    .D(\i_exotiny._0073_ ),
    .Q_N(_0061_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[16]$_SDFF_PN1_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1423),
    .D(_1179_),
    .Q_N(_0111_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1424),
    .D(\i_exotiny._0085_ ),
    .Q_N(_0084_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1425),
    .D(\i_exotiny._0062_ ),
    .Q_N(_0082_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1426),
    .D(\i_exotiny._0063_ ),
    .Q_N(_0080_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1427),
    .D(\i_exotiny._0074_ ),
    .Q_N(_0058_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[2]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1428),
    .D(\i_exotiny._0075_ ),
    .Q_N(_0055_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1429),
    .D(\i_exotiny._0076_ ),
    .Q_N(_0052_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[4]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1430),
    .D(_1180_),
    .Q_N(_5376_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[5]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1431),
    .D(\i_exotiny._0077_ ),
    .Q_N(_5377_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[6]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1432),
    .D(\i_exotiny._0079_ ),
    .Q_N(_4334_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ld_sext_o$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1433),
    .D(_1181_),
    .Q_N(_4333_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ld_sext_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1434),
    .D(_1182_),
    .Q_N(_0042_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_w_o$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1435),
    .D(_1183_),
    .Q_N(_0115_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_w_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1436),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.genblk1[3].i_fazyrv_fadd_x.c_o ),
    .Q_N(_5378_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1437),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.ex_cmp_tmp ),
    .Q_N(_0043_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.imem_stb_o$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1438),
    .D(\i_exotiny._0001_ ),
    .Q_N(_0103_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.imem_stb_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[1]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1439),
    .D(\i_exotiny._0002_ ),
    .Q_N(_0041_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1440),
    .D(\i_exotiny._0000_ ),
    .Q_N(_5379_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1441),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.c_o ),
    .Q_N(_4332_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1442),
    .D(_1184_),
    .Q_N(_4331_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1443),
    .D(_1185_),
    .Q_N(_4330_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1444),
    .D(_1186_),
    .Q_N(_0045_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1445),
    .D(_1187_),
    .Q_N(_0051_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1446),
    .D(_1188_),
    .Q_N(_0076_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1447),
    .D(_1189_),
    .Q_N(_0074_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1448),
    .D(_1190_),
    .Q_N(_0106_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1449),
    .D(_1191_),
    .Q_N(_0072_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1450),
    .D(_1192_),
    .Q_N(_0070_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15]$_SDFFE_PN0N_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1451),
    .D(_1193_),
    .Q_N(_0068_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1452),
    .D(_1194_),
    .Q_N(_4329_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1453),
    .D(_1195_),
    .Q_N(_0066_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1454),
    .D(_1196_),
    .Q_N(_0063_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19]$_SDFFE_PN0N_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1455),
    .D(_1197_),
    .Q_N(_4328_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1456),
    .D(_1198_),
    .Q_N(_0102_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1457),
    .D(_1199_),
    .Q_N(_0059_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1458),
    .D(_1200_),
    .Q_N(_0056_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23]$_SDFFE_PN0N_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1459),
    .D(_1201_),
    .Q_N(_0053_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1460),
    .D(_1202_),
    .Q_N(_4327_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1461),
    .D(_1203_),
    .Q_N(_4326_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1462),
    .D(_1204_),
    .Q_N(_4325_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1463),
    .D(_1205_),
    .Q_N(_4324_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[28]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1464),
    .D(_1206_),
    .Q_N(_4323_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1465),
    .D(_1207_),
    .Q_N(_4322_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1466),
    .D(_1208_),
    .Q_N(_4321_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31]$_SDFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1467),
    .D(_1209_),
    .Q_N(_4320_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1468),
    .D(_1210_),
    .Q_N(_0113_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1469),
    .D(_1211_),
    .Q_N(_0085_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6]$_SDFFE_PN0N_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1470),
    .D(_1212_),
    .Q_N(_0083_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1471),
    .D(_1213_),
    .Q_N(_0081_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1472),
    .D(_1214_),
    .Q_N(_0109_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1473),
    .D(_1215_),
    .Q_N(_0078_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1474),
    .D(_1216_),
    .Q_N(_0077_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1475),
    .D(_1217_),
    .Q_N(_0075_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1476),
    .D(_1218_),
    .Q_N(_0107_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1477),
    .D(_1219_),
    .Q_N(_0073_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1478),
    .D(_1220_),
    .Q_N(_0071_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1479),
    .D(_1221_),
    .Q_N(_0069_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1480),
    .D(_1222_),
    .Q_N(_4319_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1481),
    .D(_1223_),
    .Q_N(_0067_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1482),
    .D(_1224_),
    .Q_N(_0064_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1483),
    .D(_1225_),
    .Q_N(_4318_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1484),
    .D(_1226_),
    .Q_N(_0101_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1485),
    .D(_1227_),
    .Q_N(_0060_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1486),
    .D(_1228_),
    .Q_N(_0057_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1487),
    .D(_1229_),
    .Q_N(_0054_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1488),
    .D(_1230_),
    .Q_N(_4317_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1489),
    .D(_1231_),
    .Q_N(_4316_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1490),
    .D(_1232_),
    .Q_N(_4315_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1491),
    .D(_1233_),
    .Q_N(_4314_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1492),
    .D(_1234_),
    .Q_N(_4313_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1493),
    .D(_1235_),
    .Q_N(_4312_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1494),
    .D(_1236_),
    .Q_N(_0088_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1495),
    .D(_1237_),
    .Q_N(_4311_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1496),
    .D(_1238_),
    .Q_N(_4310_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1497),
    .D(_1239_),
    .Q_N(_0087_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1498),
    .D(_1240_),
    .Q_N(_0112_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1499),
    .D(_1241_),
    .Q_N(_0086_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1500),
    .D(_1242_),
    .Q_N(_0031_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[7]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1501),
    .D(_1243_),
    .Q_N(_0024_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[8]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1502),
    .D(_1244_),
    .Q_N(_0110_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1503),
    .D(_1245_),
    .Q_N(_0079_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1504),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[0] ),
    .Q_N(_0044_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1505),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[1] ),
    .Q_N(_5380_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2]$_DFF_P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1506),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[2] ),
    .Q_N(_5381_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3]$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1507),
    .D(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_n[3] ),
    .Q_N(_4309_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1508),
    .D(_1246_),
    .Q_N(_0008_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[10]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1509),
    .D(_1247_),
    .Q_N(_4308_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1510),
    .D(_1248_),
    .Q_N(_4307_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1511),
    .D(_1249_),
    .Q_N(_4306_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1512),
    .D(_1250_),
    .Q_N(_4305_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1513),
    .D(_1251_),
    .Q_N(_4304_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1514),
    .D(_1252_),
    .Q_N(_4303_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[16]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1515),
    .D(_1253_),
    .Q_N(_4302_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[17]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1516),
    .D(_1254_),
    .Q_N(_4301_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1517),
    .D(_1255_),
    .Q_N(_4300_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1518),
    .D(_1256_),
    .Q_N(_4299_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1519),
    .D(_1257_),
    .Q_N(_0007_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1520),
    .D(_1258_),
    .Q_N(_4298_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1521),
    .D(_1259_),
    .Q_N(_4297_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1522),
    .D(_1260_),
    .Q_N(_4296_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1523),
    .D(_1261_),
    .Q_N(_4295_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1524),
    .D(_1262_),
    .Q_N(_4294_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1525),
    .D(_1263_),
    .Q_N(_4293_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1526),
    .D(_1264_),
    .Q_N(_4292_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1527),
    .D(_1265_),
    .Q_N(_4291_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1528),
    .D(_1266_),
    .Q_N(_4290_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1529),
    .D(_1267_),
    .Q_N(_4289_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1530),
    .D(_1268_),
    .Q_N(_0006_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1531),
    .D(_1269_),
    .Q_N(_4288_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1532),
    .D(_1270_),
    .Q_N(_4287_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1533),
    .D(_1271_),
    .Q_N(_0004_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1534),
    .D(_1272_),
    .Q_N(_0035_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[5]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1535),
    .D(_1273_),
    .Q_N(_0034_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1536),
    .D(_1274_),
    .Q_N(_0033_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1537),
    .D(_1275_),
    .Q_N(_4286_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1538),
    .D(_1276_),
    .Q_N(_4285_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1539),
    .D(_1277_),
    .Q_N(_4284_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1540),
    .D(_1278_),
    .Q_N(_4283_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1541),
    .D(_1279_),
    .Q_N(_4282_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1542),
    .D(_1280_),
    .Q_N(_4281_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1543),
    .D(_1281_),
    .Q_N(_0036_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1544),
    .D(_1282_),
    .Q_N(_4280_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.cnt_r[0]$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1545),
    .D(_1283_),
    .Q_N(_0098_),
    .Q(\i_exotiny.i_wb_qspi_mem.cnt_r[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.cnt_r[1]$_SDFF_PN0_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1546),
    .D(_1284_),
    .Q_N(_0005_),
    .Q(\i_exotiny.i_wb_qspi_mem.cnt_r[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.cnt_r[2]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1547),
    .D(_1285_),
    .Q_N(_0097_),
    .Q(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.crm_r$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1548),
    .D(_1286_),
    .Q_N(_5382_),
    .Q(\i_exotiny.i_wb_qspi_mem.crm_r ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[0]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1549),
    .D(\i_exotiny._0006_ ),
    .Q_N(_0001_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[1]$_DFF_P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1550),
    .D(\i_exotiny._0007_ ),
    .Q_N(_5383_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[2]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1551),
    .D(\i_exotiny._0008_ ),
    .Q_N(_0104_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1552),
    .D(\i_exotiny._0009_ ),
    .Q_N(_5384_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[4]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1553),
    .D(\i_exotiny._0010_ ),
    .Q_N(_0099_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[5]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1554),
    .D(\i_exotiny._0011_ ),
    .Q_N(_5385_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.state_r_reg[6]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1555),
    .D(\i_exotiny._0012_ ),
    .Q_N(_5386_),
    .Q(\i_exotiny.i_wb_qspi_mem.state_r_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_qspi_mem.wb_mem_ack_o$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1556),
    .D(\i_exotiny._0013_ ),
    .Q_N(_4279_),
    .Q(\i_exotiny.i_wb_qspi_mem.wb_mem_ack_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_auto_cs_o$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1557),
    .D(_1287_),
    .Q_N(_4278_),
    .Q(\i_exotiny.i_wb_regs.spi_auto_cs_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_cpol_o$_SDFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1558),
    .D(_1288_),
    .Q_N(_4277_),
    .Q(\i_exotiny.i_wb_regs.spi_cpol_o ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_presc_o[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1559),
    .D(_1289_),
    .Q_N(_0095_),
    .Q(\i_exotiny.i_wb_regs.spi_presc_o[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_presc_o[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1560),
    .D(_1290_),
    .Q_N(_0094_),
    .Q(\i_exotiny.i_wb_regs.spi_presc_o[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_presc_o[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1561),
    .D(_1291_),
    .Q_N(_0093_),
    .Q(\i_exotiny.i_wb_regs.spi_presc_o[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_presc_o[3]$_SDFFE_PN1P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1562),
    .D(_1292_),
    .Q_N(_5387_),
    .Q(\i_exotiny.i_wb_regs.spi_presc_o[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_rdy_i$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1563),
    .D(\i_exotiny._0014_ ),
    .Q_N(_4276_),
    .Q(\i_exotiny.i_wb_regs.spi_rdy_i ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_size_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1564),
    .D(_1293_),
    .Q_N(_0003_),
    .Q(\i_exotiny.i_wb_regs.spi_size_o[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_regs.spi_size_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1565),
    .D(_1294_),
    .Q_N(_4275_),
    .Q(\i_exotiny.i_wb_regs.spi_size_o[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1566),
    .D(_1295_),
    .Q_N(\i_exotiny._2358_[0] ),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1567),
    .D(_1296_),
    .Q_N(_4274_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1568),
    .D(_1297_),
    .Q_N(_0050_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1569),
    .D(_1298_),
    .Q_N(_4273_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1570),
    .D(_1299_),
    .Q_N(_4272_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1571),
    .D(_1300_),
    .Q_N(_4271_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_hbit_r[6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1572),
    .D(_1301_),
    .Q_N(_5388_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[0]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1573),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[0] ),
    .Q_N(_0096_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[1]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1574),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[1] ),
    .Q_N(_5389_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[2]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1575),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[2] ),
    .Q_N(_5390_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[3]$_DFF_P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1576),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[3] ),
    .Q_N(_5391_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[4]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1577),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[4] ),
    .Q_N(_5392_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[5]$_DFF_P_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1578),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[5] ),
    .Q_N(_5393_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.cnt_presc_r[6]$_DFF_P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1579),
    .D(\i_exotiny.i_wb_spi.cnt_presc_n[6] ),
    .Q_N(_4270_),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1580),
    .D(_1302_),
    .Q_N(_4269_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[10]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1581),
    .D(_1303_),
    .Q_N(_4268_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[11]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1582),
    .D(_1304_),
    .Q_N(_4267_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[12]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1583),
    .D(_1305_),
    .Q_N(_4266_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1584),
    .D(_1306_),
    .Q_N(_4265_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[14]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1585),
    .D(_1307_),
    .Q_N(_4264_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[15]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1586),
    .D(_1308_),
    .Q_N(_4263_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[16]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1587),
    .D(_1309_),
    .Q_N(_4262_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[17]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1588),
    .D(_1310_),
    .Q_N(_4261_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[18]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1589),
    .D(_1311_),
    .Q_N(_4260_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[19]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1590),
    .D(_1312_),
    .Q_N(_4259_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1591),
    .D(_1313_),
    .Q_N(_4258_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[20]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1592),
    .D(_1314_),
    .Q_N(_4257_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[21]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1593),
    .D(_1315_),
    .Q_N(_4256_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[22]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1594),
    .D(_1316_),
    .Q_N(_4255_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[23]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1595),
    .D(_1317_),
    .Q_N(_4254_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[24]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1596),
    .D(_1318_),
    .Q_N(_4253_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[25]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1597),
    .D(_1319_),
    .Q_N(_4252_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[26]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1598),
    .D(_1320_),
    .Q_N(_4251_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[27]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1599),
    .D(_1321_),
    .Q_N(_4250_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1600),
    .D(_1322_),
    .Q_N(_4249_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1601),
    .D(_1323_),
    .Q_N(_4248_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1602),
    .D(_1324_),
    .Q_N(_4247_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1603),
    .D(_1325_),
    .Q_N(_4246_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[31]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1604),
    .D(_1326_),
    .Q_N(_4245_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[31] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[3]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1605),
    .D(_1327_),
    .Q_N(_4244_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[4]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1606),
    .D(_1328_),
    .Q_N(_4243_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[5]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1607),
    .D(_1329_),
    .Q_N(_4242_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[6]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1608),
    .D(_1330_),
    .Q_N(_4241_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[7]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1609),
    .D(_1331_),
    .Q_N(_4240_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[8]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1610),
    .D(_1332_),
    .Q_N(_4239_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_rx_r[9]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1611),
    .D(_1333_),
    .Q_N(_4238_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1612),
    .D(_1334_),
    .Q_N(_4237_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[0] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1613),
    .D(_1335_),
    .Q_N(_4236_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[10] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1614),
    .D(_1336_),
    .Q_N(_4235_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[11] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[12]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1615),
    .D(_1337_),
    .Q_N(_4234_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[12] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[13]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1616),
    .D(_1338_),
    .Q_N(_4233_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[13] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[14]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1617),
    .D(_1339_),
    .Q_N(_4232_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[14] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[15]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1618),
    .D(_1340_),
    .Q_N(_4231_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[15] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[16]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1619),
    .D(_1341_),
    .Q_N(_4230_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[16] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[17]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1620),
    .D(_1342_),
    .Q_N(_4229_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[17] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[18]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1621),
    .D(_1343_),
    .Q_N(_4228_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[18] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[19]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1622),
    .D(_1344_),
    .Q_N(_4227_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[19] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[1]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1623),
    .D(_1345_),
    .Q_N(_4226_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[20]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1624),
    .D(_1346_),
    .Q_N(_4225_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[20] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[21]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1625),
    .D(_1347_),
    .Q_N(_4224_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[21] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[22]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1626),
    .D(_1348_),
    .Q_N(_4223_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[22] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[23]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1627),
    .D(_1349_),
    .Q_N(_4222_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[23] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[24]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1628),
    .D(_1350_),
    .Q_N(_4221_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[24] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1629),
    .D(_1351_),
    .Q_N(_4220_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[25] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1630),
    .D(_1352_),
    .Q_N(_4219_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[26] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1631),
    .D(_1353_),
    .Q_N(_4218_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[27] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[28]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1632),
    .D(_1354_),
    .Q_N(_4217_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[28] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[29]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1633),
    .D(_1355_),
    .Q_N(_4216_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[29] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1634),
    .D(_1356_),
    .Q_N(_4215_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[2] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[30]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1635),
    .D(_1357_),
    .Q_N(_4214_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[30] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1636),
    .D(_1358_),
    .Q_N(_4213_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[3] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[4]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1637),
    .D(_1359_),
    .Q_N(_4212_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[4] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[5]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1638),
    .D(_1360_),
    .Q_N(_4211_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[5] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[6]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1639),
    .D(_1361_),
    .Q_N(_4210_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[6] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1640),
    .D(_1362_),
    .Q_N(_4209_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[7] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[8]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1641),
    .D(_1363_),
    .Q_N(_4208_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[8] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.dat_tx_r_reg[9]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1642),
    .D(_1364_),
    .Q_N(_5394_),
    .Q(\i_exotiny.i_wb_spi.dat_tx_r_reg[9] ));
 sg13g2_dfrbp_1 \i_exotiny.i_wb_spi.state_r_reg[1]$_DFF_P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1643),
    .D(\i_exotiny._0015_ ),
    .Q_N(_0092_),
    .Q(\i_exotiny.i_wb_spi.state_r_reg[1] ));
 sg13g2_dfrbp_1 \i_exotiny.spi_sck_o$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1644),
    .D(_1365_),
    .Q_N(_0002_),
    .Q(\i_exotiny.spi_sck_o ));
 sg13g2_dfrbp_1 \i_exotiny.spi_sdo_o$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1645),
    .D(_1366_),
    .Q_N(_4207_),
    .Q(\i_exotiny.spi_sdo_o ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[4]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[5]),
    .X(net12));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_oe[0]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_oe[1]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_oe[2]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_oe[3]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_oe[4]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[5]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[6]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[0]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uo_out[1]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uo_out[2]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uo_out[3]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uo_out[4]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uo_out[5]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uo_out[6]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout35 (.A(_3559_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_3423_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_3347_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_3278_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_3244_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_3223_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_3556_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_3420_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_3238_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_3540_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_3326_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_3234_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_3348_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_3258_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_3229_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2288_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2283_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2390_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2743_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2715_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2702_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2633_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2781_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_2701_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_4015_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_3007_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_3002_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_2973_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2968_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_2939_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_2937_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2936_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_4005_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_2910_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2762_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2666_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2630_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_1685_));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_1684_));
 sg13g2_buf_2 fanout74 (.A(_1496_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1493_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_3781_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2763_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2706_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_2695_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_2447_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_4168_),
    .X(net81));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(_2934_));
 sg13g2_buf_4 fanout83 (.X(net83),
    .A(_2933_));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(_2932_));
 sg13g2_buf_2 fanout85 (.A(_2705_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_2109_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1642_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1630_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1580_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1560_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1539_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1525_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_3682_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_2728_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_2717_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_2294_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_1994_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_1613_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_3734_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1507_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_4022_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_3713_),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(_3585_));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_3562_));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_3548_));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(_3545_));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(_3535_));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(_3534_));
 sg13g2_buf_4 fanout109 (.X(net109),
    .A(_3533_));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_3524_));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(_3523_));
 sg13g2_buf_4 fanout112 (.X(net112),
    .A(_3522_));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(_3512_));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_3510_));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_3495_));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_3494_));
 sg13g2_buf_4 fanout117 (.X(net117),
    .A(_3493_));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(_3481_));
 sg13g2_buf_4 fanout119 (.X(net119),
    .A(_3480_));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_3465_));
 sg13g2_buf_4 fanout121 (.X(net121),
    .A(_3464_));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(_3463_));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_3453_));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(_3452_));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(_3450_));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(_3438_));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_3437_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_3428_));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_3427_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_3426_));
 sg13g2_buf_4 fanout131 (.X(net131),
    .A(_3407_));
 sg13g2_buf_4 fanout132 (.X(net132),
    .A(_3402_));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(_3395_));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_3394_));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(_3390_));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_3384_));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(_3383_));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(_3365_));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(_3362_));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(_3346_));
 sg13g2_buf_4 fanout141 (.X(net141),
    .A(_3344_));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_3343_));
 sg13g2_buf_4 fanout143 (.X(net143),
    .A(_3332_));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(_3331_));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(_3318_));
 sg13g2_buf_4 fanout146 (.X(net146),
    .A(_3317_));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(_3316_));
 sg13g2_buf_4 fanout148 (.X(net148),
    .A(_3298_));
 sg13g2_buf_4 fanout149 (.X(net149),
    .A(_3295_));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(_3293_));
 sg13g2_buf_4 fanout151 (.X(net151),
    .A(_3277_));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_3276_));
 sg13g2_buf_2 fanout153 (.A(_3257_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_3253_),
    .X(net154));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_3250_));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_3249_));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(_3247_));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_3124_));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_3123_));
 sg13g2_buf_4 fanout160 (.X(net160),
    .A(_3116_));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(_3106_));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_3105_));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_3095_));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_3087_));
 sg13g2_buf_4 fanout165 (.X(net165),
    .A(_3084_));
 sg13g2_buf_2 fanout166 (.A(_3080_),
    .X(net166));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_3076_));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_3071_));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(_3064_));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_3059_));
 sg13g2_buf_2 fanout171 (.A(_3058_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_3055_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_2001_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_1843_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_1461_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_3830_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_3823_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_3807_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_3800_),
    .X(net179));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_3662_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_3653_));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(_3652_));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_3651_));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_3642_));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_3641_));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(_3640_));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_3631_));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_3630_));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(_3621_));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_3620_));
 sg13g2_buf_4 fanout191 (.X(net191),
    .A(_3619_));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_3610_));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_3609_));
 sg13g2_buf_4 fanout194 (.X(net194),
    .A(_3600_));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(_3598_));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_3597_));
 sg13g2_buf_2 fanout197 (.A(_3591_),
    .X(net197));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_3587_));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(_3586_));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_3576_));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_3575_));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_3565_));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_3564_));
 sg13g2_buf_2 fanout204 (.A(_3520_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_3474_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_3399_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_3380_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_3279_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_3265_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_3255_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_3252_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_3248_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_3245_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_3224_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_3113_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_3104_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_3089_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_3068_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_3056_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_3054_),
    .X(net220));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(_2707_));
 sg13g2_buf_2 fanout222 (.A(_1792_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_1710_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_1694_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_1567_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_1550_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_1526_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_1401_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_1394_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_1383_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_4033_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_3672_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_3321_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_3286_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_3133_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_3103_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_3053_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_2755_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_2673_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_2671_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_2324_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_2067_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_1986_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_1703_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_1693_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_1403_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_1400_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_1382_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_4016_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_3802_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_3786_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_3755_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_3671_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_3008_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_2974_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_2940_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_2672_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_2244_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_2019_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_1915_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_1914_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_1584_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_1556_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_1424_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_1413_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_3901_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_3825_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_3742_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_3696_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_3685_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_3566_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_3484_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_3351_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_3127_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_2880_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_2270_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_2120_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_2078_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_2018_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_1924_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_1913_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_1891_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_1436_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_1432_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_1427_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_1423_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_1416_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_1412_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_1390_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_1369_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_4159_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_4032_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_3914_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_3757_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_3741_),
    .X(net295));
 sg13g2_buf_1 fanout296 (.A(_3015_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_2981_),
    .X(net297));
 sg13g2_buf_1 fanout298 (.A(_2947_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_2905_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_2010_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_2004_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_1921_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_1896_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_1890_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_1797_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_1714_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_1495_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_1481_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_1451_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_1435_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_1426_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_1422_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_1419_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_1415_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_1411_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_1406_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_1396_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_1389_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_1368_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_3718_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_2878_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_1764_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_1757_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_1688_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_1515_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_1504_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_1500_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_1498_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_1485_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_1477_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_1446_),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(_1441_),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(_1438_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_1405_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_1377_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_1374_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_1371_),
    .X(net337));
 sg13g2_tielo _9559__338 (.L_LO(net338));
 sg13g2_tielo _9563__339 (.L_LO(net339));
 sg13g2_tiehi \i_exotiny.gpo_o[1]$_SDFFE_PN0P__341  (.L_HI(net341));
 sg13g2_tiehi \i_exotiny.gpo_o[2]$_SDFFE_PN0P__342  (.L_HI(net342));
 sg13g2_tiehi \i_exotiny.gpo_o[3]$_SDFFE_PN0P__343  (.L_HI(net343));
 sg13g2_tiehi \i_exotiny.gpo_o[4]$_SDFFE_PN0P__344  (.L_HI(net344));
 sg13g2_tiehi \i_exotiny.gpo_o[5]$_SDFFE_PN0P__345  (.L_HI(net345));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[0]$_DFFE_PN__346  (.L_HI(net346));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[1]$_DFFE_PN__347  (.L_HI(net347));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[2]$_DFFE_PN__348  (.L_HI(net348));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].dout[3]$_DFFE_PN__349  (.L_HI(net349));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[0]$_DFFE_PN__350  (.L_HI(net350));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[1]$_DFFE_PN__351  (.L_HI(net351));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[2]$_DFFE_PN__352  (.L_HI(net352));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].dout[3]$_DFFE_PN__353  (.L_HI(net353));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[0]$_DFFE_PN__354  (.L_HI(net354));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[1]$_DFFE_PN__355  (.L_HI(net355));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[2]$_DFFE_PN__356  (.L_HI(net356));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].dout[3]$_DFFE_PN__357  (.L_HI(net357));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[0]$_DFFE_PN__358  (.L_HI(net358));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[1]$_DFFE_PN__359  (.L_HI(net359));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[2]$_DFFE_PN__360  (.L_HI(net360));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].dout[3]$_DFFE_PN__361  (.L_HI(net361));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[0]$_DFFE_PN__362  (.L_HI(net362));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[1]$_DFFE_PN__363  (.L_HI(net363));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[2]$_DFFE_PN__364  (.L_HI(net364));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].dout[3]$_DFFE_PN__365  (.L_HI(net365));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[0]$_DFFE_PN__366  (.L_HI(net366));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[1]$_DFFE_PN__367  (.L_HI(net367));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[2]$_DFFE_PN__368  (.L_HI(net368));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].dout[3]$_DFFE_PN__369  (.L_HI(net369));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[0]$_DFFE_PN__370  (.L_HI(net370));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[1]$_DFFE_PN__371  (.L_HI(net371));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[2]$_DFFE_PN__372  (.L_HI(net372));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].dout[3]$_DFFE_PN__373  (.L_HI(net373));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[0]$_DFFE_PN__374  (.L_HI(net374));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[1]$_DFFE_PN__375  (.L_HI(net375));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[2]$_DFFE_PN__376  (.L_HI(net376));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].dout[3]$_DFFE_PN__377  (.L_HI(net377));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[0]$_DFFE_PN__378  (.L_HI(net378));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[1]$_DFFE_PN__379  (.L_HI(net379));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[2]$_DFFE_PN__380  (.L_HI(net380));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].dout[3]$_DFFE_PN__381  (.L_HI(net381));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[0]$_DFFE_PN__382  (.L_HI(net382));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[1]$_DFFE_PN__383  (.L_HI(net383));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[2]$_DFFE_PN__384  (.L_HI(net384));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].dout[3]$_DFFE_PN__385  (.L_HI(net385));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[0]$_DFFE_PN__386  (.L_HI(net386));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[1]$_DFFE_PN__387  (.L_HI(net387));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[2]$_DFFE_PN__388  (.L_HI(net388));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].dout[3]$_DFFE_PN__389  (.L_HI(net389));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[0]$_DFFE_PN__390  (.L_HI(net390));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[1]$_DFFE_PN__391  (.L_HI(net391));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[2]$_DFFE_PN__392  (.L_HI(net392));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].dout[3]$_DFFE_PN__393  (.L_HI(net393));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[0]$_DFFE_PN__394  (.L_HI(net394));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[1]$_DFFE_PN__395  (.L_HI(net395));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[2]$_DFFE_PN__396  (.L_HI(net396));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].dout[3]$_DFFE_PN__397  (.L_HI(net397));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[0]$_DFFE_PN__398  (.L_HI(net398));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[1]$_DFFE_PN__399  (.L_HI(net399));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[2]$_DFFE_PN__400  (.L_HI(net400));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].dout[3]$_DFFE_PN__401  (.L_HI(net401));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[0]$_DFFE_PN__402  (.L_HI(net402));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[1]$_DFFE_PN__403  (.L_HI(net403));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[2]$_DFFE_PN__404  (.L_HI(net404));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].dout[3]$_DFFE_PN__405  (.L_HI(net405));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[0]$_DFFE_PN__406  (.L_HI(net406));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[1]$_DFFE_PN__407  (.L_HI(net407));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[2]$_DFFE_PN__408  (.L_HI(net408));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].dout[3]$_DFFE_PN__409  (.L_HI(net409));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[0]$_DFFE_PN__410  (.L_HI(net410));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[1]$_DFFE_PN__411  (.L_HI(net411));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[2]$_DFFE_PN__412  (.L_HI(net412));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].dout[3]$_DFFE_PN__413  (.L_HI(net413));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[0]$_DFFE_PN__414  (.L_HI(net414));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[1]$_DFFE_PN__415  (.L_HI(net415));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[2]$_DFFE_PN__416  (.L_HI(net416));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].dout[3]$_DFFE_PN__417  (.L_HI(net417));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[0]$_DFFE_PN__418  (.L_HI(net418));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[1]$_DFFE_PN__419  (.L_HI(net419));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[2]$_DFFE_PN__420  (.L_HI(net420));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].dout[3]$_DFFE_PN__421  (.L_HI(net421));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[0]$_DFFE_PN__422  (.L_HI(net422));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[1]$_DFFE_PN__423  (.L_HI(net423));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[2]$_DFFE_PN__424  (.L_HI(net424));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].dout[3]$_DFFE_PN__425  (.L_HI(net425));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[0]$_DFFE_PN__426  (.L_HI(net426));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[1]$_DFFE_PN__427  (.L_HI(net427));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[2]$_DFFE_PN__428  (.L_HI(net428));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].dout[3]$_DFFE_PN__429  (.L_HI(net429));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[0]$_DFFE_PN__430  (.L_HI(net430));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[1]$_DFFE_PN__431  (.L_HI(net431));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[2]$_DFFE_PN__432  (.L_HI(net432));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].dout[3]$_DFFE_PN__433  (.L_HI(net433));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[0]$_DFFE_PN__434  (.L_HI(net434));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[1]$_DFFE_PN__435  (.L_HI(net435));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[2]$_DFFE_PN__436  (.L_HI(net436));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].dout[3]$_DFFE_PN__437  (.L_HI(net437));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[0]$_DFFE_PN__438  (.L_HI(net438));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[1]$_DFFE_PN__439  (.L_HI(net439));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[2]$_DFFE_PN__440  (.L_HI(net440));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].dout[3]$_DFFE_PN__441  (.L_HI(net441));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[0]$_DFFE_PN__442  (.L_HI(net442));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[1]$_DFFE_PN__443  (.L_HI(net443));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[2]$_DFFE_PN__444  (.L_HI(net444));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].dout[3]$_DFFE_PN__445  (.L_HI(net445));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[0]$_DFFE_PN__446  (.L_HI(net446));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[1]$_DFFE_PN__447  (.L_HI(net447));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[2]$_DFFE_PN__448  (.L_HI(net448));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].dout[3]$_DFFE_PN__449  (.L_HI(net449));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[0]$_DFFE_PN__450  (.L_HI(net450));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[1]$_DFFE_PN__451  (.L_HI(net451));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[2]$_DFFE_PN__452  (.L_HI(net452));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].dout[3]$_DFFE_PN__453  (.L_HI(net453));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[0]$_DFFE_PN__454  (.L_HI(net454));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[1]$_DFFE_PN__455  (.L_HI(net455));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[2]$_DFFE_PN__456  (.L_HI(net456));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].dout[3]$_DFFE_PN__457  (.L_HI(net457));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[0]$_DFFE_PN__458  (.L_HI(net458));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[1]$_DFFE_PN__459  (.L_HI(net459));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[2]$_DFFE_PN__460  (.L_HI(net460));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].dout[3]$_DFFE_PN__461  (.L_HI(net461));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[0]$_DFFE_PN__462  (.L_HI(net462));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[1]$_DFFE_PN__463  (.L_HI(net463));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[2]$_DFFE_PN__464  (.L_HI(net464));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].dout[3]$_DFFE_PN__465  (.L_HI(net465));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[0]$_DFFE_PN__466  (.L_HI(net466));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[1]$_DFFE_PN__467  (.L_HI(net467));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[2]$_DFFE_PN__468  (.L_HI(net468));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].dout[3]$_DFFE_PN__469  (.L_HI(net469));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[10]$_DFFE_PN__470  (.L_HI(net470));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[11]$_DFFE_PN__471  (.L_HI(net471));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[12]$_DFFE_PN__472  (.L_HI(net472));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[13]$_DFFE_PN__473  (.L_HI(net473));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[14]$_DFFE_PN__474  (.L_HI(net474));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[15]$_DFFE_PN__475  (.L_HI(net475));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[16]$_DFFE_PN__476  (.L_HI(net476));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[17]$_DFFE_PN__477  (.L_HI(net477));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[18]$_DFFE_PN__478  (.L_HI(net478));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[19]$_DFFE_PN__479  (.L_HI(net479));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[20]$_DFFE_PN__480  (.L_HI(net480));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[21]$_DFFE_PN__481  (.L_HI(net481));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[22]$_DFFE_PN__482  (.L_HI(net482));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[23]$_DFFE_PN__483  (.L_HI(net483));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[24]$_DFFE_PN__484  (.L_HI(net484));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[25]$_DFFE_PN__485  (.L_HI(net485));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[26]$_DFFE_PN__486  (.L_HI(net486));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[27]$_DFFE_PN__487  (.L_HI(net487));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[28]$_DFFE_PN__488  (.L_HI(net488));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[29]$_DFFE_PN__489  (.L_HI(net489));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[30]$_DFFE_PN__490  (.L_HI(net490));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[31]$_DFFE_PN__491  (.L_HI(net491));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[4]$_DFFE_PN__492  (.L_HI(net492));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[5]$_DFFE_PN__493  (.L_HI(net493));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[6]$_DFFE_PN__494  (.L_HI(net494));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[7]$_DFFE_PN__495  (.L_HI(net495));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[8]$_DFFE_PN__496  (.L_HI(net496));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[10].i_reg.reg_r[9]$_DFFE_PN__497  (.L_HI(net497));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[10]$_DFFE_PN__498  (.L_HI(net498));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[11]$_DFFE_PN__499  (.L_HI(net499));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[12]$_DFFE_PN__500  (.L_HI(net500));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[13]$_DFFE_PN__501  (.L_HI(net501));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[14]$_DFFE_PN__502  (.L_HI(net502));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[15]$_DFFE_PN__503  (.L_HI(net503));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[16]$_DFFE_PN__504  (.L_HI(net504));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[17]$_DFFE_PN__505  (.L_HI(net505));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[18]$_DFFE_PN__506  (.L_HI(net506));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[19]$_DFFE_PN__507  (.L_HI(net507));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[20]$_DFFE_PN__508  (.L_HI(net508));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[21]$_DFFE_PN__509  (.L_HI(net509));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[22]$_DFFE_PN__510  (.L_HI(net510));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[23]$_DFFE_PN__511  (.L_HI(net511));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[24]$_DFFE_PN__512  (.L_HI(net512));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[25]$_DFFE_PN__513  (.L_HI(net513));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[26]$_DFFE_PN__514  (.L_HI(net514));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[27]$_DFFE_PN__515  (.L_HI(net515));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[28]$_DFFE_PN__516  (.L_HI(net516));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[29]$_DFFE_PN__517  (.L_HI(net517));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[30]$_DFFE_PN__518  (.L_HI(net518));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[31]$_DFFE_PN__519  (.L_HI(net519));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[4]$_DFFE_PN__520  (.L_HI(net520));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[5]$_DFFE_PN__521  (.L_HI(net521));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[6]$_DFFE_PN__522  (.L_HI(net522));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[7]$_DFFE_PN__523  (.L_HI(net523));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[8]$_DFFE_PN__524  (.L_HI(net524));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[11].i_reg.reg_r[9]$_DFFE_PN__525  (.L_HI(net525));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[10]$_DFFE_PN__526  (.L_HI(net526));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[11]$_DFFE_PN__527  (.L_HI(net527));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[12]$_DFFE_PN__528  (.L_HI(net528));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[13]$_DFFE_PN__529  (.L_HI(net529));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[14]$_DFFE_PN__530  (.L_HI(net530));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[15]$_DFFE_PN__531  (.L_HI(net531));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[16]$_DFFE_PN__532  (.L_HI(net532));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[17]$_DFFE_PN__533  (.L_HI(net533));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[18]$_DFFE_PN__534  (.L_HI(net534));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[19]$_DFFE_PN__535  (.L_HI(net535));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[20]$_DFFE_PN__536  (.L_HI(net536));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[21]$_DFFE_PN__537  (.L_HI(net537));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[22]$_DFFE_PN__538  (.L_HI(net538));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[23]$_DFFE_PN__539  (.L_HI(net539));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[24]$_DFFE_PN__540  (.L_HI(net540));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[25]$_DFFE_PN__541  (.L_HI(net541));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[26]$_DFFE_PN__542  (.L_HI(net542));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[27]$_DFFE_PN__543  (.L_HI(net543));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[28]$_DFFE_PN__544  (.L_HI(net544));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[29]$_DFFE_PN__545  (.L_HI(net545));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[30]$_DFFE_PN__546  (.L_HI(net546));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[31]$_DFFE_PN__547  (.L_HI(net547));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[4]$_DFFE_PN__548  (.L_HI(net548));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[5]$_DFFE_PN__549  (.L_HI(net549));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[6]$_DFFE_PN__550  (.L_HI(net550));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[7]$_DFFE_PN__551  (.L_HI(net551));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[8]$_DFFE_PN__552  (.L_HI(net552));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[12].i_reg.reg_r[9]$_DFFE_PN__553  (.L_HI(net553));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[10]$_DFFE_PN__554  (.L_HI(net554));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[11]$_DFFE_PN__555  (.L_HI(net555));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[12]$_DFFE_PN__556  (.L_HI(net556));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[13]$_DFFE_PN__557  (.L_HI(net557));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[14]$_DFFE_PN__558  (.L_HI(net558));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[15]$_DFFE_PN__559  (.L_HI(net559));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[16]$_DFFE_PN__560  (.L_HI(net560));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[17]$_DFFE_PN__561  (.L_HI(net561));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[18]$_DFFE_PN__562  (.L_HI(net562));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[19]$_DFFE_PN__563  (.L_HI(net563));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[20]$_DFFE_PN__564  (.L_HI(net564));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[21]$_DFFE_PN__565  (.L_HI(net565));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[22]$_DFFE_PN__566  (.L_HI(net566));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[23]$_DFFE_PN__567  (.L_HI(net567));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[24]$_DFFE_PN__568  (.L_HI(net568));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[25]$_DFFE_PN__569  (.L_HI(net569));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[26]$_DFFE_PN__570  (.L_HI(net570));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[27]$_DFFE_PN__571  (.L_HI(net571));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[28]$_DFFE_PN__572  (.L_HI(net572));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[29]$_DFFE_PN__573  (.L_HI(net573));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[30]$_DFFE_PN__574  (.L_HI(net574));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[31]$_DFFE_PN__575  (.L_HI(net575));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[4]$_DFFE_PN__576  (.L_HI(net576));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[5]$_DFFE_PN__577  (.L_HI(net577));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[6]$_DFFE_PN__578  (.L_HI(net578));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[7]$_DFFE_PN__579  (.L_HI(net579));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[8]$_DFFE_PN__580  (.L_HI(net580));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[13].i_reg.reg_r[9]$_DFFE_PN__581  (.L_HI(net581));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[10]$_DFFE_PN__582  (.L_HI(net582));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[11]$_DFFE_PN__583  (.L_HI(net583));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[12]$_DFFE_PN__584  (.L_HI(net584));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[13]$_DFFE_PN__585  (.L_HI(net585));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[14]$_DFFE_PN__586  (.L_HI(net586));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[15]$_DFFE_PN__587  (.L_HI(net587));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[16]$_DFFE_PN__588  (.L_HI(net588));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[17]$_DFFE_PN__589  (.L_HI(net589));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[18]$_DFFE_PN__590  (.L_HI(net590));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[19]$_DFFE_PN__591  (.L_HI(net591));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[20]$_DFFE_PN__592  (.L_HI(net592));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[21]$_DFFE_PN__593  (.L_HI(net593));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[22]$_DFFE_PN__594  (.L_HI(net594));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[23]$_DFFE_PN__595  (.L_HI(net595));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[24]$_DFFE_PN__596  (.L_HI(net596));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[25]$_DFFE_PN__597  (.L_HI(net597));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[26]$_DFFE_PN__598  (.L_HI(net598));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[27]$_DFFE_PN__599  (.L_HI(net599));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[28]$_DFFE_PN__600  (.L_HI(net600));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[29]$_DFFE_PN__601  (.L_HI(net601));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[30]$_DFFE_PN__602  (.L_HI(net602));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[31]$_DFFE_PN__603  (.L_HI(net603));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[4]$_DFFE_PN__604  (.L_HI(net604));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[5]$_DFFE_PN__605  (.L_HI(net605));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[6]$_DFFE_PN__606  (.L_HI(net606));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[7]$_DFFE_PN__607  (.L_HI(net607));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[8]$_DFFE_PN__608  (.L_HI(net608));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[14].i_reg.reg_r[9]$_DFFE_PN__609  (.L_HI(net609));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[10]$_DFFE_PN__610  (.L_HI(net610));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[11]$_DFFE_PN__611  (.L_HI(net611));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[12]$_DFFE_PN__612  (.L_HI(net612));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[13]$_DFFE_PN__613  (.L_HI(net613));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[14]$_DFFE_PN__614  (.L_HI(net614));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[15]$_DFFE_PN__615  (.L_HI(net615));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[16]$_DFFE_PN__616  (.L_HI(net616));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[17]$_DFFE_PN__617  (.L_HI(net617));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[18]$_DFFE_PN__618  (.L_HI(net618));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[19]$_DFFE_PN__619  (.L_HI(net619));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[20]$_DFFE_PN__620  (.L_HI(net620));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[21]$_DFFE_PN__621  (.L_HI(net621));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[22]$_DFFE_PN__622  (.L_HI(net622));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[23]$_DFFE_PN__623  (.L_HI(net623));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[24]$_DFFE_PN__624  (.L_HI(net624));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[25]$_DFFE_PN__625  (.L_HI(net625));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[26]$_DFFE_PN__626  (.L_HI(net626));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[27]$_DFFE_PN__627  (.L_HI(net627));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[28]$_DFFE_PN__628  (.L_HI(net628));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[29]$_DFFE_PN__629  (.L_HI(net629));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[30]$_DFFE_PN__630  (.L_HI(net630));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[31]$_DFFE_PN__631  (.L_HI(net631));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[4]$_DFFE_PN__632  (.L_HI(net632));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[5]$_DFFE_PN__633  (.L_HI(net633));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[6]$_DFFE_PN__634  (.L_HI(net634));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[7]$_DFFE_PN__635  (.L_HI(net635));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[8]$_DFFE_PN__636  (.L_HI(net636));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[15].i_reg.reg_r[9]$_DFFE_PN__637  (.L_HI(net637));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[10]$_DFFE_PN__638  (.L_HI(net638));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[11]$_DFFE_PN__639  (.L_HI(net639));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[12]$_DFFE_PN__640  (.L_HI(net640));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[13]$_DFFE_PN__641  (.L_HI(net641));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[14]$_DFFE_PN__642  (.L_HI(net642));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[15]$_DFFE_PN__643  (.L_HI(net643));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[16]$_DFFE_PN__644  (.L_HI(net644));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[17]$_DFFE_PN__645  (.L_HI(net645));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[18]$_DFFE_PN__646  (.L_HI(net646));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[19]$_DFFE_PN__647  (.L_HI(net647));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[20]$_DFFE_PN__648  (.L_HI(net648));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[21]$_DFFE_PN__649  (.L_HI(net649));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[22]$_DFFE_PN__650  (.L_HI(net650));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[23]$_DFFE_PN__651  (.L_HI(net651));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[24]$_DFFE_PN__652  (.L_HI(net652));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[25]$_DFFE_PN__653  (.L_HI(net653));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[26]$_DFFE_PN__654  (.L_HI(net654));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[27]$_DFFE_PN__655  (.L_HI(net655));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[28]$_DFFE_PN__656  (.L_HI(net656));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[29]$_DFFE_PN__657  (.L_HI(net657));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[30]$_DFFE_PN__658  (.L_HI(net658));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[31]$_DFFE_PN__659  (.L_HI(net659));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[4]$_DFFE_PN__660  (.L_HI(net660));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[5]$_DFFE_PN__661  (.L_HI(net661));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[6]$_DFFE_PN__662  (.L_HI(net662));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[7]$_DFFE_PN__663  (.L_HI(net663));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[8]$_DFFE_PN__664  (.L_HI(net664));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[16].i_reg.reg_r[9]$_DFFE_PN__665  (.L_HI(net665));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[10]$_DFFE_PN__666  (.L_HI(net666));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[11]$_DFFE_PN__667  (.L_HI(net667));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[12]$_DFFE_PN__668  (.L_HI(net668));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[13]$_DFFE_PN__669  (.L_HI(net669));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[14]$_DFFE_PN__670  (.L_HI(net670));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[15]$_DFFE_PN__671  (.L_HI(net671));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[16]$_DFFE_PN__672  (.L_HI(net672));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[17]$_DFFE_PN__673  (.L_HI(net673));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[18]$_DFFE_PN__674  (.L_HI(net674));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[19]$_DFFE_PN__675  (.L_HI(net675));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[20]$_DFFE_PN__676  (.L_HI(net676));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[21]$_DFFE_PN__677  (.L_HI(net677));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[22]$_DFFE_PN__678  (.L_HI(net678));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[23]$_DFFE_PN__679  (.L_HI(net679));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[24]$_DFFE_PN__680  (.L_HI(net680));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[25]$_DFFE_PN__681  (.L_HI(net681));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[26]$_DFFE_PN__682  (.L_HI(net682));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[27]$_DFFE_PN__683  (.L_HI(net683));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[28]$_DFFE_PN__684  (.L_HI(net684));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[29]$_DFFE_PN__685  (.L_HI(net685));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[30]$_DFFE_PN__686  (.L_HI(net686));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[31]$_DFFE_PN__687  (.L_HI(net687));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[4]$_DFFE_PN__688  (.L_HI(net688));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[5]$_DFFE_PN__689  (.L_HI(net689));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[6]$_DFFE_PN__690  (.L_HI(net690));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[7]$_DFFE_PN__691  (.L_HI(net691));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[8]$_DFFE_PN__692  (.L_HI(net692));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[17].i_reg.reg_r[9]$_DFFE_PN__693  (.L_HI(net693));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[10]$_DFFE_PN__694  (.L_HI(net694));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[11]$_DFFE_PN__695  (.L_HI(net695));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[12]$_DFFE_PN__696  (.L_HI(net696));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[13]$_DFFE_PN__697  (.L_HI(net697));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[14]$_DFFE_PN__698  (.L_HI(net698));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[15]$_DFFE_PN__699  (.L_HI(net699));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[16]$_DFFE_PN__700  (.L_HI(net700));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[17]$_DFFE_PN__701  (.L_HI(net701));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[18]$_DFFE_PN__702  (.L_HI(net702));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[19]$_DFFE_PN__703  (.L_HI(net703));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[20]$_DFFE_PN__704  (.L_HI(net704));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[21]$_DFFE_PN__705  (.L_HI(net705));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[22]$_DFFE_PN__706  (.L_HI(net706));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[23]$_DFFE_PN__707  (.L_HI(net707));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[24]$_DFFE_PN__708  (.L_HI(net708));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[25]$_DFFE_PN__709  (.L_HI(net709));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[26]$_DFFE_PN__710  (.L_HI(net710));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[27]$_DFFE_PN__711  (.L_HI(net711));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[28]$_DFFE_PN__712  (.L_HI(net712));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[29]$_DFFE_PN__713  (.L_HI(net713));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[30]$_DFFE_PN__714  (.L_HI(net714));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[31]$_DFFE_PN__715  (.L_HI(net715));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[4]$_DFFE_PN__716  (.L_HI(net716));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[5]$_DFFE_PN__717  (.L_HI(net717));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[6]$_DFFE_PN__718  (.L_HI(net718));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[7]$_DFFE_PN__719  (.L_HI(net719));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[8]$_DFFE_PN__720  (.L_HI(net720));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[18].i_reg.reg_r[9]$_DFFE_PN__721  (.L_HI(net721));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[10]$_DFFE_PN__722  (.L_HI(net722));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[11]$_DFFE_PN__723  (.L_HI(net723));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[12]$_DFFE_PN__724  (.L_HI(net724));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[13]$_DFFE_PN__725  (.L_HI(net725));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[14]$_DFFE_PN__726  (.L_HI(net726));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[15]$_DFFE_PN__727  (.L_HI(net727));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[16]$_DFFE_PN__728  (.L_HI(net728));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[17]$_DFFE_PN__729  (.L_HI(net729));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[18]$_DFFE_PN__730  (.L_HI(net730));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[19]$_DFFE_PN__731  (.L_HI(net731));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[20]$_DFFE_PN__732  (.L_HI(net732));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[21]$_DFFE_PN__733  (.L_HI(net733));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[22]$_DFFE_PN__734  (.L_HI(net734));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[23]$_DFFE_PN__735  (.L_HI(net735));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[24]$_DFFE_PN__736  (.L_HI(net736));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[25]$_DFFE_PN__737  (.L_HI(net737));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[26]$_DFFE_PN__738  (.L_HI(net738));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[27]$_DFFE_PN__739  (.L_HI(net739));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[28]$_DFFE_PN__740  (.L_HI(net740));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[29]$_DFFE_PN__741  (.L_HI(net741));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[30]$_DFFE_PN__742  (.L_HI(net742));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[31]$_DFFE_PN__743  (.L_HI(net743));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[4]$_DFFE_PN__744  (.L_HI(net744));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[5]$_DFFE_PN__745  (.L_HI(net745));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[6]$_DFFE_PN__746  (.L_HI(net746));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[7]$_DFFE_PN__747  (.L_HI(net747));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[8]$_DFFE_PN__748  (.L_HI(net748));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[19].i_reg.reg_r[9]$_DFFE_PN__749  (.L_HI(net749));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[10]$_DFFE_PN__750  (.L_HI(net750));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[11]$_DFFE_PN__751  (.L_HI(net751));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[12]$_DFFE_PN__752  (.L_HI(net752));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[13]$_DFFE_PN__753  (.L_HI(net753));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[14]$_DFFE_PN__754  (.L_HI(net754));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[15]$_DFFE_PN__755  (.L_HI(net755));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[16]$_DFFE_PN__756  (.L_HI(net756));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[17]$_DFFE_PN__757  (.L_HI(net757));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[18]$_DFFE_PN__758  (.L_HI(net758));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[19]$_DFFE_PN__759  (.L_HI(net759));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[20]$_DFFE_PN__760  (.L_HI(net760));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[21]$_DFFE_PN__761  (.L_HI(net761));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[22]$_DFFE_PN__762  (.L_HI(net762));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[23]$_DFFE_PN__763  (.L_HI(net763));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[24]$_DFFE_PN__764  (.L_HI(net764));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[25]$_DFFE_PN__765  (.L_HI(net765));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[26]$_DFFE_PN__766  (.L_HI(net766));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[27]$_DFFE_PN__767  (.L_HI(net767));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[28]$_DFFE_PN__768  (.L_HI(net768));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[29]$_DFFE_PN__769  (.L_HI(net769));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[30]$_DFFE_PN__770  (.L_HI(net770));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[31]$_DFFE_PN__771  (.L_HI(net771));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[4]$_DFFE_PN__772  (.L_HI(net772));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[5]$_DFFE_PN__773  (.L_HI(net773));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[6]$_DFFE_PN__774  (.L_HI(net774));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[7]$_DFFE_PN__775  (.L_HI(net775));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[8]$_DFFE_PN__776  (.L_HI(net776));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[1].i_reg.reg_r[9]$_DFFE_PN__777  (.L_HI(net777));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[10]$_DFFE_PN__778  (.L_HI(net778));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[11]$_DFFE_PN__779  (.L_HI(net779));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[12]$_DFFE_PN__780  (.L_HI(net780));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[13]$_DFFE_PN__781  (.L_HI(net781));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[14]$_DFFE_PN__782  (.L_HI(net782));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[15]$_DFFE_PN__783  (.L_HI(net783));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[16]$_DFFE_PN__784  (.L_HI(net784));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[17]$_DFFE_PN__785  (.L_HI(net785));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[18]$_DFFE_PN__786  (.L_HI(net786));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[19]$_DFFE_PN__787  (.L_HI(net787));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[20]$_DFFE_PN__788  (.L_HI(net788));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[21]$_DFFE_PN__789  (.L_HI(net789));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[22]$_DFFE_PN__790  (.L_HI(net790));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[23]$_DFFE_PN__791  (.L_HI(net791));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[24]$_DFFE_PN__792  (.L_HI(net792));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[25]$_DFFE_PN__793  (.L_HI(net793));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[26]$_DFFE_PN__794  (.L_HI(net794));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[27]$_DFFE_PN__795  (.L_HI(net795));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[28]$_DFFE_PN__796  (.L_HI(net796));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[29]$_DFFE_PN__797  (.L_HI(net797));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[30]$_DFFE_PN__798  (.L_HI(net798));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[31]$_DFFE_PN__799  (.L_HI(net799));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[4]$_DFFE_PN__800  (.L_HI(net800));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[5]$_DFFE_PN__801  (.L_HI(net801));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[6]$_DFFE_PN__802  (.L_HI(net802));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[7]$_DFFE_PN__803  (.L_HI(net803));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[8]$_DFFE_PN__804  (.L_HI(net804));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[20].i_reg.reg_r[9]$_DFFE_PN__805  (.L_HI(net805));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[10]$_DFFE_PN__806  (.L_HI(net806));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[11]$_DFFE_PN__807  (.L_HI(net807));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[12]$_DFFE_PN__808  (.L_HI(net808));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[13]$_DFFE_PN__809  (.L_HI(net809));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[14]$_DFFE_PN__810  (.L_HI(net810));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[15]$_DFFE_PN__811  (.L_HI(net811));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[16]$_DFFE_PN__812  (.L_HI(net812));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[17]$_DFFE_PN__813  (.L_HI(net813));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[18]$_DFFE_PN__814  (.L_HI(net814));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[19]$_DFFE_PN__815  (.L_HI(net815));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[20]$_DFFE_PN__816  (.L_HI(net816));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[21]$_DFFE_PN__817  (.L_HI(net817));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[22]$_DFFE_PN__818  (.L_HI(net818));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[23]$_DFFE_PN__819  (.L_HI(net819));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[24]$_DFFE_PN__820  (.L_HI(net820));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[25]$_DFFE_PN__821  (.L_HI(net821));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[26]$_DFFE_PN__822  (.L_HI(net822));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[27]$_DFFE_PN__823  (.L_HI(net823));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[28]$_DFFE_PN__824  (.L_HI(net824));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[29]$_DFFE_PN__825  (.L_HI(net825));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[30]$_DFFE_PN__826  (.L_HI(net826));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[31]$_DFFE_PN__827  (.L_HI(net827));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[4]$_DFFE_PN__828  (.L_HI(net828));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[5]$_DFFE_PN__829  (.L_HI(net829));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[6]$_DFFE_PN__830  (.L_HI(net830));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[7]$_DFFE_PN__831  (.L_HI(net831));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[8]$_DFFE_PN__832  (.L_HI(net832));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[21].i_reg.reg_r[9]$_DFFE_PN__833  (.L_HI(net833));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[10]$_DFFE_PN__834  (.L_HI(net834));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[11]$_DFFE_PN__835  (.L_HI(net835));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[12]$_DFFE_PN__836  (.L_HI(net836));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[13]$_DFFE_PN__837  (.L_HI(net837));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[14]$_DFFE_PN__838  (.L_HI(net838));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[15]$_DFFE_PN__839  (.L_HI(net839));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[16]$_DFFE_PN__840  (.L_HI(net840));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[17]$_DFFE_PN__841  (.L_HI(net841));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[18]$_DFFE_PN__842  (.L_HI(net842));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[19]$_DFFE_PN__843  (.L_HI(net843));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[20]$_DFFE_PN__844  (.L_HI(net844));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[21]$_DFFE_PN__845  (.L_HI(net845));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[22]$_DFFE_PN__846  (.L_HI(net846));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[23]$_DFFE_PN__847  (.L_HI(net847));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[24]$_DFFE_PN__848  (.L_HI(net848));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[25]$_DFFE_PN__849  (.L_HI(net849));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[26]$_DFFE_PN__850  (.L_HI(net850));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[27]$_DFFE_PN__851  (.L_HI(net851));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[28]$_DFFE_PN__852  (.L_HI(net852));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[29]$_DFFE_PN__853  (.L_HI(net853));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[30]$_DFFE_PN__854  (.L_HI(net854));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[31]$_DFFE_PN__855  (.L_HI(net855));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[4]$_DFFE_PN__856  (.L_HI(net856));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[5]$_DFFE_PN__857  (.L_HI(net857));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[6]$_DFFE_PN__858  (.L_HI(net858));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[7]$_DFFE_PN__859  (.L_HI(net859));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[8]$_DFFE_PN__860  (.L_HI(net860));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[22].i_reg.reg_r[9]$_DFFE_PN__861  (.L_HI(net861));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[10]$_DFFE_PN__862  (.L_HI(net862));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[11]$_DFFE_PN__863  (.L_HI(net863));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[12]$_DFFE_PN__864  (.L_HI(net864));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[13]$_DFFE_PN__865  (.L_HI(net865));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[14]$_DFFE_PN__866  (.L_HI(net866));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[15]$_DFFE_PN__867  (.L_HI(net867));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[16]$_DFFE_PN__868  (.L_HI(net868));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[17]$_DFFE_PN__869  (.L_HI(net869));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[18]$_DFFE_PN__870  (.L_HI(net870));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[19]$_DFFE_PN__871  (.L_HI(net871));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[20]$_DFFE_PN__872  (.L_HI(net872));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[21]$_DFFE_PN__873  (.L_HI(net873));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[22]$_DFFE_PN__874  (.L_HI(net874));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[23]$_DFFE_PN__875  (.L_HI(net875));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[24]$_DFFE_PN__876  (.L_HI(net876));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[25]$_DFFE_PN__877  (.L_HI(net877));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[26]$_DFFE_PN__878  (.L_HI(net878));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[27]$_DFFE_PN__879  (.L_HI(net879));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[28]$_DFFE_PN__880  (.L_HI(net880));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[29]$_DFFE_PN__881  (.L_HI(net881));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[30]$_DFFE_PN__882  (.L_HI(net882));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[31]$_DFFE_PN__883  (.L_HI(net883));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[4]$_DFFE_PN__884  (.L_HI(net884));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[5]$_DFFE_PN__885  (.L_HI(net885));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[6]$_DFFE_PN__886  (.L_HI(net886));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[7]$_DFFE_PN__887  (.L_HI(net887));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[8]$_DFFE_PN__888  (.L_HI(net888));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[23].i_reg.reg_r[9]$_DFFE_PN__889  (.L_HI(net889));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[10]$_DFFE_PN__890  (.L_HI(net890));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[11]$_DFFE_PN__891  (.L_HI(net891));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[12]$_DFFE_PN__892  (.L_HI(net892));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[13]$_DFFE_PN__893  (.L_HI(net893));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[14]$_DFFE_PN__894  (.L_HI(net894));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[15]$_DFFE_PN__895  (.L_HI(net895));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[16]$_DFFE_PN__896  (.L_HI(net896));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[17]$_DFFE_PN__897  (.L_HI(net897));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[18]$_DFFE_PN__898  (.L_HI(net898));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[19]$_DFFE_PN__899  (.L_HI(net899));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[20]$_DFFE_PN__900  (.L_HI(net900));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[21]$_DFFE_PN__901  (.L_HI(net901));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[22]$_DFFE_PN__902  (.L_HI(net902));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[23]$_DFFE_PN__903  (.L_HI(net903));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[24]$_DFFE_PN__904  (.L_HI(net904));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[25]$_DFFE_PN__905  (.L_HI(net905));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[26]$_DFFE_PN__906  (.L_HI(net906));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[27]$_DFFE_PN__907  (.L_HI(net907));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[28]$_DFFE_PN__908  (.L_HI(net908));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[29]$_DFFE_PN__909  (.L_HI(net909));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[30]$_DFFE_PN__910  (.L_HI(net910));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[31]$_DFFE_PN__911  (.L_HI(net911));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[4]$_DFFE_PN__912  (.L_HI(net912));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[5]$_DFFE_PN__913  (.L_HI(net913));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[6]$_DFFE_PN__914  (.L_HI(net914));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[7]$_DFFE_PN__915  (.L_HI(net915));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[8]$_DFFE_PN__916  (.L_HI(net916));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[24].i_reg.reg_r[9]$_DFFE_PN__917  (.L_HI(net917));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[10]$_DFFE_PN__918  (.L_HI(net918));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[11]$_DFFE_PN__919  (.L_HI(net919));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[12]$_DFFE_PN__920  (.L_HI(net920));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[13]$_DFFE_PN__921  (.L_HI(net921));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[14]$_DFFE_PN__922  (.L_HI(net922));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[15]$_DFFE_PN__923  (.L_HI(net923));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[16]$_DFFE_PN__924  (.L_HI(net924));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[17]$_DFFE_PN__925  (.L_HI(net925));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[18]$_DFFE_PN__926  (.L_HI(net926));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[19]$_DFFE_PN__927  (.L_HI(net927));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[20]$_DFFE_PN__928  (.L_HI(net928));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[21]$_DFFE_PN__929  (.L_HI(net929));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[22]$_DFFE_PN__930  (.L_HI(net930));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[23]$_DFFE_PN__931  (.L_HI(net931));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[24]$_DFFE_PN__932  (.L_HI(net932));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[25]$_DFFE_PN__933  (.L_HI(net933));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[26]$_DFFE_PN__934  (.L_HI(net934));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[27]$_DFFE_PN__935  (.L_HI(net935));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[28]$_DFFE_PN__936  (.L_HI(net936));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[29]$_DFFE_PN__937  (.L_HI(net937));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[30]$_DFFE_PN__938  (.L_HI(net938));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[31]$_DFFE_PN__939  (.L_HI(net939));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[4]$_DFFE_PN__940  (.L_HI(net940));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[5]$_DFFE_PN__941  (.L_HI(net941));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[6]$_DFFE_PN__942  (.L_HI(net942));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[7]$_DFFE_PN__943  (.L_HI(net943));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[8]$_DFFE_PN__944  (.L_HI(net944));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[25].i_reg.reg_r[9]$_DFFE_PN__945  (.L_HI(net945));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[10]$_DFFE_PN__946  (.L_HI(net946));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[11]$_DFFE_PN__947  (.L_HI(net947));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[12]$_DFFE_PN__948  (.L_HI(net948));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[13]$_DFFE_PN__949  (.L_HI(net949));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[14]$_DFFE_PN__950  (.L_HI(net950));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[15]$_DFFE_PN__951  (.L_HI(net951));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[16]$_DFFE_PN__952  (.L_HI(net952));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[17]$_DFFE_PN__953  (.L_HI(net953));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[18]$_DFFE_PN__954  (.L_HI(net954));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[19]$_DFFE_PN__955  (.L_HI(net955));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[20]$_DFFE_PN__956  (.L_HI(net956));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[21]$_DFFE_PN__957  (.L_HI(net957));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[22]$_DFFE_PN__958  (.L_HI(net958));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[23]$_DFFE_PN__959  (.L_HI(net959));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[24]$_DFFE_PN__960  (.L_HI(net960));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[25]$_DFFE_PN__961  (.L_HI(net961));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[26]$_DFFE_PN__962  (.L_HI(net962));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[27]$_DFFE_PN__963  (.L_HI(net963));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[28]$_DFFE_PN__964  (.L_HI(net964));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[29]$_DFFE_PN__965  (.L_HI(net965));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[30]$_DFFE_PN__966  (.L_HI(net966));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[31]$_DFFE_PN__967  (.L_HI(net967));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[4]$_DFFE_PN__968  (.L_HI(net968));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[5]$_DFFE_PN__969  (.L_HI(net969));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[6]$_DFFE_PN__970  (.L_HI(net970));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[7]$_DFFE_PN__971  (.L_HI(net971));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[8]$_DFFE_PN__972  (.L_HI(net972));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[26].i_reg.reg_r[9]$_DFFE_PN__973  (.L_HI(net973));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[10]$_DFFE_PN__974  (.L_HI(net974));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[11]$_DFFE_PN__975  (.L_HI(net975));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[12]$_DFFE_PN__976  (.L_HI(net976));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[13]$_DFFE_PN__977  (.L_HI(net977));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[14]$_DFFE_PN__978  (.L_HI(net978));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[15]$_DFFE_PN__979  (.L_HI(net979));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[16]$_DFFE_PN__980  (.L_HI(net980));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[17]$_DFFE_PN__981  (.L_HI(net981));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[18]$_DFFE_PN__982  (.L_HI(net982));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[19]$_DFFE_PN__983  (.L_HI(net983));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[20]$_DFFE_PN__984  (.L_HI(net984));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[21]$_DFFE_PN__985  (.L_HI(net985));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[22]$_DFFE_PN__986  (.L_HI(net986));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[23]$_DFFE_PN__987  (.L_HI(net987));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[24]$_DFFE_PN__988  (.L_HI(net988));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[25]$_DFFE_PN__989  (.L_HI(net989));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[26]$_DFFE_PN__990  (.L_HI(net990));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[27]$_DFFE_PN__991  (.L_HI(net991));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[28]$_DFFE_PN__992  (.L_HI(net992));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[29]$_DFFE_PN__993  (.L_HI(net993));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[30]$_DFFE_PN__994  (.L_HI(net994));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[31]$_DFFE_PN__995  (.L_HI(net995));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[4]$_DFFE_PN__996  (.L_HI(net996));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[5]$_DFFE_PN__997  (.L_HI(net997));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[6]$_DFFE_PN__998  (.L_HI(net998));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[7]$_DFFE_PN__999  (.L_HI(net999));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[8]$_DFFE_PN__1000  (.L_HI(net1000));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[27].i_reg.reg_r[9]$_DFFE_PN__1001  (.L_HI(net1001));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[10]$_DFFE_PN__1002  (.L_HI(net1002));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[11]$_DFFE_PN__1003  (.L_HI(net1003));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[12]$_DFFE_PN__1004  (.L_HI(net1004));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[13]$_DFFE_PN__1005  (.L_HI(net1005));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[14]$_DFFE_PN__1006  (.L_HI(net1006));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[15]$_DFFE_PN__1007  (.L_HI(net1007));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[16]$_DFFE_PN__1008  (.L_HI(net1008));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[17]$_DFFE_PN__1009  (.L_HI(net1009));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[18]$_DFFE_PN__1010  (.L_HI(net1010));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[19]$_DFFE_PN__1011  (.L_HI(net1011));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[20]$_DFFE_PN__1012  (.L_HI(net1012));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[21]$_DFFE_PN__1013  (.L_HI(net1013));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[22]$_DFFE_PN__1014  (.L_HI(net1014));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[23]$_DFFE_PN__1015  (.L_HI(net1015));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[24]$_DFFE_PN__1016  (.L_HI(net1016));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[25]$_DFFE_PN__1017  (.L_HI(net1017));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[26]$_DFFE_PN__1018  (.L_HI(net1018));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[27]$_DFFE_PN__1019  (.L_HI(net1019));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[28]$_DFFE_PN__1020  (.L_HI(net1020));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[29]$_DFFE_PN__1021  (.L_HI(net1021));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[30]$_DFFE_PN__1022  (.L_HI(net1022));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[31]$_DFFE_PN__1023  (.L_HI(net1023));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[4]$_DFFE_PN__1024  (.L_HI(net1024));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[5]$_DFFE_PN__1025  (.L_HI(net1025));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[6]$_DFFE_PN__1026  (.L_HI(net1026));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[7]$_DFFE_PN__1027  (.L_HI(net1027));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[8]$_DFFE_PN__1028  (.L_HI(net1028));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[28].i_reg.reg_r[9]$_DFFE_PN__1029  (.L_HI(net1029));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[10]$_DFFE_PN__1030  (.L_HI(net1030));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[11]$_DFFE_PN__1031  (.L_HI(net1031));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[12]$_DFFE_PN__1032  (.L_HI(net1032));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[13]$_DFFE_PN__1033  (.L_HI(net1033));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[14]$_DFFE_PN__1034  (.L_HI(net1034));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[15]$_DFFE_PN__1035  (.L_HI(net1035));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[16]$_DFFE_PN__1036  (.L_HI(net1036));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[17]$_DFFE_PN__1037  (.L_HI(net1037));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[18]$_DFFE_PN__1038  (.L_HI(net1038));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[19]$_DFFE_PN__1039  (.L_HI(net1039));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[20]$_DFFE_PN__1040  (.L_HI(net1040));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[21]$_DFFE_PN__1041  (.L_HI(net1041));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[22]$_DFFE_PN__1042  (.L_HI(net1042));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[23]$_DFFE_PN__1043  (.L_HI(net1043));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[24]$_DFFE_PN__1044  (.L_HI(net1044));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[25]$_DFFE_PN__1045  (.L_HI(net1045));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[26]$_DFFE_PN__1046  (.L_HI(net1046));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[27]$_DFFE_PN__1047  (.L_HI(net1047));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[28]$_DFFE_PN__1048  (.L_HI(net1048));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[29]$_DFFE_PN__1049  (.L_HI(net1049));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[30]$_DFFE_PN__1050  (.L_HI(net1050));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[31]$_DFFE_PN__1051  (.L_HI(net1051));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[4]$_DFFE_PN__1052  (.L_HI(net1052));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[5]$_DFFE_PN__1053  (.L_HI(net1053));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[6]$_DFFE_PN__1054  (.L_HI(net1054));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[7]$_DFFE_PN__1055  (.L_HI(net1055));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[8]$_DFFE_PN__1056  (.L_HI(net1056));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[29].i_reg.reg_r[9]$_DFFE_PN__1057  (.L_HI(net1057));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[10]$_DFFE_PN__1058  (.L_HI(net1058));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[11]$_DFFE_PN__1059  (.L_HI(net1059));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[12]$_DFFE_PN__1060  (.L_HI(net1060));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[13]$_DFFE_PN__1061  (.L_HI(net1061));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[14]$_DFFE_PN__1062  (.L_HI(net1062));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[15]$_DFFE_PN__1063  (.L_HI(net1063));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[16]$_DFFE_PN__1064  (.L_HI(net1064));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[17]$_DFFE_PN__1065  (.L_HI(net1065));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[18]$_DFFE_PN__1066  (.L_HI(net1066));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[19]$_DFFE_PN__1067  (.L_HI(net1067));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[20]$_DFFE_PN__1068  (.L_HI(net1068));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[21]$_DFFE_PN__1069  (.L_HI(net1069));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[22]$_DFFE_PN__1070  (.L_HI(net1070));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[23]$_DFFE_PN__1071  (.L_HI(net1071));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[24]$_DFFE_PN__1072  (.L_HI(net1072));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[25]$_DFFE_PN__1073  (.L_HI(net1073));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[26]$_DFFE_PN__1074  (.L_HI(net1074));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[27]$_DFFE_PN__1075  (.L_HI(net1075));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[28]$_DFFE_PN__1076  (.L_HI(net1076));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[29]$_DFFE_PN__1077  (.L_HI(net1077));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[30]$_DFFE_PN__1078  (.L_HI(net1078));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[31]$_DFFE_PN__1079  (.L_HI(net1079));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[4]$_DFFE_PN__1080  (.L_HI(net1080));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[5]$_DFFE_PN__1081  (.L_HI(net1081));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[6]$_DFFE_PN__1082  (.L_HI(net1082));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[7]$_DFFE_PN__1083  (.L_HI(net1083));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[8]$_DFFE_PN__1084  (.L_HI(net1084));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[2].i_reg.reg_r[9]$_DFFE_PN__1085  (.L_HI(net1085));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[10]$_DFFE_PN__1086  (.L_HI(net1086));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[11]$_DFFE_PN__1087  (.L_HI(net1087));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[12]$_DFFE_PN__1088  (.L_HI(net1088));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[13]$_DFFE_PN__1089  (.L_HI(net1089));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[14]$_DFFE_PN__1090  (.L_HI(net1090));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[15]$_DFFE_PN__1091  (.L_HI(net1091));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[16]$_DFFE_PN__1092  (.L_HI(net1092));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[17]$_DFFE_PN__1093  (.L_HI(net1093));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[18]$_DFFE_PN__1094  (.L_HI(net1094));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[19]$_DFFE_PN__1095  (.L_HI(net1095));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[20]$_DFFE_PN__1096  (.L_HI(net1096));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[21]$_DFFE_PN__1097  (.L_HI(net1097));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[22]$_DFFE_PN__1098  (.L_HI(net1098));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[23]$_DFFE_PN__1099  (.L_HI(net1099));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[24]$_DFFE_PN__1100  (.L_HI(net1100));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[25]$_DFFE_PN__1101  (.L_HI(net1101));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[26]$_DFFE_PN__1102  (.L_HI(net1102));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[27]$_DFFE_PN__1103  (.L_HI(net1103));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[28]$_DFFE_PN__1104  (.L_HI(net1104));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[29]$_DFFE_PN__1105  (.L_HI(net1105));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[30]$_DFFE_PN__1106  (.L_HI(net1106));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[31]$_DFFE_PN__1107  (.L_HI(net1107));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[4]$_DFFE_PN__1108  (.L_HI(net1108));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[5]$_DFFE_PN__1109  (.L_HI(net1109));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[6]$_DFFE_PN__1110  (.L_HI(net1110));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[7]$_DFFE_PN__1111  (.L_HI(net1111));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[8]$_DFFE_PN__1112  (.L_HI(net1112));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[30].i_reg.reg_r[9]$_DFFE_PN__1113  (.L_HI(net1113));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[10]$_DFFE_PN__1114  (.L_HI(net1114));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[11]$_DFFE_PN__1115  (.L_HI(net1115));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[12]$_DFFE_PN__1116  (.L_HI(net1116));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[13]$_DFFE_PN__1117  (.L_HI(net1117));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[14]$_DFFE_PN__1118  (.L_HI(net1118));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[15]$_DFFE_PN__1119  (.L_HI(net1119));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[16]$_DFFE_PN__1120  (.L_HI(net1120));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[17]$_DFFE_PN__1121  (.L_HI(net1121));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[18]$_DFFE_PN__1122  (.L_HI(net1122));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[19]$_DFFE_PN__1123  (.L_HI(net1123));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[20]$_DFFE_PN__1124  (.L_HI(net1124));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[21]$_DFFE_PN__1125  (.L_HI(net1125));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[22]$_DFFE_PN__1126  (.L_HI(net1126));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[23]$_DFFE_PN__1127  (.L_HI(net1127));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[24]$_DFFE_PN__1128  (.L_HI(net1128));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[25]$_DFFE_PN__1129  (.L_HI(net1129));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[26]$_DFFE_PN__1130  (.L_HI(net1130));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[27]$_DFFE_PN__1131  (.L_HI(net1131));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[28]$_DFFE_PN__1132  (.L_HI(net1132));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[29]$_DFFE_PN__1133  (.L_HI(net1133));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[30]$_DFFE_PN__1134  (.L_HI(net1134));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[31]$_DFFE_PN__1135  (.L_HI(net1135));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[4]$_DFFE_PN__1136  (.L_HI(net1136));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[5]$_DFFE_PN__1137  (.L_HI(net1137));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[6]$_DFFE_PN__1138  (.L_HI(net1138));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[7]$_DFFE_PN__1139  (.L_HI(net1139));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[8]$_DFFE_PN__1140  (.L_HI(net1140));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[31].i_reg.reg_r[9]$_DFFE_PN__1141  (.L_HI(net1141));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[10]$_DFFE_PN__1142  (.L_HI(net1142));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[11]$_DFFE_PN__1143  (.L_HI(net1143));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[12]$_DFFE_PN__1144  (.L_HI(net1144));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[13]$_DFFE_PN__1145  (.L_HI(net1145));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[14]$_DFFE_PN__1146  (.L_HI(net1146));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[15]$_DFFE_PN__1147  (.L_HI(net1147));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[16]$_DFFE_PN__1148  (.L_HI(net1148));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[17]$_DFFE_PN__1149  (.L_HI(net1149));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[18]$_DFFE_PN__1150  (.L_HI(net1150));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[19]$_DFFE_PN__1151  (.L_HI(net1151));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[20]$_DFFE_PN__1152  (.L_HI(net1152));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[21]$_DFFE_PN__1153  (.L_HI(net1153));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[22]$_DFFE_PN__1154  (.L_HI(net1154));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[23]$_DFFE_PN__1155  (.L_HI(net1155));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[24]$_DFFE_PN__1156  (.L_HI(net1156));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[25]$_DFFE_PN__1157  (.L_HI(net1157));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[26]$_DFFE_PN__1158  (.L_HI(net1158));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[27]$_DFFE_PN__1159  (.L_HI(net1159));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[28]$_DFFE_PN__1160  (.L_HI(net1160));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[29]$_DFFE_PN__1161  (.L_HI(net1161));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[30]$_DFFE_PN__1162  (.L_HI(net1162));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[31]$_DFFE_PN__1163  (.L_HI(net1163));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[4]$_DFFE_PN__1164  (.L_HI(net1164));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[5]$_DFFE_PN__1165  (.L_HI(net1165));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[6]$_DFFE_PN__1166  (.L_HI(net1166));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[7]$_DFFE_PN__1167  (.L_HI(net1167));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[8]$_DFFE_PN__1168  (.L_HI(net1168));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[3].i_reg.reg_r[9]$_DFFE_PN__1169  (.L_HI(net1169));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[10]$_DFFE_PN__1170  (.L_HI(net1170));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[11]$_DFFE_PN__1171  (.L_HI(net1171));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[12]$_DFFE_PN__1172  (.L_HI(net1172));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[13]$_DFFE_PN__1173  (.L_HI(net1173));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[14]$_DFFE_PN__1174  (.L_HI(net1174));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[15]$_DFFE_PN__1175  (.L_HI(net1175));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[16]$_DFFE_PN__1176  (.L_HI(net1176));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[17]$_DFFE_PN__1177  (.L_HI(net1177));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[18]$_DFFE_PN__1178  (.L_HI(net1178));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[19]$_DFFE_PN__1179  (.L_HI(net1179));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[20]$_DFFE_PN__1180  (.L_HI(net1180));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[21]$_DFFE_PN__1181  (.L_HI(net1181));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[22]$_DFFE_PN__1182  (.L_HI(net1182));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[23]$_DFFE_PN__1183  (.L_HI(net1183));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[24]$_DFFE_PN__1184  (.L_HI(net1184));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[25]$_DFFE_PN__1185  (.L_HI(net1185));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[26]$_DFFE_PN__1186  (.L_HI(net1186));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[27]$_DFFE_PN__1187  (.L_HI(net1187));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[28]$_DFFE_PN__1188  (.L_HI(net1188));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[29]$_DFFE_PN__1189  (.L_HI(net1189));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[30]$_DFFE_PN__1190  (.L_HI(net1190));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[31]$_DFFE_PN__1191  (.L_HI(net1191));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[4]$_DFFE_PN__1192  (.L_HI(net1192));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[5]$_DFFE_PN__1193  (.L_HI(net1193));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[6]$_DFFE_PN__1194  (.L_HI(net1194));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[7]$_DFFE_PN__1195  (.L_HI(net1195));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[8]$_DFFE_PN__1196  (.L_HI(net1196));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[4].i_reg.reg_r[9]$_DFFE_PN__1197  (.L_HI(net1197));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[10]$_DFFE_PN__1198  (.L_HI(net1198));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[11]$_DFFE_PN__1199  (.L_HI(net1199));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[12]$_DFFE_PN__1200  (.L_HI(net1200));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[13]$_DFFE_PN__1201  (.L_HI(net1201));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[14]$_DFFE_PN__1202  (.L_HI(net1202));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[15]$_DFFE_PN__1203  (.L_HI(net1203));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[16]$_DFFE_PN__1204  (.L_HI(net1204));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[17]$_DFFE_PN__1205  (.L_HI(net1205));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[18]$_DFFE_PN__1206  (.L_HI(net1206));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[19]$_DFFE_PN__1207  (.L_HI(net1207));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[20]$_DFFE_PN__1208  (.L_HI(net1208));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[21]$_DFFE_PN__1209  (.L_HI(net1209));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[22]$_DFFE_PN__1210  (.L_HI(net1210));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[23]$_DFFE_PN__1211  (.L_HI(net1211));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[24]$_DFFE_PN__1212  (.L_HI(net1212));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[25]$_DFFE_PN__1213  (.L_HI(net1213));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[26]$_DFFE_PN__1214  (.L_HI(net1214));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[27]$_DFFE_PN__1215  (.L_HI(net1215));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[28]$_DFFE_PN__1216  (.L_HI(net1216));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[29]$_DFFE_PN__1217  (.L_HI(net1217));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[30]$_DFFE_PN__1218  (.L_HI(net1218));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[31]$_DFFE_PN__1219  (.L_HI(net1219));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[4]$_DFFE_PN__1220  (.L_HI(net1220));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[5]$_DFFE_PN__1221  (.L_HI(net1221));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[6]$_DFFE_PN__1222  (.L_HI(net1222));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[7]$_DFFE_PN__1223  (.L_HI(net1223));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[8]$_DFFE_PN__1224  (.L_HI(net1224));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[5].i_reg.reg_r[9]$_DFFE_PN__1225  (.L_HI(net1225));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[10]$_DFFE_PN__1226  (.L_HI(net1226));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[11]$_DFFE_PN__1227  (.L_HI(net1227));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[12]$_DFFE_PN__1228  (.L_HI(net1228));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[13]$_DFFE_PN__1229  (.L_HI(net1229));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[14]$_DFFE_PN__1230  (.L_HI(net1230));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[15]$_DFFE_PN__1231  (.L_HI(net1231));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[16]$_DFFE_PN__1232  (.L_HI(net1232));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[17]$_DFFE_PN__1233  (.L_HI(net1233));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[18]$_DFFE_PN__1234  (.L_HI(net1234));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[19]$_DFFE_PN__1235  (.L_HI(net1235));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[20]$_DFFE_PN__1236  (.L_HI(net1236));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[21]$_DFFE_PN__1237  (.L_HI(net1237));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[22]$_DFFE_PN__1238  (.L_HI(net1238));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[23]$_DFFE_PN__1239  (.L_HI(net1239));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[24]$_DFFE_PN__1240  (.L_HI(net1240));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[25]$_DFFE_PN__1241  (.L_HI(net1241));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[26]$_DFFE_PN__1242  (.L_HI(net1242));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[27]$_DFFE_PN__1243  (.L_HI(net1243));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[28]$_DFFE_PN__1244  (.L_HI(net1244));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[29]$_DFFE_PN__1245  (.L_HI(net1245));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[30]$_DFFE_PN__1246  (.L_HI(net1246));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[31]$_DFFE_PN__1247  (.L_HI(net1247));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[4]$_DFFE_PN__1248  (.L_HI(net1248));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[5]$_DFFE_PN__1249  (.L_HI(net1249));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[6]$_DFFE_PN__1250  (.L_HI(net1250));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[7]$_DFFE_PN__1251  (.L_HI(net1251));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[8]$_DFFE_PN__1252  (.L_HI(net1252));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[6].i_reg.reg_r[9]$_DFFE_PN__1253  (.L_HI(net1253));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[10]$_DFFE_PN__1254  (.L_HI(net1254));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[11]$_DFFE_PN__1255  (.L_HI(net1255));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[12]$_DFFE_PN__1256  (.L_HI(net1256));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[13]$_DFFE_PN__1257  (.L_HI(net1257));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[14]$_DFFE_PN__1258  (.L_HI(net1258));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[15]$_DFFE_PN__1259  (.L_HI(net1259));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[16]$_DFFE_PN__1260  (.L_HI(net1260));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[17]$_DFFE_PN__1261  (.L_HI(net1261));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[18]$_DFFE_PN__1262  (.L_HI(net1262));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[19]$_DFFE_PN__1263  (.L_HI(net1263));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[20]$_DFFE_PN__1264  (.L_HI(net1264));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[21]$_DFFE_PN__1265  (.L_HI(net1265));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[22]$_DFFE_PN__1266  (.L_HI(net1266));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[23]$_DFFE_PN__1267  (.L_HI(net1267));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[24]$_DFFE_PN__1268  (.L_HI(net1268));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[25]$_DFFE_PN__1269  (.L_HI(net1269));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[26]$_DFFE_PN__1270  (.L_HI(net1270));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[27]$_DFFE_PN__1271  (.L_HI(net1271));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[28]$_DFFE_PN__1272  (.L_HI(net1272));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[29]$_DFFE_PN__1273  (.L_HI(net1273));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[30]$_DFFE_PN__1274  (.L_HI(net1274));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[31]$_DFFE_PN__1275  (.L_HI(net1275));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[4]$_DFFE_PN__1276  (.L_HI(net1276));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[5]$_DFFE_PN__1277  (.L_HI(net1277));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[6]$_DFFE_PN__1278  (.L_HI(net1278));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[7]$_DFFE_PN__1279  (.L_HI(net1279));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[8]$_DFFE_PN__1280  (.L_HI(net1280));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[7].i_reg.reg_r[9]$_DFFE_PN__1281  (.L_HI(net1281));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[10]$_DFFE_PN__1282  (.L_HI(net1282));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[11]$_DFFE_PN__1283  (.L_HI(net1283));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[12]$_DFFE_PN__1284  (.L_HI(net1284));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[13]$_DFFE_PN__1285  (.L_HI(net1285));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[14]$_DFFE_PN__1286  (.L_HI(net1286));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[15]$_DFFE_PN__1287  (.L_HI(net1287));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[16]$_DFFE_PN__1288  (.L_HI(net1288));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[17]$_DFFE_PN__1289  (.L_HI(net1289));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[18]$_DFFE_PN__1290  (.L_HI(net1290));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[19]$_DFFE_PN__1291  (.L_HI(net1291));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[20]$_DFFE_PN__1292  (.L_HI(net1292));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[21]$_DFFE_PN__1293  (.L_HI(net1293));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[22]$_DFFE_PN__1294  (.L_HI(net1294));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[23]$_DFFE_PN__1295  (.L_HI(net1295));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[24]$_DFFE_PN__1296  (.L_HI(net1296));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[25]$_DFFE_PN__1297  (.L_HI(net1297));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[26]$_DFFE_PN__1298  (.L_HI(net1298));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[27]$_DFFE_PN__1299  (.L_HI(net1299));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[28]$_DFFE_PN__1300  (.L_HI(net1300));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[29]$_DFFE_PN__1301  (.L_HI(net1301));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[30]$_DFFE_PN__1302  (.L_HI(net1302));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[31]$_DFFE_PN__1303  (.L_HI(net1303));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[4]$_DFFE_PN__1304  (.L_HI(net1304));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[5]$_DFFE_PN__1305  (.L_HI(net1305));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[6]$_DFFE_PN__1306  (.L_HI(net1306));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[7]$_DFFE_PN__1307  (.L_HI(net1307));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[8]$_DFFE_PN__1308  (.L_HI(net1308));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[8].i_reg.reg_r[9]$_DFFE_PN__1309  (.L_HI(net1309));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[10]$_DFFE_PN__1310  (.L_HI(net1310));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[11]$_DFFE_PN__1311  (.L_HI(net1311));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[12]$_DFFE_PN__1312  (.L_HI(net1312));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[13]$_DFFE_PN__1313  (.L_HI(net1313));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[14]$_DFFE_PN__1314  (.L_HI(net1314));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[15]$_DFFE_PN__1315  (.L_HI(net1315));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[16]$_DFFE_PN__1316  (.L_HI(net1316));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[17]$_DFFE_PN__1317  (.L_HI(net1317));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[18]$_DFFE_PN__1318  (.L_HI(net1318));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[19]$_DFFE_PN__1319  (.L_HI(net1319));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[20]$_DFFE_PN__1320  (.L_HI(net1320));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[21]$_DFFE_PN__1321  (.L_HI(net1321));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[22]$_DFFE_PN__1322  (.L_HI(net1322));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[23]$_DFFE_PN__1323  (.L_HI(net1323));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[24]$_DFFE_PN__1324  (.L_HI(net1324));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[25]$_DFFE_PN__1325  (.L_HI(net1325));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[26]$_DFFE_PN__1326  (.L_HI(net1326));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[27]$_DFFE_PN__1327  (.L_HI(net1327));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[28]$_DFFE_PN__1328  (.L_HI(net1328));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[29]$_DFFE_PN__1329  (.L_HI(net1329));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[30]$_DFFE_PN__1330  (.L_HI(net1330));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[31]$_DFFE_PN__1331  (.L_HI(net1331));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[4]$_DFFE_PN__1332  (.L_HI(net1332));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[5]$_DFFE_PN__1333  (.L_HI(net1333));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[6]$_DFFE_PN__1334  (.L_HI(net1334));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[7]$_DFFE_PN__1335  (.L_HI(net1335));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[8]$_DFFE_PN__1336  (.L_HI(net1336));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1_reg[9].i_reg.reg_r[9]$_DFFE_PN__1337  (.L_HI(net1337));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[0]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[1]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[2]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[3]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs1_i[4]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[0]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[1]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[2]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[3]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rs2_i[4]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_ack$_DFF_P__1353  (.L_HI(net1353));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_shft$_DFF_P__1354  (.L_HI(net1354));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_cyc_two$_DFF_P__1355  (.L_HI(net1355));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0]$_SDFF_PP0__1356  (.L_HI(net1356));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1]$_SDFF_PP0__1357  (.L_HI(net1357));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2]$_SDFF_PP0__1358  (.L_HI(net1358));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_lsb$_DFF_P__1359  (.L_HI(net1359));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[0]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.adr_lsbs_i[1]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[10]$_DFF_P__1362  (.L_HI(net1362));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[11]$_DFF_P__1363  (.L_HI(net1363));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[1]$_SDFF_PN1__1364  (.L_HI(net1364));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[2]$_DFF_P__1365  (.L_HI(net1365));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[31]$_DFF_P__1366  (.L_HI(net1366));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[3]$_DFF_P__1367  (.L_HI(net1367));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[4]$_DFF_P__1368  (.L_HI(net1368));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[5]$_DFF_P__1369  (.L_HI(net1369));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[6]$_DFF_P__1370  (.L_HI(net1370));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[7]$_DFF_P__1371  (.L_HI(net1371));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[8]$_SDFF_PN0__1372  (.L_HI(net1372));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.b_imm_reg[9]$_DFF_P__1373  (.L_HI(net1373));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[0]$_SDFF_PN0__1374  (.L_HI(net1374));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[1]$_DFF_P__1375  (.L_HI(net1375));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[2]$_DFF_P__1376  (.L_HI(net1376));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[3]$_DFF_P__1377  (.L_HI(net1377));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_imm_reg[4]$_SDFF_PN1__1378  (.L_HI(net1378));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[29]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[2]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[30]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[3]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[4]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[5]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r_reg[6]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[10]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[11]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[12]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[13]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[14]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[15]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[16]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[17]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[18]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[19]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[20]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[21]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[22]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[23]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[24]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[25]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[26]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[27]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[28]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[29]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[30]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[31]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[4]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[5]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[6]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[7]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[8]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_r_reg[9]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[0]$_SDFF_PN0__1418  (.L_HI(net1418));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[12]$_SDFF_PN1__1419  (.L_HI(net1419));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[13]$_DFF_P__1420  (.L_HI(net1420));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[14]$_DFF_P__1421  (.L_HI(net1421));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[15]$_DFF_P__1422  (.L_HI(net1422));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[16]$_SDFF_PN1__1423  (.L_HI(net1423));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[17]$_DFF_P__1424  (.L_HI(net1424));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[18]$_DFF_P__1425  (.L_HI(net1425));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[19]$_DFF_P__1426  (.L_HI(net1426));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[1]$_DFF_P__1427  (.L_HI(net1427));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[2]$_DFF_P__1428  (.L_HI(net1428));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[3]$_DFF_P__1429  (.L_HI(net1429));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[4]$_SDFF_PN0__1430  (.L_HI(net1430));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[5]$_DFF_P__1431  (.L_HI(net1431));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.instr_i_reg[6]$_DFF_P__1432  (.L_HI(net1432));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ld_sext_o$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_h_o$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.ls_w_o$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r$_DFF_P__1436  (.L_HI(net1436));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r$_DFF_P__1437  (.L_HI(net1437));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.imem_stb_o$_DFF_P__1438  (.L_HI(net1438));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[1]$_DFF_P__1439  (.L_HI(net1439));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_cntrl.state_r_reg[3]$_DFF_P__1440  (.L_HI(net1440));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r$_DFF_P__1441  (.L_HI(net1441));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i$_SDFFE_PN0N__1442  (.L_HI(net1442));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i$_SDFFE_PN0N__1443  (.L_HI(net1443));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[2].i_hadd.a_i$_SDFFE_PN0N__1444  (.L_HI(net1444));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[3].i_hadd.a_i$_SDFFE_PN0N__1445  (.L_HI(net1445));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[10]$_SDFFE_PN0N__1446  (.L_HI(net1446));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[11]$_SDFFE_PN0N__1447  (.L_HI(net1447));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[12]$_SDFFE_PN0N__1448  (.L_HI(net1448));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[13]$_SDFFE_PN0N__1449  (.L_HI(net1449));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[14]$_SDFFE_PN0N__1450  (.L_HI(net1450));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[15]$_SDFFE_PN0N__1451  (.L_HI(net1451));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[16]$_SDFFE_PN0N__1452  (.L_HI(net1452));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[17]$_SDFFE_PN0N__1453  (.L_HI(net1453));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[18]$_SDFFE_PN0N__1454  (.L_HI(net1454));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[19]$_SDFFE_PN0N__1455  (.L_HI(net1455));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[20]$_SDFFE_PN0N__1456  (.L_HI(net1456));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[21]$_SDFFE_PN0N__1457  (.L_HI(net1457));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[22]$_SDFFE_PN0N__1458  (.L_HI(net1458));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[23]$_SDFFE_PN0N__1459  (.L_HI(net1459));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[24]$_SDFFE_PN0N__1460  (.L_HI(net1460));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[25]$_SDFFE_PN0N__1461  (.L_HI(net1461));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[26]$_SDFFE_PN0N__1462  (.L_HI(net1462));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[27]$_SDFFE_PN0N__1463  (.L_HI(net1463));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[28]$_SDFFE_PN0N__1464  (.L_HI(net1464));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[29]$_SDFFE_PN0N__1465  (.L_HI(net1465));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[30]$_SDFFE_PN0N__1466  (.L_HI(net1466));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[31]$_SDFFE_PN0N__1467  (.L_HI(net1467));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[4]$_SDFFE_PN0N__1468  (.L_HI(net1468));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[5]$_SDFFE_PN0N__1469  (.L_HI(net1469));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[6]$_SDFFE_PN0N__1470  (.L_HI(net1470));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[7]$_SDFFE_PN0N__1471  (.L_HI(net1471));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[8]$_SDFFE_PN0N__1472  (.L_HI(net1472));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.pc_o_reg[9]$_SDFFE_PN0N__1473  (.L_HI(net1473));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[10]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[11]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[12]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[13]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[14]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[15]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[16]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[17]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[18]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[19]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[20]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[21]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[22]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[23]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[24]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[25]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[26]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[27]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[28]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[29]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[2]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[30]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[31]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[3]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[4]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[5]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[6]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[7]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[8]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_a.par_o_reg[9]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0]$_DFF_P__1504  (.L_HI(net1504));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1]$_DFF_P__1505  (.L_HI(net1505));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2]$_DFF_P__1506  (.L_HI(net1506));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3]$_DFF_P__1507  (.L_HI(net1507));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[0]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[10]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[11]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[12]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[13]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[14]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[15]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[16]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[17]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[18]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[19]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[1]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[20]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[21]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[22]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[23]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[24]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[25]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[26]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[27]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[28]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[29]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[2]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[30]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[31]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[3]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[4]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[5]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[6]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[7]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[8]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.pdout_o[9]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[0]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[1]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[2]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.reg_r_reg[3]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r$_SDFFE_PN0P__1544  (.L_HI(net1544));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.cnt_r[0]$_SDFF_PN0__1545  (.L_HI(net1545));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.cnt_r[1]$_SDFF_PN0__1546  (.L_HI(net1546));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.cnt_r[2]$_SDFF_PN0__1547  (.L_HI(net1547));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.crm_r$_SDFFE_PN0P__1548  (.L_HI(net1548));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[0]$_DFF_P__1549  (.L_HI(net1549));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[1]$_DFF_P__1550  (.L_HI(net1550));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[2]$_DFF_P__1551  (.L_HI(net1551));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[3]$_DFF_P__1552  (.L_HI(net1552));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[4]$_DFF_P__1553  (.L_HI(net1553));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[5]$_DFF_P__1554  (.L_HI(net1554));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.state_r_reg[6]$_DFF_P__1555  (.L_HI(net1555));
 sg13g2_tiehi \i_exotiny.i_wb_qspi_mem.wb_mem_ack_o$_DFF_P__1556  (.L_HI(net1556));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_auto_cs_o$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_cpol_o$_SDFFE_PN0P__1558  (.L_HI(net1558));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_presc_o[0]$_SDFFE_PN1P__1559  (.L_HI(net1559));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_presc_o[1]$_SDFFE_PN1P__1560  (.L_HI(net1560));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_presc_o[2]$_SDFFE_PN0P__1561  (.L_HI(net1561));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_presc_o[3]$_SDFFE_PN1P__1562  (.L_HI(net1562));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_rdy_i$_DFF_P__1563  (.L_HI(net1563));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_size_o[0]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \i_exotiny.i_wb_regs.spi_size_o[1]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[0]$_SDFFCE_PN0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[1]$_SDFFCE_PN0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[2]$_SDFFCE_PN0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[3]$_SDFFCE_PN0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[4]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[5]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_hbit_r[6]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[0]$_DFF_P__1573  (.L_HI(net1573));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[1]$_DFF_P__1574  (.L_HI(net1574));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[2]$_DFF_P__1575  (.L_HI(net1575));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[3]$_DFF_P__1576  (.L_HI(net1576));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[4]$_DFF_P__1577  (.L_HI(net1577));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[5]$_DFF_P__1578  (.L_HI(net1578));
 sg13g2_tiehi \i_exotiny.i_wb_spi.cnt_presc_r[6]$_DFF_P__1579  (.L_HI(net1579));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[0]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[10]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[11]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[12]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[13]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[14]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[15]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[16]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[17]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[18]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[19]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[1]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[20]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[21]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[22]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[23]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[24]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[25]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[26]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[27]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[28]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[29]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[2]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[30]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[31]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[3]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[4]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[5]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[6]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[7]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[8]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_rx_r[9]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[0]$_SDFFCE_PP0P__1612  (.L_HI(net1612));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[10]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[11]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[12]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[13]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[14]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[15]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[16]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[17]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[18]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[19]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[1]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[20]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[21]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[22]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[23]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[24]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[25]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[26]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[27]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[28]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[29]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[2]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[30]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[3]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[4]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[5]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[6]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[7]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[8]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \i_exotiny.i_wb_spi.dat_tx_r_reg[9]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \i_exotiny.i_wb_spi.state_r_reg[1]$_DFF_P__1643  (.L_HI(net1643));
 sg13g2_tiehi \i_exotiny.spi_sck_o$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \i_exotiny.spi_sdo_o$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_buf_4 clkbuf_leaf_1_clk (.X(clknet_leaf_1_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_2_clk (.X(clknet_leaf_2_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_3_clk (.X(clknet_leaf_3_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_4_clk (.X(clknet_leaf_4_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_5_clk (.X(clknet_leaf_5_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_6_clk (.X(clknet_leaf_6_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_7_clk (.X(clknet_leaf_7_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_8_clk (.X(clknet_leaf_8_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_9_clk (.X(clknet_leaf_9_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_10_clk (.X(clknet_leaf_10_clk),
    .A(clknet_5_2__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_11_clk (.X(clknet_leaf_11_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_12_clk (.X(clknet_leaf_12_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_13_clk (.X(clknet_leaf_13_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_14_clk (.X(clknet_leaf_14_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_15_clk (.X(clknet_leaf_15_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_16_clk (.X(clknet_leaf_16_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_17_clk (.X(clknet_leaf_17_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_18_clk (.X(clknet_leaf_18_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_19_clk (.X(clknet_leaf_19_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_20_clk (.X(clknet_leaf_20_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_21_clk (.X(clknet_leaf_21_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_22_clk (.X(clknet_leaf_22_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_23_clk (.X(clknet_leaf_23_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_24_clk (.X(clknet_leaf_24_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_25_clk (.X(clknet_leaf_25_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_26_clk (.X(clknet_leaf_26_clk),
    .A(clknet_5_8__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_27_clk (.X(clknet_leaf_27_clk),
    .A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_28_clk (.X(clknet_leaf_28_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_29_clk (.X(clknet_leaf_29_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_30_clk (.X(clknet_leaf_30_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_31_clk (.X(clknet_leaf_31_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_32_clk (.X(clknet_leaf_32_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_33_clk (.X(clknet_leaf_33_clk),
    .A(clknet_5_10__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_34_clk (.X(clknet_leaf_34_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_35_clk (.X(clknet_leaf_35_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_36_clk (.X(clknet_leaf_36_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_37_clk (.X(clknet_leaf_37_clk),
    .A(clknet_5_11__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_38_clk (.X(clknet_leaf_38_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_39_clk (.X(clknet_leaf_39_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_40_clk (.X(clknet_leaf_40_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_41_clk (.X(clknet_leaf_41_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_42_clk (.X(clknet_leaf_42_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_43_clk (.X(clknet_leaf_43_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_44_clk (.X(clknet_leaf_44_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_45_clk (.X(clknet_leaf_45_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_46_clk (.X(clknet_leaf_46_clk),
    .A(clknet_5_15__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_47_clk (.X(clknet_leaf_47_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_48_clk (.X(clknet_leaf_48_clk),
    .A(clknet_5_14__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_49_clk (.X(clknet_leaf_49_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_50_clk (.X(clknet_leaf_50_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_51_clk (.X(clknet_leaf_51_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_52_clk (.X(clknet_leaf_52_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_53_clk (.X(clknet_leaf_53_clk),
    .A(clknet_5_12__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_54_clk (.X(clknet_leaf_54_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_55_clk (.X(clknet_leaf_55_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_56_clk (.X(clknet_leaf_56_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_57_clk (.X(clknet_leaf_57_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_58_clk (.X(clknet_leaf_58_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_59_clk (.X(clknet_leaf_59_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_60_clk (.X(clknet_leaf_60_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_61_clk (.X(clknet_leaf_61_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_62_clk (.X(clknet_leaf_62_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_63_clk (.X(clknet_leaf_63_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_64_clk (.X(clknet_leaf_64_clk),
    .A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_65_clk (.X(clknet_leaf_65_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_66_clk (.X(clknet_leaf_66_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_67_clk (.X(clknet_leaf_67_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_68_clk (.X(clknet_leaf_68_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_69_clk (.X(clknet_leaf_69_clk),
    .A(clknet_5_26__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_70_clk (.X(clknet_leaf_70_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_71_clk (.X(clknet_leaf_71_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_72_clk (.X(clknet_leaf_72_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_73_clk (.X(clknet_leaf_73_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_74_clk (.X(clknet_leaf_74_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_75_clk (.X(clknet_leaf_75_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_76_clk (.X(clknet_leaf_76_clk),
    .A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_78_clk (.X(clknet_leaf_78_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_79_clk (.X(clknet_leaf_79_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_80_clk (.X(clknet_leaf_80_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_81_clk (.X(clknet_leaf_81_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_82_clk (.X(clknet_leaf_82_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_83_clk (.X(clknet_leaf_83_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_84_clk (.X(clknet_leaf_84_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_85_clk (.X(clknet_leaf_85_clk),
    .A(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_86_clk (.X(clknet_leaf_86_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_87_clk (.X(clknet_leaf_87_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_88_clk (.X(clknet_leaf_88_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_89_clk (.X(clknet_leaf_89_clk),
    .A(clknet_5_30__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_90_clk (.X(clknet_leaf_90_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_91_clk (.X(clknet_leaf_91_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_92_clk (.X(clknet_leaf_92_clk),
    .A(clknet_5_25__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_93_clk (.X(clknet_leaf_93_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_94_clk (.X(clknet_leaf_94_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_95_clk (.X(clknet_leaf_95_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_96_clk (.X(clknet_leaf_96_clk),
    .A(clknet_5_24__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_97_clk (.X(clknet_leaf_97_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_98_clk (.X(clknet_leaf_98_clk),
    .A(clknet_5_28__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_99_clk (.X(clknet_leaf_99_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_100_clk (.X(clknet_leaf_100_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_101_clk (.X(clknet_leaf_101_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_102_clk (.X(clknet_leaf_102_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_103_clk (.X(clknet_leaf_103_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_104_clk (.X(clknet_leaf_104_clk),
    .A(clknet_5_29__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_105_clk (.X(clknet_leaf_105_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_106_clk (.X(clknet_leaf_106_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_107_clk (.X(clknet_leaf_107_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_108_clk (.X(clknet_leaf_108_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_109_clk (.X(clknet_leaf_109_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_110_clk (.X(clknet_leaf_110_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_111_clk (.X(clknet_leaf_111_clk),
    .A(clknet_5_23__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_112_clk (.X(clknet_leaf_112_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_113_clk (.X(clknet_leaf_113_clk),
    .A(clknet_5_22__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_114_clk (.X(clknet_leaf_114_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_115_clk (.X(clknet_leaf_115_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_116_clk (.X(clknet_leaf_116_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_117_clk (.X(clknet_leaf_117_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_118_clk (.X(clknet_leaf_118_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_119_clk (.X(clknet_leaf_119_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_120_clk (.X(clknet_leaf_120_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_121_clk (.X(clknet_leaf_121_clk),
    .A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_122_clk (.X(clknet_leaf_122_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_123_clk (.X(clknet_leaf_123_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_124_clk (.X(clknet_leaf_124_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_125_clk (.X(clknet_leaf_125_clk),
    .A(clknet_5_20__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_126_clk (.X(clknet_leaf_126_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_127_clk (.X(clknet_leaf_127_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_128_clk (.X(clknet_leaf_128_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_129_clk (.X(clknet_leaf_129_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_130_clk (.X(clknet_leaf_130_clk),
    .A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_131_clk (.X(clknet_leaf_131_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_132_clk (.X(clknet_leaf_132_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_133_clk (.X(clknet_leaf_133_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_134_clk (.X(clknet_leaf_134_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_135_clk (.X(clknet_leaf_135_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_136_clk (.X(clknet_leaf_136_clk),
    .A(clknet_5_16__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_137_clk (.X(clknet_leaf_137_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_138_clk (.X(clknet_leaf_138_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_139_clk (.X(clknet_leaf_139_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_140_clk (.X(clknet_leaf_140_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_141_clk (.X(clknet_leaf_141_clk),
    .A(clknet_5_19__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_142_clk (.X(clknet_leaf_142_clk),
    .A(clknet_5_18__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_143_clk (.X(clknet_leaf_143_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_144_clk (.X(clknet_leaf_144_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_145_clk (.X(clknet_leaf_145_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_146_clk (.X(clknet_leaf_146_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_147_clk (.X(clknet_leaf_147_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_148_clk (.X(clknet_leaf_148_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_149_clk (.X(clknet_leaf_149_clk),
    .A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_150_clk (.X(clknet_leaf_150_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_151_clk (.X(clknet_leaf_151_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_152_clk (.X(clknet_leaf_152_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_153_clk (.X(clknet_leaf_153_clk),
    .A(clknet_5_6__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_154_clk (.X(clknet_leaf_154_clk),
    .A(clknet_5_7__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_155_clk (.X(clknet_leaf_155_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_156_clk (.X(clknet_leaf_156_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_157_clk (.X(clknet_leaf_157_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_158_clk (.X(clknet_leaf_158_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_159_clk (.X(clknet_leaf_159_clk),
    .A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_160_clk (.X(clknet_leaf_160_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_161_clk (.X(clknet_leaf_161_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_162_clk (.X(clknet_leaf_162_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_163_clk (.X(clknet_leaf_163_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_164_clk (.X(clknet_leaf_164_clk),
    .A(clknet_5_4__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_165_clk (.X(clknet_leaf_165_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_166_clk (.X(clknet_leaf_166_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_167_clk (.X(clknet_leaf_167_clk),
    .A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkbuf_leaf_168_clk (.X(clknet_leaf_168_clk),
    .A(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_0_0_clk (.X(clknet_4_0_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_1_0_clk (.X(clknet_4_1_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_2_0_clk (.X(clknet_4_2_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_3_0_clk (.X(clknet_4_3_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_4_0_clk (.X(clknet_4_4_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_5_0_clk (.X(clknet_4_5_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_6_0_clk (.X(clknet_4_6_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_7_0_clk (.X(clknet_4_7_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_8_0_clk (.X(clknet_4_8_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_9_0_clk (.X(clknet_4_9_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_10_0_clk (.X(clknet_4_10_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_11_0_clk (.X(clknet_4_11_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_12_0_clk (.X(clknet_4_12_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_13_0_clk (.X(clknet_4_13_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_14_0_clk (.X(clknet_4_14_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_4 clkbuf_4_15_0_clk (.X(clknet_4_15_0_clk),
    .A(clknet_0_clk));
 sg13g2_buf_2 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_2 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_2 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_2 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_2 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_2 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_2 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_2 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_2 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_2 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_2 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_2 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_2 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_2 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_2 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_2 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_2 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_2 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_2 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_2 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_2 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_2 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_2 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_2 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_2 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_2 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_2 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_2 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_2 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_2 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_2 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_2 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_4 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_buf_4 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_buf_4 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_buf_4 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_buf_4 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_buf_4 clkload5 (.A(clknet_5_17__leaf_clk));
 sg13g2_buf_4 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_buf_4 clkload7 (.A(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_4 clkload9 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_16 clkload10 (.A(clknet_leaf_168_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_167_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_15_clk));
 sg13g2_inv_4 clkload13 (.A(clknet_leaf_16_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_leaf_143_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_17_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_leaf_18_clk));
 sg13g2_inv_1 clkload17 (.A(clknet_leaf_20_clk));
 sg13g2_buf_16 clkload18 (.A(clknet_leaf_49_clk));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_53_clk));
 sg13g2_buf_16 clkload20 (.A(clknet_leaf_96_clk));
 sg13g2_inv_1 clkload21 (.A(clknet_leaf_76_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_3238_));
 sg13g2_antennanp ANTENNA_2 (.A(_3238_));
 sg13g2_antennanp ANTENNA_3 (.A(_3238_));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_4 FILLER_0_259 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_fill_2 FILLER_0_347 ();
 sg13g2_fill_1 FILLER_0_349 ();
 sg13g2_fill_1 FILLER_0_380 ();
 sg13g2_fill_1 FILLER_0_469 ();
 sg13g2_fill_2 FILLER_0_500 ();
 sg13g2_fill_1 FILLER_0_536 ();
 sg13g2_fill_2 FILLER_0_567 ();
 sg13g2_fill_1 FILLER_0_569 ();
 sg13g2_fill_2 FILLER_0_604 ();
 sg13g2_fill_2 FILLER_0_690 ();
 sg13g2_fill_2 FILLER_0_736 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_884 ();
 sg13g2_decap_8 FILLER_0_891 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_905 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_8 FILLER_0_926 ();
 sg13g2_decap_8 FILLER_0_933 ();
 sg13g2_decap_8 FILLER_0_940 ();
 sg13g2_decap_8 FILLER_0_947 ();
 sg13g2_decap_8 FILLER_0_954 ();
 sg13g2_decap_8 FILLER_0_961 ();
 sg13g2_decap_8 FILLER_0_968 ();
 sg13g2_decap_8 FILLER_0_975 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_8 FILLER_0_1024 ();
 sg13g2_decap_8 FILLER_0_1031 ();
 sg13g2_decap_8 FILLER_0_1038 ();
 sg13g2_decap_8 FILLER_0_1045 ();
 sg13g2_decap_8 FILLER_0_1052 ();
 sg13g2_decap_8 FILLER_0_1059 ();
 sg13g2_decap_8 FILLER_0_1066 ();
 sg13g2_decap_8 FILLER_0_1073 ();
 sg13g2_decap_8 FILLER_0_1080 ();
 sg13g2_decap_8 FILLER_0_1087 ();
 sg13g2_decap_8 FILLER_0_1094 ();
 sg13g2_decap_8 FILLER_0_1101 ();
 sg13g2_decap_8 FILLER_0_1108 ();
 sg13g2_decap_8 FILLER_0_1115 ();
 sg13g2_decap_8 FILLER_0_1122 ();
 sg13g2_decap_8 FILLER_0_1129 ();
 sg13g2_decap_8 FILLER_0_1136 ();
 sg13g2_decap_8 FILLER_0_1143 ();
 sg13g2_decap_8 FILLER_0_1150 ();
 sg13g2_decap_8 FILLER_0_1157 ();
 sg13g2_decap_8 FILLER_0_1164 ();
 sg13g2_decap_8 FILLER_0_1171 ();
 sg13g2_decap_8 FILLER_0_1178 ();
 sg13g2_decap_8 FILLER_0_1185 ();
 sg13g2_decap_8 FILLER_0_1192 ();
 sg13g2_decap_8 FILLER_0_1199 ();
 sg13g2_decap_8 FILLER_0_1206 ();
 sg13g2_decap_8 FILLER_0_1213 ();
 sg13g2_decap_8 FILLER_0_1220 ();
 sg13g2_decap_8 FILLER_0_1227 ();
 sg13g2_decap_8 FILLER_0_1234 ();
 sg13g2_decap_8 FILLER_0_1241 ();
 sg13g2_decap_8 FILLER_0_1248 ();
 sg13g2_decap_8 FILLER_0_1255 ();
 sg13g2_decap_8 FILLER_0_1262 ();
 sg13g2_decap_8 FILLER_0_1269 ();
 sg13g2_decap_8 FILLER_0_1276 ();
 sg13g2_decap_8 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1290 ();
 sg13g2_decap_8 FILLER_0_1297 ();
 sg13g2_decap_8 FILLER_0_1304 ();
 sg13g2_decap_8 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1318 ();
 sg13g2_fill_1 FILLER_0_1325 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_414 ();
 sg13g2_fill_2 FILLER_1_451 ();
 sg13g2_fill_1 FILLER_1_453 ();
 sg13g2_fill_2 FILLER_1_536 ();
 sg13g2_fill_2 FILLER_1_628 ();
 sg13g2_fill_1 FILLER_1_660 ();
 sg13g2_fill_1 FILLER_1_665 ();
 sg13g2_fill_2 FILLER_1_692 ();
 sg13g2_fill_1 FILLER_1_694 ();
 sg13g2_fill_2 FILLER_1_825 ();
 sg13g2_fill_1 FILLER_1_827 ();
 sg13g2_decap_4 FILLER_1_866 ();
 sg13g2_fill_1 FILLER_1_870 ();
 sg13g2_decap_4 FILLER_1_875 ();
 sg13g2_fill_2 FILLER_1_879 ();
 sg13g2_decap_4 FILLER_1_885 ();
 sg13g2_fill_1 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_894 ();
 sg13g2_decap_8 FILLER_1_901 ();
 sg13g2_decap_8 FILLER_1_908 ();
 sg13g2_decap_8 FILLER_1_915 ();
 sg13g2_decap_8 FILLER_1_922 ();
 sg13g2_decap_8 FILLER_1_929 ();
 sg13g2_decap_8 FILLER_1_936 ();
 sg13g2_decap_8 FILLER_1_943 ();
 sg13g2_decap_8 FILLER_1_950 ();
 sg13g2_decap_8 FILLER_1_957 ();
 sg13g2_decap_8 FILLER_1_964 ();
 sg13g2_decap_8 FILLER_1_971 ();
 sg13g2_decap_8 FILLER_1_978 ();
 sg13g2_decap_8 FILLER_1_985 ();
 sg13g2_decap_8 FILLER_1_992 ();
 sg13g2_decap_8 FILLER_1_999 ();
 sg13g2_decap_8 FILLER_1_1006 ();
 sg13g2_decap_8 FILLER_1_1013 ();
 sg13g2_decap_8 FILLER_1_1020 ();
 sg13g2_decap_8 FILLER_1_1027 ();
 sg13g2_decap_8 FILLER_1_1034 ();
 sg13g2_decap_8 FILLER_1_1041 ();
 sg13g2_decap_8 FILLER_1_1048 ();
 sg13g2_decap_8 FILLER_1_1055 ();
 sg13g2_decap_8 FILLER_1_1062 ();
 sg13g2_decap_8 FILLER_1_1069 ();
 sg13g2_decap_8 FILLER_1_1076 ();
 sg13g2_decap_8 FILLER_1_1083 ();
 sg13g2_decap_8 FILLER_1_1090 ();
 sg13g2_decap_8 FILLER_1_1097 ();
 sg13g2_decap_8 FILLER_1_1104 ();
 sg13g2_decap_8 FILLER_1_1111 ();
 sg13g2_decap_8 FILLER_1_1118 ();
 sg13g2_decap_8 FILLER_1_1125 ();
 sg13g2_decap_8 FILLER_1_1132 ();
 sg13g2_decap_8 FILLER_1_1139 ();
 sg13g2_decap_8 FILLER_1_1146 ();
 sg13g2_decap_8 FILLER_1_1153 ();
 sg13g2_decap_8 FILLER_1_1160 ();
 sg13g2_decap_8 FILLER_1_1167 ();
 sg13g2_decap_8 FILLER_1_1174 ();
 sg13g2_decap_8 FILLER_1_1181 ();
 sg13g2_decap_8 FILLER_1_1188 ();
 sg13g2_decap_8 FILLER_1_1195 ();
 sg13g2_decap_8 FILLER_1_1202 ();
 sg13g2_decap_8 FILLER_1_1209 ();
 sg13g2_decap_8 FILLER_1_1216 ();
 sg13g2_decap_8 FILLER_1_1223 ();
 sg13g2_decap_8 FILLER_1_1230 ();
 sg13g2_decap_8 FILLER_1_1237 ();
 sg13g2_decap_8 FILLER_1_1244 ();
 sg13g2_decap_8 FILLER_1_1251 ();
 sg13g2_decap_8 FILLER_1_1258 ();
 sg13g2_decap_8 FILLER_1_1265 ();
 sg13g2_decap_8 FILLER_1_1272 ();
 sg13g2_decap_8 FILLER_1_1279 ();
 sg13g2_decap_8 FILLER_1_1286 ();
 sg13g2_decap_8 FILLER_1_1293 ();
 sg13g2_decap_8 FILLER_1_1300 ();
 sg13g2_decap_8 FILLER_1_1307 ();
 sg13g2_decap_8 FILLER_1_1314 ();
 sg13g2_decap_4 FILLER_1_1321 ();
 sg13g2_fill_1 FILLER_1_1325 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_fill_1 FILLER_2_259 ();
 sg13g2_fill_1 FILLER_2_300 ();
 sg13g2_fill_2 FILLER_2_343 ();
 sg13g2_fill_1 FILLER_2_435 ();
 sg13g2_fill_2 FILLER_2_472 ();
 sg13g2_fill_1 FILLER_2_474 ();
 sg13g2_fill_2 FILLER_2_493 ();
 sg13g2_fill_1 FILLER_2_495 ();
 sg13g2_fill_2 FILLER_2_526 ();
 sg13g2_fill_1 FILLER_2_554 ();
 sg13g2_fill_1 FILLER_2_621 ();
 sg13g2_fill_1 FILLER_2_658 ();
 sg13g2_fill_2 FILLER_2_757 ();
 sg13g2_fill_1 FILLER_2_773 ();
 sg13g2_fill_1 FILLER_2_800 ();
 sg13g2_fill_1 FILLER_2_811 ();
 sg13g2_fill_2 FILLER_2_846 ();
 sg13g2_fill_2 FILLER_2_862 ();
 sg13g2_fill_2 FILLER_2_898 ();
 sg13g2_fill_1 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_905 ();
 sg13g2_decap_8 FILLER_2_912 ();
 sg13g2_decap_8 FILLER_2_919 ();
 sg13g2_decap_8 FILLER_2_926 ();
 sg13g2_decap_8 FILLER_2_933 ();
 sg13g2_decap_8 FILLER_2_940 ();
 sg13g2_decap_8 FILLER_2_947 ();
 sg13g2_decap_8 FILLER_2_954 ();
 sg13g2_decap_8 FILLER_2_961 ();
 sg13g2_decap_8 FILLER_2_968 ();
 sg13g2_decap_8 FILLER_2_975 ();
 sg13g2_decap_8 FILLER_2_982 ();
 sg13g2_decap_8 FILLER_2_989 ();
 sg13g2_decap_8 FILLER_2_996 ();
 sg13g2_decap_8 FILLER_2_1003 ();
 sg13g2_decap_8 FILLER_2_1010 ();
 sg13g2_decap_8 FILLER_2_1017 ();
 sg13g2_decap_8 FILLER_2_1024 ();
 sg13g2_decap_8 FILLER_2_1031 ();
 sg13g2_decap_8 FILLER_2_1038 ();
 sg13g2_decap_8 FILLER_2_1045 ();
 sg13g2_decap_8 FILLER_2_1052 ();
 sg13g2_decap_8 FILLER_2_1059 ();
 sg13g2_decap_8 FILLER_2_1066 ();
 sg13g2_decap_8 FILLER_2_1073 ();
 sg13g2_decap_8 FILLER_2_1080 ();
 sg13g2_decap_8 FILLER_2_1087 ();
 sg13g2_decap_8 FILLER_2_1094 ();
 sg13g2_decap_8 FILLER_2_1101 ();
 sg13g2_decap_8 FILLER_2_1108 ();
 sg13g2_decap_8 FILLER_2_1115 ();
 sg13g2_decap_8 FILLER_2_1122 ();
 sg13g2_decap_8 FILLER_2_1129 ();
 sg13g2_decap_8 FILLER_2_1136 ();
 sg13g2_decap_8 FILLER_2_1143 ();
 sg13g2_decap_8 FILLER_2_1150 ();
 sg13g2_decap_8 FILLER_2_1157 ();
 sg13g2_decap_8 FILLER_2_1164 ();
 sg13g2_decap_8 FILLER_2_1171 ();
 sg13g2_decap_8 FILLER_2_1178 ();
 sg13g2_decap_8 FILLER_2_1185 ();
 sg13g2_decap_8 FILLER_2_1192 ();
 sg13g2_decap_8 FILLER_2_1199 ();
 sg13g2_decap_8 FILLER_2_1206 ();
 sg13g2_decap_8 FILLER_2_1213 ();
 sg13g2_decap_8 FILLER_2_1220 ();
 sg13g2_decap_8 FILLER_2_1227 ();
 sg13g2_decap_8 FILLER_2_1234 ();
 sg13g2_decap_8 FILLER_2_1241 ();
 sg13g2_decap_8 FILLER_2_1248 ();
 sg13g2_decap_8 FILLER_2_1255 ();
 sg13g2_decap_8 FILLER_2_1262 ();
 sg13g2_decap_8 FILLER_2_1269 ();
 sg13g2_decap_8 FILLER_2_1276 ();
 sg13g2_decap_8 FILLER_2_1283 ();
 sg13g2_decap_8 FILLER_2_1290 ();
 sg13g2_decap_8 FILLER_2_1297 ();
 sg13g2_decap_8 FILLER_2_1304 ();
 sg13g2_decap_8 FILLER_2_1311 ();
 sg13g2_decap_8 FILLER_2_1318 ();
 sg13g2_fill_1 FILLER_2_1325 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_359 ();
 sg13g2_fill_1 FILLER_3_453 ();
 sg13g2_fill_1 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_507 ();
 sg13g2_fill_1 FILLER_3_519 ();
 sg13g2_fill_2 FILLER_3_554 ();
 sg13g2_fill_2 FILLER_3_592 ();
 sg13g2_fill_2 FILLER_3_634 ();
 sg13g2_fill_1 FILLER_3_706 ();
 sg13g2_fill_2 FILLER_3_769 ();
 sg13g2_fill_2 FILLER_3_801 ();
 sg13g2_fill_2 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_8 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_decap_8 FILLER_3_1029 ();
 sg13g2_decap_8 FILLER_3_1036 ();
 sg13g2_decap_8 FILLER_3_1043 ();
 sg13g2_decap_8 FILLER_3_1050 ();
 sg13g2_decap_8 FILLER_3_1057 ();
 sg13g2_decap_8 FILLER_3_1064 ();
 sg13g2_decap_8 FILLER_3_1071 ();
 sg13g2_decap_8 FILLER_3_1078 ();
 sg13g2_decap_8 FILLER_3_1085 ();
 sg13g2_decap_8 FILLER_3_1092 ();
 sg13g2_decap_8 FILLER_3_1099 ();
 sg13g2_decap_8 FILLER_3_1106 ();
 sg13g2_decap_8 FILLER_3_1113 ();
 sg13g2_decap_8 FILLER_3_1120 ();
 sg13g2_decap_8 FILLER_3_1127 ();
 sg13g2_decap_8 FILLER_3_1134 ();
 sg13g2_decap_8 FILLER_3_1141 ();
 sg13g2_decap_8 FILLER_3_1148 ();
 sg13g2_decap_8 FILLER_3_1155 ();
 sg13g2_decap_8 FILLER_3_1162 ();
 sg13g2_decap_8 FILLER_3_1169 ();
 sg13g2_decap_8 FILLER_3_1176 ();
 sg13g2_decap_8 FILLER_3_1183 ();
 sg13g2_decap_8 FILLER_3_1190 ();
 sg13g2_decap_8 FILLER_3_1197 ();
 sg13g2_decap_8 FILLER_3_1204 ();
 sg13g2_decap_8 FILLER_3_1211 ();
 sg13g2_decap_8 FILLER_3_1218 ();
 sg13g2_decap_8 FILLER_3_1225 ();
 sg13g2_decap_8 FILLER_3_1232 ();
 sg13g2_decap_8 FILLER_3_1239 ();
 sg13g2_decap_8 FILLER_3_1246 ();
 sg13g2_decap_8 FILLER_3_1253 ();
 sg13g2_decap_8 FILLER_3_1260 ();
 sg13g2_decap_8 FILLER_3_1267 ();
 sg13g2_decap_8 FILLER_3_1274 ();
 sg13g2_decap_8 FILLER_3_1281 ();
 sg13g2_decap_8 FILLER_3_1288 ();
 sg13g2_decap_8 FILLER_3_1295 ();
 sg13g2_decap_8 FILLER_3_1302 ();
 sg13g2_decap_8 FILLER_3_1309 ();
 sg13g2_decap_8 FILLER_3_1316 ();
 sg13g2_fill_2 FILLER_3_1323 ();
 sg13g2_fill_1 FILLER_3_1325 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_245 ();
 sg13g2_fill_2 FILLER_4_340 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_451 ();
 sg13g2_fill_2 FILLER_4_480 ();
 sg13g2_fill_1 FILLER_4_534 ();
 sg13g2_fill_2 FILLER_4_575 ();
 sg13g2_fill_1 FILLER_4_577 ();
 sg13g2_fill_2 FILLER_4_632 ();
 sg13g2_fill_2 FILLER_4_670 ();
 sg13g2_fill_1 FILLER_4_672 ();
 sg13g2_fill_2 FILLER_4_749 ();
 sg13g2_fill_2 FILLER_4_787 ();
 sg13g2_fill_1 FILLER_4_853 ();
 sg13g2_fill_2 FILLER_4_904 ();
 sg13g2_fill_2 FILLER_4_928 ();
 sg13g2_fill_1 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_decap_8 FILLER_4_1026 ();
 sg13g2_decap_8 FILLER_4_1033 ();
 sg13g2_decap_8 FILLER_4_1040 ();
 sg13g2_decap_8 FILLER_4_1047 ();
 sg13g2_decap_8 FILLER_4_1054 ();
 sg13g2_decap_8 FILLER_4_1061 ();
 sg13g2_decap_8 FILLER_4_1068 ();
 sg13g2_decap_8 FILLER_4_1075 ();
 sg13g2_decap_8 FILLER_4_1082 ();
 sg13g2_decap_8 FILLER_4_1089 ();
 sg13g2_decap_8 FILLER_4_1096 ();
 sg13g2_decap_8 FILLER_4_1103 ();
 sg13g2_decap_8 FILLER_4_1110 ();
 sg13g2_decap_8 FILLER_4_1117 ();
 sg13g2_decap_8 FILLER_4_1124 ();
 sg13g2_decap_8 FILLER_4_1131 ();
 sg13g2_decap_8 FILLER_4_1138 ();
 sg13g2_decap_8 FILLER_4_1145 ();
 sg13g2_decap_8 FILLER_4_1152 ();
 sg13g2_decap_8 FILLER_4_1159 ();
 sg13g2_decap_8 FILLER_4_1166 ();
 sg13g2_decap_8 FILLER_4_1173 ();
 sg13g2_decap_8 FILLER_4_1180 ();
 sg13g2_decap_8 FILLER_4_1187 ();
 sg13g2_decap_8 FILLER_4_1194 ();
 sg13g2_decap_8 FILLER_4_1201 ();
 sg13g2_decap_8 FILLER_4_1208 ();
 sg13g2_decap_8 FILLER_4_1215 ();
 sg13g2_decap_8 FILLER_4_1222 ();
 sg13g2_decap_8 FILLER_4_1229 ();
 sg13g2_decap_8 FILLER_4_1236 ();
 sg13g2_decap_8 FILLER_4_1243 ();
 sg13g2_decap_8 FILLER_4_1250 ();
 sg13g2_decap_8 FILLER_4_1257 ();
 sg13g2_decap_8 FILLER_4_1264 ();
 sg13g2_decap_8 FILLER_4_1271 ();
 sg13g2_decap_8 FILLER_4_1278 ();
 sg13g2_decap_8 FILLER_4_1285 ();
 sg13g2_decap_8 FILLER_4_1292 ();
 sg13g2_decap_8 FILLER_4_1299 ();
 sg13g2_decap_8 FILLER_4_1306 ();
 sg13g2_decap_8 FILLER_4_1313 ();
 sg13g2_decap_4 FILLER_4_1320 ();
 sg13g2_fill_2 FILLER_4_1324 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_fill_2 FILLER_5_382 ();
 sg13g2_fill_1 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_425 ();
 sg13g2_fill_2 FILLER_5_452 ();
 sg13g2_fill_1 FILLER_5_454 ();
 sg13g2_fill_2 FILLER_5_511 ();
 sg13g2_fill_2 FILLER_5_563 ();
 sg13g2_fill_1 FILLER_5_565 ();
 sg13g2_fill_2 FILLER_5_584 ();
 sg13g2_fill_1 FILLER_5_586 ();
 sg13g2_fill_1 FILLER_5_705 ();
 sg13g2_fill_1 FILLER_5_710 ();
 sg13g2_fill_2 FILLER_5_730 ();
 sg13g2_fill_1 FILLER_5_732 ();
 sg13g2_fill_1 FILLER_5_759 ();
 sg13g2_fill_2 FILLER_5_866 ();
 sg13g2_fill_2 FILLER_5_904 ();
 sg13g2_decap_8 FILLER_5_944 ();
 sg13g2_decap_8 FILLER_5_951 ();
 sg13g2_decap_8 FILLER_5_958 ();
 sg13g2_decap_8 FILLER_5_965 ();
 sg13g2_decap_8 FILLER_5_972 ();
 sg13g2_decap_8 FILLER_5_979 ();
 sg13g2_decap_8 FILLER_5_986 ();
 sg13g2_decap_8 FILLER_5_993 ();
 sg13g2_decap_8 FILLER_5_1000 ();
 sg13g2_decap_8 FILLER_5_1007 ();
 sg13g2_decap_8 FILLER_5_1014 ();
 sg13g2_decap_8 FILLER_5_1021 ();
 sg13g2_decap_8 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_5_1035 ();
 sg13g2_decap_8 FILLER_5_1042 ();
 sg13g2_decap_8 FILLER_5_1049 ();
 sg13g2_decap_8 FILLER_5_1056 ();
 sg13g2_decap_8 FILLER_5_1063 ();
 sg13g2_decap_8 FILLER_5_1070 ();
 sg13g2_decap_8 FILLER_5_1077 ();
 sg13g2_decap_8 FILLER_5_1084 ();
 sg13g2_decap_8 FILLER_5_1091 ();
 sg13g2_decap_8 FILLER_5_1098 ();
 sg13g2_decap_8 FILLER_5_1105 ();
 sg13g2_decap_8 FILLER_5_1112 ();
 sg13g2_decap_8 FILLER_5_1119 ();
 sg13g2_decap_8 FILLER_5_1126 ();
 sg13g2_decap_8 FILLER_5_1133 ();
 sg13g2_decap_8 FILLER_5_1140 ();
 sg13g2_decap_8 FILLER_5_1147 ();
 sg13g2_decap_8 FILLER_5_1154 ();
 sg13g2_decap_8 FILLER_5_1161 ();
 sg13g2_decap_8 FILLER_5_1168 ();
 sg13g2_decap_8 FILLER_5_1175 ();
 sg13g2_decap_8 FILLER_5_1182 ();
 sg13g2_decap_8 FILLER_5_1189 ();
 sg13g2_decap_8 FILLER_5_1196 ();
 sg13g2_decap_8 FILLER_5_1203 ();
 sg13g2_decap_8 FILLER_5_1210 ();
 sg13g2_decap_8 FILLER_5_1217 ();
 sg13g2_decap_8 FILLER_5_1224 ();
 sg13g2_decap_8 FILLER_5_1231 ();
 sg13g2_decap_8 FILLER_5_1238 ();
 sg13g2_decap_8 FILLER_5_1245 ();
 sg13g2_decap_8 FILLER_5_1252 ();
 sg13g2_decap_8 FILLER_5_1259 ();
 sg13g2_decap_8 FILLER_5_1266 ();
 sg13g2_decap_8 FILLER_5_1273 ();
 sg13g2_decap_8 FILLER_5_1280 ();
 sg13g2_decap_8 FILLER_5_1287 ();
 sg13g2_decap_8 FILLER_5_1294 ();
 sg13g2_decap_8 FILLER_5_1301 ();
 sg13g2_decap_8 FILLER_5_1308 ();
 sg13g2_decap_8 FILLER_5_1315 ();
 sg13g2_decap_4 FILLER_5_1322 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_231 ();
 sg13g2_fill_2 FILLER_6_240 ();
 sg13g2_fill_1 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_364 ();
 sg13g2_fill_1 FILLER_6_375 ();
 sg13g2_fill_1 FILLER_6_424 ();
 sg13g2_fill_1 FILLER_6_447 ();
 sg13g2_fill_1 FILLER_6_514 ();
 sg13g2_fill_2 FILLER_6_662 ();
 sg13g2_fill_1 FILLER_6_664 ();
 sg13g2_fill_1 FILLER_6_675 ();
 sg13g2_fill_1 FILLER_6_702 ();
 sg13g2_fill_2 FILLER_6_729 ();
 sg13g2_fill_2 FILLER_6_771 ();
 sg13g2_fill_1 FILLER_6_773 ();
 sg13g2_fill_2 FILLER_6_826 ();
 sg13g2_fill_2 FILLER_6_866 ();
 sg13g2_fill_2 FILLER_6_878 ();
 sg13g2_fill_2 FILLER_6_902 ();
 sg13g2_fill_1 FILLER_6_904 ();
 sg13g2_decap_8 FILLER_6_955 ();
 sg13g2_decap_8 FILLER_6_962 ();
 sg13g2_decap_8 FILLER_6_969 ();
 sg13g2_decap_8 FILLER_6_976 ();
 sg13g2_decap_8 FILLER_6_983 ();
 sg13g2_decap_8 FILLER_6_990 ();
 sg13g2_decap_8 FILLER_6_997 ();
 sg13g2_decap_8 FILLER_6_1004 ();
 sg13g2_decap_8 FILLER_6_1011 ();
 sg13g2_decap_8 FILLER_6_1018 ();
 sg13g2_decap_8 FILLER_6_1025 ();
 sg13g2_decap_8 FILLER_6_1032 ();
 sg13g2_decap_8 FILLER_6_1039 ();
 sg13g2_decap_8 FILLER_6_1046 ();
 sg13g2_decap_8 FILLER_6_1053 ();
 sg13g2_decap_8 FILLER_6_1060 ();
 sg13g2_decap_8 FILLER_6_1067 ();
 sg13g2_decap_8 FILLER_6_1074 ();
 sg13g2_decap_8 FILLER_6_1081 ();
 sg13g2_decap_8 FILLER_6_1088 ();
 sg13g2_decap_8 FILLER_6_1095 ();
 sg13g2_decap_8 FILLER_6_1102 ();
 sg13g2_decap_8 FILLER_6_1109 ();
 sg13g2_decap_8 FILLER_6_1116 ();
 sg13g2_decap_8 FILLER_6_1123 ();
 sg13g2_decap_8 FILLER_6_1130 ();
 sg13g2_decap_8 FILLER_6_1137 ();
 sg13g2_decap_8 FILLER_6_1144 ();
 sg13g2_decap_8 FILLER_6_1151 ();
 sg13g2_decap_8 FILLER_6_1158 ();
 sg13g2_decap_8 FILLER_6_1165 ();
 sg13g2_decap_8 FILLER_6_1172 ();
 sg13g2_decap_8 FILLER_6_1179 ();
 sg13g2_decap_8 FILLER_6_1186 ();
 sg13g2_decap_8 FILLER_6_1193 ();
 sg13g2_decap_8 FILLER_6_1200 ();
 sg13g2_decap_8 FILLER_6_1207 ();
 sg13g2_decap_8 FILLER_6_1214 ();
 sg13g2_decap_8 FILLER_6_1221 ();
 sg13g2_decap_8 FILLER_6_1228 ();
 sg13g2_decap_8 FILLER_6_1235 ();
 sg13g2_decap_8 FILLER_6_1242 ();
 sg13g2_decap_8 FILLER_6_1249 ();
 sg13g2_decap_8 FILLER_6_1256 ();
 sg13g2_decap_8 FILLER_6_1263 ();
 sg13g2_decap_8 FILLER_6_1270 ();
 sg13g2_decap_8 FILLER_6_1277 ();
 sg13g2_decap_8 FILLER_6_1284 ();
 sg13g2_decap_8 FILLER_6_1291 ();
 sg13g2_decap_8 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1305 ();
 sg13g2_decap_8 FILLER_6_1312 ();
 sg13g2_decap_8 FILLER_6_1319 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_293 ();
 sg13g2_fill_1 FILLER_7_440 ();
 sg13g2_fill_1 FILLER_7_467 ();
 sg13g2_fill_2 FILLER_7_478 ();
 sg13g2_fill_2 FILLER_7_488 ();
 sg13g2_fill_1 FILLER_7_490 ();
 sg13g2_fill_2 FILLER_7_537 ();
 sg13g2_fill_1 FILLER_7_539 ();
 sg13g2_fill_1 FILLER_7_644 ();
 sg13g2_fill_2 FILLER_7_681 ();
 sg13g2_fill_2 FILLER_7_745 ();
 sg13g2_fill_1 FILLER_7_805 ();
 sg13g2_fill_2 FILLER_7_832 ();
 sg13g2_fill_2 FILLER_7_844 ();
 sg13g2_fill_2 FILLER_7_856 ();
 sg13g2_fill_1 FILLER_7_858 ();
 sg13g2_fill_2 FILLER_7_927 ();
 sg13g2_fill_1 FILLER_7_939 ();
 sg13g2_fill_2 FILLER_7_962 ();
 sg13g2_decap_8 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_993 ();
 sg13g2_decap_8 FILLER_7_1000 ();
 sg13g2_decap_8 FILLER_7_1007 ();
 sg13g2_decap_8 FILLER_7_1014 ();
 sg13g2_decap_8 FILLER_7_1021 ();
 sg13g2_decap_8 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_7_1035 ();
 sg13g2_decap_8 FILLER_7_1042 ();
 sg13g2_decap_8 FILLER_7_1049 ();
 sg13g2_decap_8 FILLER_7_1056 ();
 sg13g2_decap_8 FILLER_7_1063 ();
 sg13g2_decap_8 FILLER_7_1070 ();
 sg13g2_decap_8 FILLER_7_1077 ();
 sg13g2_decap_8 FILLER_7_1084 ();
 sg13g2_decap_8 FILLER_7_1091 ();
 sg13g2_decap_8 FILLER_7_1098 ();
 sg13g2_decap_8 FILLER_7_1105 ();
 sg13g2_decap_8 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1119 ();
 sg13g2_decap_8 FILLER_7_1126 ();
 sg13g2_decap_8 FILLER_7_1133 ();
 sg13g2_decap_8 FILLER_7_1140 ();
 sg13g2_decap_8 FILLER_7_1147 ();
 sg13g2_decap_8 FILLER_7_1154 ();
 sg13g2_decap_8 FILLER_7_1161 ();
 sg13g2_decap_8 FILLER_7_1168 ();
 sg13g2_decap_8 FILLER_7_1175 ();
 sg13g2_decap_8 FILLER_7_1182 ();
 sg13g2_decap_8 FILLER_7_1189 ();
 sg13g2_decap_8 FILLER_7_1196 ();
 sg13g2_decap_8 FILLER_7_1203 ();
 sg13g2_decap_8 FILLER_7_1210 ();
 sg13g2_decap_8 FILLER_7_1217 ();
 sg13g2_decap_8 FILLER_7_1224 ();
 sg13g2_decap_8 FILLER_7_1231 ();
 sg13g2_decap_8 FILLER_7_1238 ();
 sg13g2_decap_8 FILLER_7_1245 ();
 sg13g2_decap_8 FILLER_7_1252 ();
 sg13g2_decap_8 FILLER_7_1259 ();
 sg13g2_decap_8 FILLER_7_1266 ();
 sg13g2_decap_8 FILLER_7_1273 ();
 sg13g2_decap_8 FILLER_7_1280 ();
 sg13g2_decap_8 FILLER_7_1287 ();
 sg13g2_decap_8 FILLER_7_1294 ();
 sg13g2_decap_8 FILLER_7_1301 ();
 sg13g2_decap_8 FILLER_7_1308 ();
 sg13g2_decap_8 FILLER_7_1315 ();
 sg13g2_decap_4 FILLER_7_1322 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_1 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_fill_1 FILLER_8_275 ();
 sg13g2_fill_2 FILLER_8_286 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_fill_1 FILLER_8_386 ();
 sg13g2_fill_1 FILLER_8_445 ();
 sg13g2_fill_1 FILLER_8_456 ();
 sg13g2_fill_1 FILLER_8_507 ();
 sg13g2_fill_1 FILLER_8_584 ();
 sg13g2_fill_2 FILLER_8_657 ();
 sg13g2_fill_1 FILLER_8_729 ();
 sg13g2_fill_2 FILLER_8_793 ();
 sg13g2_fill_2 FILLER_8_831 ();
 sg13g2_fill_1 FILLER_8_833 ();
 sg13g2_fill_1 FILLER_8_860 ();
 sg13g2_fill_2 FILLER_8_891 ();
 sg13g2_fill_1 FILLER_8_893 ();
 sg13g2_fill_2 FILLER_8_920 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_decap_8 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_8_1035 ();
 sg13g2_decap_8 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1049 ();
 sg13g2_decap_8 FILLER_8_1056 ();
 sg13g2_decap_8 FILLER_8_1063 ();
 sg13g2_decap_8 FILLER_8_1070 ();
 sg13g2_decap_8 FILLER_8_1077 ();
 sg13g2_decap_8 FILLER_8_1084 ();
 sg13g2_decap_8 FILLER_8_1091 ();
 sg13g2_decap_8 FILLER_8_1098 ();
 sg13g2_decap_8 FILLER_8_1105 ();
 sg13g2_decap_8 FILLER_8_1112 ();
 sg13g2_decap_8 FILLER_8_1119 ();
 sg13g2_decap_8 FILLER_8_1126 ();
 sg13g2_decap_8 FILLER_8_1133 ();
 sg13g2_decap_8 FILLER_8_1140 ();
 sg13g2_decap_8 FILLER_8_1147 ();
 sg13g2_decap_8 FILLER_8_1154 ();
 sg13g2_decap_8 FILLER_8_1161 ();
 sg13g2_decap_8 FILLER_8_1168 ();
 sg13g2_decap_8 FILLER_8_1175 ();
 sg13g2_decap_8 FILLER_8_1182 ();
 sg13g2_decap_8 FILLER_8_1189 ();
 sg13g2_decap_8 FILLER_8_1196 ();
 sg13g2_decap_8 FILLER_8_1203 ();
 sg13g2_decap_8 FILLER_8_1210 ();
 sg13g2_decap_8 FILLER_8_1217 ();
 sg13g2_decap_8 FILLER_8_1224 ();
 sg13g2_decap_8 FILLER_8_1231 ();
 sg13g2_decap_8 FILLER_8_1238 ();
 sg13g2_decap_8 FILLER_8_1245 ();
 sg13g2_decap_8 FILLER_8_1252 ();
 sg13g2_decap_8 FILLER_8_1259 ();
 sg13g2_decap_8 FILLER_8_1266 ();
 sg13g2_decap_8 FILLER_8_1273 ();
 sg13g2_decap_8 FILLER_8_1280 ();
 sg13g2_decap_8 FILLER_8_1287 ();
 sg13g2_decap_8 FILLER_8_1294 ();
 sg13g2_decap_8 FILLER_8_1301 ();
 sg13g2_decap_8 FILLER_8_1308 ();
 sg13g2_decap_8 FILLER_8_1315 ();
 sg13g2_decap_4 FILLER_8_1322 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_4 FILLER_9_203 ();
 sg13g2_fill_2 FILLER_9_211 ();
 sg13g2_fill_1 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_334 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_fill_1 FILLER_9_348 ();
 sg13g2_fill_1 FILLER_9_430 ();
 sg13g2_fill_1 FILLER_9_441 ();
 sg13g2_fill_1 FILLER_9_468 ();
 sg13g2_fill_2 FILLER_9_503 ();
 sg13g2_fill_2 FILLER_9_551 ();
 sg13g2_fill_2 FILLER_9_605 ();
 sg13g2_fill_1 FILLER_9_607 ();
 sg13g2_fill_2 FILLER_9_680 ();
 sg13g2_fill_1 FILLER_9_682 ();
 sg13g2_fill_2 FILLER_9_717 ();
 sg13g2_fill_1 FILLER_9_745 ();
 sg13g2_fill_2 FILLER_9_831 ();
 sg13g2_fill_2 FILLER_9_841 ();
 sg13g2_fill_2 FILLER_9_861 ();
 sg13g2_fill_1 FILLER_9_863 ();
 sg13g2_fill_1 FILLER_9_904 ();
 sg13g2_fill_2 FILLER_9_961 ();
 sg13g2_decap_8 FILLER_9_1003 ();
 sg13g2_decap_8 FILLER_9_1010 ();
 sg13g2_decap_8 FILLER_9_1017 ();
 sg13g2_decap_8 FILLER_9_1024 ();
 sg13g2_decap_8 FILLER_9_1031 ();
 sg13g2_decap_8 FILLER_9_1038 ();
 sg13g2_decap_8 FILLER_9_1045 ();
 sg13g2_decap_8 FILLER_9_1052 ();
 sg13g2_decap_8 FILLER_9_1059 ();
 sg13g2_decap_8 FILLER_9_1066 ();
 sg13g2_decap_8 FILLER_9_1073 ();
 sg13g2_decap_8 FILLER_9_1080 ();
 sg13g2_decap_8 FILLER_9_1087 ();
 sg13g2_decap_8 FILLER_9_1094 ();
 sg13g2_decap_8 FILLER_9_1101 ();
 sg13g2_decap_8 FILLER_9_1108 ();
 sg13g2_decap_8 FILLER_9_1115 ();
 sg13g2_decap_8 FILLER_9_1122 ();
 sg13g2_decap_8 FILLER_9_1129 ();
 sg13g2_decap_8 FILLER_9_1136 ();
 sg13g2_decap_8 FILLER_9_1143 ();
 sg13g2_decap_8 FILLER_9_1150 ();
 sg13g2_decap_8 FILLER_9_1157 ();
 sg13g2_decap_8 FILLER_9_1164 ();
 sg13g2_decap_8 FILLER_9_1171 ();
 sg13g2_decap_8 FILLER_9_1178 ();
 sg13g2_decap_8 FILLER_9_1185 ();
 sg13g2_decap_8 FILLER_9_1192 ();
 sg13g2_decap_8 FILLER_9_1199 ();
 sg13g2_decap_8 FILLER_9_1206 ();
 sg13g2_decap_8 FILLER_9_1213 ();
 sg13g2_decap_8 FILLER_9_1220 ();
 sg13g2_decap_8 FILLER_9_1227 ();
 sg13g2_decap_8 FILLER_9_1234 ();
 sg13g2_decap_8 FILLER_9_1241 ();
 sg13g2_decap_8 FILLER_9_1248 ();
 sg13g2_decap_8 FILLER_9_1255 ();
 sg13g2_decap_8 FILLER_9_1262 ();
 sg13g2_decap_8 FILLER_9_1269 ();
 sg13g2_decap_8 FILLER_9_1276 ();
 sg13g2_decap_8 FILLER_9_1283 ();
 sg13g2_decap_8 FILLER_9_1290 ();
 sg13g2_decap_8 FILLER_9_1297 ();
 sg13g2_decap_8 FILLER_9_1304 ();
 sg13g2_decap_8 FILLER_9_1311 ();
 sg13g2_decap_8 FILLER_9_1318 ();
 sg13g2_fill_1 FILLER_9_1325 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_4 FILLER_10_189 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_2 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_379 ();
 sg13g2_fill_1 FILLER_10_436 ();
 sg13g2_fill_2 FILLER_10_477 ();
 sg13g2_fill_2 FILLER_10_489 ();
 sg13g2_fill_1 FILLER_10_491 ();
 sg13g2_fill_1 FILLER_10_518 ();
 sg13g2_fill_2 FILLER_10_568 ();
 sg13g2_fill_1 FILLER_10_570 ();
 sg13g2_fill_2 FILLER_10_591 ();
 sg13g2_fill_1 FILLER_10_593 ();
 sg13g2_fill_1 FILLER_10_650 ();
 sg13g2_fill_2 FILLER_10_749 ();
 sg13g2_fill_2 FILLER_10_769 ();
 sg13g2_fill_1 FILLER_10_775 ();
 sg13g2_fill_1 FILLER_10_790 ();
 sg13g2_fill_2 FILLER_10_805 ();
 sg13g2_fill_2 FILLER_10_821 ();
 sg13g2_fill_1 FILLER_10_849 ();
 sg13g2_fill_2 FILLER_10_888 ();
 sg13g2_fill_1 FILLER_10_890 ();
 sg13g2_fill_1 FILLER_10_905 ();
 sg13g2_fill_2 FILLER_10_924 ();
 sg13g2_fill_1 FILLER_10_978 ();
 sg13g2_decap_8 FILLER_10_1009 ();
 sg13g2_decap_8 FILLER_10_1016 ();
 sg13g2_decap_8 FILLER_10_1023 ();
 sg13g2_decap_8 FILLER_10_1030 ();
 sg13g2_decap_8 FILLER_10_1037 ();
 sg13g2_decap_8 FILLER_10_1044 ();
 sg13g2_decap_8 FILLER_10_1051 ();
 sg13g2_decap_8 FILLER_10_1058 ();
 sg13g2_decap_8 FILLER_10_1065 ();
 sg13g2_decap_8 FILLER_10_1072 ();
 sg13g2_decap_8 FILLER_10_1079 ();
 sg13g2_decap_8 FILLER_10_1086 ();
 sg13g2_decap_8 FILLER_10_1093 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_8 FILLER_10_1107 ();
 sg13g2_decap_8 FILLER_10_1114 ();
 sg13g2_decap_8 FILLER_10_1121 ();
 sg13g2_decap_8 FILLER_10_1128 ();
 sg13g2_decap_8 FILLER_10_1135 ();
 sg13g2_decap_8 FILLER_10_1142 ();
 sg13g2_decap_8 FILLER_10_1149 ();
 sg13g2_decap_8 FILLER_10_1156 ();
 sg13g2_decap_8 FILLER_10_1163 ();
 sg13g2_decap_8 FILLER_10_1170 ();
 sg13g2_decap_8 FILLER_10_1177 ();
 sg13g2_decap_8 FILLER_10_1184 ();
 sg13g2_decap_8 FILLER_10_1191 ();
 sg13g2_decap_8 FILLER_10_1198 ();
 sg13g2_decap_8 FILLER_10_1205 ();
 sg13g2_decap_8 FILLER_10_1212 ();
 sg13g2_decap_8 FILLER_10_1219 ();
 sg13g2_decap_8 FILLER_10_1226 ();
 sg13g2_decap_8 FILLER_10_1233 ();
 sg13g2_decap_8 FILLER_10_1240 ();
 sg13g2_decap_8 FILLER_10_1247 ();
 sg13g2_decap_8 FILLER_10_1254 ();
 sg13g2_decap_8 FILLER_10_1261 ();
 sg13g2_decap_8 FILLER_10_1268 ();
 sg13g2_decap_8 FILLER_10_1275 ();
 sg13g2_decap_8 FILLER_10_1282 ();
 sg13g2_decap_8 FILLER_10_1289 ();
 sg13g2_decap_8 FILLER_10_1296 ();
 sg13g2_decap_8 FILLER_10_1303 ();
 sg13g2_decap_8 FILLER_10_1310 ();
 sg13g2_decap_8 FILLER_10_1317 ();
 sg13g2_fill_2 FILLER_10_1324 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_189 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_236 ();
 sg13g2_fill_2 FILLER_11_281 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_fill_2 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_11_513 ();
 sg13g2_fill_1 FILLER_11_540 ();
 sg13g2_fill_1 FILLER_11_613 ();
 sg13g2_fill_1 FILLER_11_624 ();
 sg13g2_fill_1 FILLER_11_635 ();
 sg13g2_fill_1 FILLER_11_641 ();
 sg13g2_fill_2 FILLER_11_720 ();
 sg13g2_fill_1 FILLER_11_758 ();
 sg13g2_fill_1 FILLER_11_785 ();
 sg13g2_fill_1 FILLER_11_838 ();
 sg13g2_fill_1 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_884 ();
 sg13g2_fill_1 FILLER_11_925 ();
 sg13g2_fill_2 FILLER_11_950 ();
 sg13g2_fill_2 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1004 ();
 sg13g2_decap_8 FILLER_11_1011 ();
 sg13g2_decap_8 FILLER_11_1018 ();
 sg13g2_decap_8 FILLER_11_1025 ();
 sg13g2_decap_8 FILLER_11_1032 ();
 sg13g2_decap_8 FILLER_11_1039 ();
 sg13g2_decap_8 FILLER_11_1046 ();
 sg13g2_decap_8 FILLER_11_1053 ();
 sg13g2_decap_8 FILLER_11_1060 ();
 sg13g2_decap_8 FILLER_11_1067 ();
 sg13g2_decap_8 FILLER_11_1074 ();
 sg13g2_decap_8 FILLER_11_1081 ();
 sg13g2_decap_8 FILLER_11_1088 ();
 sg13g2_decap_8 FILLER_11_1095 ();
 sg13g2_decap_8 FILLER_11_1102 ();
 sg13g2_decap_8 FILLER_11_1109 ();
 sg13g2_decap_8 FILLER_11_1116 ();
 sg13g2_decap_8 FILLER_11_1123 ();
 sg13g2_decap_8 FILLER_11_1130 ();
 sg13g2_decap_8 FILLER_11_1137 ();
 sg13g2_decap_8 FILLER_11_1144 ();
 sg13g2_decap_8 FILLER_11_1151 ();
 sg13g2_decap_8 FILLER_11_1158 ();
 sg13g2_decap_8 FILLER_11_1165 ();
 sg13g2_decap_8 FILLER_11_1172 ();
 sg13g2_decap_8 FILLER_11_1179 ();
 sg13g2_decap_8 FILLER_11_1186 ();
 sg13g2_decap_8 FILLER_11_1193 ();
 sg13g2_decap_8 FILLER_11_1200 ();
 sg13g2_decap_8 FILLER_11_1207 ();
 sg13g2_decap_8 FILLER_11_1214 ();
 sg13g2_decap_8 FILLER_11_1221 ();
 sg13g2_decap_8 FILLER_11_1228 ();
 sg13g2_decap_8 FILLER_11_1235 ();
 sg13g2_decap_8 FILLER_11_1242 ();
 sg13g2_decap_8 FILLER_11_1249 ();
 sg13g2_decap_8 FILLER_11_1256 ();
 sg13g2_decap_8 FILLER_11_1263 ();
 sg13g2_decap_8 FILLER_11_1270 ();
 sg13g2_decap_8 FILLER_11_1277 ();
 sg13g2_decap_8 FILLER_11_1284 ();
 sg13g2_decap_8 FILLER_11_1291 ();
 sg13g2_decap_8 FILLER_11_1298 ();
 sg13g2_decap_8 FILLER_11_1305 ();
 sg13g2_decap_8 FILLER_11_1312 ();
 sg13g2_decap_8 FILLER_11_1319 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_182 ();
 sg13g2_fill_1 FILLER_12_186 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_303 ();
 sg13g2_fill_2 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_422 ();
 sg13g2_fill_1 FILLER_12_540 ();
 sg13g2_fill_1 FILLER_12_549 ();
 sg13g2_fill_2 FILLER_12_600 ();
 sg13g2_fill_1 FILLER_12_602 ();
 sg13g2_fill_2 FILLER_12_677 ();
 sg13g2_fill_1 FILLER_12_705 ();
 sg13g2_fill_1 FILLER_12_716 ();
 sg13g2_fill_1 FILLER_12_743 ();
 sg13g2_fill_1 FILLER_12_756 ();
 sg13g2_fill_2 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_12_835 ();
 sg13g2_fill_2 FILLER_12_846 ();
 sg13g2_fill_2 FILLER_12_856 ();
 sg13g2_fill_1 FILLER_12_858 ();
 sg13g2_fill_1 FILLER_12_885 ();
 sg13g2_fill_2 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_1008 ();
 sg13g2_decap_8 FILLER_12_1015 ();
 sg13g2_decap_8 FILLER_12_1022 ();
 sg13g2_decap_8 FILLER_12_1029 ();
 sg13g2_decap_8 FILLER_12_1036 ();
 sg13g2_decap_8 FILLER_12_1043 ();
 sg13g2_decap_8 FILLER_12_1050 ();
 sg13g2_decap_8 FILLER_12_1057 ();
 sg13g2_decap_8 FILLER_12_1064 ();
 sg13g2_decap_8 FILLER_12_1071 ();
 sg13g2_decap_8 FILLER_12_1078 ();
 sg13g2_decap_8 FILLER_12_1085 ();
 sg13g2_decap_8 FILLER_12_1092 ();
 sg13g2_decap_8 FILLER_12_1099 ();
 sg13g2_decap_8 FILLER_12_1106 ();
 sg13g2_decap_8 FILLER_12_1113 ();
 sg13g2_decap_8 FILLER_12_1120 ();
 sg13g2_decap_8 FILLER_12_1127 ();
 sg13g2_decap_8 FILLER_12_1134 ();
 sg13g2_decap_8 FILLER_12_1141 ();
 sg13g2_decap_8 FILLER_12_1148 ();
 sg13g2_decap_8 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1162 ();
 sg13g2_decap_8 FILLER_12_1169 ();
 sg13g2_decap_8 FILLER_12_1176 ();
 sg13g2_decap_8 FILLER_12_1183 ();
 sg13g2_decap_8 FILLER_12_1190 ();
 sg13g2_decap_8 FILLER_12_1197 ();
 sg13g2_decap_8 FILLER_12_1204 ();
 sg13g2_decap_8 FILLER_12_1211 ();
 sg13g2_decap_8 FILLER_12_1218 ();
 sg13g2_decap_8 FILLER_12_1225 ();
 sg13g2_decap_8 FILLER_12_1232 ();
 sg13g2_decap_8 FILLER_12_1239 ();
 sg13g2_decap_8 FILLER_12_1246 ();
 sg13g2_decap_8 FILLER_12_1253 ();
 sg13g2_decap_8 FILLER_12_1260 ();
 sg13g2_decap_8 FILLER_12_1267 ();
 sg13g2_decap_8 FILLER_12_1274 ();
 sg13g2_decap_8 FILLER_12_1281 ();
 sg13g2_decap_8 FILLER_12_1288 ();
 sg13g2_decap_8 FILLER_12_1295 ();
 sg13g2_decap_8 FILLER_12_1302 ();
 sg13g2_decap_8 FILLER_12_1309 ();
 sg13g2_decap_8 FILLER_12_1316 ();
 sg13g2_fill_2 FILLER_12_1323 ();
 sg13g2_fill_1 FILLER_12_1325 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_4 FILLER_13_175 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_373 ();
 sg13g2_fill_1 FILLER_13_435 ();
 sg13g2_fill_2 FILLER_13_462 ();
 sg13g2_fill_1 FILLER_13_464 ();
 sg13g2_fill_2 FILLER_13_533 ();
 sg13g2_fill_1 FILLER_13_535 ();
 sg13g2_fill_2 FILLER_13_576 ();
 sg13g2_fill_1 FILLER_13_578 ();
 sg13g2_fill_1 FILLER_13_615 ();
 sg13g2_fill_1 FILLER_13_650 ();
 sg13g2_fill_2 FILLER_13_677 ();
 sg13g2_fill_2 FILLER_13_693 ();
 sg13g2_fill_1 FILLER_13_695 ();
 sg13g2_fill_2 FILLER_13_793 ();
 sg13g2_fill_1 FILLER_13_894 ();
 sg13g2_fill_1 FILLER_13_905 ();
 sg13g2_fill_2 FILLER_13_916 ();
 sg13g2_fill_1 FILLER_13_928 ();
 sg13g2_fill_2 FILLER_13_955 ();
 sg13g2_decap_8 FILLER_13_1013 ();
 sg13g2_decap_8 FILLER_13_1020 ();
 sg13g2_decap_8 FILLER_13_1027 ();
 sg13g2_decap_8 FILLER_13_1034 ();
 sg13g2_decap_8 FILLER_13_1041 ();
 sg13g2_decap_8 FILLER_13_1048 ();
 sg13g2_decap_8 FILLER_13_1055 ();
 sg13g2_decap_8 FILLER_13_1062 ();
 sg13g2_decap_8 FILLER_13_1069 ();
 sg13g2_decap_8 FILLER_13_1076 ();
 sg13g2_decap_8 FILLER_13_1083 ();
 sg13g2_decap_8 FILLER_13_1090 ();
 sg13g2_decap_8 FILLER_13_1097 ();
 sg13g2_decap_8 FILLER_13_1104 ();
 sg13g2_decap_8 FILLER_13_1111 ();
 sg13g2_decap_8 FILLER_13_1118 ();
 sg13g2_decap_8 FILLER_13_1125 ();
 sg13g2_decap_8 FILLER_13_1132 ();
 sg13g2_decap_8 FILLER_13_1139 ();
 sg13g2_decap_8 FILLER_13_1146 ();
 sg13g2_decap_8 FILLER_13_1153 ();
 sg13g2_decap_8 FILLER_13_1160 ();
 sg13g2_decap_8 FILLER_13_1167 ();
 sg13g2_decap_8 FILLER_13_1174 ();
 sg13g2_decap_8 FILLER_13_1181 ();
 sg13g2_decap_8 FILLER_13_1188 ();
 sg13g2_decap_8 FILLER_13_1195 ();
 sg13g2_decap_8 FILLER_13_1202 ();
 sg13g2_decap_8 FILLER_13_1209 ();
 sg13g2_decap_8 FILLER_13_1216 ();
 sg13g2_decap_8 FILLER_13_1223 ();
 sg13g2_decap_8 FILLER_13_1230 ();
 sg13g2_decap_8 FILLER_13_1237 ();
 sg13g2_decap_8 FILLER_13_1244 ();
 sg13g2_decap_8 FILLER_13_1251 ();
 sg13g2_decap_8 FILLER_13_1258 ();
 sg13g2_decap_8 FILLER_13_1265 ();
 sg13g2_decap_8 FILLER_13_1272 ();
 sg13g2_decap_8 FILLER_13_1279 ();
 sg13g2_decap_8 FILLER_13_1286 ();
 sg13g2_decap_8 FILLER_13_1293 ();
 sg13g2_decap_8 FILLER_13_1300 ();
 sg13g2_decap_8 FILLER_13_1307 ();
 sg13g2_decap_8 FILLER_13_1314 ();
 sg13g2_decap_4 FILLER_13_1321 ();
 sg13g2_fill_1 FILLER_13_1325 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_175 ();
 sg13g2_fill_2 FILLER_14_237 ();
 sg13g2_fill_1 FILLER_14_249 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_fill_2 FILLER_14_409 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_fill_1 FILLER_14_438 ();
 sg13g2_fill_1 FILLER_14_525 ();
 sg13g2_fill_2 FILLER_14_603 ();
 sg13g2_fill_1 FILLER_14_605 ();
 sg13g2_fill_2 FILLER_14_616 ();
 sg13g2_fill_2 FILLER_14_628 ();
 sg13g2_fill_2 FILLER_14_682 ();
 sg13g2_fill_1 FILLER_14_684 ();
 sg13g2_fill_2 FILLER_14_721 ();
 sg13g2_fill_1 FILLER_14_723 ();
 sg13g2_fill_2 FILLER_14_782 ();
 sg13g2_fill_2 FILLER_14_830 ();
 sg13g2_fill_2 FILLER_14_858 ();
 sg13g2_fill_1 FILLER_14_860 ();
 sg13g2_fill_1 FILLER_14_906 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_decap_8 FILLER_14_1026 ();
 sg13g2_decap_8 FILLER_14_1033 ();
 sg13g2_decap_8 FILLER_14_1040 ();
 sg13g2_decap_8 FILLER_14_1047 ();
 sg13g2_decap_8 FILLER_14_1054 ();
 sg13g2_decap_8 FILLER_14_1061 ();
 sg13g2_decap_8 FILLER_14_1068 ();
 sg13g2_decap_8 FILLER_14_1075 ();
 sg13g2_decap_8 FILLER_14_1082 ();
 sg13g2_decap_8 FILLER_14_1089 ();
 sg13g2_decap_8 FILLER_14_1096 ();
 sg13g2_decap_8 FILLER_14_1103 ();
 sg13g2_decap_8 FILLER_14_1110 ();
 sg13g2_decap_8 FILLER_14_1117 ();
 sg13g2_decap_8 FILLER_14_1124 ();
 sg13g2_decap_8 FILLER_14_1131 ();
 sg13g2_decap_8 FILLER_14_1138 ();
 sg13g2_decap_8 FILLER_14_1145 ();
 sg13g2_decap_8 FILLER_14_1152 ();
 sg13g2_decap_8 FILLER_14_1159 ();
 sg13g2_decap_8 FILLER_14_1166 ();
 sg13g2_decap_8 FILLER_14_1173 ();
 sg13g2_decap_8 FILLER_14_1180 ();
 sg13g2_decap_8 FILLER_14_1187 ();
 sg13g2_decap_8 FILLER_14_1194 ();
 sg13g2_decap_8 FILLER_14_1201 ();
 sg13g2_decap_8 FILLER_14_1208 ();
 sg13g2_decap_8 FILLER_14_1215 ();
 sg13g2_decap_8 FILLER_14_1222 ();
 sg13g2_decap_8 FILLER_14_1229 ();
 sg13g2_decap_8 FILLER_14_1236 ();
 sg13g2_decap_8 FILLER_14_1243 ();
 sg13g2_decap_8 FILLER_14_1250 ();
 sg13g2_decap_8 FILLER_14_1257 ();
 sg13g2_decap_8 FILLER_14_1264 ();
 sg13g2_decap_8 FILLER_14_1271 ();
 sg13g2_decap_8 FILLER_14_1278 ();
 sg13g2_decap_8 FILLER_14_1285 ();
 sg13g2_decap_8 FILLER_14_1292 ();
 sg13g2_decap_8 FILLER_14_1299 ();
 sg13g2_decap_8 FILLER_14_1306 ();
 sg13g2_decap_8 FILLER_14_1313 ();
 sg13g2_decap_4 FILLER_14_1320 ();
 sg13g2_fill_2 FILLER_14_1324 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_248 ();
 sg13g2_fill_2 FILLER_15_280 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_328 ();
 sg13g2_fill_1 FILLER_15_339 ();
 sg13g2_fill_2 FILLER_15_388 ();
 sg13g2_fill_1 FILLER_15_390 ();
 sg13g2_fill_1 FILLER_15_453 ();
 sg13g2_fill_2 FILLER_15_512 ();
 sg13g2_fill_1 FILLER_15_548 ();
 sg13g2_fill_2 FILLER_15_559 ();
 sg13g2_fill_1 FILLER_15_561 ();
 sg13g2_fill_2 FILLER_15_616 ();
 sg13g2_fill_1 FILLER_15_644 ();
 sg13g2_decap_4 FILLER_15_655 ();
 sg13g2_fill_2 FILLER_15_699 ();
 sg13g2_fill_2 FILLER_15_805 ();
 sg13g2_fill_1 FILLER_15_841 ();
 sg13g2_fill_2 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_916 ();
 sg13g2_fill_2 FILLER_15_928 ();
 sg13g2_fill_1 FILLER_15_930 ();
 sg13g2_fill_2 FILLER_15_965 ();
 sg13g2_fill_2 FILLER_15_993 ();
 sg13g2_fill_1 FILLER_15_1009 ();
 sg13g2_decap_8 FILLER_15_1036 ();
 sg13g2_decap_8 FILLER_15_1043 ();
 sg13g2_decap_8 FILLER_15_1050 ();
 sg13g2_decap_8 FILLER_15_1057 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_decap_8 FILLER_15_1071 ();
 sg13g2_decap_8 FILLER_15_1078 ();
 sg13g2_decap_8 FILLER_15_1085 ();
 sg13g2_decap_8 FILLER_15_1092 ();
 sg13g2_decap_8 FILLER_15_1099 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1134 ();
 sg13g2_decap_8 FILLER_15_1141 ();
 sg13g2_decap_8 FILLER_15_1148 ();
 sg13g2_decap_8 FILLER_15_1155 ();
 sg13g2_decap_8 FILLER_15_1162 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_decap_8 FILLER_15_1176 ();
 sg13g2_decap_8 FILLER_15_1183 ();
 sg13g2_decap_8 FILLER_15_1190 ();
 sg13g2_decap_8 FILLER_15_1197 ();
 sg13g2_decap_8 FILLER_15_1204 ();
 sg13g2_decap_8 FILLER_15_1211 ();
 sg13g2_decap_8 FILLER_15_1218 ();
 sg13g2_decap_8 FILLER_15_1225 ();
 sg13g2_decap_8 FILLER_15_1232 ();
 sg13g2_decap_8 FILLER_15_1239 ();
 sg13g2_decap_8 FILLER_15_1246 ();
 sg13g2_decap_8 FILLER_15_1253 ();
 sg13g2_decap_8 FILLER_15_1260 ();
 sg13g2_decap_8 FILLER_15_1267 ();
 sg13g2_decap_8 FILLER_15_1274 ();
 sg13g2_decap_8 FILLER_15_1281 ();
 sg13g2_decap_8 FILLER_15_1288 ();
 sg13g2_decap_8 FILLER_15_1295 ();
 sg13g2_decap_8 FILLER_15_1302 ();
 sg13g2_decap_8 FILLER_15_1309 ();
 sg13g2_decap_8 FILLER_15_1316 ();
 sg13g2_fill_2 FILLER_15_1323 ();
 sg13g2_fill_1 FILLER_15_1325 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_fill_2 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_497 ();
 sg13g2_fill_2 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_564 ();
 sg13g2_fill_1 FILLER_16_591 ();
 sg13g2_fill_2 FILLER_16_668 ();
 sg13g2_fill_1 FILLER_16_670 ();
 sg13g2_fill_1 FILLER_16_689 ();
 sg13g2_fill_1 FILLER_16_765 ();
 sg13g2_fill_1 FILLER_16_776 ();
 sg13g2_fill_2 FILLER_16_839 ();
 sg13g2_fill_1 FILLER_16_841 ();
 sg13g2_fill_1 FILLER_16_856 ();
 sg13g2_fill_1 FILLER_16_883 ();
 sg13g2_fill_1 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_1031 ();
 sg13g2_decap_8 FILLER_16_1038 ();
 sg13g2_decap_8 FILLER_16_1045 ();
 sg13g2_decap_8 FILLER_16_1052 ();
 sg13g2_decap_8 FILLER_16_1059 ();
 sg13g2_decap_8 FILLER_16_1066 ();
 sg13g2_decap_8 FILLER_16_1073 ();
 sg13g2_decap_8 FILLER_16_1080 ();
 sg13g2_decap_8 FILLER_16_1087 ();
 sg13g2_decap_8 FILLER_16_1094 ();
 sg13g2_decap_8 FILLER_16_1101 ();
 sg13g2_decap_8 FILLER_16_1108 ();
 sg13g2_decap_8 FILLER_16_1115 ();
 sg13g2_decap_8 FILLER_16_1122 ();
 sg13g2_decap_8 FILLER_16_1129 ();
 sg13g2_decap_8 FILLER_16_1136 ();
 sg13g2_decap_8 FILLER_16_1143 ();
 sg13g2_decap_8 FILLER_16_1150 ();
 sg13g2_decap_8 FILLER_16_1157 ();
 sg13g2_decap_8 FILLER_16_1164 ();
 sg13g2_decap_8 FILLER_16_1171 ();
 sg13g2_decap_8 FILLER_16_1178 ();
 sg13g2_decap_8 FILLER_16_1185 ();
 sg13g2_decap_8 FILLER_16_1192 ();
 sg13g2_decap_8 FILLER_16_1199 ();
 sg13g2_decap_8 FILLER_16_1206 ();
 sg13g2_decap_8 FILLER_16_1213 ();
 sg13g2_decap_8 FILLER_16_1220 ();
 sg13g2_decap_8 FILLER_16_1227 ();
 sg13g2_decap_8 FILLER_16_1234 ();
 sg13g2_decap_8 FILLER_16_1241 ();
 sg13g2_decap_8 FILLER_16_1248 ();
 sg13g2_decap_8 FILLER_16_1255 ();
 sg13g2_decap_8 FILLER_16_1262 ();
 sg13g2_decap_8 FILLER_16_1269 ();
 sg13g2_decap_8 FILLER_16_1276 ();
 sg13g2_decap_8 FILLER_16_1283 ();
 sg13g2_decap_8 FILLER_16_1290 ();
 sg13g2_decap_8 FILLER_16_1297 ();
 sg13g2_decap_8 FILLER_16_1304 ();
 sg13g2_decap_8 FILLER_16_1311 ();
 sg13g2_decap_8 FILLER_16_1318 ();
 sg13g2_fill_1 FILLER_16_1325 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_147 ();
 sg13g2_fill_2 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_241 ();
 sg13g2_fill_1 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_399 ();
 sg13g2_fill_1 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_440 ();
 sg13g2_fill_1 FILLER_17_462 ();
 sg13g2_fill_1 FILLER_17_468 ();
 sg13g2_fill_1 FILLER_17_500 ();
 sg13g2_fill_2 FILLER_17_571 ();
 sg13g2_fill_1 FILLER_17_573 ();
 sg13g2_fill_2 FILLER_17_631 ();
 sg13g2_fill_1 FILLER_17_633 ();
 sg13g2_decap_4 FILLER_17_638 ();
 sg13g2_fill_1 FILLER_17_642 ();
 sg13g2_fill_1 FILLER_17_690 ();
 sg13g2_fill_2 FILLER_17_697 ();
 sg13g2_fill_1 FILLER_17_733 ();
 sg13g2_fill_1 FILLER_17_812 ();
 sg13g2_fill_1 FILLER_17_839 ();
 sg13g2_fill_2 FILLER_17_898 ();
 sg13g2_fill_1 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_1033 ();
 sg13g2_decap_8 FILLER_17_1040 ();
 sg13g2_decap_8 FILLER_17_1047 ();
 sg13g2_decap_8 FILLER_17_1054 ();
 sg13g2_decap_8 FILLER_17_1061 ();
 sg13g2_decap_8 FILLER_17_1068 ();
 sg13g2_decap_8 FILLER_17_1075 ();
 sg13g2_decap_8 FILLER_17_1082 ();
 sg13g2_decap_8 FILLER_17_1089 ();
 sg13g2_decap_8 FILLER_17_1096 ();
 sg13g2_decap_8 FILLER_17_1103 ();
 sg13g2_decap_8 FILLER_17_1110 ();
 sg13g2_decap_8 FILLER_17_1117 ();
 sg13g2_decap_8 FILLER_17_1124 ();
 sg13g2_decap_8 FILLER_17_1131 ();
 sg13g2_decap_8 FILLER_17_1138 ();
 sg13g2_decap_8 FILLER_17_1145 ();
 sg13g2_decap_8 FILLER_17_1152 ();
 sg13g2_decap_8 FILLER_17_1159 ();
 sg13g2_decap_8 FILLER_17_1166 ();
 sg13g2_decap_8 FILLER_17_1173 ();
 sg13g2_decap_8 FILLER_17_1180 ();
 sg13g2_decap_8 FILLER_17_1187 ();
 sg13g2_decap_8 FILLER_17_1194 ();
 sg13g2_decap_8 FILLER_17_1201 ();
 sg13g2_decap_8 FILLER_17_1208 ();
 sg13g2_decap_8 FILLER_17_1215 ();
 sg13g2_decap_8 FILLER_17_1222 ();
 sg13g2_decap_8 FILLER_17_1229 ();
 sg13g2_decap_8 FILLER_17_1236 ();
 sg13g2_decap_8 FILLER_17_1243 ();
 sg13g2_decap_8 FILLER_17_1250 ();
 sg13g2_decap_8 FILLER_17_1257 ();
 sg13g2_decap_8 FILLER_17_1264 ();
 sg13g2_decap_8 FILLER_17_1271 ();
 sg13g2_decap_8 FILLER_17_1278 ();
 sg13g2_decap_8 FILLER_17_1285 ();
 sg13g2_decap_8 FILLER_17_1292 ();
 sg13g2_decap_8 FILLER_17_1299 ();
 sg13g2_decap_8 FILLER_17_1306 ();
 sg13g2_decap_8 FILLER_17_1313 ();
 sg13g2_decap_4 FILLER_17_1320 ();
 sg13g2_fill_2 FILLER_17_1324 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_4 FILLER_18_140 ();
 sg13g2_fill_2 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_279 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_334 ();
 sg13g2_fill_1 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_441 ();
 sg13g2_fill_1 FILLER_18_533 ();
 sg13g2_fill_2 FILLER_18_554 ();
 sg13g2_fill_2 FILLER_18_591 ();
 sg13g2_fill_2 FILLER_18_773 ();
 sg13g2_fill_2 FILLER_18_809 ();
 sg13g2_fill_1 FILLER_18_937 ();
 sg13g2_decap_8 FILLER_18_1020 ();
 sg13g2_decap_8 FILLER_18_1027 ();
 sg13g2_decap_8 FILLER_18_1034 ();
 sg13g2_decap_8 FILLER_18_1041 ();
 sg13g2_decap_8 FILLER_18_1048 ();
 sg13g2_decap_8 FILLER_18_1055 ();
 sg13g2_decap_8 FILLER_18_1062 ();
 sg13g2_decap_8 FILLER_18_1069 ();
 sg13g2_decap_8 FILLER_18_1076 ();
 sg13g2_decap_8 FILLER_18_1083 ();
 sg13g2_decap_8 FILLER_18_1090 ();
 sg13g2_decap_8 FILLER_18_1097 ();
 sg13g2_decap_8 FILLER_18_1104 ();
 sg13g2_decap_8 FILLER_18_1111 ();
 sg13g2_decap_8 FILLER_18_1118 ();
 sg13g2_decap_8 FILLER_18_1125 ();
 sg13g2_decap_8 FILLER_18_1132 ();
 sg13g2_decap_8 FILLER_18_1139 ();
 sg13g2_decap_8 FILLER_18_1146 ();
 sg13g2_decap_8 FILLER_18_1153 ();
 sg13g2_decap_8 FILLER_18_1160 ();
 sg13g2_decap_8 FILLER_18_1167 ();
 sg13g2_decap_8 FILLER_18_1174 ();
 sg13g2_decap_8 FILLER_18_1181 ();
 sg13g2_decap_8 FILLER_18_1188 ();
 sg13g2_decap_8 FILLER_18_1195 ();
 sg13g2_decap_8 FILLER_18_1202 ();
 sg13g2_decap_8 FILLER_18_1209 ();
 sg13g2_decap_8 FILLER_18_1216 ();
 sg13g2_decap_8 FILLER_18_1223 ();
 sg13g2_decap_8 FILLER_18_1230 ();
 sg13g2_decap_8 FILLER_18_1237 ();
 sg13g2_decap_8 FILLER_18_1244 ();
 sg13g2_decap_8 FILLER_18_1251 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_8 FILLER_18_1265 ();
 sg13g2_decap_8 FILLER_18_1272 ();
 sg13g2_decap_8 FILLER_18_1279 ();
 sg13g2_decap_8 FILLER_18_1286 ();
 sg13g2_decap_8 FILLER_18_1293 ();
 sg13g2_decap_8 FILLER_18_1300 ();
 sg13g2_decap_8 FILLER_18_1307 ();
 sg13g2_decap_8 FILLER_18_1314 ();
 sg13g2_decap_4 FILLER_18_1321 ();
 sg13g2_fill_1 FILLER_18_1325 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_fill_2 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_2 FILLER_19_276 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_fill_1 FILLER_19_409 ();
 sg13g2_fill_2 FILLER_19_469 ();
 sg13g2_fill_1 FILLER_19_523 ();
 sg13g2_fill_1 FILLER_19_543 ();
 sg13g2_fill_2 FILLER_19_576 ();
 sg13g2_fill_1 FILLER_19_587 ();
 sg13g2_fill_1 FILLER_19_621 ();
 sg13g2_fill_2 FILLER_19_626 ();
 sg13g2_fill_1 FILLER_19_641 ();
 sg13g2_fill_1 FILLER_19_648 ();
 sg13g2_fill_2 FILLER_19_697 ();
 sg13g2_fill_1 FILLER_19_699 ();
 sg13g2_fill_1 FILLER_19_721 ();
 sg13g2_fill_2 FILLER_19_760 ();
 sg13g2_fill_1 FILLER_19_762 ();
 sg13g2_fill_2 FILLER_19_873 ();
 sg13g2_fill_2 FILLER_19_920 ();
 sg13g2_fill_1 FILLER_19_922 ();
 sg13g2_fill_2 FILLER_19_937 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_decap_8 FILLER_19_1029 ();
 sg13g2_decap_8 FILLER_19_1036 ();
 sg13g2_decap_8 FILLER_19_1043 ();
 sg13g2_decap_8 FILLER_19_1050 ();
 sg13g2_decap_8 FILLER_19_1057 ();
 sg13g2_decap_8 FILLER_19_1064 ();
 sg13g2_decap_8 FILLER_19_1071 ();
 sg13g2_decap_8 FILLER_19_1078 ();
 sg13g2_decap_8 FILLER_19_1085 ();
 sg13g2_decap_8 FILLER_19_1092 ();
 sg13g2_decap_8 FILLER_19_1099 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_decap_8 FILLER_19_1113 ();
 sg13g2_decap_8 FILLER_19_1120 ();
 sg13g2_decap_8 FILLER_19_1127 ();
 sg13g2_decap_8 FILLER_19_1134 ();
 sg13g2_decap_8 FILLER_19_1141 ();
 sg13g2_decap_8 FILLER_19_1148 ();
 sg13g2_decap_8 FILLER_19_1155 ();
 sg13g2_decap_8 FILLER_19_1162 ();
 sg13g2_decap_8 FILLER_19_1169 ();
 sg13g2_decap_8 FILLER_19_1176 ();
 sg13g2_decap_8 FILLER_19_1183 ();
 sg13g2_decap_8 FILLER_19_1190 ();
 sg13g2_decap_8 FILLER_19_1197 ();
 sg13g2_decap_8 FILLER_19_1204 ();
 sg13g2_decap_8 FILLER_19_1211 ();
 sg13g2_decap_8 FILLER_19_1218 ();
 sg13g2_decap_8 FILLER_19_1225 ();
 sg13g2_decap_8 FILLER_19_1232 ();
 sg13g2_decap_8 FILLER_19_1239 ();
 sg13g2_decap_8 FILLER_19_1246 ();
 sg13g2_decap_8 FILLER_19_1253 ();
 sg13g2_decap_8 FILLER_19_1260 ();
 sg13g2_decap_8 FILLER_19_1267 ();
 sg13g2_decap_8 FILLER_19_1274 ();
 sg13g2_decap_8 FILLER_19_1281 ();
 sg13g2_decap_8 FILLER_19_1288 ();
 sg13g2_decap_8 FILLER_19_1295 ();
 sg13g2_decap_8 FILLER_19_1302 ();
 sg13g2_decap_8 FILLER_19_1309 ();
 sg13g2_decap_8 FILLER_19_1316 ();
 sg13g2_fill_2 FILLER_19_1323 ();
 sg13g2_fill_1 FILLER_19_1325 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_94 ();
 sg13g2_fill_1 FILLER_20_96 ();
 sg13g2_fill_2 FILLER_20_113 ();
 sg13g2_fill_1 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_122 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_fill_2 FILLER_20_356 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_468 ();
 sg13g2_fill_2 FILLER_20_505 ();
 sg13g2_fill_1 FILLER_20_512 ();
 sg13g2_fill_2 FILLER_20_566 ();
 sg13g2_fill_2 FILLER_20_584 ();
 sg13g2_fill_1 FILLER_20_626 ();
 sg13g2_fill_1 FILLER_20_658 ();
 sg13g2_fill_2 FILLER_20_689 ();
 sg13g2_fill_1 FILLER_20_691 ();
 sg13g2_fill_1 FILLER_20_697 ();
 sg13g2_fill_1 FILLER_20_703 ();
 sg13g2_fill_2 FILLER_20_815 ();
 sg13g2_fill_1 FILLER_20_905 ();
 sg13g2_fill_1 FILLER_20_932 ();
 sg13g2_fill_1 FILLER_20_963 ();
 sg13g2_decap_8 FILLER_20_1022 ();
 sg13g2_decap_8 FILLER_20_1029 ();
 sg13g2_decap_8 FILLER_20_1036 ();
 sg13g2_decap_8 FILLER_20_1043 ();
 sg13g2_decap_8 FILLER_20_1050 ();
 sg13g2_decap_8 FILLER_20_1057 ();
 sg13g2_decap_8 FILLER_20_1064 ();
 sg13g2_decap_8 FILLER_20_1071 ();
 sg13g2_decap_8 FILLER_20_1078 ();
 sg13g2_decap_8 FILLER_20_1085 ();
 sg13g2_decap_8 FILLER_20_1092 ();
 sg13g2_decap_8 FILLER_20_1099 ();
 sg13g2_decap_8 FILLER_20_1106 ();
 sg13g2_decap_8 FILLER_20_1113 ();
 sg13g2_decap_8 FILLER_20_1120 ();
 sg13g2_decap_8 FILLER_20_1127 ();
 sg13g2_decap_8 FILLER_20_1134 ();
 sg13g2_decap_8 FILLER_20_1141 ();
 sg13g2_decap_8 FILLER_20_1148 ();
 sg13g2_decap_8 FILLER_20_1155 ();
 sg13g2_decap_8 FILLER_20_1162 ();
 sg13g2_decap_8 FILLER_20_1169 ();
 sg13g2_decap_8 FILLER_20_1176 ();
 sg13g2_decap_8 FILLER_20_1183 ();
 sg13g2_decap_8 FILLER_20_1190 ();
 sg13g2_decap_8 FILLER_20_1197 ();
 sg13g2_decap_8 FILLER_20_1204 ();
 sg13g2_decap_8 FILLER_20_1211 ();
 sg13g2_decap_8 FILLER_20_1218 ();
 sg13g2_decap_8 FILLER_20_1225 ();
 sg13g2_decap_8 FILLER_20_1232 ();
 sg13g2_decap_8 FILLER_20_1239 ();
 sg13g2_decap_8 FILLER_20_1246 ();
 sg13g2_decap_8 FILLER_20_1253 ();
 sg13g2_decap_8 FILLER_20_1260 ();
 sg13g2_decap_8 FILLER_20_1267 ();
 sg13g2_decap_8 FILLER_20_1274 ();
 sg13g2_decap_8 FILLER_20_1281 ();
 sg13g2_decap_8 FILLER_20_1288 ();
 sg13g2_decap_8 FILLER_20_1295 ();
 sg13g2_decap_8 FILLER_20_1302 ();
 sg13g2_decap_8 FILLER_20_1309 ();
 sg13g2_decap_8 FILLER_20_1316 ();
 sg13g2_fill_2 FILLER_20_1323 ();
 sg13g2_fill_1 FILLER_20_1325 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_4 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_65 ();
 sg13g2_fill_1 FILLER_21_84 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_120 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_fill_2 FILLER_21_161 ();
 sg13g2_fill_1 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_253 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_308 ();
 sg13g2_fill_2 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_542 ();
 sg13g2_fill_1 FILLER_21_635 ();
 sg13g2_fill_2 FILLER_21_651 ();
 sg13g2_fill_2 FILLER_21_670 ();
 sg13g2_fill_1 FILLER_21_685 ();
 sg13g2_fill_2 FILLER_21_697 ();
 sg13g2_fill_1 FILLER_21_699 ();
 sg13g2_fill_2 FILLER_21_714 ();
 sg13g2_fill_2 FILLER_21_724 ();
 sg13g2_fill_1 FILLER_21_734 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_fill_1 FILLER_21_749 ();
 sg13g2_fill_1 FILLER_21_755 ();
 sg13g2_fill_2 FILLER_21_842 ();
 sg13g2_fill_1 FILLER_21_844 ();
 sg13g2_fill_2 FILLER_21_909 ();
 sg13g2_fill_1 FILLER_21_941 ();
 sg13g2_fill_1 FILLER_21_1000 ();
 sg13g2_decap_8 FILLER_21_1037 ();
 sg13g2_decap_8 FILLER_21_1044 ();
 sg13g2_decap_8 FILLER_21_1051 ();
 sg13g2_decap_8 FILLER_21_1058 ();
 sg13g2_decap_8 FILLER_21_1065 ();
 sg13g2_decap_8 FILLER_21_1072 ();
 sg13g2_decap_8 FILLER_21_1079 ();
 sg13g2_decap_8 FILLER_21_1086 ();
 sg13g2_decap_8 FILLER_21_1093 ();
 sg13g2_decap_8 FILLER_21_1100 ();
 sg13g2_decap_8 FILLER_21_1107 ();
 sg13g2_decap_8 FILLER_21_1114 ();
 sg13g2_decap_8 FILLER_21_1121 ();
 sg13g2_decap_8 FILLER_21_1128 ();
 sg13g2_decap_8 FILLER_21_1135 ();
 sg13g2_decap_8 FILLER_21_1142 ();
 sg13g2_decap_8 FILLER_21_1149 ();
 sg13g2_decap_8 FILLER_21_1156 ();
 sg13g2_decap_8 FILLER_21_1163 ();
 sg13g2_decap_8 FILLER_21_1170 ();
 sg13g2_decap_8 FILLER_21_1177 ();
 sg13g2_decap_8 FILLER_21_1184 ();
 sg13g2_decap_8 FILLER_21_1191 ();
 sg13g2_decap_8 FILLER_21_1198 ();
 sg13g2_decap_8 FILLER_21_1205 ();
 sg13g2_decap_8 FILLER_21_1212 ();
 sg13g2_decap_8 FILLER_21_1219 ();
 sg13g2_decap_8 FILLER_21_1226 ();
 sg13g2_decap_8 FILLER_21_1233 ();
 sg13g2_decap_8 FILLER_21_1240 ();
 sg13g2_decap_8 FILLER_21_1247 ();
 sg13g2_decap_8 FILLER_21_1254 ();
 sg13g2_decap_8 FILLER_21_1261 ();
 sg13g2_decap_8 FILLER_21_1268 ();
 sg13g2_decap_8 FILLER_21_1275 ();
 sg13g2_decap_8 FILLER_21_1282 ();
 sg13g2_decap_8 FILLER_21_1289 ();
 sg13g2_decap_8 FILLER_21_1296 ();
 sg13g2_decap_8 FILLER_21_1303 ();
 sg13g2_decap_8 FILLER_21_1310 ();
 sg13g2_decap_8 FILLER_21_1317 ();
 sg13g2_fill_2 FILLER_21_1324 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_4 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_25 ();
 sg13g2_fill_2 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_103 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_238 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_336 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_22_456 ();
 sg13g2_fill_1 FILLER_22_467 ();
 sg13g2_fill_1 FILLER_22_478 ();
 sg13g2_fill_2 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_507 ();
 sg13g2_fill_2 FILLER_22_596 ();
 sg13g2_fill_2 FILLER_22_634 ();
 sg13g2_fill_1 FILLER_22_636 ();
 sg13g2_fill_1 FILLER_22_704 ();
 sg13g2_fill_2 FILLER_22_710 ();
 sg13g2_fill_2 FILLER_22_718 ();
 sg13g2_fill_2 FILLER_22_734 ();
 sg13g2_fill_1 FILLER_22_776 ();
 sg13g2_fill_2 FILLER_22_827 ();
 sg13g2_fill_2 FILLER_22_949 ();
 sg13g2_decap_4 FILLER_22_1013 ();
 sg13g2_decap_8 FILLER_22_1021 ();
 sg13g2_decap_8 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_22_1035 ();
 sg13g2_decap_8 FILLER_22_1042 ();
 sg13g2_decap_8 FILLER_22_1049 ();
 sg13g2_decap_8 FILLER_22_1056 ();
 sg13g2_decap_8 FILLER_22_1063 ();
 sg13g2_decap_8 FILLER_22_1070 ();
 sg13g2_decap_8 FILLER_22_1077 ();
 sg13g2_decap_8 FILLER_22_1084 ();
 sg13g2_decap_8 FILLER_22_1091 ();
 sg13g2_decap_8 FILLER_22_1098 ();
 sg13g2_decap_8 FILLER_22_1105 ();
 sg13g2_decap_8 FILLER_22_1112 ();
 sg13g2_decap_8 FILLER_22_1119 ();
 sg13g2_decap_8 FILLER_22_1126 ();
 sg13g2_decap_8 FILLER_22_1133 ();
 sg13g2_decap_8 FILLER_22_1140 ();
 sg13g2_decap_8 FILLER_22_1147 ();
 sg13g2_decap_8 FILLER_22_1154 ();
 sg13g2_decap_8 FILLER_22_1161 ();
 sg13g2_decap_8 FILLER_22_1168 ();
 sg13g2_decap_8 FILLER_22_1175 ();
 sg13g2_decap_8 FILLER_22_1182 ();
 sg13g2_decap_8 FILLER_22_1189 ();
 sg13g2_decap_8 FILLER_22_1196 ();
 sg13g2_decap_8 FILLER_22_1203 ();
 sg13g2_decap_8 FILLER_22_1210 ();
 sg13g2_decap_8 FILLER_22_1217 ();
 sg13g2_decap_8 FILLER_22_1224 ();
 sg13g2_decap_8 FILLER_22_1231 ();
 sg13g2_decap_8 FILLER_22_1238 ();
 sg13g2_decap_8 FILLER_22_1245 ();
 sg13g2_decap_8 FILLER_22_1252 ();
 sg13g2_decap_8 FILLER_22_1259 ();
 sg13g2_decap_8 FILLER_22_1266 ();
 sg13g2_decap_8 FILLER_22_1273 ();
 sg13g2_decap_8 FILLER_22_1280 ();
 sg13g2_decap_8 FILLER_22_1287 ();
 sg13g2_decap_8 FILLER_22_1294 ();
 sg13g2_decap_8 FILLER_22_1301 ();
 sg13g2_decap_8 FILLER_22_1308 ();
 sg13g2_decap_8 FILLER_22_1315 ();
 sg13g2_decap_4 FILLER_22_1322 ();
 sg13g2_fill_2 FILLER_23_8 ();
 sg13g2_fill_1 FILLER_23_10 ();
 sg13g2_fill_2 FILLER_23_19 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_2 FILLER_23_172 ();
 sg13g2_fill_1 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_200 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_fill_1 FILLER_23_245 ();
 sg13g2_fill_1 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_296 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_338 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_23_444 ();
 sg13g2_fill_1 FILLER_23_450 ();
 sg13g2_fill_2 FILLER_23_469 ();
 sg13g2_fill_2 FILLER_23_498 ();
 sg13g2_fill_2 FILLER_23_558 ();
 sg13g2_fill_1 FILLER_23_570 ();
 sg13g2_fill_1 FILLER_23_597 ();
 sg13g2_fill_1 FILLER_23_624 ();
 sg13g2_fill_1 FILLER_23_630 ();
 sg13g2_fill_2 FILLER_23_695 ();
 sg13g2_fill_1 FILLER_23_697 ();
 sg13g2_fill_1 FILLER_23_732 ();
 sg13g2_fill_1 FILLER_23_759 ();
 sg13g2_fill_1 FILLER_23_774 ();
 sg13g2_fill_2 FILLER_23_805 ();
 sg13g2_fill_1 FILLER_23_817 ();
 sg13g2_fill_1 FILLER_23_828 ();
 sg13g2_fill_1 FILLER_23_855 ();
 sg13g2_fill_2 FILLER_23_866 ();
 sg13g2_fill_2 FILLER_23_922 ();
 sg13g2_fill_1 FILLER_23_924 ();
 sg13g2_fill_1 FILLER_23_929 ();
 sg13g2_fill_2 FILLER_23_956 ();
 sg13g2_fill_1 FILLER_23_988 ();
 sg13g2_decap_8 FILLER_23_1027 ();
 sg13g2_decap_8 FILLER_23_1034 ();
 sg13g2_decap_8 FILLER_23_1041 ();
 sg13g2_decap_8 FILLER_23_1048 ();
 sg13g2_decap_8 FILLER_23_1055 ();
 sg13g2_decap_8 FILLER_23_1062 ();
 sg13g2_decap_8 FILLER_23_1069 ();
 sg13g2_decap_8 FILLER_23_1076 ();
 sg13g2_decap_8 FILLER_23_1083 ();
 sg13g2_decap_8 FILLER_23_1090 ();
 sg13g2_decap_8 FILLER_23_1097 ();
 sg13g2_decap_8 FILLER_23_1104 ();
 sg13g2_decap_8 FILLER_23_1111 ();
 sg13g2_decap_8 FILLER_23_1118 ();
 sg13g2_decap_8 FILLER_23_1125 ();
 sg13g2_decap_8 FILLER_23_1132 ();
 sg13g2_decap_8 FILLER_23_1139 ();
 sg13g2_decap_8 FILLER_23_1146 ();
 sg13g2_decap_8 FILLER_23_1153 ();
 sg13g2_decap_8 FILLER_23_1160 ();
 sg13g2_decap_8 FILLER_23_1167 ();
 sg13g2_decap_8 FILLER_23_1174 ();
 sg13g2_decap_8 FILLER_23_1181 ();
 sg13g2_decap_8 FILLER_23_1188 ();
 sg13g2_decap_8 FILLER_23_1195 ();
 sg13g2_decap_8 FILLER_23_1202 ();
 sg13g2_decap_8 FILLER_23_1209 ();
 sg13g2_decap_8 FILLER_23_1216 ();
 sg13g2_decap_8 FILLER_23_1223 ();
 sg13g2_decap_8 FILLER_23_1230 ();
 sg13g2_decap_8 FILLER_23_1237 ();
 sg13g2_decap_8 FILLER_23_1244 ();
 sg13g2_decap_8 FILLER_23_1251 ();
 sg13g2_decap_8 FILLER_23_1258 ();
 sg13g2_decap_8 FILLER_23_1265 ();
 sg13g2_decap_8 FILLER_23_1272 ();
 sg13g2_decap_8 FILLER_23_1279 ();
 sg13g2_decap_8 FILLER_23_1286 ();
 sg13g2_decap_8 FILLER_23_1293 ();
 sg13g2_decap_8 FILLER_23_1300 ();
 sg13g2_decap_8 FILLER_23_1307 ();
 sg13g2_decap_8 FILLER_23_1314 ();
 sg13g2_decap_4 FILLER_23_1321 ();
 sg13g2_fill_1 FILLER_23_1325 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_2 FILLER_24_51 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_62 ();
 sg13g2_fill_2 FILLER_24_77 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_140 ();
 sg13g2_fill_1 FILLER_24_146 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_214 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_320 ();
 sg13g2_fill_1 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_592 ();
 sg13g2_fill_1 FILLER_24_594 ();
 sg13g2_fill_1 FILLER_24_603 ();
 sg13g2_fill_1 FILLER_24_638 ();
 sg13g2_fill_1 FILLER_24_644 ();
 sg13g2_fill_1 FILLER_24_675 ();
 sg13g2_fill_1 FILLER_24_741 ();
 sg13g2_fill_1 FILLER_24_794 ();
 sg13g2_fill_2 FILLER_24_825 ();
 sg13g2_fill_2 FILLER_24_837 ();
 sg13g2_fill_2 FILLER_24_939 ();
 sg13g2_fill_2 FILLER_24_969 ();
 sg13g2_fill_1 FILLER_24_971 ();
 sg13g2_fill_1 FILLER_24_982 ();
 sg13g2_decap_8 FILLER_24_1027 ();
 sg13g2_decap_8 FILLER_24_1034 ();
 sg13g2_decap_8 FILLER_24_1041 ();
 sg13g2_decap_8 FILLER_24_1048 ();
 sg13g2_decap_8 FILLER_24_1055 ();
 sg13g2_decap_8 FILLER_24_1062 ();
 sg13g2_decap_8 FILLER_24_1069 ();
 sg13g2_decap_8 FILLER_24_1076 ();
 sg13g2_decap_8 FILLER_24_1083 ();
 sg13g2_decap_8 FILLER_24_1090 ();
 sg13g2_decap_8 FILLER_24_1097 ();
 sg13g2_decap_8 FILLER_24_1104 ();
 sg13g2_decap_8 FILLER_24_1111 ();
 sg13g2_decap_8 FILLER_24_1118 ();
 sg13g2_decap_8 FILLER_24_1125 ();
 sg13g2_decap_8 FILLER_24_1132 ();
 sg13g2_decap_8 FILLER_24_1139 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_8 FILLER_24_1153 ();
 sg13g2_decap_8 FILLER_24_1160 ();
 sg13g2_decap_8 FILLER_24_1167 ();
 sg13g2_decap_8 FILLER_24_1174 ();
 sg13g2_decap_8 FILLER_24_1181 ();
 sg13g2_decap_8 FILLER_24_1188 ();
 sg13g2_decap_8 FILLER_24_1195 ();
 sg13g2_decap_8 FILLER_24_1202 ();
 sg13g2_decap_8 FILLER_24_1209 ();
 sg13g2_decap_8 FILLER_24_1216 ();
 sg13g2_decap_8 FILLER_24_1223 ();
 sg13g2_decap_8 FILLER_24_1230 ();
 sg13g2_decap_8 FILLER_24_1237 ();
 sg13g2_decap_8 FILLER_24_1244 ();
 sg13g2_decap_8 FILLER_24_1251 ();
 sg13g2_decap_8 FILLER_24_1258 ();
 sg13g2_decap_8 FILLER_24_1265 ();
 sg13g2_decap_8 FILLER_24_1272 ();
 sg13g2_decap_8 FILLER_24_1279 ();
 sg13g2_decap_8 FILLER_24_1286 ();
 sg13g2_decap_8 FILLER_24_1293 ();
 sg13g2_decap_8 FILLER_24_1300 ();
 sg13g2_decap_8 FILLER_24_1307 ();
 sg13g2_decap_8 FILLER_24_1314 ();
 sg13g2_decap_4 FILLER_24_1321 ();
 sg13g2_fill_1 FILLER_24_1325 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_88 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_201 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_fill_1 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_352 ();
 sg13g2_fill_1 FILLER_25_358 ();
 sg13g2_fill_1 FILLER_25_373 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_fill_1 FILLER_25_449 ();
 sg13g2_fill_2 FILLER_25_468 ();
 sg13g2_fill_2 FILLER_25_515 ();
 sg13g2_fill_1 FILLER_25_576 ();
 sg13g2_fill_2 FILLER_25_584 ();
 sg13g2_decap_4 FILLER_25_661 ();
 sg13g2_fill_2 FILLER_25_665 ();
 sg13g2_fill_1 FILLER_25_684 ();
 sg13g2_fill_2 FILLER_25_709 ();
 sg13g2_fill_2 FILLER_25_757 ();
 sg13g2_fill_1 FILLER_25_773 ();
 sg13g2_fill_2 FILLER_25_800 ();
 sg13g2_fill_1 FILLER_25_810 ();
 sg13g2_fill_2 FILLER_25_837 ();
 sg13g2_fill_1 FILLER_25_905 ();
 sg13g2_fill_2 FILLER_25_916 ();
 sg13g2_fill_1 FILLER_25_980 ();
 sg13g2_fill_1 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_1030 ();
 sg13g2_decap_8 FILLER_25_1037 ();
 sg13g2_decap_8 FILLER_25_1044 ();
 sg13g2_decap_8 FILLER_25_1051 ();
 sg13g2_decap_8 FILLER_25_1058 ();
 sg13g2_decap_8 FILLER_25_1065 ();
 sg13g2_decap_8 FILLER_25_1072 ();
 sg13g2_decap_8 FILLER_25_1079 ();
 sg13g2_decap_8 FILLER_25_1086 ();
 sg13g2_decap_8 FILLER_25_1093 ();
 sg13g2_decap_8 FILLER_25_1100 ();
 sg13g2_decap_8 FILLER_25_1107 ();
 sg13g2_decap_8 FILLER_25_1114 ();
 sg13g2_decap_8 FILLER_25_1121 ();
 sg13g2_decap_8 FILLER_25_1128 ();
 sg13g2_decap_8 FILLER_25_1135 ();
 sg13g2_decap_8 FILLER_25_1142 ();
 sg13g2_decap_8 FILLER_25_1149 ();
 sg13g2_decap_8 FILLER_25_1156 ();
 sg13g2_decap_8 FILLER_25_1163 ();
 sg13g2_decap_8 FILLER_25_1170 ();
 sg13g2_decap_8 FILLER_25_1177 ();
 sg13g2_decap_8 FILLER_25_1184 ();
 sg13g2_decap_8 FILLER_25_1191 ();
 sg13g2_decap_8 FILLER_25_1198 ();
 sg13g2_decap_8 FILLER_25_1205 ();
 sg13g2_decap_8 FILLER_25_1212 ();
 sg13g2_decap_8 FILLER_25_1219 ();
 sg13g2_decap_8 FILLER_25_1226 ();
 sg13g2_decap_8 FILLER_25_1233 ();
 sg13g2_decap_8 FILLER_25_1240 ();
 sg13g2_decap_8 FILLER_25_1247 ();
 sg13g2_decap_8 FILLER_25_1254 ();
 sg13g2_decap_8 FILLER_25_1261 ();
 sg13g2_decap_8 FILLER_25_1268 ();
 sg13g2_decap_8 FILLER_25_1275 ();
 sg13g2_decap_8 FILLER_25_1282 ();
 sg13g2_decap_8 FILLER_25_1289 ();
 sg13g2_decap_8 FILLER_25_1296 ();
 sg13g2_decap_8 FILLER_25_1303 ();
 sg13g2_decap_8 FILLER_25_1310 ();
 sg13g2_decap_8 FILLER_25_1317 ();
 sg13g2_fill_2 FILLER_25_1324 ();
 sg13g2_fill_2 FILLER_26_34 ();
 sg13g2_fill_1 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_122 ();
 sg13g2_fill_1 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_161 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_2 FILLER_26_183 ();
 sg13g2_fill_1 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_412 ();
 sg13g2_fill_1 FILLER_26_498 ();
 sg13g2_fill_1 FILLER_26_532 ();
 sg13g2_fill_2 FILLER_26_542 ();
 sg13g2_fill_1 FILLER_26_544 ();
 sg13g2_fill_2 FILLER_26_580 ();
 sg13g2_fill_1 FILLER_26_582 ();
 sg13g2_fill_2 FILLER_26_588 ();
 sg13g2_fill_1 FILLER_26_618 ();
 sg13g2_fill_1 FILLER_26_626 ();
 sg13g2_fill_1 FILLER_26_632 ();
 sg13g2_fill_1 FILLER_26_638 ();
 sg13g2_fill_1 FILLER_26_644 ();
 sg13g2_fill_1 FILLER_26_650 ();
 sg13g2_fill_1 FILLER_26_729 ();
 sg13g2_fill_1 FILLER_26_756 ();
 sg13g2_fill_1 FILLER_26_761 ();
 sg13g2_fill_2 FILLER_26_792 ();
 sg13g2_fill_2 FILLER_26_838 ();
 sg13g2_fill_2 FILLER_26_870 ();
 sg13g2_fill_1 FILLER_26_884 ();
 sg13g2_fill_2 FILLER_26_963 ();
 sg13g2_decap_8 FILLER_26_1017 ();
 sg13g2_decap_8 FILLER_26_1024 ();
 sg13g2_decap_8 FILLER_26_1031 ();
 sg13g2_decap_8 FILLER_26_1038 ();
 sg13g2_decap_8 FILLER_26_1045 ();
 sg13g2_decap_8 FILLER_26_1052 ();
 sg13g2_decap_8 FILLER_26_1059 ();
 sg13g2_decap_8 FILLER_26_1066 ();
 sg13g2_decap_8 FILLER_26_1073 ();
 sg13g2_decap_8 FILLER_26_1080 ();
 sg13g2_decap_8 FILLER_26_1087 ();
 sg13g2_decap_8 FILLER_26_1094 ();
 sg13g2_decap_8 FILLER_26_1101 ();
 sg13g2_decap_8 FILLER_26_1108 ();
 sg13g2_decap_8 FILLER_26_1115 ();
 sg13g2_decap_8 FILLER_26_1122 ();
 sg13g2_decap_8 FILLER_26_1129 ();
 sg13g2_decap_8 FILLER_26_1136 ();
 sg13g2_decap_8 FILLER_26_1143 ();
 sg13g2_decap_8 FILLER_26_1150 ();
 sg13g2_decap_8 FILLER_26_1157 ();
 sg13g2_decap_8 FILLER_26_1164 ();
 sg13g2_decap_8 FILLER_26_1171 ();
 sg13g2_decap_8 FILLER_26_1178 ();
 sg13g2_decap_8 FILLER_26_1185 ();
 sg13g2_decap_8 FILLER_26_1192 ();
 sg13g2_decap_8 FILLER_26_1199 ();
 sg13g2_decap_8 FILLER_26_1206 ();
 sg13g2_decap_8 FILLER_26_1213 ();
 sg13g2_decap_8 FILLER_26_1220 ();
 sg13g2_decap_8 FILLER_26_1227 ();
 sg13g2_decap_8 FILLER_26_1234 ();
 sg13g2_decap_8 FILLER_26_1241 ();
 sg13g2_decap_8 FILLER_26_1248 ();
 sg13g2_decap_8 FILLER_26_1255 ();
 sg13g2_decap_8 FILLER_26_1262 ();
 sg13g2_decap_8 FILLER_26_1269 ();
 sg13g2_decap_8 FILLER_26_1276 ();
 sg13g2_decap_8 FILLER_26_1283 ();
 sg13g2_decap_8 FILLER_26_1290 ();
 sg13g2_decap_8 FILLER_26_1297 ();
 sg13g2_decap_8 FILLER_26_1304 ();
 sg13g2_decap_8 FILLER_26_1311 ();
 sg13g2_decap_8 FILLER_26_1318 ();
 sg13g2_fill_1 FILLER_26_1325 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_67 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_213 ();
 sg13g2_fill_2 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_268 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_312 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_fill_2 FILLER_27_389 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_fill_1 FILLER_27_462 ();
 sg13g2_fill_1 FILLER_27_473 ();
 sg13g2_fill_1 FILLER_27_478 ();
 sg13g2_fill_1 FILLER_27_535 ();
 sg13g2_fill_1 FILLER_27_546 ();
 sg13g2_fill_1 FILLER_27_552 ();
 sg13g2_fill_1 FILLER_27_560 ();
 sg13g2_fill_1 FILLER_27_571 ();
 sg13g2_fill_1 FILLER_27_593 ();
 sg13g2_fill_1 FILLER_27_618 ();
 sg13g2_fill_1 FILLER_27_634 ();
 sg13g2_fill_1 FILLER_27_640 ();
 sg13g2_fill_1 FILLER_27_647 ();
 sg13g2_fill_1 FILLER_27_658 ();
 sg13g2_decap_4 FILLER_27_669 ();
 sg13g2_fill_2 FILLER_27_673 ();
 sg13g2_fill_1 FILLER_27_680 ();
 sg13g2_fill_2 FILLER_27_685 ();
 sg13g2_fill_2 FILLER_27_692 ();
 sg13g2_decap_4 FILLER_27_701 ();
 sg13g2_fill_1 FILLER_27_709 ();
 sg13g2_fill_2 FILLER_27_740 ();
 sg13g2_fill_2 FILLER_27_772 ();
 sg13g2_fill_1 FILLER_27_774 ();
 sg13g2_fill_2 FILLER_27_809 ();
 sg13g2_fill_1 FILLER_27_873 ();
 sg13g2_fill_1 FILLER_27_892 ();
 sg13g2_fill_2 FILLER_27_985 ();
 sg13g2_decap_8 FILLER_27_1025 ();
 sg13g2_decap_8 FILLER_27_1032 ();
 sg13g2_decap_8 FILLER_27_1039 ();
 sg13g2_decap_8 FILLER_27_1046 ();
 sg13g2_decap_8 FILLER_27_1053 ();
 sg13g2_decap_8 FILLER_27_1060 ();
 sg13g2_decap_8 FILLER_27_1067 ();
 sg13g2_decap_8 FILLER_27_1074 ();
 sg13g2_decap_8 FILLER_27_1081 ();
 sg13g2_decap_8 FILLER_27_1088 ();
 sg13g2_decap_8 FILLER_27_1095 ();
 sg13g2_decap_8 FILLER_27_1102 ();
 sg13g2_decap_8 FILLER_27_1109 ();
 sg13g2_decap_8 FILLER_27_1116 ();
 sg13g2_decap_8 FILLER_27_1123 ();
 sg13g2_decap_8 FILLER_27_1130 ();
 sg13g2_decap_8 FILLER_27_1137 ();
 sg13g2_decap_8 FILLER_27_1144 ();
 sg13g2_decap_8 FILLER_27_1151 ();
 sg13g2_decap_8 FILLER_27_1158 ();
 sg13g2_decap_8 FILLER_27_1165 ();
 sg13g2_decap_8 FILLER_27_1172 ();
 sg13g2_decap_8 FILLER_27_1179 ();
 sg13g2_decap_8 FILLER_27_1186 ();
 sg13g2_decap_8 FILLER_27_1193 ();
 sg13g2_decap_8 FILLER_27_1200 ();
 sg13g2_decap_8 FILLER_27_1207 ();
 sg13g2_decap_8 FILLER_27_1214 ();
 sg13g2_decap_8 FILLER_27_1221 ();
 sg13g2_decap_8 FILLER_27_1228 ();
 sg13g2_decap_8 FILLER_27_1235 ();
 sg13g2_decap_8 FILLER_27_1242 ();
 sg13g2_decap_8 FILLER_27_1249 ();
 sg13g2_decap_8 FILLER_27_1256 ();
 sg13g2_decap_8 FILLER_27_1263 ();
 sg13g2_decap_8 FILLER_27_1270 ();
 sg13g2_decap_8 FILLER_27_1277 ();
 sg13g2_decap_8 FILLER_27_1284 ();
 sg13g2_decap_8 FILLER_27_1291 ();
 sg13g2_decap_8 FILLER_27_1298 ();
 sg13g2_decap_8 FILLER_27_1305 ();
 sg13g2_decap_8 FILLER_27_1312 ();
 sg13g2_decap_8 FILLER_27_1319 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_fill_2 FILLER_28_172 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_261 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_385 ();
 sg13g2_fill_1 FILLER_28_412 ();
 sg13g2_fill_2 FILLER_28_512 ();
 sg13g2_fill_1 FILLER_28_559 ();
 sg13g2_fill_1 FILLER_28_566 ();
 sg13g2_fill_1 FILLER_28_619 ();
 sg13g2_fill_2 FILLER_28_668 ();
 sg13g2_fill_2 FILLER_28_717 ();
 sg13g2_fill_1 FILLER_28_737 ();
 sg13g2_fill_2 FILLER_28_752 ();
 sg13g2_fill_1 FILLER_28_768 ();
 sg13g2_fill_1 FILLER_28_795 ();
 sg13g2_fill_1 FILLER_28_822 ();
 sg13g2_fill_1 FILLER_28_827 ();
 sg13g2_fill_1 FILLER_28_920 ();
 sg13g2_fill_2 FILLER_28_931 ();
 sg13g2_fill_1 FILLER_28_933 ();
 sg13g2_decap_8 FILLER_28_1020 ();
 sg13g2_decap_8 FILLER_28_1027 ();
 sg13g2_decap_8 FILLER_28_1034 ();
 sg13g2_decap_8 FILLER_28_1041 ();
 sg13g2_decap_8 FILLER_28_1048 ();
 sg13g2_decap_8 FILLER_28_1055 ();
 sg13g2_decap_8 FILLER_28_1062 ();
 sg13g2_decap_8 FILLER_28_1069 ();
 sg13g2_decap_8 FILLER_28_1076 ();
 sg13g2_decap_8 FILLER_28_1083 ();
 sg13g2_decap_8 FILLER_28_1090 ();
 sg13g2_decap_8 FILLER_28_1097 ();
 sg13g2_decap_8 FILLER_28_1104 ();
 sg13g2_decap_8 FILLER_28_1111 ();
 sg13g2_decap_8 FILLER_28_1118 ();
 sg13g2_decap_8 FILLER_28_1125 ();
 sg13g2_decap_8 FILLER_28_1132 ();
 sg13g2_decap_8 FILLER_28_1139 ();
 sg13g2_decap_8 FILLER_28_1146 ();
 sg13g2_decap_8 FILLER_28_1153 ();
 sg13g2_decap_8 FILLER_28_1160 ();
 sg13g2_decap_8 FILLER_28_1167 ();
 sg13g2_decap_8 FILLER_28_1174 ();
 sg13g2_decap_8 FILLER_28_1181 ();
 sg13g2_decap_8 FILLER_28_1188 ();
 sg13g2_decap_8 FILLER_28_1195 ();
 sg13g2_decap_8 FILLER_28_1202 ();
 sg13g2_decap_8 FILLER_28_1209 ();
 sg13g2_decap_8 FILLER_28_1216 ();
 sg13g2_decap_8 FILLER_28_1223 ();
 sg13g2_decap_8 FILLER_28_1230 ();
 sg13g2_decap_8 FILLER_28_1237 ();
 sg13g2_decap_8 FILLER_28_1244 ();
 sg13g2_decap_8 FILLER_28_1251 ();
 sg13g2_decap_8 FILLER_28_1258 ();
 sg13g2_decap_8 FILLER_28_1265 ();
 sg13g2_decap_8 FILLER_28_1272 ();
 sg13g2_decap_8 FILLER_28_1279 ();
 sg13g2_decap_8 FILLER_28_1286 ();
 sg13g2_decap_8 FILLER_28_1293 ();
 sg13g2_decap_8 FILLER_28_1300 ();
 sg13g2_decap_8 FILLER_28_1307 ();
 sg13g2_decap_8 FILLER_28_1314 ();
 sg13g2_decap_4 FILLER_28_1321 ();
 sg13g2_fill_1 FILLER_28_1325 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_106 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_fill_1 FILLER_29_187 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_238 ();
 sg13g2_fill_1 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_315 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_391 ();
 sg13g2_fill_2 FILLER_29_412 ();
 sg13g2_fill_1 FILLER_29_447 ();
 sg13g2_fill_1 FILLER_29_453 ();
 sg13g2_fill_1 FILLER_29_480 ();
 sg13g2_fill_1 FILLER_29_592 ();
 sg13g2_fill_1 FILLER_29_602 ();
 sg13g2_fill_1 FILLER_29_620 ();
 sg13g2_fill_1 FILLER_29_628 ();
 sg13g2_fill_1 FILLER_29_634 ();
 sg13g2_fill_2 FILLER_29_640 ();
 sg13g2_fill_2 FILLER_29_648 ();
 sg13g2_fill_1 FILLER_29_672 ();
 sg13g2_fill_2 FILLER_29_686 ();
 sg13g2_fill_2 FILLER_29_692 ();
 sg13g2_fill_1 FILLER_29_699 ();
 sg13g2_fill_1 FILLER_29_787 ();
 sg13g2_fill_2 FILLER_29_822 ();
 sg13g2_fill_2 FILLER_29_838 ();
 sg13g2_fill_1 FILLER_29_840 ();
 sg13g2_fill_2 FILLER_29_901 ();
 sg13g2_fill_1 FILLER_29_989 ();
 sg13g2_decap_8 FILLER_29_1020 ();
 sg13g2_decap_8 FILLER_29_1027 ();
 sg13g2_decap_8 FILLER_29_1034 ();
 sg13g2_decap_8 FILLER_29_1041 ();
 sg13g2_decap_8 FILLER_29_1048 ();
 sg13g2_decap_8 FILLER_29_1055 ();
 sg13g2_decap_8 FILLER_29_1062 ();
 sg13g2_decap_8 FILLER_29_1069 ();
 sg13g2_decap_8 FILLER_29_1076 ();
 sg13g2_decap_8 FILLER_29_1083 ();
 sg13g2_decap_8 FILLER_29_1090 ();
 sg13g2_decap_8 FILLER_29_1097 ();
 sg13g2_decap_8 FILLER_29_1104 ();
 sg13g2_decap_8 FILLER_29_1111 ();
 sg13g2_decap_8 FILLER_29_1118 ();
 sg13g2_decap_8 FILLER_29_1125 ();
 sg13g2_decap_8 FILLER_29_1132 ();
 sg13g2_decap_8 FILLER_29_1139 ();
 sg13g2_decap_8 FILLER_29_1146 ();
 sg13g2_decap_8 FILLER_29_1153 ();
 sg13g2_decap_8 FILLER_29_1160 ();
 sg13g2_decap_8 FILLER_29_1167 ();
 sg13g2_decap_8 FILLER_29_1174 ();
 sg13g2_decap_8 FILLER_29_1181 ();
 sg13g2_decap_8 FILLER_29_1188 ();
 sg13g2_decap_8 FILLER_29_1195 ();
 sg13g2_decap_8 FILLER_29_1202 ();
 sg13g2_decap_8 FILLER_29_1209 ();
 sg13g2_decap_8 FILLER_29_1216 ();
 sg13g2_decap_8 FILLER_29_1223 ();
 sg13g2_decap_8 FILLER_29_1230 ();
 sg13g2_decap_8 FILLER_29_1237 ();
 sg13g2_decap_8 FILLER_29_1244 ();
 sg13g2_decap_8 FILLER_29_1251 ();
 sg13g2_decap_8 FILLER_29_1258 ();
 sg13g2_decap_8 FILLER_29_1265 ();
 sg13g2_decap_8 FILLER_29_1272 ();
 sg13g2_decap_8 FILLER_29_1279 ();
 sg13g2_decap_8 FILLER_29_1286 ();
 sg13g2_decap_8 FILLER_29_1293 ();
 sg13g2_decap_8 FILLER_29_1300 ();
 sg13g2_decap_8 FILLER_29_1307 ();
 sg13g2_decap_8 FILLER_29_1314 ();
 sg13g2_decap_4 FILLER_29_1321 ();
 sg13g2_fill_1 FILLER_29_1325 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_5 ();
 sg13g2_fill_2 FILLER_30_16 ();
 sg13g2_fill_1 FILLER_30_33 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_fill_1 FILLER_30_152 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_fill_1 FILLER_30_308 ();
 sg13g2_fill_2 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_379 ();
 sg13g2_fill_2 FILLER_30_483 ();
 sg13g2_fill_2 FILLER_30_490 ();
 sg13g2_fill_2 FILLER_30_533 ();
 sg13g2_fill_2 FILLER_30_550 ();
 sg13g2_fill_2 FILLER_30_585 ();
 sg13g2_fill_1 FILLER_30_593 ();
 sg13g2_fill_2 FILLER_30_625 ();
 sg13g2_fill_1 FILLER_30_632 ();
 sg13g2_fill_1 FILLER_30_676 ();
 sg13g2_fill_1 FILLER_30_681 ();
 sg13g2_fill_2 FILLER_30_687 ();
 sg13g2_fill_1 FILLER_30_715 ();
 sg13g2_fill_2 FILLER_30_742 ();
 sg13g2_decap_4 FILLER_30_748 ();
 sg13g2_fill_1 FILLER_30_752 ();
 sg13g2_fill_2 FILLER_30_809 ();
 sg13g2_fill_2 FILLER_30_933 ();
 sg13g2_fill_2 FILLER_30_965 ();
 sg13g2_fill_1 FILLER_30_967 ();
 sg13g2_fill_2 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1026 ();
 sg13g2_decap_8 FILLER_30_1033 ();
 sg13g2_decap_8 FILLER_30_1040 ();
 sg13g2_decap_8 FILLER_30_1047 ();
 sg13g2_decap_8 FILLER_30_1054 ();
 sg13g2_decap_8 FILLER_30_1061 ();
 sg13g2_decap_8 FILLER_30_1068 ();
 sg13g2_decap_8 FILLER_30_1075 ();
 sg13g2_decap_8 FILLER_30_1082 ();
 sg13g2_decap_8 FILLER_30_1089 ();
 sg13g2_decap_8 FILLER_30_1096 ();
 sg13g2_decap_8 FILLER_30_1103 ();
 sg13g2_decap_8 FILLER_30_1110 ();
 sg13g2_decap_8 FILLER_30_1117 ();
 sg13g2_decap_8 FILLER_30_1124 ();
 sg13g2_decap_8 FILLER_30_1131 ();
 sg13g2_decap_8 FILLER_30_1138 ();
 sg13g2_decap_8 FILLER_30_1145 ();
 sg13g2_decap_8 FILLER_30_1152 ();
 sg13g2_decap_8 FILLER_30_1159 ();
 sg13g2_decap_8 FILLER_30_1166 ();
 sg13g2_decap_8 FILLER_30_1173 ();
 sg13g2_decap_8 FILLER_30_1180 ();
 sg13g2_decap_8 FILLER_30_1187 ();
 sg13g2_decap_8 FILLER_30_1194 ();
 sg13g2_decap_8 FILLER_30_1201 ();
 sg13g2_decap_8 FILLER_30_1208 ();
 sg13g2_decap_8 FILLER_30_1215 ();
 sg13g2_decap_8 FILLER_30_1222 ();
 sg13g2_decap_8 FILLER_30_1229 ();
 sg13g2_decap_8 FILLER_30_1236 ();
 sg13g2_decap_8 FILLER_30_1243 ();
 sg13g2_decap_8 FILLER_30_1250 ();
 sg13g2_decap_8 FILLER_30_1257 ();
 sg13g2_decap_8 FILLER_30_1264 ();
 sg13g2_decap_8 FILLER_30_1271 ();
 sg13g2_decap_8 FILLER_30_1278 ();
 sg13g2_decap_8 FILLER_30_1285 ();
 sg13g2_decap_8 FILLER_30_1292 ();
 sg13g2_decap_8 FILLER_30_1299 ();
 sg13g2_decap_8 FILLER_30_1306 ();
 sg13g2_decap_8 FILLER_30_1313 ();
 sg13g2_decap_4 FILLER_30_1320 ();
 sg13g2_fill_2 FILLER_30_1324 ();
 sg13g2_fill_2 FILLER_31_72 ();
 sg13g2_fill_1 FILLER_31_79 ();
 sg13g2_fill_2 FILLER_31_85 ();
 sg13g2_fill_1 FILLER_31_110 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_fill_1 FILLER_31_166 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_fill_2 FILLER_31_432 ();
 sg13g2_fill_2 FILLER_31_494 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_1 FILLER_31_551 ();
 sg13g2_fill_1 FILLER_31_570 ();
 sg13g2_fill_1 FILLER_31_576 ();
 sg13g2_fill_1 FILLER_31_583 ();
 sg13g2_fill_1 FILLER_31_618 ();
 sg13g2_fill_2 FILLER_31_629 ();
 sg13g2_fill_1 FILLER_31_653 ();
 sg13g2_fill_1 FILLER_31_660 ();
 sg13g2_fill_1 FILLER_31_670 ();
 sg13g2_fill_1 FILLER_31_690 ();
 sg13g2_fill_1 FILLER_31_695 ();
 sg13g2_fill_1 FILLER_31_786 ();
 sg13g2_fill_1 FILLER_31_813 ();
 sg13g2_fill_1 FILLER_31_840 ();
 sg13g2_fill_2 FILLER_31_859 ();
 sg13g2_fill_1 FILLER_31_869 ();
 sg13g2_fill_1 FILLER_31_883 ();
 sg13g2_fill_2 FILLER_31_950 ();
 sg13g2_decap_8 FILLER_31_1034 ();
 sg13g2_decap_8 FILLER_31_1041 ();
 sg13g2_decap_8 FILLER_31_1048 ();
 sg13g2_decap_8 FILLER_31_1055 ();
 sg13g2_decap_8 FILLER_31_1062 ();
 sg13g2_decap_8 FILLER_31_1069 ();
 sg13g2_decap_8 FILLER_31_1076 ();
 sg13g2_decap_8 FILLER_31_1083 ();
 sg13g2_decap_8 FILLER_31_1090 ();
 sg13g2_decap_8 FILLER_31_1097 ();
 sg13g2_decap_8 FILLER_31_1104 ();
 sg13g2_decap_8 FILLER_31_1111 ();
 sg13g2_decap_8 FILLER_31_1118 ();
 sg13g2_decap_8 FILLER_31_1125 ();
 sg13g2_decap_8 FILLER_31_1132 ();
 sg13g2_decap_8 FILLER_31_1139 ();
 sg13g2_decap_8 FILLER_31_1146 ();
 sg13g2_decap_8 FILLER_31_1153 ();
 sg13g2_decap_8 FILLER_31_1160 ();
 sg13g2_decap_8 FILLER_31_1167 ();
 sg13g2_decap_8 FILLER_31_1174 ();
 sg13g2_decap_8 FILLER_31_1181 ();
 sg13g2_decap_8 FILLER_31_1188 ();
 sg13g2_decap_8 FILLER_31_1195 ();
 sg13g2_decap_8 FILLER_31_1202 ();
 sg13g2_decap_8 FILLER_31_1209 ();
 sg13g2_decap_8 FILLER_31_1216 ();
 sg13g2_decap_8 FILLER_31_1223 ();
 sg13g2_decap_8 FILLER_31_1230 ();
 sg13g2_decap_8 FILLER_31_1237 ();
 sg13g2_decap_8 FILLER_31_1244 ();
 sg13g2_decap_8 FILLER_31_1251 ();
 sg13g2_decap_8 FILLER_31_1258 ();
 sg13g2_decap_8 FILLER_31_1265 ();
 sg13g2_decap_8 FILLER_31_1272 ();
 sg13g2_decap_8 FILLER_31_1279 ();
 sg13g2_decap_8 FILLER_31_1286 ();
 sg13g2_decap_8 FILLER_31_1293 ();
 sg13g2_decap_8 FILLER_31_1300 ();
 sg13g2_decap_8 FILLER_31_1307 ();
 sg13g2_decap_8 FILLER_31_1314 ();
 sg13g2_decap_4 FILLER_31_1321 ();
 sg13g2_fill_1 FILLER_31_1325 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_367 ();
 sg13g2_fill_1 FILLER_32_488 ();
 sg13g2_fill_1 FILLER_32_523 ();
 sg13g2_fill_2 FILLER_32_553 ();
 sg13g2_fill_1 FILLER_32_613 ();
 sg13g2_fill_2 FILLER_32_631 ();
 sg13g2_fill_2 FILLER_32_674 ();
 sg13g2_fill_1 FILLER_32_681 ();
 sg13g2_fill_2 FILLER_32_687 ();
 sg13g2_fill_2 FILLER_32_694 ();
 sg13g2_fill_1 FILLER_32_696 ();
 sg13g2_fill_1 FILLER_32_701 ();
 sg13g2_fill_2 FILLER_32_814 ();
 sg13g2_fill_1 FILLER_32_842 ();
 sg13g2_fill_2 FILLER_32_935 ();
 sg13g2_fill_1 FILLER_32_937 ();
 sg13g2_fill_2 FILLER_32_968 ();
 sg13g2_fill_2 FILLER_32_980 ();
 sg13g2_decap_8 FILLER_32_1022 ();
 sg13g2_decap_8 FILLER_32_1029 ();
 sg13g2_decap_8 FILLER_32_1036 ();
 sg13g2_decap_8 FILLER_32_1043 ();
 sg13g2_decap_8 FILLER_32_1050 ();
 sg13g2_decap_8 FILLER_32_1057 ();
 sg13g2_decap_8 FILLER_32_1064 ();
 sg13g2_decap_8 FILLER_32_1071 ();
 sg13g2_decap_8 FILLER_32_1078 ();
 sg13g2_decap_8 FILLER_32_1085 ();
 sg13g2_decap_8 FILLER_32_1092 ();
 sg13g2_decap_8 FILLER_32_1099 ();
 sg13g2_decap_8 FILLER_32_1106 ();
 sg13g2_decap_8 FILLER_32_1113 ();
 sg13g2_decap_8 FILLER_32_1120 ();
 sg13g2_decap_8 FILLER_32_1127 ();
 sg13g2_decap_8 FILLER_32_1134 ();
 sg13g2_decap_8 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1148 ();
 sg13g2_decap_8 FILLER_32_1155 ();
 sg13g2_decap_8 FILLER_32_1162 ();
 sg13g2_decap_8 FILLER_32_1169 ();
 sg13g2_decap_8 FILLER_32_1176 ();
 sg13g2_decap_8 FILLER_32_1183 ();
 sg13g2_decap_8 FILLER_32_1190 ();
 sg13g2_decap_8 FILLER_32_1197 ();
 sg13g2_decap_8 FILLER_32_1204 ();
 sg13g2_decap_8 FILLER_32_1211 ();
 sg13g2_decap_8 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1225 ();
 sg13g2_decap_8 FILLER_32_1232 ();
 sg13g2_decap_8 FILLER_32_1239 ();
 sg13g2_decap_8 FILLER_32_1246 ();
 sg13g2_decap_8 FILLER_32_1253 ();
 sg13g2_decap_8 FILLER_32_1260 ();
 sg13g2_decap_8 FILLER_32_1267 ();
 sg13g2_decap_8 FILLER_32_1274 ();
 sg13g2_decap_8 FILLER_32_1281 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1302 ();
 sg13g2_decap_8 FILLER_32_1309 ();
 sg13g2_decap_8 FILLER_32_1316 ();
 sg13g2_fill_2 FILLER_32_1323 ();
 sg13g2_fill_1 FILLER_32_1325 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_90 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_309 ();
 sg13g2_decap_4 FILLER_33_348 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_365 ();
 sg13g2_fill_2 FILLER_33_421 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_2 FILLER_33_439 ();
 sg13g2_fill_2 FILLER_33_451 ();
 sg13g2_fill_1 FILLER_33_453 ();
 sg13g2_fill_1 FILLER_33_467 ();
 sg13g2_fill_2 FILLER_33_503 ();
 sg13g2_fill_1 FILLER_33_513 ();
 sg13g2_fill_1 FILLER_33_519 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_2 FILLER_33_559 ();
 sg13g2_fill_2 FILLER_33_607 ();
 sg13g2_fill_1 FILLER_33_619 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_fill_1 FILLER_33_632 ();
 sg13g2_fill_2 FILLER_33_639 ();
 sg13g2_fill_1 FILLER_33_641 ();
 sg13g2_fill_2 FILLER_33_680 ();
 sg13g2_fill_2 FILLER_33_745 ();
 sg13g2_fill_1 FILLER_33_747 ();
 sg13g2_fill_1 FILLER_33_774 ();
 sg13g2_fill_1 FILLER_33_805 ();
 sg13g2_fill_1 FILLER_33_832 ();
 sg13g2_fill_1 FILLER_33_843 ();
 sg13g2_fill_2 FILLER_33_914 ();
 sg13g2_fill_1 FILLER_33_983 ();
 sg13g2_decap_8 FILLER_33_1024 ();
 sg13g2_decap_8 FILLER_33_1031 ();
 sg13g2_decap_8 FILLER_33_1038 ();
 sg13g2_decap_8 FILLER_33_1045 ();
 sg13g2_decap_8 FILLER_33_1052 ();
 sg13g2_decap_8 FILLER_33_1059 ();
 sg13g2_decap_8 FILLER_33_1066 ();
 sg13g2_decap_8 FILLER_33_1073 ();
 sg13g2_decap_8 FILLER_33_1080 ();
 sg13g2_decap_8 FILLER_33_1087 ();
 sg13g2_decap_8 FILLER_33_1094 ();
 sg13g2_decap_8 FILLER_33_1101 ();
 sg13g2_decap_8 FILLER_33_1108 ();
 sg13g2_decap_8 FILLER_33_1115 ();
 sg13g2_decap_8 FILLER_33_1122 ();
 sg13g2_decap_8 FILLER_33_1129 ();
 sg13g2_decap_8 FILLER_33_1136 ();
 sg13g2_decap_8 FILLER_33_1143 ();
 sg13g2_decap_8 FILLER_33_1150 ();
 sg13g2_decap_8 FILLER_33_1157 ();
 sg13g2_decap_8 FILLER_33_1164 ();
 sg13g2_decap_8 FILLER_33_1171 ();
 sg13g2_decap_8 FILLER_33_1178 ();
 sg13g2_decap_8 FILLER_33_1185 ();
 sg13g2_decap_8 FILLER_33_1192 ();
 sg13g2_decap_8 FILLER_33_1199 ();
 sg13g2_decap_8 FILLER_33_1206 ();
 sg13g2_decap_8 FILLER_33_1213 ();
 sg13g2_decap_8 FILLER_33_1220 ();
 sg13g2_decap_8 FILLER_33_1227 ();
 sg13g2_decap_8 FILLER_33_1234 ();
 sg13g2_decap_8 FILLER_33_1241 ();
 sg13g2_decap_8 FILLER_33_1248 ();
 sg13g2_decap_8 FILLER_33_1255 ();
 sg13g2_decap_8 FILLER_33_1262 ();
 sg13g2_decap_8 FILLER_33_1269 ();
 sg13g2_decap_8 FILLER_33_1276 ();
 sg13g2_decap_8 FILLER_33_1283 ();
 sg13g2_decap_8 FILLER_33_1290 ();
 sg13g2_decap_8 FILLER_33_1297 ();
 sg13g2_decap_8 FILLER_33_1304 ();
 sg13g2_decap_8 FILLER_33_1311 ();
 sg13g2_decap_8 FILLER_33_1318 ();
 sg13g2_fill_1 FILLER_33_1325 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_36 ();
 sg13g2_fill_2 FILLER_34_89 ();
 sg13g2_fill_1 FILLER_34_96 ();
 sg13g2_fill_1 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_151 ();
 sg13g2_fill_2 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_180 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_fill_2 FILLER_34_192 ();
 sg13g2_fill_1 FILLER_34_223 ();
 sg13g2_fill_1 FILLER_34_234 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_2 FILLER_34_439 ();
 sg13g2_fill_2 FILLER_34_477 ();
 sg13g2_fill_1 FILLER_34_479 ();
 sg13g2_fill_1 FILLER_34_522 ();
 sg13g2_fill_1 FILLER_34_572 ();
 sg13g2_fill_2 FILLER_34_578 ();
 sg13g2_fill_2 FILLER_34_590 ();
 sg13g2_fill_1 FILLER_34_604 ();
 sg13g2_fill_2 FILLER_34_645 ();
 sg13g2_fill_2 FILLER_34_667 ();
 sg13g2_fill_2 FILLER_34_679 ();
 sg13g2_fill_1 FILLER_34_681 ();
 sg13g2_decap_4 FILLER_34_686 ();
 sg13g2_fill_1 FILLER_34_690 ();
 sg13g2_fill_2 FILLER_34_703 ();
 sg13g2_decap_4 FILLER_34_710 ();
 sg13g2_fill_1 FILLER_34_714 ();
 sg13g2_fill_2 FILLER_34_786 ();
 sg13g2_fill_2 FILLER_34_822 ();
 sg13g2_fill_1 FILLER_34_886 ();
 sg13g2_fill_1 FILLER_34_913 ();
 sg13g2_fill_1 FILLER_34_924 ();
 sg13g2_fill_1 FILLER_34_935 ();
 sg13g2_fill_2 FILLER_34_966 ();
 sg13g2_fill_1 FILLER_34_968 ();
 sg13g2_fill_2 FILLER_34_979 ();
 sg13g2_decap_8 FILLER_34_1021 ();
 sg13g2_decap_8 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_34_1035 ();
 sg13g2_decap_8 FILLER_34_1042 ();
 sg13g2_decap_8 FILLER_34_1049 ();
 sg13g2_decap_8 FILLER_34_1056 ();
 sg13g2_decap_8 FILLER_34_1063 ();
 sg13g2_decap_8 FILLER_34_1070 ();
 sg13g2_decap_8 FILLER_34_1077 ();
 sg13g2_decap_8 FILLER_34_1084 ();
 sg13g2_decap_8 FILLER_34_1091 ();
 sg13g2_decap_8 FILLER_34_1098 ();
 sg13g2_decap_8 FILLER_34_1105 ();
 sg13g2_decap_8 FILLER_34_1112 ();
 sg13g2_decap_8 FILLER_34_1119 ();
 sg13g2_decap_8 FILLER_34_1126 ();
 sg13g2_decap_8 FILLER_34_1133 ();
 sg13g2_decap_8 FILLER_34_1140 ();
 sg13g2_decap_8 FILLER_34_1147 ();
 sg13g2_decap_8 FILLER_34_1154 ();
 sg13g2_decap_8 FILLER_34_1161 ();
 sg13g2_decap_8 FILLER_34_1168 ();
 sg13g2_decap_8 FILLER_34_1175 ();
 sg13g2_decap_8 FILLER_34_1182 ();
 sg13g2_decap_8 FILLER_34_1189 ();
 sg13g2_decap_8 FILLER_34_1196 ();
 sg13g2_decap_8 FILLER_34_1203 ();
 sg13g2_decap_8 FILLER_34_1210 ();
 sg13g2_decap_8 FILLER_34_1217 ();
 sg13g2_decap_8 FILLER_34_1224 ();
 sg13g2_decap_8 FILLER_34_1231 ();
 sg13g2_decap_8 FILLER_34_1238 ();
 sg13g2_decap_8 FILLER_34_1245 ();
 sg13g2_decap_8 FILLER_34_1252 ();
 sg13g2_decap_8 FILLER_34_1259 ();
 sg13g2_decap_8 FILLER_34_1266 ();
 sg13g2_decap_8 FILLER_34_1273 ();
 sg13g2_decap_8 FILLER_34_1280 ();
 sg13g2_decap_8 FILLER_34_1287 ();
 sg13g2_decap_8 FILLER_34_1294 ();
 sg13g2_decap_8 FILLER_34_1301 ();
 sg13g2_decap_8 FILLER_34_1308 ();
 sg13g2_decap_8 FILLER_34_1315 ();
 sg13g2_decap_4 FILLER_34_1322 ();
 sg13g2_fill_2 FILLER_35_31 ();
 sg13g2_fill_1 FILLER_35_33 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_fill_2 FILLER_35_94 ();
 sg13g2_fill_2 FILLER_35_122 ();
 sg13g2_fill_1 FILLER_35_124 ();
 sg13g2_fill_1 FILLER_35_142 ();
 sg13g2_fill_2 FILLER_35_178 ();
 sg13g2_fill_2 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_300 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_fill_1 FILLER_35_484 ();
 sg13g2_fill_2 FILLER_35_521 ();
 sg13g2_fill_2 FILLER_35_528 ();
 sg13g2_fill_2 FILLER_35_547 ();
 sg13g2_fill_1 FILLER_35_559 ();
 sg13g2_fill_1 FILLER_35_581 ();
 sg13g2_fill_1 FILLER_35_618 ();
 sg13g2_fill_1 FILLER_35_634 ();
 sg13g2_fill_2 FILLER_35_646 ();
 sg13g2_fill_1 FILLER_35_653 ();
 sg13g2_fill_1 FILLER_35_661 ();
 sg13g2_fill_1 FILLER_35_667 ();
 sg13g2_fill_1 FILLER_35_672 ();
 sg13g2_fill_1 FILLER_35_694 ();
 sg13g2_fill_1 FILLER_35_699 ();
 sg13g2_fill_2 FILLER_35_715 ();
 sg13g2_fill_1 FILLER_35_717 ();
 sg13g2_decap_4 FILLER_35_724 ();
 sg13g2_fill_2 FILLER_35_883 ();
 sg13g2_fill_2 FILLER_35_895 ();
 sg13g2_fill_1 FILLER_35_897 ();
 sg13g2_fill_2 FILLER_35_950 ();
 sg13g2_fill_1 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_1017 ();
 sg13g2_decap_8 FILLER_35_1024 ();
 sg13g2_decap_8 FILLER_35_1031 ();
 sg13g2_decap_8 FILLER_35_1038 ();
 sg13g2_decap_8 FILLER_35_1045 ();
 sg13g2_decap_8 FILLER_35_1052 ();
 sg13g2_decap_8 FILLER_35_1059 ();
 sg13g2_decap_8 FILLER_35_1066 ();
 sg13g2_decap_8 FILLER_35_1073 ();
 sg13g2_decap_8 FILLER_35_1080 ();
 sg13g2_decap_8 FILLER_35_1087 ();
 sg13g2_decap_8 FILLER_35_1094 ();
 sg13g2_decap_8 FILLER_35_1101 ();
 sg13g2_decap_8 FILLER_35_1108 ();
 sg13g2_decap_8 FILLER_35_1115 ();
 sg13g2_decap_8 FILLER_35_1122 ();
 sg13g2_decap_8 FILLER_35_1129 ();
 sg13g2_decap_8 FILLER_35_1136 ();
 sg13g2_decap_8 FILLER_35_1143 ();
 sg13g2_decap_8 FILLER_35_1150 ();
 sg13g2_decap_8 FILLER_35_1157 ();
 sg13g2_decap_8 FILLER_35_1164 ();
 sg13g2_decap_8 FILLER_35_1171 ();
 sg13g2_decap_8 FILLER_35_1178 ();
 sg13g2_decap_8 FILLER_35_1185 ();
 sg13g2_decap_8 FILLER_35_1192 ();
 sg13g2_decap_8 FILLER_35_1199 ();
 sg13g2_decap_8 FILLER_35_1206 ();
 sg13g2_decap_8 FILLER_35_1213 ();
 sg13g2_decap_8 FILLER_35_1220 ();
 sg13g2_decap_8 FILLER_35_1227 ();
 sg13g2_decap_8 FILLER_35_1234 ();
 sg13g2_decap_8 FILLER_35_1241 ();
 sg13g2_decap_8 FILLER_35_1248 ();
 sg13g2_decap_8 FILLER_35_1255 ();
 sg13g2_decap_8 FILLER_35_1262 ();
 sg13g2_decap_8 FILLER_35_1269 ();
 sg13g2_decap_8 FILLER_35_1276 ();
 sg13g2_decap_8 FILLER_35_1283 ();
 sg13g2_decap_8 FILLER_35_1290 ();
 sg13g2_decap_8 FILLER_35_1297 ();
 sg13g2_decap_8 FILLER_35_1304 ();
 sg13g2_decap_8 FILLER_35_1311 ();
 sg13g2_decap_8 FILLER_35_1318 ();
 sg13g2_fill_1 FILLER_35_1325 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_80 ();
 sg13g2_fill_1 FILLER_36_87 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_111 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_157 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_207 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_fill_1 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_313 ();
 sg13g2_fill_1 FILLER_36_328 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_387 ();
 sg13g2_fill_2 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_427 ();
 sg13g2_fill_2 FILLER_36_464 ();
 sg13g2_fill_1 FILLER_36_466 ();
 sg13g2_fill_2 FILLER_36_506 ();
 sg13g2_fill_1 FILLER_36_508 ();
 sg13g2_fill_2 FILLER_36_575 ();
 sg13g2_fill_1 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_594 ();
 sg13g2_fill_2 FILLER_36_604 ();
 sg13g2_fill_1 FILLER_36_636 ();
 sg13g2_fill_1 FILLER_36_686 ();
 sg13g2_fill_2 FILLER_36_748 ();
 sg13g2_fill_2 FILLER_36_836 ();
 sg13g2_fill_1 FILLER_36_838 ();
 sg13g2_fill_1 FILLER_36_899 ();
 sg13g2_fill_1 FILLER_36_910 ();
 sg13g2_fill_2 FILLER_36_965 ();
 sg13g2_fill_1 FILLER_36_967 ();
 sg13g2_decap_8 FILLER_36_1012 ();
 sg13g2_decap_8 FILLER_36_1019 ();
 sg13g2_decap_8 FILLER_36_1026 ();
 sg13g2_decap_8 FILLER_36_1033 ();
 sg13g2_decap_8 FILLER_36_1040 ();
 sg13g2_decap_8 FILLER_36_1047 ();
 sg13g2_decap_8 FILLER_36_1054 ();
 sg13g2_decap_8 FILLER_36_1061 ();
 sg13g2_decap_8 FILLER_36_1068 ();
 sg13g2_decap_8 FILLER_36_1075 ();
 sg13g2_decap_8 FILLER_36_1082 ();
 sg13g2_decap_8 FILLER_36_1089 ();
 sg13g2_decap_8 FILLER_36_1096 ();
 sg13g2_decap_8 FILLER_36_1103 ();
 sg13g2_decap_8 FILLER_36_1110 ();
 sg13g2_decap_8 FILLER_36_1117 ();
 sg13g2_decap_8 FILLER_36_1124 ();
 sg13g2_decap_8 FILLER_36_1131 ();
 sg13g2_decap_8 FILLER_36_1138 ();
 sg13g2_decap_8 FILLER_36_1145 ();
 sg13g2_decap_8 FILLER_36_1152 ();
 sg13g2_decap_8 FILLER_36_1159 ();
 sg13g2_decap_8 FILLER_36_1166 ();
 sg13g2_decap_8 FILLER_36_1173 ();
 sg13g2_decap_8 FILLER_36_1180 ();
 sg13g2_decap_8 FILLER_36_1187 ();
 sg13g2_decap_8 FILLER_36_1194 ();
 sg13g2_decap_8 FILLER_36_1201 ();
 sg13g2_decap_8 FILLER_36_1208 ();
 sg13g2_decap_8 FILLER_36_1215 ();
 sg13g2_decap_8 FILLER_36_1222 ();
 sg13g2_decap_8 FILLER_36_1229 ();
 sg13g2_decap_8 FILLER_36_1236 ();
 sg13g2_decap_8 FILLER_36_1243 ();
 sg13g2_decap_8 FILLER_36_1250 ();
 sg13g2_decap_8 FILLER_36_1257 ();
 sg13g2_decap_8 FILLER_36_1264 ();
 sg13g2_decap_8 FILLER_36_1271 ();
 sg13g2_decap_8 FILLER_36_1278 ();
 sg13g2_decap_8 FILLER_36_1285 ();
 sg13g2_decap_8 FILLER_36_1292 ();
 sg13g2_decap_8 FILLER_36_1299 ();
 sg13g2_decap_8 FILLER_36_1306 ();
 sg13g2_decap_8 FILLER_36_1313 ();
 sg13g2_decap_4 FILLER_36_1320 ();
 sg13g2_fill_2 FILLER_36_1324 ();
 sg13g2_fill_1 FILLER_37_26 ();
 sg13g2_fill_1 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_136 ();
 sg13g2_fill_1 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_175 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_2 FILLER_37_246 ();
 sg13g2_fill_1 FILLER_37_256 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_decap_4 FILLER_37_317 ();
 sg13g2_fill_2 FILLER_37_388 ();
 sg13g2_fill_2 FILLER_37_400 ();
 sg13g2_fill_1 FILLER_37_402 ();
 sg13g2_fill_2 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_430 ();
 sg13g2_decap_4 FILLER_37_437 ();
 sg13g2_fill_2 FILLER_37_481 ();
 sg13g2_fill_1 FILLER_37_542 ();
 sg13g2_fill_2 FILLER_37_582 ();
 sg13g2_fill_2 FILLER_37_620 ();
 sg13g2_fill_2 FILLER_37_651 ();
 sg13g2_fill_2 FILLER_37_659 ();
 sg13g2_fill_1 FILLER_37_667 ();
 sg13g2_fill_1 FILLER_37_673 ();
 sg13g2_fill_1 FILLER_37_682 ();
 sg13g2_fill_1 FILLER_37_689 ();
 sg13g2_fill_1 FILLER_37_695 ();
 sg13g2_fill_1 FILLER_37_700 ();
 sg13g2_fill_1 FILLER_37_704 ();
 sg13g2_fill_1 FILLER_37_715 ();
 sg13g2_fill_1 FILLER_37_720 ();
 sg13g2_fill_1 FILLER_37_725 ();
 sg13g2_fill_1 FILLER_37_744 ();
 sg13g2_fill_2 FILLER_37_755 ();
 sg13g2_fill_1 FILLER_37_757 ();
 sg13g2_fill_2 FILLER_37_762 ();
 sg13g2_decap_4 FILLER_37_774 ();
 sg13g2_fill_1 FILLER_37_792 ();
 sg13g2_fill_1 FILLER_37_803 ();
 sg13g2_fill_1 FILLER_37_814 ();
 sg13g2_fill_1 FILLER_37_819 ();
 sg13g2_fill_1 FILLER_37_830 ();
 sg13g2_fill_1 FILLER_37_841 ();
 sg13g2_fill_2 FILLER_37_868 ();
 sg13g2_fill_1 FILLER_37_870 ();
 sg13g2_fill_2 FILLER_37_961 ();
 sg13g2_fill_1 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_1000 ();
 sg13g2_decap_8 FILLER_37_1007 ();
 sg13g2_decap_8 FILLER_37_1014 ();
 sg13g2_decap_8 FILLER_37_1021 ();
 sg13g2_decap_8 FILLER_37_1028 ();
 sg13g2_decap_8 FILLER_37_1035 ();
 sg13g2_decap_8 FILLER_37_1042 ();
 sg13g2_decap_8 FILLER_37_1049 ();
 sg13g2_decap_8 FILLER_37_1056 ();
 sg13g2_decap_8 FILLER_37_1063 ();
 sg13g2_decap_8 FILLER_37_1070 ();
 sg13g2_decap_8 FILLER_37_1077 ();
 sg13g2_decap_8 FILLER_37_1084 ();
 sg13g2_decap_8 FILLER_37_1091 ();
 sg13g2_decap_8 FILLER_37_1098 ();
 sg13g2_decap_8 FILLER_37_1105 ();
 sg13g2_decap_8 FILLER_37_1112 ();
 sg13g2_decap_8 FILLER_37_1119 ();
 sg13g2_decap_8 FILLER_37_1126 ();
 sg13g2_decap_8 FILLER_37_1133 ();
 sg13g2_decap_8 FILLER_37_1140 ();
 sg13g2_decap_8 FILLER_37_1147 ();
 sg13g2_decap_8 FILLER_37_1154 ();
 sg13g2_decap_8 FILLER_37_1161 ();
 sg13g2_decap_8 FILLER_37_1168 ();
 sg13g2_decap_8 FILLER_37_1175 ();
 sg13g2_decap_8 FILLER_37_1182 ();
 sg13g2_decap_8 FILLER_37_1189 ();
 sg13g2_decap_8 FILLER_37_1196 ();
 sg13g2_decap_8 FILLER_37_1203 ();
 sg13g2_decap_8 FILLER_37_1210 ();
 sg13g2_decap_8 FILLER_37_1217 ();
 sg13g2_decap_8 FILLER_37_1224 ();
 sg13g2_decap_8 FILLER_37_1231 ();
 sg13g2_decap_8 FILLER_37_1238 ();
 sg13g2_decap_8 FILLER_37_1245 ();
 sg13g2_decap_8 FILLER_37_1252 ();
 sg13g2_decap_8 FILLER_37_1259 ();
 sg13g2_decap_8 FILLER_37_1266 ();
 sg13g2_decap_8 FILLER_37_1273 ();
 sg13g2_decap_8 FILLER_37_1280 ();
 sg13g2_decap_8 FILLER_37_1287 ();
 sg13g2_decap_8 FILLER_37_1294 ();
 sg13g2_decap_8 FILLER_37_1301 ();
 sg13g2_decap_8 FILLER_37_1308 ();
 sg13g2_decap_8 FILLER_37_1315 ();
 sg13g2_decap_4 FILLER_37_1322 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_41 ();
 sg13g2_decap_4 FILLER_38_54 ();
 sg13g2_fill_1 FILLER_38_117 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_fill_1 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_366 ();
 sg13g2_fill_1 FILLER_38_378 ();
 sg13g2_fill_1 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_440 ();
 sg13g2_fill_1 FILLER_38_447 ();
 sg13g2_fill_2 FILLER_38_453 ();
 sg13g2_fill_1 FILLER_38_459 ();
 sg13g2_fill_2 FILLER_38_473 ();
 sg13g2_fill_1 FILLER_38_506 ();
 sg13g2_fill_2 FILLER_38_535 ();
 sg13g2_fill_1 FILLER_38_542 ();
 sg13g2_fill_1 FILLER_38_552 ();
 sg13g2_fill_1 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_573 ();
 sg13g2_fill_2 FILLER_38_626 ();
 sg13g2_fill_1 FILLER_38_628 ();
 sg13g2_fill_1 FILLER_38_652 ();
 sg13g2_fill_2 FILLER_38_658 ();
 sg13g2_fill_2 FILLER_38_665 ();
 sg13g2_fill_1 FILLER_38_667 ();
 sg13g2_fill_1 FILLER_38_711 ();
 sg13g2_fill_2 FILLER_38_738 ();
 sg13g2_fill_1 FILLER_38_750 ();
 sg13g2_fill_2 FILLER_38_755 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_fill_2 FILLER_38_902 ();
 sg13g2_fill_1 FILLER_38_912 ();
 sg13g2_decap_8 FILLER_38_995 ();
 sg13g2_decap_8 FILLER_38_1002 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_decap_8 FILLER_38_1016 ();
 sg13g2_decap_8 FILLER_38_1023 ();
 sg13g2_decap_8 FILLER_38_1030 ();
 sg13g2_decap_8 FILLER_38_1037 ();
 sg13g2_decap_8 FILLER_38_1044 ();
 sg13g2_decap_8 FILLER_38_1051 ();
 sg13g2_decap_8 FILLER_38_1058 ();
 sg13g2_decap_8 FILLER_38_1065 ();
 sg13g2_decap_8 FILLER_38_1072 ();
 sg13g2_decap_8 FILLER_38_1079 ();
 sg13g2_decap_8 FILLER_38_1086 ();
 sg13g2_decap_8 FILLER_38_1093 ();
 sg13g2_decap_8 FILLER_38_1100 ();
 sg13g2_decap_8 FILLER_38_1107 ();
 sg13g2_decap_8 FILLER_38_1114 ();
 sg13g2_decap_8 FILLER_38_1121 ();
 sg13g2_decap_8 FILLER_38_1128 ();
 sg13g2_decap_8 FILLER_38_1135 ();
 sg13g2_decap_8 FILLER_38_1142 ();
 sg13g2_decap_8 FILLER_38_1149 ();
 sg13g2_decap_8 FILLER_38_1156 ();
 sg13g2_decap_8 FILLER_38_1163 ();
 sg13g2_decap_8 FILLER_38_1170 ();
 sg13g2_decap_8 FILLER_38_1177 ();
 sg13g2_decap_8 FILLER_38_1184 ();
 sg13g2_decap_8 FILLER_38_1191 ();
 sg13g2_decap_8 FILLER_38_1198 ();
 sg13g2_decap_8 FILLER_38_1205 ();
 sg13g2_decap_8 FILLER_38_1212 ();
 sg13g2_decap_8 FILLER_38_1219 ();
 sg13g2_decap_8 FILLER_38_1226 ();
 sg13g2_decap_8 FILLER_38_1233 ();
 sg13g2_decap_8 FILLER_38_1240 ();
 sg13g2_decap_8 FILLER_38_1247 ();
 sg13g2_decap_8 FILLER_38_1254 ();
 sg13g2_decap_8 FILLER_38_1261 ();
 sg13g2_decap_8 FILLER_38_1268 ();
 sg13g2_decap_8 FILLER_38_1275 ();
 sg13g2_decap_8 FILLER_38_1282 ();
 sg13g2_decap_8 FILLER_38_1289 ();
 sg13g2_decap_8 FILLER_38_1296 ();
 sg13g2_decap_8 FILLER_38_1303 ();
 sg13g2_decap_8 FILLER_38_1310 ();
 sg13g2_decap_8 FILLER_38_1317 ();
 sg13g2_fill_2 FILLER_38_1324 ();
 sg13g2_fill_1 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_39 ();
 sg13g2_fill_1 FILLER_39_79 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_2 FILLER_39_163 ();
 sg13g2_fill_1 FILLER_39_173 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_fill_2 FILLER_39_211 ();
 sg13g2_fill_2 FILLER_39_218 ();
 sg13g2_fill_1 FILLER_39_220 ();
 sg13g2_fill_1 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_280 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_336 ();
 sg13g2_decap_4 FILLER_39_349 ();
 sg13g2_fill_1 FILLER_39_353 ();
 sg13g2_fill_2 FILLER_39_361 ();
 sg13g2_fill_1 FILLER_39_363 ();
 sg13g2_fill_1 FILLER_39_392 ();
 sg13g2_fill_1 FILLER_39_401 ();
 sg13g2_fill_2 FILLER_39_415 ();
 sg13g2_fill_1 FILLER_39_439 ();
 sg13g2_fill_2 FILLER_39_445 ();
 sg13g2_decap_4 FILLER_39_452 ();
 sg13g2_decap_4 FILLER_39_461 ();
 sg13g2_fill_2 FILLER_39_470 ();
 sg13g2_fill_1 FILLER_39_472 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_fill_2 FILLER_39_491 ();
 sg13g2_fill_1 FILLER_39_548 ();
 sg13g2_fill_2 FILLER_39_557 ();
 sg13g2_fill_1 FILLER_39_559 ();
 sg13g2_fill_2 FILLER_39_595 ();
 sg13g2_fill_1 FILLER_39_610 ();
 sg13g2_fill_1 FILLER_39_621 ();
 sg13g2_fill_2 FILLER_39_630 ();
 sg13g2_fill_1 FILLER_39_671 ();
 sg13g2_fill_2 FILLER_39_691 ();
 sg13g2_fill_1 FILLER_39_693 ();
 sg13g2_decap_4 FILLER_39_698 ();
 sg13g2_fill_1 FILLER_39_702 ();
 sg13g2_fill_1 FILLER_39_860 ();
 sg13g2_fill_2 FILLER_39_947 ();
 sg13g2_decap_8 FILLER_39_1001 ();
 sg13g2_decap_8 FILLER_39_1008 ();
 sg13g2_decap_8 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1022 ();
 sg13g2_decap_8 FILLER_39_1029 ();
 sg13g2_decap_8 FILLER_39_1036 ();
 sg13g2_decap_8 FILLER_39_1043 ();
 sg13g2_decap_8 FILLER_39_1050 ();
 sg13g2_decap_8 FILLER_39_1057 ();
 sg13g2_decap_8 FILLER_39_1064 ();
 sg13g2_decap_8 FILLER_39_1071 ();
 sg13g2_decap_8 FILLER_39_1078 ();
 sg13g2_decap_8 FILLER_39_1085 ();
 sg13g2_decap_8 FILLER_39_1092 ();
 sg13g2_decap_8 FILLER_39_1099 ();
 sg13g2_decap_8 FILLER_39_1106 ();
 sg13g2_decap_8 FILLER_39_1113 ();
 sg13g2_decap_8 FILLER_39_1120 ();
 sg13g2_decap_8 FILLER_39_1127 ();
 sg13g2_decap_8 FILLER_39_1134 ();
 sg13g2_decap_8 FILLER_39_1141 ();
 sg13g2_decap_8 FILLER_39_1148 ();
 sg13g2_decap_8 FILLER_39_1155 ();
 sg13g2_decap_8 FILLER_39_1162 ();
 sg13g2_decap_8 FILLER_39_1169 ();
 sg13g2_decap_8 FILLER_39_1176 ();
 sg13g2_decap_8 FILLER_39_1183 ();
 sg13g2_decap_8 FILLER_39_1190 ();
 sg13g2_decap_8 FILLER_39_1197 ();
 sg13g2_decap_8 FILLER_39_1204 ();
 sg13g2_decap_8 FILLER_39_1211 ();
 sg13g2_decap_8 FILLER_39_1218 ();
 sg13g2_decap_8 FILLER_39_1225 ();
 sg13g2_decap_8 FILLER_39_1232 ();
 sg13g2_decap_8 FILLER_39_1239 ();
 sg13g2_decap_8 FILLER_39_1246 ();
 sg13g2_decap_8 FILLER_39_1253 ();
 sg13g2_decap_8 FILLER_39_1260 ();
 sg13g2_decap_8 FILLER_39_1267 ();
 sg13g2_decap_8 FILLER_39_1274 ();
 sg13g2_decap_8 FILLER_39_1281 ();
 sg13g2_decap_8 FILLER_39_1288 ();
 sg13g2_decap_8 FILLER_39_1295 ();
 sg13g2_decap_8 FILLER_39_1302 ();
 sg13g2_decap_8 FILLER_39_1309 ();
 sg13g2_decap_8 FILLER_39_1316 ();
 sg13g2_fill_2 FILLER_39_1323 ();
 sg13g2_fill_1 FILLER_39_1325 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_5 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_decap_4 FILLER_40_68 ();
 sg13g2_fill_1 FILLER_40_105 ();
 sg13g2_fill_1 FILLER_40_161 ();
 sg13g2_fill_2 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_fill_1 FILLER_40_203 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_fill_1 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_fill_1 FILLER_40_249 ();
 sg13g2_fill_2 FILLER_40_259 ();
 sg13g2_fill_2 FILLER_40_266 ();
 sg13g2_decap_4 FILLER_40_278 ();
 sg13g2_decap_4 FILLER_40_286 ();
 sg13g2_fill_2 FILLER_40_294 ();
 sg13g2_fill_1 FILLER_40_296 ();
 sg13g2_fill_1 FILLER_40_328 ();
 sg13g2_fill_1 FILLER_40_338 ();
 sg13g2_fill_2 FILLER_40_399 ();
 sg13g2_fill_1 FILLER_40_416 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_fill_2 FILLER_40_464 ();
 sg13g2_fill_1 FILLER_40_486 ();
 sg13g2_fill_1 FILLER_40_513 ();
 sg13g2_fill_1 FILLER_40_519 ();
 sg13g2_fill_2 FILLER_40_530 ();
 sg13g2_fill_1 FILLER_40_541 ();
 sg13g2_fill_1 FILLER_40_556 ();
 sg13g2_fill_1 FILLER_40_585 ();
 sg13g2_fill_1 FILLER_40_591 ();
 sg13g2_fill_2 FILLER_40_643 ();
 sg13g2_fill_1 FILLER_40_650 ();
 sg13g2_fill_1 FILLER_40_658 ();
 sg13g2_fill_1 FILLER_40_663 ();
 sg13g2_fill_2 FILLER_40_668 ();
 sg13g2_fill_1 FILLER_40_675 ();
 sg13g2_fill_1 FILLER_40_680 ();
 sg13g2_fill_1 FILLER_40_687 ();
 sg13g2_fill_1 FILLER_40_714 ();
 sg13g2_fill_1 FILLER_40_719 ();
 sg13g2_fill_2 FILLER_40_724 ();
 sg13g2_fill_2 FILLER_40_730 ();
 sg13g2_fill_2 FILLER_40_742 ();
 sg13g2_fill_1 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_823 ();
 sg13g2_fill_1 FILLER_40_833 ();
 sg13g2_fill_2 FILLER_40_892 ();
 sg13g2_fill_2 FILLER_40_930 ();
 sg13g2_fill_1 FILLER_40_932 ();
 sg13g2_fill_2 FILLER_40_969 ();
 sg13g2_fill_1 FILLER_40_981 ();
 sg13g2_fill_2 FILLER_40_986 ();
 sg13g2_fill_1 FILLER_40_988 ();
 sg13g2_decap_8 FILLER_40_993 ();
 sg13g2_decap_8 FILLER_40_1000 ();
 sg13g2_decap_8 FILLER_40_1007 ();
 sg13g2_decap_8 FILLER_40_1014 ();
 sg13g2_decap_8 FILLER_40_1021 ();
 sg13g2_decap_8 FILLER_40_1028 ();
 sg13g2_decap_8 FILLER_40_1035 ();
 sg13g2_decap_8 FILLER_40_1042 ();
 sg13g2_decap_8 FILLER_40_1049 ();
 sg13g2_decap_8 FILLER_40_1056 ();
 sg13g2_decap_8 FILLER_40_1063 ();
 sg13g2_decap_8 FILLER_40_1070 ();
 sg13g2_decap_8 FILLER_40_1077 ();
 sg13g2_decap_8 FILLER_40_1084 ();
 sg13g2_decap_8 FILLER_40_1091 ();
 sg13g2_decap_8 FILLER_40_1098 ();
 sg13g2_decap_8 FILLER_40_1105 ();
 sg13g2_decap_8 FILLER_40_1112 ();
 sg13g2_decap_8 FILLER_40_1119 ();
 sg13g2_decap_8 FILLER_40_1126 ();
 sg13g2_decap_8 FILLER_40_1133 ();
 sg13g2_decap_8 FILLER_40_1140 ();
 sg13g2_decap_8 FILLER_40_1147 ();
 sg13g2_decap_8 FILLER_40_1154 ();
 sg13g2_decap_8 FILLER_40_1161 ();
 sg13g2_decap_8 FILLER_40_1168 ();
 sg13g2_decap_8 FILLER_40_1175 ();
 sg13g2_decap_8 FILLER_40_1182 ();
 sg13g2_decap_8 FILLER_40_1189 ();
 sg13g2_decap_8 FILLER_40_1196 ();
 sg13g2_decap_8 FILLER_40_1203 ();
 sg13g2_decap_8 FILLER_40_1210 ();
 sg13g2_decap_8 FILLER_40_1217 ();
 sg13g2_decap_8 FILLER_40_1224 ();
 sg13g2_decap_8 FILLER_40_1231 ();
 sg13g2_decap_8 FILLER_40_1238 ();
 sg13g2_decap_8 FILLER_40_1245 ();
 sg13g2_decap_8 FILLER_40_1252 ();
 sg13g2_decap_8 FILLER_40_1259 ();
 sg13g2_decap_8 FILLER_40_1266 ();
 sg13g2_decap_8 FILLER_40_1273 ();
 sg13g2_decap_8 FILLER_40_1280 ();
 sg13g2_decap_8 FILLER_40_1287 ();
 sg13g2_decap_8 FILLER_40_1294 ();
 sg13g2_decap_8 FILLER_40_1301 ();
 sg13g2_decap_8 FILLER_40_1308 ();
 sg13g2_decap_8 FILLER_40_1315 ();
 sg13g2_decap_4 FILLER_40_1322 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_11 ();
 sg13g2_fill_2 FILLER_41_16 ();
 sg13g2_fill_2 FILLER_41_22 ();
 sg13g2_fill_1 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_112 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_fill_2 FILLER_41_152 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_fill_2 FILLER_41_218 ();
 sg13g2_fill_1 FILLER_41_239 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_fill_2 FILLER_41_296 ();
 sg13g2_fill_1 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_320 ();
 sg13g2_fill_1 FILLER_41_325 ();
 sg13g2_fill_1 FILLER_41_331 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_fill_2 FILLER_41_347 ();
 sg13g2_fill_2 FILLER_41_354 ();
 sg13g2_fill_2 FILLER_41_360 ();
 sg13g2_fill_1 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_373 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_392 ();
 sg13g2_fill_2 FILLER_41_398 ();
 sg13g2_fill_2 FILLER_41_422 ();
 sg13g2_decap_8 FILLER_41_430 ();
 sg13g2_decap_4 FILLER_41_448 ();
 sg13g2_decap_4 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_466 ();
 sg13g2_fill_1 FILLER_41_477 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_fill_1 FILLER_41_508 ();
 sg13g2_fill_2 FILLER_41_524 ();
 sg13g2_fill_2 FILLER_41_544 ();
 sg13g2_fill_2 FILLER_41_550 ();
 sg13g2_fill_1 FILLER_41_561 ();
 sg13g2_fill_1 FILLER_41_616 ();
 sg13g2_fill_1 FILLER_41_631 ();
 sg13g2_fill_1 FILLER_41_648 ();
 sg13g2_fill_2 FILLER_41_654 ();
 sg13g2_fill_2 FILLER_41_665 ();
 sg13g2_fill_2 FILLER_41_671 ();
 sg13g2_fill_1 FILLER_41_673 ();
 sg13g2_fill_1 FILLER_41_678 ();
 sg13g2_fill_2 FILLER_41_683 ();
 sg13g2_decap_4 FILLER_41_699 ();
 sg13g2_fill_1 FILLER_41_703 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_739 ();
 sg13g2_fill_2 FILLER_41_766 ();
 sg13g2_fill_1 FILLER_41_794 ();
 sg13g2_fill_2 FILLER_41_799 ();
 sg13g2_fill_1 FILLER_41_811 ();
 sg13g2_fill_1 FILLER_41_838 ();
 sg13g2_fill_1 FILLER_41_865 ();
 sg13g2_fill_1 FILLER_41_876 ();
 sg13g2_fill_2 FILLER_41_923 ();
 sg13g2_fill_1 FILLER_41_925 ();
 sg13g2_fill_2 FILLER_41_940 ();
 sg13g2_fill_2 FILLER_41_950 ();
 sg13g2_decap_4 FILLER_41_978 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_41_1029 ();
 sg13g2_decap_8 FILLER_41_1036 ();
 sg13g2_decap_8 FILLER_41_1043 ();
 sg13g2_decap_8 FILLER_41_1050 ();
 sg13g2_decap_8 FILLER_41_1057 ();
 sg13g2_decap_8 FILLER_41_1064 ();
 sg13g2_decap_8 FILLER_41_1071 ();
 sg13g2_decap_8 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1085 ();
 sg13g2_decap_8 FILLER_41_1092 ();
 sg13g2_decap_8 FILLER_41_1099 ();
 sg13g2_decap_8 FILLER_41_1106 ();
 sg13g2_decap_8 FILLER_41_1113 ();
 sg13g2_decap_8 FILLER_41_1120 ();
 sg13g2_decap_8 FILLER_41_1127 ();
 sg13g2_decap_8 FILLER_41_1134 ();
 sg13g2_decap_8 FILLER_41_1141 ();
 sg13g2_decap_8 FILLER_41_1148 ();
 sg13g2_decap_8 FILLER_41_1155 ();
 sg13g2_decap_8 FILLER_41_1162 ();
 sg13g2_decap_8 FILLER_41_1169 ();
 sg13g2_decap_8 FILLER_41_1176 ();
 sg13g2_decap_8 FILLER_41_1183 ();
 sg13g2_decap_8 FILLER_41_1190 ();
 sg13g2_decap_8 FILLER_41_1197 ();
 sg13g2_decap_8 FILLER_41_1204 ();
 sg13g2_decap_8 FILLER_41_1211 ();
 sg13g2_decap_8 FILLER_41_1218 ();
 sg13g2_decap_8 FILLER_41_1225 ();
 sg13g2_decap_8 FILLER_41_1232 ();
 sg13g2_decap_8 FILLER_41_1239 ();
 sg13g2_decap_8 FILLER_41_1246 ();
 sg13g2_decap_8 FILLER_41_1253 ();
 sg13g2_decap_8 FILLER_41_1260 ();
 sg13g2_decap_8 FILLER_41_1267 ();
 sg13g2_decap_8 FILLER_41_1274 ();
 sg13g2_decap_8 FILLER_41_1281 ();
 sg13g2_decap_8 FILLER_41_1288 ();
 sg13g2_decap_8 FILLER_41_1295 ();
 sg13g2_decap_8 FILLER_41_1302 ();
 sg13g2_decap_8 FILLER_41_1309 ();
 sg13g2_decap_8 FILLER_41_1316 ();
 sg13g2_fill_2 FILLER_41_1323 ();
 sg13g2_fill_1 FILLER_41_1325 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_6 ();
 sg13g2_fill_1 FILLER_42_8 ();
 sg13g2_fill_1 FILLER_42_35 ();
 sg13g2_fill_2 FILLER_42_40 ();
 sg13g2_fill_1 FILLER_42_42 ();
 sg13g2_decap_4 FILLER_42_53 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_fill_1 FILLER_42_62 ();
 sg13g2_fill_1 FILLER_42_87 ();
 sg13g2_fill_1 FILLER_42_135 ();
 sg13g2_fill_1 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_173 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_fill_2 FILLER_42_230 ();
 sg13g2_fill_1 FILLER_42_232 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_248 ();
 sg13g2_fill_1 FILLER_42_259 ();
 sg13g2_fill_2 FILLER_42_270 ();
 sg13g2_fill_1 FILLER_42_272 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_284 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_decap_4 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_42_361 ();
 sg13g2_fill_2 FILLER_42_381 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_419 ();
 sg13g2_fill_2 FILLER_42_425 ();
 sg13g2_fill_2 FILLER_42_448 ();
 sg13g2_fill_2 FILLER_42_525 ();
 sg13g2_fill_1 FILLER_42_532 ();
 sg13g2_fill_2 FILLER_42_547 ();
 sg13g2_fill_2 FILLER_42_577 ();
 sg13g2_fill_2 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_699 ();
 sg13g2_fill_1 FILLER_42_707 ();
 sg13g2_fill_2 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_fill_1 FILLER_42_737 ();
 sg13g2_fill_1 FILLER_42_752 ();
 sg13g2_fill_1 FILLER_42_783 ();
 sg13g2_fill_2 FILLER_42_848 ();
 sg13g2_fill_2 FILLER_42_876 ();
 sg13g2_fill_1 FILLER_42_878 ();
 sg13g2_fill_2 FILLER_42_893 ();
 sg13g2_fill_1 FILLER_42_895 ();
 sg13g2_fill_1 FILLER_42_958 ();
 sg13g2_decap_8 FILLER_42_995 ();
 sg13g2_decap_8 FILLER_42_1002 ();
 sg13g2_decap_8 FILLER_42_1009 ();
 sg13g2_decap_8 FILLER_42_1016 ();
 sg13g2_decap_8 FILLER_42_1023 ();
 sg13g2_decap_8 FILLER_42_1030 ();
 sg13g2_decap_8 FILLER_42_1037 ();
 sg13g2_decap_8 FILLER_42_1044 ();
 sg13g2_decap_8 FILLER_42_1051 ();
 sg13g2_decap_8 FILLER_42_1058 ();
 sg13g2_decap_8 FILLER_42_1065 ();
 sg13g2_decap_8 FILLER_42_1072 ();
 sg13g2_decap_8 FILLER_42_1079 ();
 sg13g2_decap_8 FILLER_42_1086 ();
 sg13g2_decap_8 FILLER_42_1093 ();
 sg13g2_decap_8 FILLER_42_1100 ();
 sg13g2_decap_8 FILLER_42_1107 ();
 sg13g2_decap_8 FILLER_42_1114 ();
 sg13g2_decap_8 FILLER_42_1121 ();
 sg13g2_decap_8 FILLER_42_1128 ();
 sg13g2_decap_8 FILLER_42_1135 ();
 sg13g2_decap_8 FILLER_42_1142 ();
 sg13g2_decap_8 FILLER_42_1149 ();
 sg13g2_decap_8 FILLER_42_1156 ();
 sg13g2_decap_8 FILLER_42_1163 ();
 sg13g2_decap_8 FILLER_42_1170 ();
 sg13g2_decap_8 FILLER_42_1177 ();
 sg13g2_decap_8 FILLER_42_1184 ();
 sg13g2_decap_8 FILLER_42_1191 ();
 sg13g2_decap_8 FILLER_42_1198 ();
 sg13g2_decap_8 FILLER_42_1205 ();
 sg13g2_decap_8 FILLER_42_1212 ();
 sg13g2_decap_8 FILLER_42_1219 ();
 sg13g2_decap_8 FILLER_42_1226 ();
 sg13g2_decap_8 FILLER_42_1233 ();
 sg13g2_decap_8 FILLER_42_1240 ();
 sg13g2_decap_8 FILLER_42_1247 ();
 sg13g2_decap_8 FILLER_42_1254 ();
 sg13g2_decap_8 FILLER_42_1261 ();
 sg13g2_decap_8 FILLER_42_1268 ();
 sg13g2_decap_8 FILLER_42_1275 ();
 sg13g2_decap_8 FILLER_42_1282 ();
 sg13g2_decap_8 FILLER_42_1289 ();
 sg13g2_decap_8 FILLER_42_1296 ();
 sg13g2_decap_8 FILLER_42_1303 ();
 sg13g2_decap_8 FILLER_42_1310 ();
 sg13g2_decap_8 FILLER_42_1317 ();
 sg13g2_fill_2 FILLER_42_1324 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_13 ();
 sg13g2_fill_2 FILLER_43_18 ();
 sg13g2_fill_1 FILLER_43_20 ();
 sg13g2_fill_1 FILLER_43_25 ();
 sg13g2_fill_1 FILLER_43_40 ();
 sg13g2_fill_1 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_104 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_fill_1 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_205 ();
 sg13g2_fill_1 FILLER_43_250 ();
 sg13g2_fill_1 FILLER_43_255 ();
 sg13g2_fill_1 FILLER_43_337 ();
 sg13g2_fill_1 FILLER_43_346 ();
 sg13g2_decap_4 FILLER_43_351 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_fill_1 FILLER_43_366 ();
 sg13g2_fill_1 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_382 ();
 sg13g2_fill_1 FILLER_43_411 ();
 sg13g2_decap_4 FILLER_43_428 ();
 sg13g2_fill_1 FILLER_43_432 ();
 sg13g2_fill_1 FILLER_43_441 ();
 sg13g2_decap_4 FILLER_43_452 ();
 sg13g2_fill_2 FILLER_43_456 ();
 sg13g2_fill_2 FILLER_43_462 ();
 sg13g2_fill_2 FILLER_43_504 ();
 sg13g2_fill_2 FILLER_43_558 ();
 sg13g2_fill_1 FILLER_43_560 ();
 sg13g2_fill_2 FILLER_43_584 ();
 sg13g2_fill_2 FILLER_43_607 ();
 sg13g2_fill_2 FILLER_43_614 ();
 sg13g2_fill_2 FILLER_43_626 ();
 sg13g2_fill_2 FILLER_43_677 ();
 sg13g2_fill_2 FILLER_43_771 ();
 sg13g2_fill_1 FILLER_43_773 ();
 sg13g2_fill_1 FILLER_43_782 ();
 sg13g2_fill_1 FILLER_43_793 ();
 sg13g2_fill_2 FILLER_43_817 ();
 sg13g2_fill_2 FILLER_43_941 ();
 sg13g2_fill_1 FILLER_43_943 ();
 sg13g2_fill_1 FILLER_43_962 ();
 sg13g2_decap_8 FILLER_43_1003 ();
 sg13g2_decap_8 FILLER_43_1010 ();
 sg13g2_decap_8 FILLER_43_1017 ();
 sg13g2_decap_8 FILLER_43_1024 ();
 sg13g2_decap_8 FILLER_43_1031 ();
 sg13g2_decap_8 FILLER_43_1038 ();
 sg13g2_decap_8 FILLER_43_1045 ();
 sg13g2_decap_8 FILLER_43_1052 ();
 sg13g2_decap_8 FILLER_43_1059 ();
 sg13g2_decap_8 FILLER_43_1066 ();
 sg13g2_decap_8 FILLER_43_1073 ();
 sg13g2_decap_8 FILLER_43_1080 ();
 sg13g2_decap_8 FILLER_43_1087 ();
 sg13g2_decap_8 FILLER_43_1094 ();
 sg13g2_decap_8 FILLER_43_1101 ();
 sg13g2_decap_8 FILLER_43_1108 ();
 sg13g2_decap_8 FILLER_43_1115 ();
 sg13g2_decap_8 FILLER_43_1122 ();
 sg13g2_decap_8 FILLER_43_1129 ();
 sg13g2_decap_8 FILLER_43_1136 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1150 ();
 sg13g2_decap_8 FILLER_43_1157 ();
 sg13g2_decap_8 FILLER_43_1164 ();
 sg13g2_decap_8 FILLER_43_1171 ();
 sg13g2_decap_8 FILLER_43_1178 ();
 sg13g2_decap_8 FILLER_43_1185 ();
 sg13g2_decap_8 FILLER_43_1192 ();
 sg13g2_decap_8 FILLER_43_1199 ();
 sg13g2_decap_8 FILLER_43_1206 ();
 sg13g2_decap_8 FILLER_43_1213 ();
 sg13g2_decap_8 FILLER_43_1220 ();
 sg13g2_decap_8 FILLER_43_1227 ();
 sg13g2_decap_8 FILLER_43_1234 ();
 sg13g2_decap_8 FILLER_43_1241 ();
 sg13g2_decap_8 FILLER_43_1248 ();
 sg13g2_decap_8 FILLER_43_1255 ();
 sg13g2_decap_8 FILLER_43_1262 ();
 sg13g2_decap_8 FILLER_43_1269 ();
 sg13g2_decap_8 FILLER_43_1276 ();
 sg13g2_decap_8 FILLER_43_1283 ();
 sg13g2_decap_8 FILLER_43_1290 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_8 FILLER_43_1304 ();
 sg13g2_decap_8 FILLER_43_1311 ();
 sg13g2_decap_8 FILLER_43_1318 ();
 sg13g2_fill_1 FILLER_43_1325 ();
 sg13g2_fill_1 FILLER_44_44 ();
 sg13g2_fill_2 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_99 ();
 sg13g2_fill_1 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_166 ();
 sg13g2_fill_2 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_357 ();
 sg13g2_fill_1 FILLER_44_363 ();
 sg13g2_fill_2 FILLER_44_376 ();
 sg13g2_fill_1 FILLER_44_396 ();
 sg13g2_fill_1 FILLER_44_415 ();
 sg13g2_fill_1 FILLER_44_420 ();
 sg13g2_fill_1 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_430 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_decap_8 FILLER_44_450 ();
 sg13g2_decap_8 FILLER_44_461 ();
 sg13g2_fill_1 FILLER_44_473 ();
 sg13g2_fill_1 FILLER_44_478 ();
 sg13g2_fill_2 FILLER_44_544 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_decap_4 FILLER_44_555 ();
 sg13g2_fill_1 FILLER_44_559 ();
 sg13g2_fill_1 FILLER_44_575 ();
 sg13g2_fill_2 FILLER_44_586 ();
 sg13g2_decap_4 FILLER_44_591 ();
 sg13g2_fill_1 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_601 ();
 sg13g2_fill_2 FILLER_44_608 ();
 sg13g2_fill_1 FILLER_44_610 ();
 sg13g2_fill_2 FILLER_44_614 ();
 sg13g2_fill_1 FILLER_44_665 ();
 sg13g2_fill_2 FILLER_44_707 ();
 sg13g2_fill_2 FILLER_44_715 ();
 sg13g2_fill_1 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_726 ();
 sg13g2_fill_1 FILLER_44_818 ();
 sg13g2_fill_2 FILLER_44_881 ();
 sg13g2_fill_1 FILLER_44_883 ();
 sg13g2_fill_2 FILLER_44_920 ();
 sg13g2_fill_1 FILLER_44_922 ();
 sg13g2_fill_2 FILLER_44_989 ();
 sg13g2_decap_8 FILLER_44_995 ();
 sg13g2_decap_8 FILLER_44_1002 ();
 sg13g2_decap_8 FILLER_44_1009 ();
 sg13g2_decap_8 FILLER_44_1016 ();
 sg13g2_decap_8 FILLER_44_1023 ();
 sg13g2_decap_8 FILLER_44_1030 ();
 sg13g2_decap_8 FILLER_44_1037 ();
 sg13g2_decap_8 FILLER_44_1044 ();
 sg13g2_decap_8 FILLER_44_1051 ();
 sg13g2_decap_8 FILLER_44_1058 ();
 sg13g2_decap_8 FILLER_44_1065 ();
 sg13g2_decap_8 FILLER_44_1072 ();
 sg13g2_decap_8 FILLER_44_1079 ();
 sg13g2_decap_8 FILLER_44_1086 ();
 sg13g2_decap_8 FILLER_44_1093 ();
 sg13g2_decap_8 FILLER_44_1100 ();
 sg13g2_decap_8 FILLER_44_1107 ();
 sg13g2_decap_8 FILLER_44_1114 ();
 sg13g2_decap_8 FILLER_44_1121 ();
 sg13g2_decap_8 FILLER_44_1128 ();
 sg13g2_decap_8 FILLER_44_1135 ();
 sg13g2_decap_8 FILLER_44_1142 ();
 sg13g2_decap_8 FILLER_44_1149 ();
 sg13g2_decap_8 FILLER_44_1156 ();
 sg13g2_decap_8 FILLER_44_1163 ();
 sg13g2_decap_8 FILLER_44_1170 ();
 sg13g2_decap_8 FILLER_44_1177 ();
 sg13g2_decap_8 FILLER_44_1184 ();
 sg13g2_decap_8 FILLER_44_1191 ();
 sg13g2_decap_8 FILLER_44_1198 ();
 sg13g2_decap_8 FILLER_44_1205 ();
 sg13g2_decap_8 FILLER_44_1212 ();
 sg13g2_decap_8 FILLER_44_1219 ();
 sg13g2_decap_8 FILLER_44_1226 ();
 sg13g2_decap_8 FILLER_44_1233 ();
 sg13g2_decap_8 FILLER_44_1240 ();
 sg13g2_decap_8 FILLER_44_1247 ();
 sg13g2_decap_8 FILLER_44_1254 ();
 sg13g2_decap_8 FILLER_44_1261 ();
 sg13g2_decap_8 FILLER_44_1268 ();
 sg13g2_decap_8 FILLER_44_1275 ();
 sg13g2_decap_8 FILLER_44_1282 ();
 sg13g2_decap_8 FILLER_44_1289 ();
 sg13g2_decap_8 FILLER_44_1296 ();
 sg13g2_decap_8 FILLER_44_1303 ();
 sg13g2_decap_8 FILLER_44_1310 ();
 sg13g2_decap_8 FILLER_44_1317 ();
 sg13g2_fill_2 FILLER_44_1324 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_34 ();
 sg13g2_fill_1 FILLER_45_36 ();
 sg13g2_fill_2 FILLER_45_57 ();
 sg13g2_fill_2 FILLER_45_85 ();
 sg13g2_fill_1 FILLER_45_87 ();
 sg13g2_fill_1 FILLER_45_92 ();
 sg13g2_fill_1 FILLER_45_139 ();
 sg13g2_fill_1 FILLER_45_153 ();
 sg13g2_fill_2 FILLER_45_217 ();
 sg13g2_decap_4 FILLER_45_223 ();
 sg13g2_decap_8 FILLER_45_235 ();
 sg13g2_fill_1 FILLER_45_242 ();
 sg13g2_fill_2 FILLER_45_257 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_fill_2 FILLER_45_281 ();
 sg13g2_fill_1 FILLER_45_283 ();
 sg13g2_fill_1 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_fill_1 FILLER_45_344 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_2 FILLER_45_355 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_368 ();
 sg13g2_fill_2 FILLER_45_415 ();
 sg13g2_fill_2 FILLER_45_422 ();
 sg13g2_fill_1 FILLER_45_424 ();
 sg13g2_decap_4 FILLER_45_462 ();
 sg13g2_fill_1 FILLER_45_466 ();
 sg13g2_fill_2 FILLER_45_534 ();
 sg13g2_fill_1 FILLER_45_585 ();
 sg13g2_fill_1 FILLER_45_612 ();
 sg13g2_fill_1 FILLER_45_647 ();
 sg13g2_fill_1 FILLER_45_666 ();
 sg13g2_fill_2 FILLER_45_672 ();
 sg13g2_fill_2 FILLER_45_678 ();
 sg13g2_fill_1 FILLER_45_706 ();
 sg13g2_fill_2 FILLER_45_780 ();
 sg13g2_fill_1 FILLER_45_796 ();
 sg13g2_fill_2 FILLER_45_917 ();
 sg13g2_fill_1 FILLER_45_919 ();
 sg13g2_fill_2 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_45_1029 ();
 sg13g2_decap_8 FILLER_45_1036 ();
 sg13g2_decap_8 FILLER_45_1043 ();
 sg13g2_decap_8 FILLER_45_1050 ();
 sg13g2_decap_8 FILLER_45_1057 ();
 sg13g2_decap_8 FILLER_45_1064 ();
 sg13g2_decap_8 FILLER_45_1071 ();
 sg13g2_decap_8 FILLER_45_1078 ();
 sg13g2_decap_8 FILLER_45_1085 ();
 sg13g2_decap_8 FILLER_45_1092 ();
 sg13g2_decap_8 FILLER_45_1099 ();
 sg13g2_decap_8 FILLER_45_1106 ();
 sg13g2_decap_8 FILLER_45_1113 ();
 sg13g2_decap_8 FILLER_45_1120 ();
 sg13g2_decap_8 FILLER_45_1127 ();
 sg13g2_decap_8 FILLER_45_1134 ();
 sg13g2_decap_8 FILLER_45_1141 ();
 sg13g2_decap_8 FILLER_45_1148 ();
 sg13g2_decap_8 FILLER_45_1155 ();
 sg13g2_decap_8 FILLER_45_1162 ();
 sg13g2_decap_8 FILLER_45_1169 ();
 sg13g2_decap_8 FILLER_45_1176 ();
 sg13g2_decap_8 FILLER_45_1183 ();
 sg13g2_decap_8 FILLER_45_1190 ();
 sg13g2_decap_8 FILLER_45_1197 ();
 sg13g2_decap_8 FILLER_45_1204 ();
 sg13g2_decap_8 FILLER_45_1211 ();
 sg13g2_decap_8 FILLER_45_1218 ();
 sg13g2_decap_8 FILLER_45_1225 ();
 sg13g2_decap_8 FILLER_45_1232 ();
 sg13g2_decap_8 FILLER_45_1239 ();
 sg13g2_decap_8 FILLER_45_1246 ();
 sg13g2_decap_8 FILLER_45_1253 ();
 sg13g2_decap_8 FILLER_45_1260 ();
 sg13g2_decap_8 FILLER_45_1267 ();
 sg13g2_decap_8 FILLER_45_1274 ();
 sg13g2_decap_8 FILLER_45_1281 ();
 sg13g2_decap_8 FILLER_45_1288 ();
 sg13g2_decap_8 FILLER_45_1295 ();
 sg13g2_decap_8 FILLER_45_1302 ();
 sg13g2_decap_8 FILLER_45_1309 ();
 sg13g2_decap_8 FILLER_45_1316 ();
 sg13g2_fill_2 FILLER_45_1323 ();
 sg13g2_fill_1 FILLER_45_1325 ();
 sg13g2_fill_1 FILLER_46_30 ();
 sg13g2_fill_1 FILLER_46_100 ();
 sg13g2_fill_2 FILLER_46_137 ();
 sg13g2_fill_2 FILLER_46_168 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_190 ();
 sg13g2_decap_4 FILLER_46_206 ();
 sg13g2_fill_1 FILLER_46_210 ();
 sg13g2_fill_1 FILLER_46_308 ();
 sg13g2_fill_1 FILLER_46_313 ();
 sg13g2_fill_2 FILLER_46_319 ();
 sg13g2_fill_1 FILLER_46_326 ();
 sg13g2_fill_2 FILLER_46_331 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_344 ();
 sg13g2_fill_1 FILLER_46_349 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_fill_1 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_410 ();
 sg13g2_fill_2 FILLER_46_432 ();
 sg13g2_fill_1 FILLER_46_434 ();
 sg13g2_fill_1 FILLER_46_445 ();
 sg13g2_fill_1 FILLER_46_453 ();
 sg13g2_fill_1 FILLER_46_467 ();
 sg13g2_fill_1 FILLER_46_472 ();
 sg13g2_fill_2 FILLER_46_477 ();
 sg13g2_fill_1 FILLER_46_483 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_1 FILLER_46_500 ();
 sg13g2_fill_1 FILLER_46_506 ();
 sg13g2_fill_1 FILLER_46_518 ();
 sg13g2_fill_1 FILLER_46_528 ();
 sg13g2_fill_2 FILLER_46_533 ();
 sg13g2_fill_1 FILLER_46_556 ();
 sg13g2_fill_1 FILLER_46_640 ();
 sg13g2_fill_2 FILLER_46_740 ();
 sg13g2_fill_2 FILLER_46_760 ();
 sg13g2_fill_1 FILLER_46_762 ();
 sg13g2_fill_1 FILLER_46_833 ();
 sg13g2_fill_2 FILLER_46_957 ();
 sg13g2_decap_8 FILLER_46_985 ();
 sg13g2_decap_8 FILLER_46_992 ();
 sg13g2_decap_8 FILLER_46_999 ();
 sg13g2_decap_8 FILLER_46_1006 ();
 sg13g2_decap_8 FILLER_46_1013 ();
 sg13g2_decap_8 FILLER_46_1020 ();
 sg13g2_decap_8 FILLER_46_1027 ();
 sg13g2_decap_8 FILLER_46_1034 ();
 sg13g2_decap_8 FILLER_46_1041 ();
 sg13g2_decap_8 FILLER_46_1048 ();
 sg13g2_decap_8 FILLER_46_1055 ();
 sg13g2_decap_8 FILLER_46_1062 ();
 sg13g2_decap_8 FILLER_46_1069 ();
 sg13g2_decap_8 FILLER_46_1076 ();
 sg13g2_decap_8 FILLER_46_1083 ();
 sg13g2_decap_8 FILLER_46_1090 ();
 sg13g2_decap_8 FILLER_46_1097 ();
 sg13g2_decap_8 FILLER_46_1104 ();
 sg13g2_decap_8 FILLER_46_1111 ();
 sg13g2_decap_8 FILLER_46_1118 ();
 sg13g2_decap_8 FILLER_46_1125 ();
 sg13g2_decap_8 FILLER_46_1132 ();
 sg13g2_decap_8 FILLER_46_1139 ();
 sg13g2_decap_8 FILLER_46_1146 ();
 sg13g2_decap_8 FILLER_46_1153 ();
 sg13g2_decap_8 FILLER_46_1160 ();
 sg13g2_decap_8 FILLER_46_1167 ();
 sg13g2_decap_8 FILLER_46_1174 ();
 sg13g2_decap_8 FILLER_46_1181 ();
 sg13g2_decap_8 FILLER_46_1188 ();
 sg13g2_decap_8 FILLER_46_1195 ();
 sg13g2_decap_8 FILLER_46_1202 ();
 sg13g2_decap_8 FILLER_46_1209 ();
 sg13g2_decap_8 FILLER_46_1216 ();
 sg13g2_decap_8 FILLER_46_1223 ();
 sg13g2_decap_8 FILLER_46_1230 ();
 sg13g2_decap_8 FILLER_46_1237 ();
 sg13g2_decap_8 FILLER_46_1244 ();
 sg13g2_decap_8 FILLER_46_1251 ();
 sg13g2_decap_8 FILLER_46_1258 ();
 sg13g2_decap_8 FILLER_46_1265 ();
 sg13g2_decap_8 FILLER_46_1272 ();
 sg13g2_decap_8 FILLER_46_1279 ();
 sg13g2_decap_8 FILLER_46_1286 ();
 sg13g2_decap_8 FILLER_46_1293 ();
 sg13g2_decap_8 FILLER_46_1300 ();
 sg13g2_decap_8 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1314 ();
 sg13g2_decap_4 FILLER_46_1321 ();
 sg13g2_fill_1 FILLER_46_1325 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_134 ();
 sg13g2_fill_2 FILLER_47_196 ();
 sg13g2_fill_1 FILLER_47_198 ();
 sg13g2_decap_4 FILLER_47_225 ();
 sg13g2_decap_8 FILLER_47_233 ();
 sg13g2_decap_8 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_decap_4 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_decap_4 FILLER_47_380 ();
 sg13g2_fill_1 FILLER_47_384 ();
 sg13g2_fill_2 FILLER_47_469 ();
 sg13g2_fill_1 FILLER_47_493 ();
 sg13g2_fill_1 FILLER_47_498 ();
 sg13g2_fill_1 FILLER_47_515 ();
 sg13g2_fill_1 FILLER_47_560 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_607 ();
 sg13g2_fill_2 FILLER_47_621 ();
 sg13g2_fill_1 FILLER_47_645 ();
 sg13g2_fill_2 FILLER_47_704 ();
 sg13g2_fill_1 FILLER_47_711 ();
 sg13g2_fill_2 FILLER_47_739 ();
 sg13g2_fill_2 FILLER_47_775 ();
 sg13g2_fill_1 FILLER_47_777 ();
 sg13g2_fill_2 FILLER_47_788 ();
 sg13g2_fill_1 FILLER_47_790 ();
 sg13g2_fill_2 FILLER_47_855 ();
 sg13g2_fill_2 FILLER_47_871 ();
 sg13g2_fill_1 FILLER_47_873 ();
 sg13g2_decap_8 FILLER_47_990 ();
 sg13g2_decap_8 FILLER_47_997 ();
 sg13g2_decap_8 FILLER_47_1004 ();
 sg13g2_decap_8 FILLER_47_1011 ();
 sg13g2_decap_8 FILLER_47_1018 ();
 sg13g2_decap_8 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_47_1032 ();
 sg13g2_decap_8 FILLER_47_1039 ();
 sg13g2_decap_8 FILLER_47_1046 ();
 sg13g2_decap_8 FILLER_47_1053 ();
 sg13g2_decap_8 FILLER_47_1060 ();
 sg13g2_decap_8 FILLER_47_1067 ();
 sg13g2_decap_8 FILLER_47_1074 ();
 sg13g2_decap_8 FILLER_47_1081 ();
 sg13g2_decap_8 FILLER_47_1088 ();
 sg13g2_decap_8 FILLER_47_1095 ();
 sg13g2_decap_8 FILLER_47_1102 ();
 sg13g2_decap_8 FILLER_47_1109 ();
 sg13g2_decap_8 FILLER_47_1116 ();
 sg13g2_decap_8 FILLER_47_1123 ();
 sg13g2_decap_8 FILLER_47_1130 ();
 sg13g2_decap_8 FILLER_47_1137 ();
 sg13g2_decap_8 FILLER_47_1144 ();
 sg13g2_decap_8 FILLER_47_1151 ();
 sg13g2_decap_8 FILLER_47_1158 ();
 sg13g2_decap_8 FILLER_47_1165 ();
 sg13g2_decap_8 FILLER_47_1172 ();
 sg13g2_decap_8 FILLER_47_1179 ();
 sg13g2_decap_8 FILLER_47_1186 ();
 sg13g2_decap_8 FILLER_47_1193 ();
 sg13g2_decap_8 FILLER_47_1200 ();
 sg13g2_decap_8 FILLER_47_1207 ();
 sg13g2_decap_8 FILLER_47_1214 ();
 sg13g2_decap_8 FILLER_47_1221 ();
 sg13g2_decap_8 FILLER_47_1228 ();
 sg13g2_decap_8 FILLER_47_1235 ();
 sg13g2_decap_8 FILLER_47_1242 ();
 sg13g2_decap_8 FILLER_47_1249 ();
 sg13g2_decap_8 FILLER_47_1256 ();
 sg13g2_decap_8 FILLER_47_1263 ();
 sg13g2_decap_8 FILLER_47_1270 ();
 sg13g2_decap_8 FILLER_47_1277 ();
 sg13g2_decap_8 FILLER_47_1284 ();
 sg13g2_decap_8 FILLER_47_1291 ();
 sg13g2_decap_8 FILLER_47_1298 ();
 sg13g2_decap_8 FILLER_47_1305 ();
 sg13g2_decap_8 FILLER_47_1312 ();
 sg13g2_decap_8 FILLER_47_1319 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_60 ();
 sg13g2_fill_2 FILLER_48_97 ();
 sg13g2_fill_1 FILLER_48_150 ();
 sg13g2_fill_1 FILLER_48_155 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_202 ();
 sg13g2_fill_2 FILLER_48_207 ();
 sg13g2_fill_1 FILLER_48_235 ();
 sg13g2_fill_2 FILLER_48_240 ();
 sg13g2_fill_2 FILLER_48_247 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_280 ();
 sg13g2_fill_2 FILLER_48_290 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_355 ();
 sg13g2_fill_1 FILLER_48_357 ();
 sg13g2_fill_2 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_376 ();
 sg13g2_fill_1 FILLER_48_414 ();
 sg13g2_fill_1 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_443 ();
 sg13g2_fill_1 FILLER_48_448 ();
 sg13g2_fill_2 FILLER_48_453 ();
 sg13g2_fill_1 FILLER_48_602 ();
 sg13g2_fill_1 FILLER_48_608 ();
 sg13g2_fill_1 FILLER_48_635 ();
 sg13g2_fill_1 FILLER_48_737 ();
 sg13g2_fill_1 FILLER_48_764 ();
 sg13g2_fill_1 FILLER_48_791 ();
 sg13g2_fill_1 FILLER_48_800 ();
 sg13g2_fill_2 FILLER_48_815 ();
 sg13g2_fill_1 FILLER_48_817 ();
 sg13g2_fill_2 FILLER_48_880 ();
 sg13g2_fill_1 FILLER_48_926 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_48_1029 ();
 sg13g2_decap_8 FILLER_48_1036 ();
 sg13g2_decap_8 FILLER_48_1043 ();
 sg13g2_decap_8 FILLER_48_1050 ();
 sg13g2_decap_8 FILLER_48_1057 ();
 sg13g2_decap_8 FILLER_48_1064 ();
 sg13g2_decap_8 FILLER_48_1071 ();
 sg13g2_decap_8 FILLER_48_1078 ();
 sg13g2_decap_8 FILLER_48_1085 ();
 sg13g2_decap_8 FILLER_48_1092 ();
 sg13g2_decap_8 FILLER_48_1099 ();
 sg13g2_decap_8 FILLER_48_1106 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_decap_8 FILLER_48_1120 ();
 sg13g2_decap_8 FILLER_48_1127 ();
 sg13g2_decap_8 FILLER_48_1134 ();
 sg13g2_decap_8 FILLER_48_1141 ();
 sg13g2_decap_8 FILLER_48_1148 ();
 sg13g2_decap_8 FILLER_48_1155 ();
 sg13g2_decap_8 FILLER_48_1162 ();
 sg13g2_decap_8 FILLER_48_1169 ();
 sg13g2_decap_8 FILLER_48_1176 ();
 sg13g2_decap_8 FILLER_48_1183 ();
 sg13g2_decap_8 FILLER_48_1190 ();
 sg13g2_decap_8 FILLER_48_1197 ();
 sg13g2_decap_8 FILLER_48_1204 ();
 sg13g2_decap_8 FILLER_48_1211 ();
 sg13g2_decap_8 FILLER_48_1218 ();
 sg13g2_decap_8 FILLER_48_1225 ();
 sg13g2_decap_8 FILLER_48_1232 ();
 sg13g2_decap_8 FILLER_48_1239 ();
 sg13g2_decap_8 FILLER_48_1246 ();
 sg13g2_decap_8 FILLER_48_1253 ();
 sg13g2_decap_8 FILLER_48_1260 ();
 sg13g2_decap_8 FILLER_48_1267 ();
 sg13g2_decap_8 FILLER_48_1274 ();
 sg13g2_decap_8 FILLER_48_1281 ();
 sg13g2_decap_8 FILLER_48_1288 ();
 sg13g2_decap_8 FILLER_48_1295 ();
 sg13g2_decap_8 FILLER_48_1302 ();
 sg13g2_decap_8 FILLER_48_1309 ();
 sg13g2_decap_8 FILLER_48_1316 ();
 sg13g2_fill_2 FILLER_48_1323 ();
 sg13g2_fill_1 FILLER_48_1325 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_11 ();
 sg13g2_fill_1 FILLER_49_16 ();
 sg13g2_fill_2 FILLER_49_43 ();
 sg13g2_fill_1 FILLER_49_55 ();
 sg13g2_fill_2 FILLER_49_82 ();
 sg13g2_fill_1 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_222 ();
 sg13g2_fill_2 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_230 ();
 sg13g2_decap_4 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_fill_1 FILLER_49_296 ();
 sg13g2_fill_2 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_399 ();
 sg13g2_fill_1 FILLER_49_401 ();
 sg13g2_fill_1 FILLER_49_540 ();
 sg13g2_fill_2 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_fill_1 FILLER_49_648 ();
 sg13g2_fill_1 FILLER_49_663 ();
 sg13g2_fill_1 FILLER_49_669 ();
 sg13g2_fill_2 FILLER_49_745 ();
 sg13g2_fill_1 FILLER_49_747 ();
 sg13g2_fill_2 FILLER_49_792 ();
 sg13g2_fill_1 FILLER_49_820 ();
 sg13g2_fill_1 FILLER_49_847 ();
 sg13g2_fill_2 FILLER_49_919 ();
 sg13g2_fill_1 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_988 ();
 sg13g2_decap_8 FILLER_49_995 ();
 sg13g2_decap_8 FILLER_49_1002 ();
 sg13g2_decap_8 FILLER_49_1009 ();
 sg13g2_decap_8 FILLER_49_1016 ();
 sg13g2_decap_8 FILLER_49_1023 ();
 sg13g2_decap_8 FILLER_49_1030 ();
 sg13g2_decap_8 FILLER_49_1037 ();
 sg13g2_decap_8 FILLER_49_1044 ();
 sg13g2_decap_8 FILLER_49_1051 ();
 sg13g2_decap_8 FILLER_49_1058 ();
 sg13g2_decap_8 FILLER_49_1065 ();
 sg13g2_decap_8 FILLER_49_1072 ();
 sg13g2_decap_8 FILLER_49_1079 ();
 sg13g2_decap_8 FILLER_49_1086 ();
 sg13g2_decap_8 FILLER_49_1093 ();
 sg13g2_decap_8 FILLER_49_1100 ();
 sg13g2_decap_8 FILLER_49_1107 ();
 sg13g2_decap_8 FILLER_49_1114 ();
 sg13g2_decap_8 FILLER_49_1121 ();
 sg13g2_decap_8 FILLER_49_1128 ();
 sg13g2_decap_8 FILLER_49_1135 ();
 sg13g2_decap_8 FILLER_49_1142 ();
 sg13g2_decap_8 FILLER_49_1149 ();
 sg13g2_decap_8 FILLER_49_1156 ();
 sg13g2_decap_8 FILLER_49_1163 ();
 sg13g2_decap_8 FILLER_49_1170 ();
 sg13g2_decap_8 FILLER_49_1177 ();
 sg13g2_decap_8 FILLER_49_1184 ();
 sg13g2_decap_8 FILLER_49_1191 ();
 sg13g2_decap_8 FILLER_49_1198 ();
 sg13g2_decap_8 FILLER_49_1205 ();
 sg13g2_decap_8 FILLER_49_1212 ();
 sg13g2_decap_8 FILLER_49_1219 ();
 sg13g2_decap_8 FILLER_49_1226 ();
 sg13g2_decap_8 FILLER_49_1233 ();
 sg13g2_decap_8 FILLER_49_1240 ();
 sg13g2_decap_8 FILLER_49_1247 ();
 sg13g2_decap_8 FILLER_49_1254 ();
 sg13g2_decap_8 FILLER_49_1261 ();
 sg13g2_decap_8 FILLER_49_1268 ();
 sg13g2_decap_8 FILLER_49_1275 ();
 sg13g2_decap_8 FILLER_49_1282 ();
 sg13g2_decap_8 FILLER_49_1289 ();
 sg13g2_decap_8 FILLER_49_1296 ();
 sg13g2_decap_8 FILLER_49_1303 ();
 sg13g2_decap_8 FILLER_49_1310 ();
 sg13g2_decap_8 FILLER_49_1317 ();
 sg13g2_fill_2 FILLER_49_1324 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_40 ();
 sg13g2_fill_1 FILLER_50_51 ();
 sg13g2_fill_2 FILLER_50_62 ();
 sg13g2_fill_2 FILLER_50_115 ();
 sg13g2_fill_1 FILLER_50_122 ();
 sg13g2_fill_1 FILLER_50_127 ();
 sg13g2_fill_1 FILLER_50_134 ();
 sg13g2_fill_1 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_190 ();
 sg13g2_fill_2 FILLER_50_202 ();
 sg13g2_fill_1 FILLER_50_230 ();
 sg13g2_fill_1 FILLER_50_234 ();
 sg13g2_fill_1 FILLER_50_239 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_fill_1 FILLER_50_290 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_312 ();
 sg13g2_fill_2 FILLER_50_351 ();
 sg13g2_decap_4 FILLER_50_367 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_2 FILLER_50_418 ();
 sg13g2_fill_1 FILLER_50_420 ();
 sg13g2_fill_1 FILLER_50_511 ();
 sg13g2_fill_1 FILLER_50_555 ();
 sg13g2_fill_1 FILLER_50_560 ();
 sg13g2_fill_2 FILLER_50_589 ();
 sg13g2_fill_1 FILLER_50_662 ();
 sg13g2_fill_1 FILLER_50_689 ();
 sg13g2_fill_1 FILLER_50_716 ();
 sg13g2_fill_2 FILLER_50_745 ();
 sg13g2_fill_2 FILLER_50_783 ();
 sg13g2_fill_1 FILLER_50_795 ();
 sg13g2_fill_1 FILLER_50_806 ();
 sg13g2_fill_1 FILLER_50_825 ();
 sg13g2_fill_2 FILLER_50_856 ();
 sg13g2_fill_1 FILLER_50_858 ();
 sg13g2_fill_1 FILLER_50_885 ();
 sg13g2_fill_2 FILLER_50_894 ();
 sg13g2_fill_1 FILLER_50_906 ();
 sg13g2_fill_1 FILLER_50_917 ();
 sg13g2_fill_2 FILLER_50_949 ();
 sg13g2_fill_2 FILLER_50_961 ();
 sg13g2_decap_8 FILLER_50_989 ();
 sg13g2_decap_8 FILLER_50_996 ();
 sg13g2_decap_8 FILLER_50_1003 ();
 sg13g2_decap_8 FILLER_50_1010 ();
 sg13g2_decap_8 FILLER_50_1017 ();
 sg13g2_decap_8 FILLER_50_1024 ();
 sg13g2_decap_8 FILLER_50_1031 ();
 sg13g2_decap_8 FILLER_50_1038 ();
 sg13g2_decap_8 FILLER_50_1045 ();
 sg13g2_decap_8 FILLER_50_1052 ();
 sg13g2_decap_8 FILLER_50_1059 ();
 sg13g2_decap_8 FILLER_50_1066 ();
 sg13g2_decap_8 FILLER_50_1073 ();
 sg13g2_decap_8 FILLER_50_1080 ();
 sg13g2_decap_8 FILLER_50_1087 ();
 sg13g2_decap_8 FILLER_50_1094 ();
 sg13g2_decap_8 FILLER_50_1101 ();
 sg13g2_decap_8 FILLER_50_1108 ();
 sg13g2_decap_8 FILLER_50_1115 ();
 sg13g2_decap_8 FILLER_50_1122 ();
 sg13g2_decap_8 FILLER_50_1129 ();
 sg13g2_decap_8 FILLER_50_1136 ();
 sg13g2_decap_8 FILLER_50_1143 ();
 sg13g2_decap_8 FILLER_50_1150 ();
 sg13g2_decap_8 FILLER_50_1157 ();
 sg13g2_decap_8 FILLER_50_1164 ();
 sg13g2_decap_8 FILLER_50_1171 ();
 sg13g2_decap_8 FILLER_50_1178 ();
 sg13g2_decap_8 FILLER_50_1185 ();
 sg13g2_decap_8 FILLER_50_1192 ();
 sg13g2_decap_8 FILLER_50_1199 ();
 sg13g2_decap_8 FILLER_50_1206 ();
 sg13g2_decap_8 FILLER_50_1213 ();
 sg13g2_decap_8 FILLER_50_1220 ();
 sg13g2_decap_8 FILLER_50_1227 ();
 sg13g2_decap_8 FILLER_50_1234 ();
 sg13g2_decap_8 FILLER_50_1241 ();
 sg13g2_decap_8 FILLER_50_1248 ();
 sg13g2_decap_8 FILLER_50_1255 ();
 sg13g2_decap_8 FILLER_50_1262 ();
 sg13g2_decap_8 FILLER_50_1269 ();
 sg13g2_decap_8 FILLER_50_1276 ();
 sg13g2_decap_8 FILLER_50_1283 ();
 sg13g2_decap_8 FILLER_50_1290 ();
 sg13g2_decap_8 FILLER_50_1297 ();
 sg13g2_decap_8 FILLER_50_1304 ();
 sg13g2_decap_8 FILLER_50_1311 ();
 sg13g2_decap_8 FILLER_50_1318 ();
 sg13g2_fill_1 FILLER_50_1325 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_139 ();
 sg13g2_fill_1 FILLER_51_185 ();
 sg13g2_fill_1 FILLER_51_200 ();
 sg13g2_fill_1 FILLER_51_206 ();
 sg13g2_fill_1 FILLER_51_216 ();
 sg13g2_fill_2 FILLER_51_221 ();
 sg13g2_fill_2 FILLER_51_227 ();
 sg13g2_fill_2 FILLER_51_242 ();
 sg13g2_fill_2 FILLER_51_257 ();
 sg13g2_fill_2 FILLER_51_282 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_fill_1 FILLER_51_306 ();
 sg13g2_fill_2 FILLER_51_423 ();
 sg13g2_fill_1 FILLER_51_425 ();
 sg13g2_fill_1 FILLER_51_435 ();
 sg13g2_fill_2 FILLER_51_448 ();
 sg13g2_fill_1 FILLER_51_450 ();
 sg13g2_fill_1 FILLER_51_485 ();
 sg13g2_fill_2 FILLER_51_496 ();
 sg13g2_fill_2 FILLER_51_550 ();
 sg13g2_fill_1 FILLER_51_565 ();
 sg13g2_fill_2 FILLER_51_596 ();
 sg13g2_fill_2 FILLER_51_602 ();
 sg13g2_fill_2 FILLER_51_608 ();
 sg13g2_fill_1 FILLER_51_619 ();
 sg13g2_fill_2 FILLER_51_656 ();
 sg13g2_fill_2 FILLER_51_677 ();
 sg13g2_fill_1 FILLER_51_684 ();
 sg13g2_decap_4 FILLER_51_703 ();
 sg13g2_fill_1 FILLER_51_869 ();
 sg13g2_fill_2 FILLER_51_942 ();
 sg13g2_decap_8 FILLER_51_984 ();
 sg13g2_decap_8 FILLER_51_991 ();
 sg13g2_decap_8 FILLER_51_998 ();
 sg13g2_decap_8 FILLER_51_1005 ();
 sg13g2_decap_8 FILLER_51_1012 ();
 sg13g2_decap_8 FILLER_51_1019 ();
 sg13g2_decap_8 FILLER_51_1026 ();
 sg13g2_decap_8 FILLER_51_1033 ();
 sg13g2_decap_8 FILLER_51_1040 ();
 sg13g2_decap_8 FILLER_51_1047 ();
 sg13g2_decap_8 FILLER_51_1054 ();
 sg13g2_decap_8 FILLER_51_1061 ();
 sg13g2_decap_8 FILLER_51_1068 ();
 sg13g2_decap_8 FILLER_51_1075 ();
 sg13g2_decap_8 FILLER_51_1082 ();
 sg13g2_decap_8 FILLER_51_1089 ();
 sg13g2_decap_8 FILLER_51_1096 ();
 sg13g2_decap_8 FILLER_51_1103 ();
 sg13g2_decap_8 FILLER_51_1110 ();
 sg13g2_decap_8 FILLER_51_1117 ();
 sg13g2_decap_8 FILLER_51_1124 ();
 sg13g2_decap_8 FILLER_51_1131 ();
 sg13g2_decap_8 FILLER_51_1138 ();
 sg13g2_decap_8 FILLER_51_1145 ();
 sg13g2_decap_8 FILLER_51_1152 ();
 sg13g2_decap_8 FILLER_51_1159 ();
 sg13g2_decap_8 FILLER_51_1166 ();
 sg13g2_decap_8 FILLER_51_1173 ();
 sg13g2_decap_8 FILLER_51_1180 ();
 sg13g2_decap_8 FILLER_51_1187 ();
 sg13g2_decap_8 FILLER_51_1194 ();
 sg13g2_decap_8 FILLER_51_1201 ();
 sg13g2_decap_8 FILLER_51_1208 ();
 sg13g2_decap_8 FILLER_51_1215 ();
 sg13g2_decap_8 FILLER_51_1222 ();
 sg13g2_decap_8 FILLER_51_1229 ();
 sg13g2_decap_8 FILLER_51_1236 ();
 sg13g2_decap_8 FILLER_51_1243 ();
 sg13g2_decap_8 FILLER_51_1250 ();
 sg13g2_decap_8 FILLER_51_1257 ();
 sg13g2_decap_8 FILLER_51_1264 ();
 sg13g2_decap_8 FILLER_51_1271 ();
 sg13g2_decap_8 FILLER_51_1278 ();
 sg13g2_decap_8 FILLER_51_1285 ();
 sg13g2_decap_8 FILLER_51_1292 ();
 sg13g2_decap_8 FILLER_51_1299 ();
 sg13g2_decap_8 FILLER_51_1306 ();
 sg13g2_decap_8 FILLER_51_1313 ();
 sg13g2_decap_4 FILLER_51_1320 ();
 sg13g2_fill_2 FILLER_51_1324 ();
 sg13g2_fill_2 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_121 ();
 sg13g2_fill_1 FILLER_52_148 ();
 sg13g2_fill_1 FILLER_52_170 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_fill_1 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_1 FILLER_52_270 ();
 sg13g2_decap_4 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_1 FILLER_52_333 ();
 sg13g2_fill_1 FILLER_52_346 ();
 sg13g2_fill_2 FILLER_52_356 ();
 sg13g2_fill_2 FILLER_52_363 ();
 sg13g2_fill_1 FILLER_52_365 ();
 sg13g2_fill_2 FILLER_52_443 ();
 sg13g2_fill_2 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_497 ();
 sg13g2_fill_1 FILLER_52_534 ();
 sg13g2_fill_2 FILLER_52_592 ();
 sg13g2_fill_1 FILLER_52_599 ();
 sg13g2_fill_2 FILLER_52_606 ();
 sg13g2_fill_1 FILLER_52_612 ();
 sg13g2_fill_1 FILLER_52_639 ();
 sg13g2_fill_1 FILLER_52_692 ();
 sg13g2_fill_2 FILLER_52_776 ();
 sg13g2_fill_2 FILLER_52_788 ();
 sg13g2_fill_1 FILLER_52_934 ();
 sg13g2_fill_1 FILLER_52_945 ();
 sg13g2_fill_1 FILLER_52_982 ();
 sg13g2_decap_8 FILLER_52_987 ();
 sg13g2_decap_8 FILLER_52_994 ();
 sg13g2_decap_8 FILLER_52_1001 ();
 sg13g2_decap_8 FILLER_52_1008 ();
 sg13g2_decap_8 FILLER_52_1015 ();
 sg13g2_decap_8 FILLER_52_1022 ();
 sg13g2_decap_8 FILLER_52_1029 ();
 sg13g2_decap_8 FILLER_52_1036 ();
 sg13g2_decap_8 FILLER_52_1043 ();
 sg13g2_decap_8 FILLER_52_1050 ();
 sg13g2_decap_8 FILLER_52_1057 ();
 sg13g2_decap_8 FILLER_52_1064 ();
 sg13g2_decap_8 FILLER_52_1071 ();
 sg13g2_decap_8 FILLER_52_1078 ();
 sg13g2_decap_8 FILLER_52_1085 ();
 sg13g2_decap_8 FILLER_52_1092 ();
 sg13g2_decap_8 FILLER_52_1099 ();
 sg13g2_decap_8 FILLER_52_1106 ();
 sg13g2_decap_8 FILLER_52_1113 ();
 sg13g2_decap_8 FILLER_52_1120 ();
 sg13g2_decap_8 FILLER_52_1127 ();
 sg13g2_decap_8 FILLER_52_1134 ();
 sg13g2_decap_8 FILLER_52_1141 ();
 sg13g2_decap_8 FILLER_52_1148 ();
 sg13g2_decap_8 FILLER_52_1155 ();
 sg13g2_decap_8 FILLER_52_1162 ();
 sg13g2_decap_8 FILLER_52_1169 ();
 sg13g2_decap_8 FILLER_52_1176 ();
 sg13g2_decap_8 FILLER_52_1183 ();
 sg13g2_decap_8 FILLER_52_1190 ();
 sg13g2_decap_8 FILLER_52_1197 ();
 sg13g2_decap_8 FILLER_52_1204 ();
 sg13g2_decap_8 FILLER_52_1211 ();
 sg13g2_decap_8 FILLER_52_1218 ();
 sg13g2_decap_8 FILLER_52_1225 ();
 sg13g2_decap_8 FILLER_52_1232 ();
 sg13g2_decap_8 FILLER_52_1239 ();
 sg13g2_decap_8 FILLER_52_1246 ();
 sg13g2_decap_8 FILLER_52_1253 ();
 sg13g2_decap_8 FILLER_52_1260 ();
 sg13g2_decap_8 FILLER_52_1267 ();
 sg13g2_decap_8 FILLER_52_1274 ();
 sg13g2_decap_8 FILLER_52_1281 ();
 sg13g2_decap_8 FILLER_52_1288 ();
 sg13g2_decap_8 FILLER_52_1295 ();
 sg13g2_decap_8 FILLER_52_1302 ();
 sg13g2_decap_8 FILLER_52_1309 ();
 sg13g2_decap_8 FILLER_52_1316 ();
 sg13g2_fill_2 FILLER_52_1323 ();
 sg13g2_fill_1 FILLER_52_1325 ();
 sg13g2_fill_2 FILLER_53_124 ();
 sg13g2_fill_1 FILLER_53_144 ();
 sg13g2_fill_1 FILLER_53_173 ();
 sg13g2_fill_2 FILLER_53_184 ();
 sg13g2_fill_2 FILLER_53_195 ();
 sg13g2_fill_1 FILLER_53_216 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_227 ();
 sg13g2_decap_8 FILLER_53_233 ();
 sg13g2_decap_4 FILLER_53_240 ();
 sg13g2_decap_4 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_272 ();
 sg13g2_fill_2 FILLER_53_279 ();
 sg13g2_decap_4 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_295 ();
 sg13g2_fill_1 FILLER_53_319 ();
 sg13g2_fill_1 FILLER_53_337 ();
 sg13g2_fill_2 FILLER_53_364 ();
 sg13g2_fill_2 FILLER_53_370 ();
 sg13g2_fill_1 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_405 ();
 sg13g2_fill_2 FILLER_53_416 ();
 sg13g2_fill_2 FILLER_53_422 ();
 sg13g2_fill_2 FILLER_53_472 ();
 sg13g2_fill_1 FILLER_53_474 ();
 sg13g2_fill_2 FILLER_53_513 ();
 sg13g2_fill_1 FILLER_53_541 ();
 sg13g2_fill_1 FILLER_53_569 ();
 sg13g2_fill_1 FILLER_53_647 ();
 sg13g2_fill_2 FILLER_53_652 ();
 sg13g2_fill_1 FILLER_53_658 ();
 sg13g2_fill_2 FILLER_53_669 ();
 sg13g2_fill_1 FILLER_53_675 ();
 sg13g2_fill_1 FILLER_53_702 ();
 sg13g2_fill_1 FILLER_53_708 ();
 sg13g2_fill_2 FILLER_53_713 ();
 sg13g2_fill_1 FILLER_53_719 ();
 sg13g2_fill_1 FILLER_53_746 ();
 sg13g2_fill_2 FILLER_53_751 ();
 sg13g2_fill_2 FILLER_53_763 ();
 sg13g2_fill_2 FILLER_53_791 ();
 sg13g2_fill_2 FILLER_53_859 ();
 sg13g2_fill_1 FILLER_53_961 ();
 sg13g2_decap_8 FILLER_53_988 ();
 sg13g2_decap_8 FILLER_53_995 ();
 sg13g2_decap_8 FILLER_53_1002 ();
 sg13g2_decap_8 FILLER_53_1009 ();
 sg13g2_decap_8 FILLER_53_1016 ();
 sg13g2_decap_8 FILLER_53_1023 ();
 sg13g2_decap_8 FILLER_53_1030 ();
 sg13g2_decap_8 FILLER_53_1037 ();
 sg13g2_decap_8 FILLER_53_1044 ();
 sg13g2_decap_8 FILLER_53_1051 ();
 sg13g2_decap_8 FILLER_53_1058 ();
 sg13g2_decap_8 FILLER_53_1065 ();
 sg13g2_decap_8 FILLER_53_1072 ();
 sg13g2_decap_8 FILLER_53_1079 ();
 sg13g2_decap_8 FILLER_53_1086 ();
 sg13g2_decap_8 FILLER_53_1093 ();
 sg13g2_decap_8 FILLER_53_1100 ();
 sg13g2_decap_8 FILLER_53_1107 ();
 sg13g2_decap_8 FILLER_53_1114 ();
 sg13g2_decap_8 FILLER_53_1121 ();
 sg13g2_decap_8 FILLER_53_1128 ();
 sg13g2_decap_8 FILLER_53_1135 ();
 sg13g2_decap_8 FILLER_53_1142 ();
 sg13g2_decap_8 FILLER_53_1149 ();
 sg13g2_decap_8 FILLER_53_1156 ();
 sg13g2_decap_8 FILLER_53_1163 ();
 sg13g2_decap_8 FILLER_53_1170 ();
 sg13g2_decap_8 FILLER_53_1177 ();
 sg13g2_decap_8 FILLER_53_1184 ();
 sg13g2_decap_8 FILLER_53_1191 ();
 sg13g2_decap_8 FILLER_53_1198 ();
 sg13g2_decap_8 FILLER_53_1205 ();
 sg13g2_decap_8 FILLER_53_1212 ();
 sg13g2_decap_8 FILLER_53_1219 ();
 sg13g2_decap_8 FILLER_53_1226 ();
 sg13g2_decap_8 FILLER_53_1233 ();
 sg13g2_decap_8 FILLER_53_1240 ();
 sg13g2_decap_8 FILLER_53_1247 ();
 sg13g2_decap_8 FILLER_53_1254 ();
 sg13g2_decap_8 FILLER_53_1261 ();
 sg13g2_decap_8 FILLER_53_1268 ();
 sg13g2_decap_8 FILLER_53_1275 ();
 sg13g2_decap_8 FILLER_53_1282 ();
 sg13g2_decap_8 FILLER_53_1289 ();
 sg13g2_decap_8 FILLER_53_1296 ();
 sg13g2_decap_8 FILLER_53_1303 ();
 sg13g2_decap_8 FILLER_53_1310 ();
 sg13g2_decap_8 FILLER_53_1317 ();
 sg13g2_fill_2 FILLER_53_1324 ();
 sg13g2_fill_1 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_fill_2 FILLER_54_109 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_fill_2 FILLER_54_138 ();
 sg13g2_fill_2 FILLER_54_196 ();
 sg13g2_decap_4 FILLER_54_218 ();
 sg13g2_fill_2 FILLER_54_291 ();
 sg13g2_fill_1 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_298 ();
 sg13g2_fill_1 FILLER_54_304 ();
 sg13g2_fill_2 FILLER_54_310 ();
 sg13g2_fill_1 FILLER_54_318 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_fill_1 FILLER_54_335 ();
 sg13g2_fill_1 FILLER_54_414 ();
 sg13g2_fill_2 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_427 ();
 sg13g2_fill_1 FILLER_54_510 ();
 sg13g2_fill_1 FILLER_54_541 ();
 sg13g2_fill_2 FILLER_54_577 ();
 sg13g2_fill_1 FILLER_54_579 ();
 sg13g2_fill_1 FILLER_54_606 ();
 sg13g2_fill_1 FILLER_54_617 ();
 sg13g2_fill_1 FILLER_54_623 ();
 sg13g2_fill_2 FILLER_54_704 ();
 sg13g2_fill_1 FILLER_54_710 ();
 sg13g2_fill_1 FILLER_54_721 ();
 sg13g2_fill_1 FILLER_54_758 ();
 sg13g2_fill_2 FILLER_54_769 ();
 sg13g2_fill_2 FILLER_54_807 ();
 sg13g2_fill_1 FILLER_54_809 ();
 sg13g2_fill_2 FILLER_54_947 ();
 sg13g2_fill_1 FILLER_54_959 ();
 sg13g2_decap_8 FILLER_54_982 ();
 sg13g2_decap_8 FILLER_54_989 ();
 sg13g2_decap_8 FILLER_54_996 ();
 sg13g2_decap_8 FILLER_54_1003 ();
 sg13g2_decap_8 FILLER_54_1010 ();
 sg13g2_decap_8 FILLER_54_1017 ();
 sg13g2_decap_8 FILLER_54_1024 ();
 sg13g2_decap_8 FILLER_54_1031 ();
 sg13g2_decap_8 FILLER_54_1038 ();
 sg13g2_decap_8 FILLER_54_1045 ();
 sg13g2_decap_8 FILLER_54_1052 ();
 sg13g2_decap_8 FILLER_54_1059 ();
 sg13g2_decap_8 FILLER_54_1066 ();
 sg13g2_decap_8 FILLER_54_1073 ();
 sg13g2_decap_8 FILLER_54_1080 ();
 sg13g2_decap_8 FILLER_54_1087 ();
 sg13g2_decap_8 FILLER_54_1094 ();
 sg13g2_decap_8 FILLER_54_1101 ();
 sg13g2_decap_8 FILLER_54_1108 ();
 sg13g2_decap_8 FILLER_54_1115 ();
 sg13g2_decap_8 FILLER_54_1122 ();
 sg13g2_decap_8 FILLER_54_1129 ();
 sg13g2_decap_8 FILLER_54_1136 ();
 sg13g2_decap_8 FILLER_54_1143 ();
 sg13g2_decap_8 FILLER_54_1150 ();
 sg13g2_decap_8 FILLER_54_1157 ();
 sg13g2_decap_8 FILLER_54_1164 ();
 sg13g2_decap_8 FILLER_54_1171 ();
 sg13g2_decap_8 FILLER_54_1178 ();
 sg13g2_decap_8 FILLER_54_1185 ();
 sg13g2_decap_8 FILLER_54_1192 ();
 sg13g2_decap_8 FILLER_54_1199 ();
 sg13g2_decap_8 FILLER_54_1206 ();
 sg13g2_decap_8 FILLER_54_1213 ();
 sg13g2_decap_8 FILLER_54_1220 ();
 sg13g2_decap_8 FILLER_54_1227 ();
 sg13g2_decap_8 FILLER_54_1234 ();
 sg13g2_decap_8 FILLER_54_1241 ();
 sg13g2_decap_8 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1255 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_decap_8 FILLER_54_1269 ();
 sg13g2_decap_8 FILLER_54_1276 ();
 sg13g2_decap_8 FILLER_54_1283 ();
 sg13g2_decap_8 FILLER_54_1290 ();
 sg13g2_decap_8 FILLER_54_1297 ();
 sg13g2_decap_8 FILLER_54_1304 ();
 sg13g2_decap_8 FILLER_54_1311 ();
 sg13g2_decap_8 FILLER_54_1318 ();
 sg13g2_fill_1 FILLER_54_1325 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_52 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_124 ();
 sg13g2_fill_2 FILLER_55_171 ();
 sg13g2_fill_1 FILLER_55_173 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_fill_1 FILLER_55_212 ();
 sg13g2_fill_2 FILLER_55_218 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_decap_4 FILLER_55_292 ();
 sg13g2_fill_1 FILLER_55_312 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_365 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_fill_2 FILLER_55_390 ();
 sg13g2_fill_1 FILLER_55_405 ();
 sg13g2_fill_1 FILLER_55_450 ();
 sg13g2_fill_2 FILLER_55_507 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_fill_1 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_652 ();
 sg13g2_fill_1 FILLER_55_679 ();
 sg13g2_fill_1 FILLER_55_684 ();
 sg13g2_fill_1 FILLER_55_689 ();
 sg13g2_fill_2 FILLER_55_818 ();
 sg13g2_fill_1 FILLER_55_820 ();
 sg13g2_fill_2 FILLER_55_925 ();
 sg13g2_fill_1 FILLER_55_937 ();
 sg13g2_fill_1 FILLER_55_948 ();
 sg13g2_decap_8 FILLER_55_983 ();
 sg13g2_decap_8 FILLER_55_990 ();
 sg13g2_decap_8 FILLER_55_997 ();
 sg13g2_decap_8 FILLER_55_1004 ();
 sg13g2_decap_8 FILLER_55_1011 ();
 sg13g2_decap_8 FILLER_55_1018 ();
 sg13g2_decap_8 FILLER_55_1025 ();
 sg13g2_decap_8 FILLER_55_1032 ();
 sg13g2_decap_8 FILLER_55_1039 ();
 sg13g2_decap_8 FILLER_55_1046 ();
 sg13g2_decap_8 FILLER_55_1053 ();
 sg13g2_decap_8 FILLER_55_1060 ();
 sg13g2_decap_8 FILLER_55_1067 ();
 sg13g2_decap_8 FILLER_55_1074 ();
 sg13g2_decap_8 FILLER_55_1081 ();
 sg13g2_decap_8 FILLER_55_1088 ();
 sg13g2_decap_8 FILLER_55_1095 ();
 sg13g2_decap_8 FILLER_55_1102 ();
 sg13g2_decap_8 FILLER_55_1109 ();
 sg13g2_decap_8 FILLER_55_1116 ();
 sg13g2_decap_8 FILLER_55_1123 ();
 sg13g2_decap_8 FILLER_55_1130 ();
 sg13g2_decap_8 FILLER_55_1137 ();
 sg13g2_decap_8 FILLER_55_1144 ();
 sg13g2_decap_8 FILLER_55_1151 ();
 sg13g2_decap_8 FILLER_55_1158 ();
 sg13g2_decap_8 FILLER_55_1165 ();
 sg13g2_decap_8 FILLER_55_1172 ();
 sg13g2_decap_8 FILLER_55_1179 ();
 sg13g2_decap_8 FILLER_55_1186 ();
 sg13g2_decap_8 FILLER_55_1193 ();
 sg13g2_decap_8 FILLER_55_1200 ();
 sg13g2_decap_8 FILLER_55_1207 ();
 sg13g2_decap_8 FILLER_55_1214 ();
 sg13g2_decap_8 FILLER_55_1221 ();
 sg13g2_decap_8 FILLER_55_1228 ();
 sg13g2_decap_8 FILLER_55_1235 ();
 sg13g2_decap_8 FILLER_55_1242 ();
 sg13g2_decap_8 FILLER_55_1249 ();
 sg13g2_decap_8 FILLER_55_1256 ();
 sg13g2_decap_8 FILLER_55_1263 ();
 sg13g2_decap_8 FILLER_55_1270 ();
 sg13g2_decap_8 FILLER_55_1277 ();
 sg13g2_decap_8 FILLER_55_1284 ();
 sg13g2_decap_8 FILLER_55_1291 ();
 sg13g2_decap_8 FILLER_55_1298 ();
 sg13g2_decap_8 FILLER_55_1305 ();
 sg13g2_decap_8 FILLER_55_1312 ();
 sg13g2_decap_8 FILLER_55_1319 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_2 ();
 sg13g2_fill_1 FILLER_56_75 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_129 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_205 ();
 sg13g2_fill_1 FILLER_56_226 ();
 sg13g2_fill_1 FILLER_56_261 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_1 FILLER_56_279 ();
 sg13g2_fill_2 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_352 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_fill_2 FILLER_56_430 ();
 sg13g2_fill_2 FILLER_56_488 ();
 sg13g2_fill_1 FILLER_56_490 ();
 sg13g2_fill_2 FILLER_56_495 ();
 sg13g2_fill_2 FILLER_56_505 ();
 sg13g2_fill_1 FILLER_56_507 ();
 sg13g2_fill_1 FILLER_56_564 ();
 sg13g2_fill_1 FILLER_56_611 ();
 sg13g2_fill_1 FILLER_56_664 ();
 sg13g2_fill_1 FILLER_56_691 ();
 sg13g2_fill_1 FILLER_56_718 ();
 sg13g2_fill_1 FILLER_56_729 ();
 sg13g2_fill_2 FILLER_56_734 ();
 sg13g2_fill_2 FILLER_56_766 ();
 sg13g2_fill_2 FILLER_56_802 ();
 sg13g2_fill_1 FILLER_56_804 ();
 sg13g2_fill_1 FILLER_56_831 ();
 sg13g2_fill_1 FILLER_56_896 ();
 sg13g2_decap_8 FILLER_56_985 ();
 sg13g2_decap_8 FILLER_56_992 ();
 sg13g2_decap_8 FILLER_56_999 ();
 sg13g2_decap_8 FILLER_56_1006 ();
 sg13g2_decap_8 FILLER_56_1013 ();
 sg13g2_decap_8 FILLER_56_1020 ();
 sg13g2_decap_8 FILLER_56_1027 ();
 sg13g2_decap_8 FILLER_56_1034 ();
 sg13g2_decap_8 FILLER_56_1041 ();
 sg13g2_decap_8 FILLER_56_1048 ();
 sg13g2_decap_8 FILLER_56_1055 ();
 sg13g2_decap_8 FILLER_56_1062 ();
 sg13g2_decap_8 FILLER_56_1069 ();
 sg13g2_decap_8 FILLER_56_1076 ();
 sg13g2_decap_8 FILLER_56_1083 ();
 sg13g2_decap_8 FILLER_56_1090 ();
 sg13g2_decap_8 FILLER_56_1097 ();
 sg13g2_decap_8 FILLER_56_1104 ();
 sg13g2_decap_8 FILLER_56_1111 ();
 sg13g2_decap_8 FILLER_56_1118 ();
 sg13g2_decap_8 FILLER_56_1125 ();
 sg13g2_decap_8 FILLER_56_1132 ();
 sg13g2_decap_8 FILLER_56_1139 ();
 sg13g2_decap_8 FILLER_56_1146 ();
 sg13g2_decap_8 FILLER_56_1153 ();
 sg13g2_decap_8 FILLER_56_1160 ();
 sg13g2_decap_8 FILLER_56_1167 ();
 sg13g2_decap_8 FILLER_56_1174 ();
 sg13g2_decap_8 FILLER_56_1181 ();
 sg13g2_decap_8 FILLER_56_1188 ();
 sg13g2_decap_8 FILLER_56_1195 ();
 sg13g2_decap_8 FILLER_56_1202 ();
 sg13g2_decap_8 FILLER_56_1209 ();
 sg13g2_decap_8 FILLER_56_1216 ();
 sg13g2_decap_8 FILLER_56_1223 ();
 sg13g2_decap_8 FILLER_56_1230 ();
 sg13g2_decap_8 FILLER_56_1237 ();
 sg13g2_decap_8 FILLER_56_1244 ();
 sg13g2_decap_8 FILLER_56_1251 ();
 sg13g2_decap_8 FILLER_56_1258 ();
 sg13g2_decap_8 FILLER_56_1265 ();
 sg13g2_decap_8 FILLER_56_1272 ();
 sg13g2_decap_8 FILLER_56_1279 ();
 sg13g2_decap_8 FILLER_56_1286 ();
 sg13g2_decap_8 FILLER_56_1293 ();
 sg13g2_decap_8 FILLER_56_1300 ();
 sg13g2_decap_8 FILLER_56_1307 ();
 sg13g2_decap_8 FILLER_56_1314 ();
 sg13g2_decap_4 FILLER_56_1321 ();
 sg13g2_fill_1 FILLER_56_1325 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_27 ();
 sg13g2_fill_1 FILLER_57_33 ();
 sg13g2_fill_1 FILLER_57_40 ();
 sg13g2_fill_1 FILLER_57_46 ();
 sg13g2_fill_1 FILLER_57_52 ();
 sg13g2_fill_1 FILLER_57_59 ();
 sg13g2_fill_2 FILLER_57_69 ();
 sg13g2_fill_2 FILLER_57_83 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_128 ();
 sg13g2_fill_1 FILLER_57_149 ();
 sg13g2_fill_2 FILLER_57_160 ();
 sg13g2_fill_1 FILLER_57_162 ();
 sg13g2_fill_2 FILLER_57_167 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_fill_2 FILLER_57_178 ();
 sg13g2_fill_2 FILLER_57_271 ();
 sg13g2_fill_1 FILLER_57_281 ();
 sg13g2_fill_1 FILLER_57_295 ();
 sg13g2_fill_1 FILLER_57_336 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_364 ();
 sg13g2_fill_1 FILLER_57_392 ();
 sg13g2_fill_2 FILLER_57_450 ();
 sg13g2_fill_1 FILLER_57_452 ();
 sg13g2_fill_2 FILLER_57_585 ();
 sg13g2_fill_1 FILLER_57_623 ();
 sg13g2_fill_1 FILLER_57_634 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_fill_1 FILLER_57_700 ();
 sg13g2_fill_1 FILLER_57_735 ();
 sg13g2_fill_1 FILLER_57_780 ();
 sg13g2_fill_1 FILLER_57_872 ();
 sg13g2_fill_2 FILLER_57_925 ();
 sg13g2_fill_1 FILLER_57_949 ();
 sg13g2_fill_2 FILLER_57_960 ();
 sg13g2_fill_1 FILLER_57_962 ();
 sg13g2_decap_8 FILLER_57_971 ();
 sg13g2_decap_8 FILLER_57_978 ();
 sg13g2_decap_8 FILLER_57_985 ();
 sg13g2_decap_8 FILLER_57_992 ();
 sg13g2_decap_8 FILLER_57_999 ();
 sg13g2_decap_8 FILLER_57_1006 ();
 sg13g2_decap_8 FILLER_57_1013 ();
 sg13g2_decap_8 FILLER_57_1020 ();
 sg13g2_decap_8 FILLER_57_1027 ();
 sg13g2_decap_8 FILLER_57_1034 ();
 sg13g2_decap_8 FILLER_57_1041 ();
 sg13g2_decap_8 FILLER_57_1048 ();
 sg13g2_decap_8 FILLER_57_1055 ();
 sg13g2_decap_8 FILLER_57_1062 ();
 sg13g2_decap_8 FILLER_57_1069 ();
 sg13g2_decap_8 FILLER_57_1076 ();
 sg13g2_decap_8 FILLER_57_1083 ();
 sg13g2_decap_8 FILLER_57_1090 ();
 sg13g2_decap_8 FILLER_57_1097 ();
 sg13g2_decap_8 FILLER_57_1104 ();
 sg13g2_decap_8 FILLER_57_1111 ();
 sg13g2_decap_8 FILLER_57_1118 ();
 sg13g2_decap_8 FILLER_57_1125 ();
 sg13g2_decap_8 FILLER_57_1132 ();
 sg13g2_decap_8 FILLER_57_1139 ();
 sg13g2_decap_8 FILLER_57_1146 ();
 sg13g2_decap_8 FILLER_57_1153 ();
 sg13g2_decap_8 FILLER_57_1160 ();
 sg13g2_decap_8 FILLER_57_1167 ();
 sg13g2_decap_8 FILLER_57_1174 ();
 sg13g2_decap_8 FILLER_57_1181 ();
 sg13g2_decap_8 FILLER_57_1188 ();
 sg13g2_decap_8 FILLER_57_1195 ();
 sg13g2_decap_8 FILLER_57_1202 ();
 sg13g2_decap_8 FILLER_57_1209 ();
 sg13g2_decap_8 FILLER_57_1216 ();
 sg13g2_decap_8 FILLER_57_1223 ();
 sg13g2_decap_8 FILLER_57_1230 ();
 sg13g2_decap_8 FILLER_57_1237 ();
 sg13g2_decap_8 FILLER_57_1244 ();
 sg13g2_decap_8 FILLER_57_1251 ();
 sg13g2_decap_8 FILLER_57_1258 ();
 sg13g2_decap_8 FILLER_57_1265 ();
 sg13g2_decap_8 FILLER_57_1272 ();
 sg13g2_decap_8 FILLER_57_1279 ();
 sg13g2_decap_8 FILLER_57_1286 ();
 sg13g2_decap_8 FILLER_57_1293 ();
 sg13g2_decap_8 FILLER_57_1300 ();
 sg13g2_decap_8 FILLER_57_1307 ();
 sg13g2_decap_8 FILLER_57_1314 ();
 sg13g2_decap_4 FILLER_57_1321 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_94 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_151 ();
 sg13g2_fill_2 FILLER_58_177 ();
 sg13g2_fill_1 FILLER_58_204 ();
 sg13g2_fill_1 FILLER_58_237 ();
 sg13g2_fill_1 FILLER_58_246 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_256 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_299 ();
 sg13g2_fill_2 FILLER_58_333 ();
 sg13g2_fill_1 FILLER_58_344 ();
 sg13g2_fill_1 FILLER_58_378 ();
 sg13g2_fill_2 FILLER_58_420 ();
 sg13g2_fill_2 FILLER_58_448 ();
 sg13g2_fill_1 FILLER_58_450 ();
 sg13g2_fill_2 FILLER_58_491 ();
 sg13g2_fill_2 FILLER_58_539 ();
 sg13g2_fill_1 FILLER_58_571 ();
 sg13g2_fill_1 FILLER_58_602 ();
 sg13g2_fill_1 FILLER_58_629 ();
 sg13g2_fill_1 FILLER_58_660 ();
 sg13g2_fill_1 FILLER_58_687 ();
 sg13g2_fill_2 FILLER_58_853 ();
 sg13g2_decap_8 FILLER_58_931 ();
 sg13g2_decap_4 FILLER_58_938 ();
 sg13g2_decap_8 FILLER_58_972 ();
 sg13g2_decap_8 FILLER_58_979 ();
 sg13g2_decap_8 FILLER_58_986 ();
 sg13g2_decap_8 FILLER_58_993 ();
 sg13g2_decap_8 FILLER_58_1000 ();
 sg13g2_decap_8 FILLER_58_1007 ();
 sg13g2_decap_8 FILLER_58_1014 ();
 sg13g2_decap_8 FILLER_58_1021 ();
 sg13g2_decap_8 FILLER_58_1028 ();
 sg13g2_decap_8 FILLER_58_1035 ();
 sg13g2_decap_8 FILLER_58_1042 ();
 sg13g2_decap_8 FILLER_58_1049 ();
 sg13g2_decap_8 FILLER_58_1056 ();
 sg13g2_decap_8 FILLER_58_1063 ();
 sg13g2_decap_8 FILLER_58_1070 ();
 sg13g2_decap_8 FILLER_58_1077 ();
 sg13g2_decap_8 FILLER_58_1084 ();
 sg13g2_decap_8 FILLER_58_1091 ();
 sg13g2_decap_8 FILLER_58_1098 ();
 sg13g2_decap_8 FILLER_58_1105 ();
 sg13g2_decap_8 FILLER_58_1112 ();
 sg13g2_decap_8 FILLER_58_1119 ();
 sg13g2_decap_8 FILLER_58_1126 ();
 sg13g2_decap_8 FILLER_58_1133 ();
 sg13g2_decap_8 FILLER_58_1140 ();
 sg13g2_decap_8 FILLER_58_1147 ();
 sg13g2_decap_8 FILLER_58_1154 ();
 sg13g2_decap_8 FILLER_58_1161 ();
 sg13g2_decap_8 FILLER_58_1168 ();
 sg13g2_decap_8 FILLER_58_1175 ();
 sg13g2_decap_8 FILLER_58_1182 ();
 sg13g2_decap_8 FILLER_58_1189 ();
 sg13g2_decap_8 FILLER_58_1196 ();
 sg13g2_decap_8 FILLER_58_1203 ();
 sg13g2_decap_8 FILLER_58_1210 ();
 sg13g2_decap_8 FILLER_58_1217 ();
 sg13g2_decap_8 FILLER_58_1224 ();
 sg13g2_decap_8 FILLER_58_1231 ();
 sg13g2_decap_8 FILLER_58_1238 ();
 sg13g2_decap_8 FILLER_58_1245 ();
 sg13g2_decap_8 FILLER_58_1252 ();
 sg13g2_decap_8 FILLER_58_1259 ();
 sg13g2_decap_8 FILLER_58_1266 ();
 sg13g2_decap_8 FILLER_58_1273 ();
 sg13g2_decap_8 FILLER_58_1280 ();
 sg13g2_decap_8 FILLER_58_1287 ();
 sg13g2_decap_8 FILLER_58_1294 ();
 sg13g2_decap_8 FILLER_58_1301 ();
 sg13g2_decap_8 FILLER_58_1308 ();
 sg13g2_decap_8 FILLER_58_1315 ();
 sg13g2_decap_4 FILLER_58_1322 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_116 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_161 ();
 sg13g2_fill_1 FILLER_59_193 ();
 sg13g2_fill_2 FILLER_59_228 ();
 sg13g2_fill_2 FILLER_59_238 ();
 sg13g2_fill_2 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_383 ();
 sg13g2_fill_2 FILLER_59_389 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_fill_2 FILLER_59_459 ();
 sg13g2_fill_1 FILLER_59_532 ();
 sg13g2_fill_1 FILLER_59_665 ();
 sg13g2_fill_2 FILLER_59_728 ();
 sg13g2_fill_1 FILLER_59_730 ();
 sg13g2_fill_2 FILLER_59_765 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_1 FILLER_59_871 ();
 sg13g2_decap_8 FILLER_59_920 ();
 sg13g2_decap_8 FILLER_59_927 ();
 sg13g2_decap_8 FILLER_59_934 ();
 sg13g2_decap_8 FILLER_59_941 ();
 sg13g2_decap_8 FILLER_59_948 ();
 sg13g2_decap_8 FILLER_59_955 ();
 sg13g2_decap_8 FILLER_59_962 ();
 sg13g2_decap_8 FILLER_59_969 ();
 sg13g2_decap_8 FILLER_59_976 ();
 sg13g2_decap_8 FILLER_59_983 ();
 sg13g2_decap_8 FILLER_59_990 ();
 sg13g2_decap_8 FILLER_59_997 ();
 sg13g2_decap_8 FILLER_59_1004 ();
 sg13g2_decap_8 FILLER_59_1011 ();
 sg13g2_decap_8 FILLER_59_1018 ();
 sg13g2_decap_8 FILLER_59_1025 ();
 sg13g2_decap_8 FILLER_59_1032 ();
 sg13g2_decap_8 FILLER_59_1039 ();
 sg13g2_decap_8 FILLER_59_1046 ();
 sg13g2_decap_8 FILLER_59_1053 ();
 sg13g2_decap_8 FILLER_59_1060 ();
 sg13g2_decap_8 FILLER_59_1067 ();
 sg13g2_decap_8 FILLER_59_1074 ();
 sg13g2_decap_8 FILLER_59_1081 ();
 sg13g2_decap_8 FILLER_59_1088 ();
 sg13g2_decap_8 FILLER_59_1095 ();
 sg13g2_decap_8 FILLER_59_1102 ();
 sg13g2_decap_8 FILLER_59_1109 ();
 sg13g2_decap_8 FILLER_59_1116 ();
 sg13g2_decap_8 FILLER_59_1123 ();
 sg13g2_decap_8 FILLER_59_1130 ();
 sg13g2_decap_8 FILLER_59_1137 ();
 sg13g2_decap_8 FILLER_59_1144 ();
 sg13g2_decap_8 FILLER_59_1151 ();
 sg13g2_decap_8 FILLER_59_1158 ();
 sg13g2_decap_8 FILLER_59_1165 ();
 sg13g2_decap_8 FILLER_59_1172 ();
 sg13g2_decap_8 FILLER_59_1179 ();
 sg13g2_decap_8 FILLER_59_1186 ();
 sg13g2_decap_8 FILLER_59_1193 ();
 sg13g2_decap_8 FILLER_59_1200 ();
 sg13g2_decap_8 FILLER_59_1207 ();
 sg13g2_decap_8 FILLER_59_1214 ();
 sg13g2_decap_8 FILLER_59_1221 ();
 sg13g2_decap_8 FILLER_59_1228 ();
 sg13g2_decap_8 FILLER_59_1235 ();
 sg13g2_decap_8 FILLER_59_1242 ();
 sg13g2_decap_8 FILLER_59_1249 ();
 sg13g2_decap_8 FILLER_59_1256 ();
 sg13g2_decap_8 FILLER_59_1263 ();
 sg13g2_decap_8 FILLER_59_1270 ();
 sg13g2_decap_8 FILLER_59_1277 ();
 sg13g2_decap_8 FILLER_59_1284 ();
 sg13g2_decap_8 FILLER_59_1291 ();
 sg13g2_decap_8 FILLER_59_1298 ();
 sg13g2_decap_8 FILLER_59_1305 ();
 sg13g2_decap_8 FILLER_59_1312 ();
 sg13g2_decap_8 FILLER_59_1319 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_1 FILLER_60_6 ();
 sg13g2_fill_1 FILLER_60_21 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_2 FILLER_60_81 ();
 sg13g2_fill_2 FILLER_60_94 ();
 sg13g2_fill_1 FILLER_60_127 ();
 sg13g2_fill_1 FILLER_60_136 ();
 sg13g2_fill_2 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_149 ();
 sg13g2_fill_1 FILLER_60_160 ();
 sg13g2_fill_2 FILLER_60_232 ();
 sg13g2_fill_2 FILLER_60_291 ();
 sg13g2_fill_2 FILLER_60_301 ();
 sg13g2_fill_2 FILLER_60_311 ();
 sg13g2_fill_1 FILLER_60_325 ();
 sg13g2_fill_1 FILLER_60_332 ();
 sg13g2_fill_1 FILLER_60_461 ();
 sg13g2_fill_2 FILLER_60_472 ();
 sg13g2_fill_2 FILLER_60_580 ();
 sg13g2_fill_1 FILLER_60_640 ();
 sg13g2_fill_1 FILLER_60_675 ();
 sg13g2_fill_2 FILLER_60_723 ();
 sg13g2_fill_1 FILLER_60_847 ();
 sg13g2_decap_8 FILLER_60_908 ();
 sg13g2_decap_8 FILLER_60_915 ();
 sg13g2_decap_8 FILLER_60_922 ();
 sg13g2_decap_8 FILLER_60_929 ();
 sg13g2_decap_8 FILLER_60_936 ();
 sg13g2_decap_8 FILLER_60_943 ();
 sg13g2_decap_8 FILLER_60_950 ();
 sg13g2_decap_8 FILLER_60_957 ();
 sg13g2_decap_8 FILLER_60_964 ();
 sg13g2_decap_8 FILLER_60_971 ();
 sg13g2_decap_8 FILLER_60_978 ();
 sg13g2_decap_8 FILLER_60_985 ();
 sg13g2_decap_8 FILLER_60_992 ();
 sg13g2_decap_8 FILLER_60_999 ();
 sg13g2_decap_8 FILLER_60_1006 ();
 sg13g2_decap_8 FILLER_60_1013 ();
 sg13g2_decap_8 FILLER_60_1020 ();
 sg13g2_decap_8 FILLER_60_1027 ();
 sg13g2_decap_8 FILLER_60_1034 ();
 sg13g2_decap_8 FILLER_60_1041 ();
 sg13g2_decap_8 FILLER_60_1048 ();
 sg13g2_decap_8 FILLER_60_1055 ();
 sg13g2_decap_8 FILLER_60_1062 ();
 sg13g2_decap_8 FILLER_60_1069 ();
 sg13g2_decap_8 FILLER_60_1076 ();
 sg13g2_decap_8 FILLER_60_1083 ();
 sg13g2_decap_8 FILLER_60_1090 ();
 sg13g2_decap_8 FILLER_60_1097 ();
 sg13g2_decap_8 FILLER_60_1104 ();
 sg13g2_decap_8 FILLER_60_1111 ();
 sg13g2_decap_8 FILLER_60_1118 ();
 sg13g2_decap_8 FILLER_60_1125 ();
 sg13g2_decap_8 FILLER_60_1132 ();
 sg13g2_decap_8 FILLER_60_1139 ();
 sg13g2_decap_8 FILLER_60_1146 ();
 sg13g2_decap_8 FILLER_60_1153 ();
 sg13g2_decap_8 FILLER_60_1160 ();
 sg13g2_decap_8 FILLER_60_1167 ();
 sg13g2_decap_8 FILLER_60_1174 ();
 sg13g2_decap_8 FILLER_60_1181 ();
 sg13g2_decap_8 FILLER_60_1188 ();
 sg13g2_decap_8 FILLER_60_1195 ();
 sg13g2_decap_8 FILLER_60_1202 ();
 sg13g2_decap_8 FILLER_60_1209 ();
 sg13g2_decap_8 FILLER_60_1216 ();
 sg13g2_decap_8 FILLER_60_1223 ();
 sg13g2_decap_8 FILLER_60_1230 ();
 sg13g2_decap_8 FILLER_60_1237 ();
 sg13g2_decap_8 FILLER_60_1244 ();
 sg13g2_decap_8 FILLER_60_1251 ();
 sg13g2_decap_8 FILLER_60_1258 ();
 sg13g2_decap_8 FILLER_60_1265 ();
 sg13g2_decap_8 FILLER_60_1272 ();
 sg13g2_decap_8 FILLER_60_1279 ();
 sg13g2_decap_8 FILLER_60_1286 ();
 sg13g2_decap_8 FILLER_60_1293 ();
 sg13g2_decap_8 FILLER_60_1300 ();
 sg13g2_decap_8 FILLER_60_1307 ();
 sg13g2_decap_8 FILLER_60_1314 ();
 sg13g2_decap_4 FILLER_60_1321 ();
 sg13g2_fill_1 FILLER_60_1325 ();
 sg13g2_fill_2 FILLER_61_107 ();
 sg13g2_fill_1 FILLER_61_161 ();
 sg13g2_fill_1 FILLER_61_166 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_176 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_fill_1 FILLER_61_220 ();
 sg13g2_fill_1 FILLER_61_330 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_2 FILLER_61_393 ();
 sg13g2_fill_2 FILLER_61_491 ();
 sg13g2_fill_2 FILLER_61_549 ();
 sg13g2_fill_1 FILLER_61_565 ();
 sg13g2_fill_2 FILLER_61_592 ();
 sg13g2_fill_2 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_606 ();
 sg13g2_fill_1 FILLER_61_627 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_fill_1 FILLER_61_673 ();
 sg13g2_fill_1 FILLER_61_734 ();
 sg13g2_fill_2 FILLER_61_782 ();
 sg13g2_fill_1 FILLER_61_824 ();
 sg13g2_decap_8 FILLER_61_907 ();
 sg13g2_decap_8 FILLER_61_914 ();
 sg13g2_decap_8 FILLER_61_921 ();
 sg13g2_decap_8 FILLER_61_928 ();
 sg13g2_decap_8 FILLER_61_935 ();
 sg13g2_decap_8 FILLER_61_942 ();
 sg13g2_decap_8 FILLER_61_949 ();
 sg13g2_decap_8 FILLER_61_956 ();
 sg13g2_decap_8 FILLER_61_963 ();
 sg13g2_decap_8 FILLER_61_970 ();
 sg13g2_decap_8 FILLER_61_977 ();
 sg13g2_decap_8 FILLER_61_984 ();
 sg13g2_decap_8 FILLER_61_991 ();
 sg13g2_decap_8 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1005 ();
 sg13g2_decap_8 FILLER_61_1012 ();
 sg13g2_decap_8 FILLER_61_1019 ();
 sg13g2_decap_8 FILLER_61_1026 ();
 sg13g2_decap_8 FILLER_61_1033 ();
 sg13g2_decap_8 FILLER_61_1040 ();
 sg13g2_decap_8 FILLER_61_1047 ();
 sg13g2_decap_8 FILLER_61_1054 ();
 sg13g2_decap_8 FILLER_61_1061 ();
 sg13g2_decap_8 FILLER_61_1068 ();
 sg13g2_decap_8 FILLER_61_1075 ();
 sg13g2_decap_8 FILLER_61_1082 ();
 sg13g2_decap_8 FILLER_61_1089 ();
 sg13g2_decap_8 FILLER_61_1096 ();
 sg13g2_decap_8 FILLER_61_1103 ();
 sg13g2_decap_8 FILLER_61_1110 ();
 sg13g2_decap_8 FILLER_61_1117 ();
 sg13g2_decap_8 FILLER_61_1124 ();
 sg13g2_decap_8 FILLER_61_1131 ();
 sg13g2_decap_8 FILLER_61_1138 ();
 sg13g2_decap_8 FILLER_61_1145 ();
 sg13g2_decap_8 FILLER_61_1152 ();
 sg13g2_decap_8 FILLER_61_1159 ();
 sg13g2_decap_8 FILLER_61_1166 ();
 sg13g2_decap_8 FILLER_61_1173 ();
 sg13g2_decap_8 FILLER_61_1180 ();
 sg13g2_decap_8 FILLER_61_1187 ();
 sg13g2_decap_8 FILLER_61_1194 ();
 sg13g2_decap_8 FILLER_61_1201 ();
 sg13g2_decap_8 FILLER_61_1208 ();
 sg13g2_decap_8 FILLER_61_1215 ();
 sg13g2_decap_8 FILLER_61_1222 ();
 sg13g2_decap_8 FILLER_61_1229 ();
 sg13g2_decap_8 FILLER_61_1236 ();
 sg13g2_decap_8 FILLER_61_1243 ();
 sg13g2_decap_8 FILLER_61_1250 ();
 sg13g2_decap_8 FILLER_61_1257 ();
 sg13g2_decap_8 FILLER_61_1264 ();
 sg13g2_decap_8 FILLER_61_1271 ();
 sg13g2_decap_8 FILLER_61_1278 ();
 sg13g2_decap_8 FILLER_61_1285 ();
 sg13g2_decap_8 FILLER_61_1292 ();
 sg13g2_decap_8 FILLER_61_1299 ();
 sg13g2_decap_8 FILLER_61_1306 ();
 sg13g2_decap_8 FILLER_61_1313 ();
 sg13g2_decap_4 FILLER_61_1320 ();
 sg13g2_fill_2 FILLER_61_1324 ();
 sg13g2_fill_2 FILLER_62_46 ();
 sg13g2_fill_1 FILLER_62_48 ();
 sg13g2_fill_1 FILLER_62_64 ();
 sg13g2_fill_2 FILLER_62_70 ();
 sg13g2_fill_2 FILLER_62_81 ();
 sg13g2_fill_1 FILLER_62_111 ();
 sg13g2_fill_2 FILLER_62_167 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_297 ();
 sg13g2_fill_1 FILLER_62_335 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_62_364 ();
 sg13g2_fill_1 FILLER_62_456 ();
 sg13g2_fill_1 FILLER_62_467 ();
 sg13g2_fill_1 FILLER_62_494 ();
 sg13g2_fill_1 FILLER_62_531 ();
 sg13g2_fill_1 FILLER_62_542 ();
 sg13g2_fill_2 FILLER_62_553 ();
 sg13g2_fill_1 FILLER_62_555 ();
 sg13g2_fill_2 FILLER_62_608 ();
 sg13g2_fill_1 FILLER_62_610 ();
 sg13g2_fill_2 FILLER_62_651 ();
 sg13g2_fill_2 FILLER_62_663 ();
 sg13g2_fill_1 FILLER_62_665 ();
 sg13g2_fill_2 FILLER_62_710 ();
 sg13g2_fill_1 FILLER_62_722 ();
 sg13g2_fill_2 FILLER_62_749 ();
 sg13g2_fill_2 FILLER_62_791 ();
 sg13g2_fill_1 FILLER_62_793 ();
 sg13g2_fill_2 FILLER_62_804 ();
 sg13g2_fill_1 FILLER_62_820 ();
 sg13g2_fill_1 FILLER_62_857 ();
 sg13g2_decap_8 FILLER_62_884 ();
 sg13g2_decap_8 FILLER_62_891 ();
 sg13g2_decap_8 FILLER_62_898 ();
 sg13g2_decap_8 FILLER_62_905 ();
 sg13g2_decap_8 FILLER_62_912 ();
 sg13g2_decap_8 FILLER_62_919 ();
 sg13g2_decap_8 FILLER_62_926 ();
 sg13g2_decap_8 FILLER_62_933 ();
 sg13g2_decap_8 FILLER_62_940 ();
 sg13g2_decap_8 FILLER_62_947 ();
 sg13g2_decap_8 FILLER_62_954 ();
 sg13g2_decap_8 FILLER_62_961 ();
 sg13g2_decap_8 FILLER_62_968 ();
 sg13g2_decap_8 FILLER_62_975 ();
 sg13g2_decap_8 FILLER_62_982 ();
 sg13g2_decap_8 FILLER_62_989 ();
 sg13g2_decap_8 FILLER_62_996 ();
 sg13g2_decap_8 FILLER_62_1003 ();
 sg13g2_decap_8 FILLER_62_1010 ();
 sg13g2_decap_8 FILLER_62_1017 ();
 sg13g2_decap_8 FILLER_62_1024 ();
 sg13g2_decap_8 FILLER_62_1031 ();
 sg13g2_decap_8 FILLER_62_1038 ();
 sg13g2_decap_8 FILLER_62_1045 ();
 sg13g2_decap_8 FILLER_62_1052 ();
 sg13g2_decap_8 FILLER_62_1059 ();
 sg13g2_decap_8 FILLER_62_1066 ();
 sg13g2_decap_8 FILLER_62_1073 ();
 sg13g2_decap_8 FILLER_62_1080 ();
 sg13g2_decap_8 FILLER_62_1087 ();
 sg13g2_decap_8 FILLER_62_1094 ();
 sg13g2_decap_8 FILLER_62_1101 ();
 sg13g2_decap_8 FILLER_62_1108 ();
 sg13g2_decap_8 FILLER_62_1115 ();
 sg13g2_decap_8 FILLER_62_1122 ();
 sg13g2_decap_8 FILLER_62_1129 ();
 sg13g2_decap_8 FILLER_62_1136 ();
 sg13g2_decap_8 FILLER_62_1143 ();
 sg13g2_decap_8 FILLER_62_1150 ();
 sg13g2_decap_8 FILLER_62_1157 ();
 sg13g2_decap_8 FILLER_62_1164 ();
 sg13g2_decap_8 FILLER_62_1171 ();
 sg13g2_decap_8 FILLER_62_1178 ();
 sg13g2_decap_8 FILLER_62_1185 ();
 sg13g2_decap_8 FILLER_62_1192 ();
 sg13g2_decap_8 FILLER_62_1199 ();
 sg13g2_decap_8 FILLER_62_1206 ();
 sg13g2_decap_8 FILLER_62_1213 ();
 sg13g2_decap_8 FILLER_62_1220 ();
 sg13g2_decap_8 FILLER_62_1227 ();
 sg13g2_decap_8 FILLER_62_1234 ();
 sg13g2_decap_8 FILLER_62_1241 ();
 sg13g2_decap_8 FILLER_62_1248 ();
 sg13g2_decap_8 FILLER_62_1255 ();
 sg13g2_decap_8 FILLER_62_1262 ();
 sg13g2_decap_8 FILLER_62_1269 ();
 sg13g2_decap_8 FILLER_62_1276 ();
 sg13g2_decap_8 FILLER_62_1283 ();
 sg13g2_decap_8 FILLER_62_1290 ();
 sg13g2_decap_8 FILLER_62_1297 ();
 sg13g2_decap_8 FILLER_62_1304 ();
 sg13g2_decap_8 FILLER_62_1311 ();
 sg13g2_decap_8 FILLER_62_1318 ();
 sg13g2_fill_1 FILLER_62_1325 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_86 ();
 sg13g2_fill_1 FILLER_63_101 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_fill_2 FILLER_63_164 ();
 sg13g2_fill_1 FILLER_63_166 ();
 sg13g2_fill_2 FILLER_63_225 ();
 sg13g2_fill_2 FILLER_63_247 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_fill_2 FILLER_63_344 ();
 sg13g2_fill_2 FILLER_63_363 ();
 sg13g2_fill_2 FILLER_63_387 ();
 sg13g2_fill_1 FILLER_63_419 ();
 sg13g2_fill_2 FILLER_63_474 ();
 sg13g2_fill_1 FILLER_63_476 ();
 sg13g2_fill_1 FILLER_63_669 ();
 sg13g2_fill_2 FILLER_63_690 ();
 sg13g2_fill_1 FILLER_63_692 ();
 sg13g2_fill_1 FILLER_63_805 ();
 sg13g2_fill_1 FILLER_63_832 ();
 sg13g2_decap_8 FILLER_63_877 ();
 sg13g2_decap_8 FILLER_63_884 ();
 sg13g2_decap_8 FILLER_63_891 ();
 sg13g2_decap_8 FILLER_63_898 ();
 sg13g2_decap_8 FILLER_63_905 ();
 sg13g2_decap_8 FILLER_63_912 ();
 sg13g2_decap_8 FILLER_63_919 ();
 sg13g2_decap_8 FILLER_63_926 ();
 sg13g2_decap_8 FILLER_63_933 ();
 sg13g2_decap_8 FILLER_63_940 ();
 sg13g2_decap_8 FILLER_63_947 ();
 sg13g2_decap_8 FILLER_63_954 ();
 sg13g2_decap_8 FILLER_63_961 ();
 sg13g2_decap_8 FILLER_63_968 ();
 sg13g2_decap_8 FILLER_63_975 ();
 sg13g2_decap_8 FILLER_63_982 ();
 sg13g2_decap_8 FILLER_63_989 ();
 sg13g2_decap_8 FILLER_63_996 ();
 sg13g2_decap_8 FILLER_63_1003 ();
 sg13g2_decap_8 FILLER_63_1010 ();
 sg13g2_decap_8 FILLER_63_1017 ();
 sg13g2_decap_8 FILLER_63_1024 ();
 sg13g2_decap_8 FILLER_63_1031 ();
 sg13g2_decap_8 FILLER_63_1038 ();
 sg13g2_decap_8 FILLER_63_1045 ();
 sg13g2_decap_8 FILLER_63_1052 ();
 sg13g2_decap_8 FILLER_63_1059 ();
 sg13g2_decap_8 FILLER_63_1066 ();
 sg13g2_decap_8 FILLER_63_1073 ();
 sg13g2_decap_8 FILLER_63_1080 ();
 sg13g2_decap_8 FILLER_63_1087 ();
 sg13g2_decap_8 FILLER_63_1094 ();
 sg13g2_decap_8 FILLER_63_1101 ();
 sg13g2_decap_8 FILLER_63_1108 ();
 sg13g2_decap_8 FILLER_63_1115 ();
 sg13g2_decap_8 FILLER_63_1122 ();
 sg13g2_decap_8 FILLER_63_1129 ();
 sg13g2_decap_8 FILLER_63_1136 ();
 sg13g2_decap_8 FILLER_63_1143 ();
 sg13g2_decap_8 FILLER_63_1150 ();
 sg13g2_decap_8 FILLER_63_1157 ();
 sg13g2_decap_8 FILLER_63_1164 ();
 sg13g2_decap_8 FILLER_63_1171 ();
 sg13g2_decap_8 FILLER_63_1178 ();
 sg13g2_decap_8 FILLER_63_1185 ();
 sg13g2_decap_8 FILLER_63_1192 ();
 sg13g2_decap_8 FILLER_63_1199 ();
 sg13g2_decap_8 FILLER_63_1206 ();
 sg13g2_decap_8 FILLER_63_1213 ();
 sg13g2_decap_8 FILLER_63_1220 ();
 sg13g2_decap_8 FILLER_63_1227 ();
 sg13g2_decap_8 FILLER_63_1234 ();
 sg13g2_decap_8 FILLER_63_1241 ();
 sg13g2_decap_8 FILLER_63_1248 ();
 sg13g2_decap_8 FILLER_63_1255 ();
 sg13g2_decap_8 FILLER_63_1262 ();
 sg13g2_decap_8 FILLER_63_1269 ();
 sg13g2_decap_8 FILLER_63_1276 ();
 sg13g2_decap_8 FILLER_63_1283 ();
 sg13g2_decap_8 FILLER_63_1290 ();
 sg13g2_decap_8 FILLER_63_1297 ();
 sg13g2_decap_8 FILLER_63_1304 ();
 sg13g2_decap_8 FILLER_63_1311 ();
 sg13g2_decap_8 FILLER_63_1318 ();
 sg13g2_fill_1 FILLER_63_1325 ();
 sg13g2_fill_1 FILLER_64_26 ();
 sg13g2_fill_2 FILLER_64_50 ();
 sg13g2_fill_1 FILLER_64_52 ();
 sg13g2_fill_2 FILLER_64_58 ();
 sg13g2_fill_1 FILLER_64_60 ();
 sg13g2_fill_2 FILLER_64_137 ();
 sg13g2_fill_2 FILLER_64_153 ();
 sg13g2_fill_2 FILLER_64_166 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_1 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_340 ();
 sg13g2_fill_1 FILLER_64_354 ();
 sg13g2_fill_2 FILLER_64_432 ();
 sg13g2_fill_1 FILLER_64_434 ();
 sg13g2_fill_1 FILLER_64_491 ();
 sg13g2_fill_2 FILLER_64_554 ();
 sg13g2_fill_2 FILLER_64_612 ();
 sg13g2_fill_1 FILLER_64_614 ();
 sg13g2_fill_2 FILLER_64_649 ();
 sg13g2_fill_2 FILLER_64_775 ();
 sg13g2_fill_1 FILLER_64_777 ();
 sg13g2_fill_1 FILLER_64_850 ();
 sg13g2_decap_8 FILLER_64_875 ();
 sg13g2_decap_8 FILLER_64_882 ();
 sg13g2_decap_8 FILLER_64_889 ();
 sg13g2_decap_8 FILLER_64_896 ();
 sg13g2_decap_8 FILLER_64_903 ();
 sg13g2_decap_8 FILLER_64_910 ();
 sg13g2_decap_8 FILLER_64_917 ();
 sg13g2_decap_8 FILLER_64_924 ();
 sg13g2_decap_8 FILLER_64_931 ();
 sg13g2_decap_8 FILLER_64_938 ();
 sg13g2_decap_8 FILLER_64_945 ();
 sg13g2_decap_8 FILLER_64_952 ();
 sg13g2_decap_8 FILLER_64_959 ();
 sg13g2_decap_8 FILLER_64_966 ();
 sg13g2_decap_8 FILLER_64_973 ();
 sg13g2_decap_8 FILLER_64_980 ();
 sg13g2_decap_8 FILLER_64_987 ();
 sg13g2_decap_8 FILLER_64_994 ();
 sg13g2_decap_8 FILLER_64_1001 ();
 sg13g2_decap_8 FILLER_64_1008 ();
 sg13g2_decap_8 FILLER_64_1015 ();
 sg13g2_decap_8 FILLER_64_1022 ();
 sg13g2_decap_8 FILLER_64_1029 ();
 sg13g2_decap_8 FILLER_64_1036 ();
 sg13g2_decap_8 FILLER_64_1043 ();
 sg13g2_decap_8 FILLER_64_1050 ();
 sg13g2_decap_8 FILLER_64_1057 ();
 sg13g2_decap_8 FILLER_64_1064 ();
 sg13g2_decap_8 FILLER_64_1071 ();
 sg13g2_decap_8 FILLER_64_1078 ();
 sg13g2_decap_8 FILLER_64_1085 ();
 sg13g2_decap_8 FILLER_64_1092 ();
 sg13g2_decap_8 FILLER_64_1099 ();
 sg13g2_decap_8 FILLER_64_1106 ();
 sg13g2_decap_8 FILLER_64_1113 ();
 sg13g2_decap_8 FILLER_64_1120 ();
 sg13g2_decap_8 FILLER_64_1127 ();
 sg13g2_decap_8 FILLER_64_1134 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_decap_8 FILLER_64_1148 ();
 sg13g2_decap_8 FILLER_64_1155 ();
 sg13g2_decap_8 FILLER_64_1162 ();
 sg13g2_decap_8 FILLER_64_1169 ();
 sg13g2_decap_8 FILLER_64_1176 ();
 sg13g2_decap_8 FILLER_64_1183 ();
 sg13g2_decap_8 FILLER_64_1190 ();
 sg13g2_decap_8 FILLER_64_1197 ();
 sg13g2_decap_8 FILLER_64_1204 ();
 sg13g2_decap_8 FILLER_64_1211 ();
 sg13g2_decap_8 FILLER_64_1218 ();
 sg13g2_decap_8 FILLER_64_1225 ();
 sg13g2_decap_8 FILLER_64_1232 ();
 sg13g2_decap_8 FILLER_64_1239 ();
 sg13g2_decap_8 FILLER_64_1246 ();
 sg13g2_decap_8 FILLER_64_1253 ();
 sg13g2_decap_8 FILLER_64_1260 ();
 sg13g2_decap_8 FILLER_64_1267 ();
 sg13g2_decap_8 FILLER_64_1274 ();
 sg13g2_decap_8 FILLER_64_1281 ();
 sg13g2_decap_8 FILLER_64_1288 ();
 sg13g2_decap_8 FILLER_64_1295 ();
 sg13g2_decap_8 FILLER_64_1302 ();
 sg13g2_decap_8 FILLER_64_1309 ();
 sg13g2_decap_8 FILLER_64_1316 ();
 sg13g2_fill_2 FILLER_64_1323 ();
 sg13g2_fill_1 FILLER_64_1325 ();
 sg13g2_fill_2 FILLER_65_65 ();
 sg13g2_fill_2 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_95 ();
 sg13g2_fill_1 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_128 ();
 sg13g2_fill_1 FILLER_65_149 ();
 sg13g2_fill_2 FILLER_65_163 ();
 sg13g2_fill_1 FILLER_65_165 ();
 sg13g2_fill_2 FILLER_65_181 ();
 sg13g2_fill_1 FILLER_65_189 ();
 sg13g2_fill_1 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_217 ();
 sg13g2_fill_1 FILLER_65_235 ();
 sg13g2_fill_1 FILLER_65_294 ();
 sg13g2_fill_2 FILLER_65_329 ();
 sg13g2_fill_1 FILLER_65_410 ();
 sg13g2_fill_1 FILLER_65_437 ();
 sg13g2_fill_2 FILLER_65_448 ();
 sg13g2_fill_1 FILLER_65_450 ();
 sg13g2_fill_1 FILLER_65_491 ();
 sg13g2_fill_2 FILLER_65_518 ();
 sg13g2_fill_1 FILLER_65_560 ();
 sg13g2_fill_1 FILLER_65_583 ();
 sg13g2_fill_2 FILLER_65_623 ();
 sg13g2_fill_2 FILLER_65_695 ();
 sg13g2_fill_1 FILLER_65_697 ();
 sg13g2_fill_1 FILLER_65_738 ();
 sg13g2_fill_2 FILLER_65_827 ();
 sg13g2_fill_1 FILLER_65_829 ();
 sg13g2_decap_8 FILLER_65_868 ();
 sg13g2_decap_8 FILLER_65_875 ();
 sg13g2_decap_8 FILLER_65_882 ();
 sg13g2_decap_8 FILLER_65_889 ();
 sg13g2_decap_8 FILLER_65_896 ();
 sg13g2_decap_8 FILLER_65_903 ();
 sg13g2_decap_8 FILLER_65_910 ();
 sg13g2_decap_8 FILLER_65_917 ();
 sg13g2_decap_8 FILLER_65_924 ();
 sg13g2_decap_8 FILLER_65_931 ();
 sg13g2_decap_8 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_945 ();
 sg13g2_decap_8 FILLER_65_952 ();
 sg13g2_decap_8 FILLER_65_959 ();
 sg13g2_decap_8 FILLER_65_966 ();
 sg13g2_decap_8 FILLER_65_973 ();
 sg13g2_decap_8 FILLER_65_980 ();
 sg13g2_decap_8 FILLER_65_987 ();
 sg13g2_decap_8 FILLER_65_994 ();
 sg13g2_decap_8 FILLER_65_1001 ();
 sg13g2_decap_8 FILLER_65_1008 ();
 sg13g2_decap_8 FILLER_65_1015 ();
 sg13g2_decap_8 FILLER_65_1022 ();
 sg13g2_decap_8 FILLER_65_1029 ();
 sg13g2_decap_8 FILLER_65_1036 ();
 sg13g2_decap_8 FILLER_65_1043 ();
 sg13g2_decap_8 FILLER_65_1050 ();
 sg13g2_decap_8 FILLER_65_1057 ();
 sg13g2_decap_8 FILLER_65_1064 ();
 sg13g2_decap_8 FILLER_65_1071 ();
 sg13g2_decap_8 FILLER_65_1078 ();
 sg13g2_decap_8 FILLER_65_1085 ();
 sg13g2_decap_8 FILLER_65_1092 ();
 sg13g2_decap_8 FILLER_65_1099 ();
 sg13g2_decap_8 FILLER_65_1106 ();
 sg13g2_decap_8 FILLER_65_1113 ();
 sg13g2_decap_8 FILLER_65_1120 ();
 sg13g2_decap_8 FILLER_65_1127 ();
 sg13g2_decap_8 FILLER_65_1134 ();
 sg13g2_decap_8 FILLER_65_1141 ();
 sg13g2_decap_8 FILLER_65_1148 ();
 sg13g2_decap_8 FILLER_65_1155 ();
 sg13g2_decap_8 FILLER_65_1162 ();
 sg13g2_decap_8 FILLER_65_1169 ();
 sg13g2_decap_8 FILLER_65_1176 ();
 sg13g2_decap_8 FILLER_65_1183 ();
 sg13g2_decap_8 FILLER_65_1190 ();
 sg13g2_decap_8 FILLER_65_1197 ();
 sg13g2_decap_8 FILLER_65_1204 ();
 sg13g2_decap_8 FILLER_65_1211 ();
 sg13g2_decap_8 FILLER_65_1218 ();
 sg13g2_decap_8 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1232 ();
 sg13g2_decap_8 FILLER_65_1239 ();
 sg13g2_decap_8 FILLER_65_1246 ();
 sg13g2_decap_8 FILLER_65_1253 ();
 sg13g2_decap_8 FILLER_65_1260 ();
 sg13g2_decap_8 FILLER_65_1267 ();
 sg13g2_decap_8 FILLER_65_1274 ();
 sg13g2_decap_8 FILLER_65_1281 ();
 sg13g2_decap_8 FILLER_65_1288 ();
 sg13g2_decap_8 FILLER_65_1295 ();
 sg13g2_decap_8 FILLER_65_1302 ();
 sg13g2_decap_8 FILLER_65_1309 ();
 sg13g2_decap_8 FILLER_65_1316 ();
 sg13g2_fill_2 FILLER_65_1323 ();
 sg13g2_fill_1 FILLER_65_1325 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_25 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_fill_1 FILLER_66_189 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_1 FILLER_66_277 ();
 sg13g2_fill_2 FILLER_66_340 ();
 sg13g2_fill_1 FILLER_66_402 ();
 sg13g2_fill_1 FILLER_66_413 ();
 sg13g2_fill_1 FILLER_66_428 ();
 sg13g2_fill_1 FILLER_66_469 ();
 sg13g2_fill_2 FILLER_66_612 ();
 sg13g2_fill_2 FILLER_66_628 ();
 sg13g2_fill_1 FILLER_66_652 ();
 sg13g2_fill_2 FILLER_66_711 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_729 ();
 sg13g2_fill_2 FILLER_66_764 ();
 sg13g2_fill_1 FILLER_66_766 ();
 sg13g2_fill_1 FILLER_66_829 ();
 sg13g2_decap_8 FILLER_66_856 ();
 sg13g2_decap_8 FILLER_66_863 ();
 sg13g2_decap_8 FILLER_66_870 ();
 sg13g2_decap_8 FILLER_66_877 ();
 sg13g2_decap_8 FILLER_66_884 ();
 sg13g2_decap_8 FILLER_66_891 ();
 sg13g2_decap_8 FILLER_66_898 ();
 sg13g2_decap_8 FILLER_66_905 ();
 sg13g2_decap_8 FILLER_66_912 ();
 sg13g2_decap_8 FILLER_66_919 ();
 sg13g2_decap_8 FILLER_66_926 ();
 sg13g2_decap_8 FILLER_66_933 ();
 sg13g2_decap_8 FILLER_66_940 ();
 sg13g2_decap_8 FILLER_66_947 ();
 sg13g2_decap_8 FILLER_66_954 ();
 sg13g2_decap_8 FILLER_66_961 ();
 sg13g2_decap_8 FILLER_66_968 ();
 sg13g2_decap_8 FILLER_66_975 ();
 sg13g2_decap_8 FILLER_66_982 ();
 sg13g2_decap_8 FILLER_66_989 ();
 sg13g2_decap_8 FILLER_66_996 ();
 sg13g2_decap_8 FILLER_66_1003 ();
 sg13g2_decap_8 FILLER_66_1010 ();
 sg13g2_decap_8 FILLER_66_1017 ();
 sg13g2_decap_8 FILLER_66_1024 ();
 sg13g2_decap_8 FILLER_66_1031 ();
 sg13g2_decap_8 FILLER_66_1038 ();
 sg13g2_decap_8 FILLER_66_1045 ();
 sg13g2_decap_8 FILLER_66_1052 ();
 sg13g2_decap_8 FILLER_66_1059 ();
 sg13g2_decap_8 FILLER_66_1066 ();
 sg13g2_decap_8 FILLER_66_1073 ();
 sg13g2_decap_8 FILLER_66_1080 ();
 sg13g2_decap_8 FILLER_66_1087 ();
 sg13g2_decap_8 FILLER_66_1094 ();
 sg13g2_decap_8 FILLER_66_1101 ();
 sg13g2_decap_8 FILLER_66_1108 ();
 sg13g2_decap_8 FILLER_66_1115 ();
 sg13g2_decap_8 FILLER_66_1122 ();
 sg13g2_decap_8 FILLER_66_1129 ();
 sg13g2_decap_8 FILLER_66_1136 ();
 sg13g2_decap_8 FILLER_66_1143 ();
 sg13g2_decap_8 FILLER_66_1150 ();
 sg13g2_decap_8 FILLER_66_1157 ();
 sg13g2_decap_8 FILLER_66_1164 ();
 sg13g2_decap_8 FILLER_66_1171 ();
 sg13g2_decap_8 FILLER_66_1178 ();
 sg13g2_decap_8 FILLER_66_1185 ();
 sg13g2_decap_8 FILLER_66_1192 ();
 sg13g2_decap_8 FILLER_66_1199 ();
 sg13g2_decap_8 FILLER_66_1206 ();
 sg13g2_decap_8 FILLER_66_1213 ();
 sg13g2_decap_8 FILLER_66_1220 ();
 sg13g2_decap_8 FILLER_66_1227 ();
 sg13g2_decap_8 FILLER_66_1234 ();
 sg13g2_decap_8 FILLER_66_1241 ();
 sg13g2_decap_8 FILLER_66_1248 ();
 sg13g2_decap_8 FILLER_66_1255 ();
 sg13g2_decap_8 FILLER_66_1262 ();
 sg13g2_decap_8 FILLER_66_1269 ();
 sg13g2_decap_8 FILLER_66_1276 ();
 sg13g2_decap_8 FILLER_66_1283 ();
 sg13g2_decap_8 FILLER_66_1290 ();
 sg13g2_decap_8 FILLER_66_1297 ();
 sg13g2_decap_8 FILLER_66_1304 ();
 sg13g2_decap_8 FILLER_66_1311 ();
 sg13g2_decap_8 FILLER_66_1318 ();
 sg13g2_fill_1 FILLER_66_1325 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_27 ();
 sg13g2_fill_1 FILLER_67_33 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_81 ();
 sg13g2_fill_1 FILLER_67_88 ();
 sg13g2_fill_2 FILLER_67_94 ();
 sg13g2_fill_1 FILLER_67_96 ();
 sg13g2_fill_2 FILLER_67_164 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_193 ();
 sg13g2_fill_1 FILLER_67_226 ();
 sg13g2_fill_2 FILLER_67_247 ();
 sg13g2_fill_2 FILLER_67_307 ();
 sg13g2_fill_2 FILLER_67_315 ();
 sg13g2_fill_1 FILLER_67_425 ();
 sg13g2_fill_2 FILLER_67_452 ();
 sg13g2_fill_1 FILLER_67_454 ();
 sg13g2_fill_2 FILLER_67_575 ();
 sg13g2_fill_1 FILLER_67_577 ();
 sg13g2_fill_1 FILLER_67_612 ();
 sg13g2_fill_1 FILLER_67_776 ();
 sg13g2_fill_2 FILLER_67_815 ();
 sg13g2_fill_2 FILLER_67_827 ();
 sg13g2_fill_2 FILLER_67_839 ();
 sg13g2_decap_8 FILLER_67_845 ();
 sg13g2_decap_8 FILLER_67_852 ();
 sg13g2_decap_8 FILLER_67_859 ();
 sg13g2_decap_8 FILLER_67_866 ();
 sg13g2_decap_8 FILLER_67_873 ();
 sg13g2_decap_8 FILLER_67_880 ();
 sg13g2_decap_8 FILLER_67_887 ();
 sg13g2_decap_8 FILLER_67_894 ();
 sg13g2_decap_8 FILLER_67_901 ();
 sg13g2_decap_8 FILLER_67_908 ();
 sg13g2_decap_8 FILLER_67_915 ();
 sg13g2_decap_8 FILLER_67_922 ();
 sg13g2_decap_8 FILLER_67_929 ();
 sg13g2_decap_8 FILLER_67_936 ();
 sg13g2_decap_8 FILLER_67_943 ();
 sg13g2_decap_8 FILLER_67_950 ();
 sg13g2_decap_8 FILLER_67_957 ();
 sg13g2_decap_8 FILLER_67_964 ();
 sg13g2_decap_8 FILLER_67_971 ();
 sg13g2_decap_8 FILLER_67_978 ();
 sg13g2_decap_8 FILLER_67_985 ();
 sg13g2_decap_8 FILLER_67_992 ();
 sg13g2_decap_8 FILLER_67_999 ();
 sg13g2_decap_8 FILLER_67_1006 ();
 sg13g2_decap_8 FILLER_67_1013 ();
 sg13g2_decap_8 FILLER_67_1020 ();
 sg13g2_decap_8 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1034 ();
 sg13g2_decap_8 FILLER_67_1041 ();
 sg13g2_decap_8 FILLER_67_1048 ();
 sg13g2_decap_8 FILLER_67_1055 ();
 sg13g2_decap_8 FILLER_67_1062 ();
 sg13g2_decap_8 FILLER_67_1069 ();
 sg13g2_decap_8 FILLER_67_1076 ();
 sg13g2_decap_8 FILLER_67_1083 ();
 sg13g2_decap_8 FILLER_67_1090 ();
 sg13g2_decap_8 FILLER_67_1097 ();
 sg13g2_decap_8 FILLER_67_1104 ();
 sg13g2_decap_8 FILLER_67_1111 ();
 sg13g2_decap_8 FILLER_67_1118 ();
 sg13g2_decap_8 FILLER_67_1125 ();
 sg13g2_decap_8 FILLER_67_1132 ();
 sg13g2_decap_8 FILLER_67_1139 ();
 sg13g2_decap_8 FILLER_67_1146 ();
 sg13g2_decap_8 FILLER_67_1153 ();
 sg13g2_decap_8 FILLER_67_1160 ();
 sg13g2_decap_8 FILLER_67_1167 ();
 sg13g2_decap_8 FILLER_67_1174 ();
 sg13g2_decap_8 FILLER_67_1181 ();
 sg13g2_decap_8 FILLER_67_1188 ();
 sg13g2_decap_8 FILLER_67_1195 ();
 sg13g2_decap_8 FILLER_67_1202 ();
 sg13g2_decap_8 FILLER_67_1209 ();
 sg13g2_decap_8 FILLER_67_1216 ();
 sg13g2_decap_8 FILLER_67_1223 ();
 sg13g2_decap_8 FILLER_67_1230 ();
 sg13g2_decap_8 FILLER_67_1237 ();
 sg13g2_decap_8 FILLER_67_1244 ();
 sg13g2_decap_8 FILLER_67_1251 ();
 sg13g2_decap_8 FILLER_67_1258 ();
 sg13g2_decap_8 FILLER_67_1265 ();
 sg13g2_decap_8 FILLER_67_1272 ();
 sg13g2_decap_8 FILLER_67_1279 ();
 sg13g2_decap_8 FILLER_67_1286 ();
 sg13g2_decap_8 FILLER_67_1293 ();
 sg13g2_decap_8 FILLER_67_1300 ();
 sg13g2_decap_8 FILLER_67_1307 ();
 sg13g2_decap_8 FILLER_67_1314 ();
 sg13g2_decap_4 FILLER_67_1321 ();
 sg13g2_fill_1 FILLER_67_1325 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_fill_2 FILLER_68_42 ();
 sg13g2_fill_1 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_85 ();
 sg13g2_fill_1 FILLER_68_99 ();
 sg13g2_fill_1 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_115 ();
 sg13g2_fill_2 FILLER_68_122 ();
 sg13g2_fill_2 FILLER_68_150 ();
 sg13g2_fill_1 FILLER_68_269 ();
 sg13g2_fill_2 FILLER_68_375 ();
 sg13g2_fill_1 FILLER_68_411 ();
 sg13g2_fill_1 FILLER_68_438 ();
 sg13g2_fill_2 FILLER_68_475 ();
 sg13g2_fill_1 FILLER_68_477 ();
 sg13g2_fill_1 FILLER_68_508 ();
 sg13g2_fill_1 FILLER_68_542 ();
 sg13g2_fill_1 FILLER_68_569 ();
 sg13g2_fill_1 FILLER_68_580 ();
 sg13g2_fill_1 FILLER_68_591 ();
 sg13g2_fill_1 FILLER_68_630 ();
 sg13g2_fill_1 FILLER_68_635 ();
 sg13g2_fill_1 FILLER_68_662 ();
 sg13g2_fill_2 FILLER_68_703 ();
 sg13g2_fill_1 FILLER_68_705 ();
 sg13g2_fill_1 FILLER_68_742 ();
 sg13g2_fill_2 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_771 ();
 sg13g2_decap_8 FILLER_68_828 ();
 sg13g2_decap_8 FILLER_68_835 ();
 sg13g2_decap_8 FILLER_68_842 ();
 sg13g2_decap_8 FILLER_68_849 ();
 sg13g2_decap_8 FILLER_68_856 ();
 sg13g2_decap_8 FILLER_68_863 ();
 sg13g2_decap_8 FILLER_68_870 ();
 sg13g2_decap_8 FILLER_68_877 ();
 sg13g2_decap_8 FILLER_68_884 ();
 sg13g2_decap_8 FILLER_68_891 ();
 sg13g2_decap_8 FILLER_68_898 ();
 sg13g2_decap_8 FILLER_68_905 ();
 sg13g2_decap_8 FILLER_68_912 ();
 sg13g2_decap_8 FILLER_68_919 ();
 sg13g2_decap_8 FILLER_68_926 ();
 sg13g2_decap_8 FILLER_68_933 ();
 sg13g2_decap_8 FILLER_68_940 ();
 sg13g2_decap_8 FILLER_68_947 ();
 sg13g2_decap_8 FILLER_68_954 ();
 sg13g2_decap_8 FILLER_68_961 ();
 sg13g2_decap_8 FILLER_68_968 ();
 sg13g2_decap_8 FILLER_68_975 ();
 sg13g2_decap_8 FILLER_68_982 ();
 sg13g2_decap_8 FILLER_68_989 ();
 sg13g2_decap_8 FILLER_68_996 ();
 sg13g2_decap_8 FILLER_68_1003 ();
 sg13g2_decap_8 FILLER_68_1010 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_decap_8 FILLER_68_1024 ();
 sg13g2_decap_8 FILLER_68_1031 ();
 sg13g2_decap_8 FILLER_68_1038 ();
 sg13g2_decap_8 FILLER_68_1045 ();
 sg13g2_decap_8 FILLER_68_1052 ();
 sg13g2_decap_8 FILLER_68_1059 ();
 sg13g2_decap_8 FILLER_68_1066 ();
 sg13g2_decap_8 FILLER_68_1073 ();
 sg13g2_decap_8 FILLER_68_1080 ();
 sg13g2_decap_8 FILLER_68_1087 ();
 sg13g2_decap_8 FILLER_68_1094 ();
 sg13g2_decap_8 FILLER_68_1101 ();
 sg13g2_decap_8 FILLER_68_1108 ();
 sg13g2_decap_8 FILLER_68_1115 ();
 sg13g2_decap_8 FILLER_68_1122 ();
 sg13g2_decap_8 FILLER_68_1129 ();
 sg13g2_decap_8 FILLER_68_1136 ();
 sg13g2_decap_8 FILLER_68_1143 ();
 sg13g2_decap_8 FILLER_68_1150 ();
 sg13g2_decap_8 FILLER_68_1157 ();
 sg13g2_decap_8 FILLER_68_1164 ();
 sg13g2_decap_8 FILLER_68_1171 ();
 sg13g2_decap_8 FILLER_68_1178 ();
 sg13g2_decap_8 FILLER_68_1185 ();
 sg13g2_decap_8 FILLER_68_1192 ();
 sg13g2_decap_8 FILLER_68_1199 ();
 sg13g2_decap_8 FILLER_68_1206 ();
 sg13g2_decap_8 FILLER_68_1213 ();
 sg13g2_decap_8 FILLER_68_1220 ();
 sg13g2_decap_8 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1234 ();
 sg13g2_decap_8 FILLER_68_1241 ();
 sg13g2_decap_8 FILLER_68_1248 ();
 sg13g2_decap_8 FILLER_68_1255 ();
 sg13g2_decap_8 FILLER_68_1262 ();
 sg13g2_decap_8 FILLER_68_1269 ();
 sg13g2_decap_8 FILLER_68_1276 ();
 sg13g2_decap_8 FILLER_68_1283 ();
 sg13g2_decap_8 FILLER_68_1290 ();
 sg13g2_decap_8 FILLER_68_1297 ();
 sg13g2_decap_8 FILLER_68_1304 ();
 sg13g2_decap_8 FILLER_68_1311 ();
 sg13g2_decap_8 FILLER_68_1318 ();
 sg13g2_fill_1 FILLER_68_1325 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_fill_2 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_9 ();
 sg13g2_fill_1 FILLER_69_64 ();
 sg13g2_fill_1 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_76 ();
 sg13g2_fill_1 FILLER_69_103 ();
 sg13g2_fill_1 FILLER_69_130 ();
 sg13g2_fill_1 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_147 ();
 sg13g2_fill_1 FILLER_69_149 ();
 sg13g2_fill_2 FILLER_69_178 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_297 ();
 sg13g2_fill_2 FILLER_69_304 ();
 sg13g2_fill_1 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_352 ();
 sg13g2_fill_2 FILLER_69_454 ();
 sg13g2_fill_2 FILLER_69_470 ();
 sg13g2_fill_2 FILLER_69_494 ();
 sg13g2_fill_1 FILLER_69_496 ();
 sg13g2_fill_1 FILLER_69_606 ();
 sg13g2_fill_1 FILLER_69_617 ();
 sg13g2_fill_1 FILLER_69_644 ();
 sg13g2_fill_2 FILLER_69_653 ();
 sg13g2_fill_2 FILLER_69_659 ();
 sg13g2_fill_2 FILLER_69_683 ();
 sg13g2_fill_1 FILLER_69_685 ();
 sg13g2_fill_1 FILLER_69_694 ();
 sg13g2_fill_1 FILLER_69_700 ();
 sg13g2_fill_2 FILLER_69_711 ();
 sg13g2_fill_1 FILLER_69_713 ();
 sg13g2_fill_2 FILLER_69_762 ();
 sg13g2_fill_2 FILLER_69_792 ();
 sg13g2_fill_1 FILLER_69_794 ();
 sg13g2_decap_8 FILLER_69_821 ();
 sg13g2_decap_8 FILLER_69_828 ();
 sg13g2_decap_8 FILLER_69_835 ();
 sg13g2_decap_8 FILLER_69_842 ();
 sg13g2_decap_8 FILLER_69_849 ();
 sg13g2_decap_8 FILLER_69_856 ();
 sg13g2_decap_8 FILLER_69_863 ();
 sg13g2_decap_8 FILLER_69_870 ();
 sg13g2_decap_8 FILLER_69_877 ();
 sg13g2_decap_8 FILLER_69_884 ();
 sg13g2_decap_8 FILLER_69_891 ();
 sg13g2_decap_8 FILLER_69_898 ();
 sg13g2_decap_8 FILLER_69_905 ();
 sg13g2_decap_8 FILLER_69_912 ();
 sg13g2_decap_8 FILLER_69_919 ();
 sg13g2_decap_8 FILLER_69_926 ();
 sg13g2_decap_8 FILLER_69_933 ();
 sg13g2_decap_8 FILLER_69_940 ();
 sg13g2_decap_8 FILLER_69_947 ();
 sg13g2_decap_8 FILLER_69_954 ();
 sg13g2_decap_8 FILLER_69_961 ();
 sg13g2_decap_8 FILLER_69_968 ();
 sg13g2_decap_8 FILLER_69_975 ();
 sg13g2_decap_8 FILLER_69_982 ();
 sg13g2_decap_8 FILLER_69_989 ();
 sg13g2_decap_8 FILLER_69_996 ();
 sg13g2_decap_8 FILLER_69_1003 ();
 sg13g2_decap_8 FILLER_69_1010 ();
 sg13g2_decap_8 FILLER_69_1017 ();
 sg13g2_decap_8 FILLER_69_1024 ();
 sg13g2_decap_8 FILLER_69_1031 ();
 sg13g2_decap_8 FILLER_69_1038 ();
 sg13g2_decap_8 FILLER_69_1045 ();
 sg13g2_decap_8 FILLER_69_1052 ();
 sg13g2_decap_8 FILLER_69_1059 ();
 sg13g2_decap_8 FILLER_69_1066 ();
 sg13g2_decap_8 FILLER_69_1073 ();
 sg13g2_decap_8 FILLER_69_1080 ();
 sg13g2_decap_8 FILLER_69_1087 ();
 sg13g2_decap_8 FILLER_69_1094 ();
 sg13g2_decap_8 FILLER_69_1101 ();
 sg13g2_decap_8 FILLER_69_1108 ();
 sg13g2_decap_8 FILLER_69_1115 ();
 sg13g2_decap_8 FILLER_69_1122 ();
 sg13g2_decap_8 FILLER_69_1129 ();
 sg13g2_decap_8 FILLER_69_1136 ();
 sg13g2_decap_8 FILLER_69_1143 ();
 sg13g2_decap_8 FILLER_69_1150 ();
 sg13g2_decap_8 FILLER_69_1157 ();
 sg13g2_decap_8 FILLER_69_1164 ();
 sg13g2_decap_8 FILLER_69_1171 ();
 sg13g2_decap_8 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1185 ();
 sg13g2_decap_8 FILLER_69_1192 ();
 sg13g2_decap_8 FILLER_69_1199 ();
 sg13g2_decap_8 FILLER_69_1206 ();
 sg13g2_decap_8 FILLER_69_1213 ();
 sg13g2_decap_8 FILLER_69_1220 ();
 sg13g2_decap_8 FILLER_69_1227 ();
 sg13g2_decap_8 FILLER_69_1234 ();
 sg13g2_decap_8 FILLER_69_1241 ();
 sg13g2_decap_8 FILLER_69_1248 ();
 sg13g2_decap_8 FILLER_69_1255 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_decap_8 FILLER_69_1269 ();
 sg13g2_decap_8 FILLER_69_1276 ();
 sg13g2_decap_8 FILLER_69_1283 ();
 sg13g2_decap_8 FILLER_69_1290 ();
 sg13g2_decap_8 FILLER_69_1297 ();
 sg13g2_decap_8 FILLER_69_1304 ();
 sg13g2_decap_8 FILLER_69_1311 ();
 sg13g2_decap_8 FILLER_69_1318 ();
 sg13g2_fill_1 FILLER_69_1325 ();
 sg13g2_fill_1 FILLER_70_100 ();
 sg13g2_fill_2 FILLER_70_106 ();
 sg13g2_fill_1 FILLER_70_108 ();
 sg13g2_fill_1 FILLER_70_149 ();
 sg13g2_fill_1 FILLER_70_160 ();
 sg13g2_fill_1 FILLER_70_187 ();
 sg13g2_fill_2 FILLER_70_218 ();
 sg13g2_fill_2 FILLER_70_237 ();
 sg13g2_fill_1 FILLER_70_244 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_256 ();
 sg13g2_fill_2 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_306 ();
 sg13g2_fill_1 FILLER_70_316 ();
 sg13g2_fill_1 FILLER_70_343 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_fill_1 FILLER_70_379 ();
 sg13g2_fill_2 FILLER_70_390 ();
 sg13g2_fill_1 FILLER_70_402 ();
 sg13g2_fill_1 FILLER_70_413 ();
 sg13g2_fill_1 FILLER_70_516 ();
 sg13g2_fill_2 FILLER_70_531 ();
 sg13g2_fill_2 FILLER_70_559 ();
 sg13g2_fill_2 FILLER_70_571 ();
 sg13g2_fill_1 FILLER_70_589 ();
 sg13g2_fill_2 FILLER_70_604 ();
 sg13g2_fill_2 FILLER_70_632 ();
 sg13g2_fill_1 FILLER_70_634 ();
 sg13g2_fill_1 FILLER_70_661 ();
 sg13g2_fill_1 FILLER_70_666 ();
 sg13g2_fill_2 FILLER_70_681 ();
 sg13g2_fill_1 FILLER_70_683 ();
 sg13g2_fill_1 FILLER_70_696 ();
 sg13g2_fill_1 FILLER_70_747 ();
 sg13g2_fill_1 FILLER_70_788 ();
 sg13g2_decap_8 FILLER_70_801 ();
 sg13g2_decap_8 FILLER_70_808 ();
 sg13g2_decap_8 FILLER_70_815 ();
 sg13g2_decap_8 FILLER_70_822 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_8 FILLER_70_836 ();
 sg13g2_decap_8 FILLER_70_843 ();
 sg13g2_decap_8 FILLER_70_850 ();
 sg13g2_decap_8 FILLER_70_857 ();
 sg13g2_decap_8 FILLER_70_864 ();
 sg13g2_decap_8 FILLER_70_871 ();
 sg13g2_decap_8 FILLER_70_878 ();
 sg13g2_decap_8 FILLER_70_885 ();
 sg13g2_decap_8 FILLER_70_892 ();
 sg13g2_decap_8 FILLER_70_899 ();
 sg13g2_decap_8 FILLER_70_906 ();
 sg13g2_decap_8 FILLER_70_913 ();
 sg13g2_decap_8 FILLER_70_920 ();
 sg13g2_decap_8 FILLER_70_927 ();
 sg13g2_decap_8 FILLER_70_934 ();
 sg13g2_decap_8 FILLER_70_941 ();
 sg13g2_decap_8 FILLER_70_948 ();
 sg13g2_decap_8 FILLER_70_955 ();
 sg13g2_decap_8 FILLER_70_962 ();
 sg13g2_decap_8 FILLER_70_969 ();
 sg13g2_decap_8 FILLER_70_976 ();
 sg13g2_decap_8 FILLER_70_983 ();
 sg13g2_decap_8 FILLER_70_990 ();
 sg13g2_decap_8 FILLER_70_997 ();
 sg13g2_decap_8 FILLER_70_1004 ();
 sg13g2_decap_8 FILLER_70_1011 ();
 sg13g2_decap_8 FILLER_70_1018 ();
 sg13g2_decap_8 FILLER_70_1025 ();
 sg13g2_decap_8 FILLER_70_1032 ();
 sg13g2_decap_8 FILLER_70_1039 ();
 sg13g2_decap_8 FILLER_70_1046 ();
 sg13g2_decap_8 FILLER_70_1053 ();
 sg13g2_decap_8 FILLER_70_1060 ();
 sg13g2_decap_8 FILLER_70_1067 ();
 sg13g2_decap_8 FILLER_70_1074 ();
 sg13g2_decap_8 FILLER_70_1081 ();
 sg13g2_decap_8 FILLER_70_1088 ();
 sg13g2_decap_8 FILLER_70_1095 ();
 sg13g2_decap_8 FILLER_70_1102 ();
 sg13g2_decap_8 FILLER_70_1109 ();
 sg13g2_decap_8 FILLER_70_1116 ();
 sg13g2_decap_8 FILLER_70_1123 ();
 sg13g2_decap_8 FILLER_70_1130 ();
 sg13g2_decap_8 FILLER_70_1137 ();
 sg13g2_decap_8 FILLER_70_1144 ();
 sg13g2_decap_8 FILLER_70_1151 ();
 sg13g2_decap_8 FILLER_70_1158 ();
 sg13g2_decap_8 FILLER_70_1165 ();
 sg13g2_decap_8 FILLER_70_1172 ();
 sg13g2_decap_8 FILLER_70_1179 ();
 sg13g2_decap_8 FILLER_70_1186 ();
 sg13g2_decap_8 FILLER_70_1193 ();
 sg13g2_decap_8 FILLER_70_1200 ();
 sg13g2_decap_8 FILLER_70_1207 ();
 sg13g2_decap_8 FILLER_70_1214 ();
 sg13g2_decap_8 FILLER_70_1221 ();
 sg13g2_decap_8 FILLER_70_1228 ();
 sg13g2_decap_8 FILLER_70_1235 ();
 sg13g2_decap_8 FILLER_70_1242 ();
 sg13g2_decap_8 FILLER_70_1249 ();
 sg13g2_decap_8 FILLER_70_1256 ();
 sg13g2_decap_8 FILLER_70_1263 ();
 sg13g2_decap_8 FILLER_70_1270 ();
 sg13g2_decap_8 FILLER_70_1277 ();
 sg13g2_decap_8 FILLER_70_1284 ();
 sg13g2_decap_8 FILLER_70_1291 ();
 sg13g2_decap_8 FILLER_70_1298 ();
 sg13g2_decap_8 FILLER_70_1305 ();
 sg13g2_decap_8 FILLER_70_1312 ();
 sg13g2_decap_8 FILLER_70_1319 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_6 ();
 sg13g2_fill_2 FILLER_71_20 ();
 sg13g2_fill_1 FILLER_71_22 ();
 sg13g2_fill_1 FILLER_71_32 ();
 sg13g2_fill_2 FILLER_71_38 ();
 sg13g2_fill_2 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_102 ();
 sg13g2_fill_2 FILLER_71_181 ();
 sg13g2_fill_1 FILLER_71_223 ();
 sg13g2_fill_2 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_284 ();
 sg13g2_fill_1 FILLER_71_352 ();
 sg13g2_fill_1 FILLER_71_450 ();
 sg13g2_fill_2 FILLER_71_547 ();
 sg13g2_fill_2 FILLER_71_601 ();
 sg13g2_fill_1 FILLER_71_705 ();
 sg13g2_decap_8 FILLER_71_810 ();
 sg13g2_decap_8 FILLER_71_817 ();
 sg13g2_decap_8 FILLER_71_824 ();
 sg13g2_decap_8 FILLER_71_831 ();
 sg13g2_decap_8 FILLER_71_838 ();
 sg13g2_decap_8 FILLER_71_845 ();
 sg13g2_decap_8 FILLER_71_852 ();
 sg13g2_decap_8 FILLER_71_859 ();
 sg13g2_decap_8 FILLER_71_866 ();
 sg13g2_decap_8 FILLER_71_873 ();
 sg13g2_decap_8 FILLER_71_880 ();
 sg13g2_decap_8 FILLER_71_887 ();
 sg13g2_decap_8 FILLER_71_894 ();
 sg13g2_decap_8 FILLER_71_901 ();
 sg13g2_decap_8 FILLER_71_908 ();
 sg13g2_decap_8 FILLER_71_915 ();
 sg13g2_decap_8 FILLER_71_922 ();
 sg13g2_decap_8 FILLER_71_929 ();
 sg13g2_decap_8 FILLER_71_936 ();
 sg13g2_decap_8 FILLER_71_943 ();
 sg13g2_decap_8 FILLER_71_950 ();
 sg13g2_decap_8 FILLER_71_957 ();
 sg13g2_decap_8 FILLER_71_964 ();
 sg13g2_decap_8 FILLER_71_971 ();
 sg13g2_decap_8 FILLER_71_978 ();
 sg13g2_decap_8 FILLER_71_985 ();
 sg13g2_decap_8 FILLER_71_992 ();
 sg13g2_decap_8 FILLER_71_999 ();
 sg13g2_decap_8 FILLER_71_1006 ();
 sg13g2_decap_8 FILLER_71_1013 ();
 sg13g2_decap_8 FILLER_71_1020 ();
 sg13g2_decap_8 FILLER_71_1027 ();
 sg13g2_decap_8 FILLER_71_1034 ();
 sg13g2_decap_8 FILLER_71_1041 ();
 sg13g2_decap_8 FILLER_71_1048 ();
 sg13g2_decap_8 FILLER_71_1055 ();
 sg13g2_decap_8 FILLER_71_1062 ();
 sg13g2_decap_8 FILLER_71_1069 ();
 sg13g2_decap_8 FILLER_71_1076 ();
 sg13g2_decap_8 FILLER_71_1083 ();
 sg13g2_decap_8 FILLER_71_1090 ();
 sg13g2_decap_8 FILLER_71_1097 ();
 sg13g2_decap_8 FILLER_71_1104 ();
 sg13g2_decap_8 FILLER_71_1111 ();
 sg13g2_decap_8 FILLER_71_1118 ();
 sg13g2_decap_8 FILLER_71_1125 ();
 sg13g2_decap_8 FILLER_71_1132 ();
 sg13g2_decap_8 FILLER_71_1139 ();
 sg13g2_decap_8 FILLER_71_1146 ();
 sg13g2_decap_8 FILLER_71_1153 ();
 sg13g2_decap_8 FILLER_71_1160 ();
 sg13g2_decap_8 FILLER_71_1167 ();
 sg13g2_decap_8 FILLER_71_1174 ();
 sg13g2_decap_8 FILLER_71_1181 ();
 sg13g2_decap_8 FILLER_71_1188 ();
 sg13g2_decap_8 FILLER_71_1195 ();
 sg13g2_decap_8 FILLER_71_1202 ();
 sg13g2_decap_8 FILLER_71_1209 ();
 sg13g2_decap_8 FILLER_71_1216 ();
 sg13g2_decap_8 FILLER_71_1223 ();
 sg13g2_decap_8 FILLER_71_1230 ();
 sg13g2_decap_8 FILLER_71_1237 ();
 sg13g2_decap_8 FILLER_71_1244 ();
 sg13g2_decap_8 FILLER_71_1251 ();
 sg13g2_decap_8 FILLER_71_1258 ();
 sg13g2_decap_8 FILLER_71_1265 ();
 sg13g2_decap_8 FILLER_71_1272 ();
 sg13g2_decap_8 FILLER_71_1279 ();
 sg13g2_decap_8 FILLER_71_1286 ();
 sg13g2_decap_8 FILLER_71_1293 ();
 sg13g2_decap_8 FILLER_71_1300 ();
 sg13g2_decap_8 FILLER_71_1307 ();
 sg13g2_decap_8 FILLER_71_1314 ();
 sg13g2_decap_4 FILLER_71_1321 ();
 sg13g2_fill_1 FILLER_71_1325 ();
 sg13g2_fill_2 FILLER_72_4 ();
 sg13g2_fill_1 FILLER_72_80 ();
 sg13g2_fill_2 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_189 ();
 sg13g2_fill_1 FILLER_72_310 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_fill_1 FILLER_72_348 ();
 sg13g2_fill_2 FILLER_72_359 ();
 sg13g2_fill_2 FILLER_72_371 ();
 sg13g2_fill_2 FILLER_72_383 ();
 sg13g2_fill_1 FILLER_72_439 ();
 sg13g2_fill_1 FILLER_72_466 ();
 sg13g2_fill_1 FILLER_72_472 ();
 sg13g2_fill_1 FILLER_72_499 ();
 sg13g2_fill_2 FILLER_72_580 ();
 sg13g2_fill_2 FILLER_72_680 ();
 sg13g2_fill_1 FILLER_72_764 ();
 sg13g2_decap_8 FILLER_72_801 ();
 sg13g2_decap_8 FILLER_72_808 ();
 sg13g2_decap_8 FILLER_72_815 ();
 sg13g2_decap_8 FILLER_72_822 ();
 sg13g2_decap_8 FILLER_72_829 ();
 sg13g2_decap_8 FILLER_72_836 ();
 sg13g2_decap_8 FILLER_72_843 ();
 sg13g2_decap_8 FILLER_72_850 ();
 sg13g2_decap_8 FILLER_72_857 ();
 sg13g2_decap_8 FILLER_72_864 ();
 sg13g2_decap_8 FILLER_72_871 ();
 sg13g2_decap_8 FILLER_72_878 ();
 sg13g2_decap_8 FILLER_72_885 ();
 sg13g2_decap_8 FILLER_72_892 ();
 sg13g2_decap_8 FILLER_72_899 ();
 sg13g2_decap_8 FILLER_72_906 ();
 sg13g2_decap_8 FILLER_72_913 ();
 sg13g2_decap_8 FILLER_72_920 ();
 sg13g2_decap_8 FILLER_72_927 ();
 sg13g2_decap_8 FILLER_72_934 ();
 sg13g2_decap_8 FILLER_72_941 ();
 sg13g2_decap_8 FILLER_72_948 ();
 sg13g2_decap_8 FILLER_72_955 ();
 sg13g2_decap_8 FILLER_72_962 ();
 sg13g2_decap_8 FILLER_72_969 ();
 sg13g2_decap_8 FILLER_72_976 ();
 sg13g2_decap_8 FILLER_72_983 ();
 sg13g2_decap_8 FILLER_72_990 ();
 sg13g2_decap_8 FILLER_72_997 ();
 sg13g2_decap_8 FILLER_72_1004 ();
 sg13g2_decap_8 FILLER_72_1011 ();
 sg13g2_decap_8 FILLER_72_1018 ();
 sg13g2_decap_8 FILLER_72_1025 ();
 sg13g2_decap_8 FILLER_72_1032 ();
 sg13g2_decap_8 FILLER_72_1039 ();
 sg13g2_decap_8 FILLER_72_1046 ();
 sg13g2_decap_8 FILLER_72_1053 ();
 sg13g2_decap_8 FILLER_72_1060 ();
 sg13g2_decap_8 FILLER_72_1067 ();
 sg13g2_decap_8 FILLER_72_1074 ();
 sg13g2_decap_8 FILLER_72_1081 ();
 sg13g2_decap_8 FILLER_72_1088 ();
 sg13g2_decap_8 FILLER_72_1095 ();
 sg13g2_decap_8 FILLER_72_1102 ();
 sg13g2_decap_8 FILLER_72_1109 ();
 sg13g2_decap_8 FILLER_72_1116 ();
 sg13g2_decap_8 FILLER_72_1123 ();
 sg13g2_decap_8 FILLER_72_1130 ();
 sg13g2_decap_8 FILLER_72_1137 ();
 sg13g2_decap_8 FILLER_72_1144 ();
 sg13g2_decap_8 FILLER_72_1151 ();
 sg13g2_decap_8 FILLER_72_1158 ();
 sg13g2_decap_8 FILLER_72_1165 ();
 sg13g2_decap_8 FILLER_72_1172 ();
 sg13g2_decap_8 FILLER_72_1179 ();
 sg13g2_decap_8 FILLER_72_1186 ();
 sg13g2_decap_8 FILLER_72_1193 ();
 sg13g2_decap_8 FILLER_72_1200 ();
 sg13g2_decap_8 FILLER_72_1207 ();
 sg13g2_decap_8 FILLER_72_1214 ();
 sg13g2_decap_8 FILLER_72_1221 ();
 sg13g2_decap_8 FILLER_72_1228 ();
 sg13g2_decap_8 FILLER_72_1235 ();
 sg13g2_decap_8 FILLER_72_1242 ();
 sg13g2_decap_8 FILLER_72_1249 ();
 sg13g2_decap_8 FILLER_72_1256 ();
 sg13g2_decap_8 FILLER_72_1263 ();
 sg13g2_decap_8 FILLER_72_1270 ();
 sg13g2_decap_8 FILLER_72_1277 ();
 sg13g2_decap_8 FILLER_72_1284 ();
 sg13g2_decap_8 FILLER_72_1291 ();
 sg13g2_decap_8 FILLER_72_1298 ();
 sg13g2_decap_8 FILLER_72_1305 ();
 sg13g2_decap_8 FILLER_72_1312 ();
 sg13g2_decap_8 FILLER_72_1319 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_1 FILLER_73_24 ();
 sg13g2_fill_2 FILLER_73_38 ();
 sg13g2_fill_1 FILLER_73_101 ();
 sg13g2_fill_1 FILLER_73_117 ();
 sg13g2_fill_1 FILLER_73_164 ();
 sg13g2_fill_2 FILLER_73_222 ();
 sg13g2_fill_1 FILLER_73_254 ();
 sg13g2_fill_2 FILLER_73_267 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_354 ();
 sg13g2_fill_1 FILLER_73_381 ();
 sg13g2_fill_1 FILLER_73_418 ();
 sg13g2_fill_2 FILLER_73_508 ();
 sg13g2_fill_1 FILLER_73_510 ();
 sg13g2_fill_2 FILLER_73_535 ();
 sg13g2_fill_2 FILLER_73_611 ();
 sg13g2_fill_2 FILLER_73_639 ();
 sg13g2_fill_1 FILLER_73_641 ();
 sg13g2_fill_1 FILLER_73_720 ();
 sg13g2_fill_2 FILLER_73_751 ();
 sg13g2_fill_1 FILLER_73_763 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_8 FILLER_73_857 ();
 sg13g2_decap_8 FILLER_73_864 ();
 sg13g2_decap_8 FILLER_73_871 ();
 sg13g2_decap_8 FILLER_73_878 ();
 sg13g2_decap_8 FILLER_73_885 ();
 sg13g2_decap_8 FILLER_73_892 ();
 sg13g2_decap_8 FILLER_73_899 ();
 sg13g2_decap_8 FILLER_73_906 ();
 sg13g2_decap_8 FILLER_73_913 ();
 sg13g2_decap_8 FILLER_73_920 ();
 sg13g2_decap_8 FILLER_73_927 ();
 sg13g2_decap_8 FILLER_73_934 ();
 sg13g2_decap_8 FILLER_73_941 ();
 sg13g2_decap_8 FILLER_73_948 ();
 sg13g2_decap_8 FILLER_73_955 ();
 sg13g2_decap_8 FILLER_73_962 ();
 sg13g2_decap_8 FILLER_73_969 ();
 sg13g2_decap_8 FILLER_73_976 ();
 sg13g2_decap_8 FILLER_73_983 ();
 sg13g2_decap_8 FILLER_73_990 ();
 sg13g2_decap_8 FILLER_73_997 ();
 sg13g2_decap_8 FILLER_73_1004 ();
 sg13g2_decap_8 FILLER_73_1011 ();
 sg13g2_decap_8 FILLER_73_1018 ();
 sg13g2_decap_8 FILLER_73_1025 ();
 sg13g2_decap_8 FILLER_73_1032 ();
 sg13g2_decap_8 FILLER_73_1039 ();
 sg13g2_decap_8 FILLER_73_1046 ();
 sg13g2_decap_8 FILLER_73_1053 ();
 sg13g2_decap_8 FILLER_73_1060 ();
 sg13g2_decap_8 FILLER_73_1067 ();
 sg13g2_decap_8 FILLER_73_1074 ();
 sg13g2_decap_8 FILLER_73_1081 ();
 sg13g2_decap_8 FILLER_73_1088 ();
 sg13g2_decap_8 FILLER_73_1095 ();
 sg13g2_decap_8 FILLER_73_1102 ();
 sg13g2_decap_8 FILLER_73_1109 ();
 sg13g2_decap_8 FILLER_73_1116 ();
 sg13g2_decap_8 FILLER_73_1123 ();
 sg13g2_decap_8 FILLER_73_1130 ();
 sg13g2_decap_8 FILLER_73_1137 ();
 sg13g2_decap_8 FILLER_73_1144 ();
 sg13g2_decap_8 FILLER_73_1151 ();
 sg13g2_decap_8 FILLER_73_1158 ();
 sg13g2_decap_8 FILLER_73_1165 ();
 sg13g2_decap_8 FILLER_73_1172 ();
 sg13g2_decap_8 FILLER_73_1179 ();
 sg13g2_decap_8 FILLER_73_1186 ();
 sg13g2_decap_8 FILLER_73_1193 ();
 sg13g2_decap_8 FILLER_73_1200 ();
 sg13g2_decap_8 FILLER_73_1207 ();
 sg13g2_decap_8 FILLER_73_1214 ();
 sg13g2_decap_8 FILLER_73_1221 ();
 sg13g2_decap_8 FILLER_73_1228 ();
 sg13g2_decap_8 FILLER_73_1235 ();
 sg13g2_decap_8 FILLER_73_1242 ();
 sg13g2_decap_8 FILLER_73_1249 ();
 sg13g2_decap_8 FILLER_73_1256 ();
 sg13g2_decap_8 FILLER_73_1263 ();
 sg13g2_decap_8 FILLER_73_1270 ();
 sg13g2_decap_8 FILLER_73_1277 ();
 sg13g2_decap_8 FILLER_73_1284 ();
 sg13g2_decap_8 FILLER_73_1291 ();
 sg13g2_decap_8 FILLER_73_1298 ();
 sg13g2_decap_8 FILLER_73_1305 ();
 sg13g2_decap_8 FILLER_73_1312 ();
 sg13g2_decap_8 FILLER_73_1319 ();
 sg13g2_fill_2 FILLER_74_8 ();
 sg13g2_fill_1 FILLER_74_18 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_74 ();
 sg13g2_fill_1 FILLER_74_110 ();
 sg13g2_fill_2 FILLER_74_149 ();
 sg13g2_fill_1 FILLER_74_312 ();
 sg13g2_fill_1 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_440 ();
 sg13g2_fill_1 FILLER_74_467 ();
 sg13g2_fill_2 FILLER_74_498 ();
 sg13g2_fill_1 FILLER_74_564 ();
 sg13g2_fill_2 FILLER_74_575 ();
 sg13g2_fill_2 FILLER_74_661 ();
 sg13g2_fill_1 FILLER_74_673 ();
 sg13g2_fill_2 FILLER_74_704 ();
 sg13g2_fill_1 FILLER_74_716 ();
 sg13g2_fill_1 FILLER_74_727 ();
 sg13g2_fill_2 FILLER_74_742 ();
 sg13g2_fill_2 FILLER_74_788 ();
 sg13g2_decap_8 FILLER_74_801 ();
 sg13g2_decap_8 FILLER_74_808 ();
 sg13g2_decap_8 FILLER_74_815 ();
 sg13g2_decap_8 FILLER_74_822 ();
 sg13g2_decap_8 FILLER_74_829 ();
 sg13g2_decap_8 FILLER_74_836 ();
 sg13g2_decap_8 FILLER_74_843 ();
 sg13g2_decap_8 FILLER_74_850 ();
 sg13g2_decap_8 FILLER_74_857 ();
 sg13g2_decap_8 FILLER_74_864 ();
 sg13g2_decap_8 FILLER_74_871 ();
 sg13g2_decap_8 FILLER_74_878 ();
 sg13g2_decap_8 FILLER_74_885 ();
 sg13g2_decap_8 FILLER_74_892 ();
 sg13g2_decap_8 FILLER_74_899 ();
 sg13g2_decap_8 FILLER_74_906 ();
 sg13g2_decap_8 FILLER_74_913 ();
 sg13g2_decap_8 FILLER_74_920 ();
 sg13g2_decap_8 FILLER_74_927 ();
 sg13g2_decap_8 FILLER_74_934 ();
 sg13g2_decap_8 FILLER_74_941 ();
 sg13g2_decap_8 FILLER_74_948 ();
 sg13g2_decap_8 FILLER_74_955 ();
 sg13g2_decap_8 FILLER_74_962 ();
 sg13g2_decap_8 FILLER_74_969 ();
 sg13g2_decap_8 FILLER_74_976 ();
 sg13g2_decap_8 FILLER_74_983 ();
 sg13g2_decap_8 FILLER_74_990 ();
 sg13g2_decap_8 FILLER_74_997 ();
 sg13g2_decap_8 FILLER_74_1004 ();
 sg13g2_decap_8 FILLER_74_1011 ();
 sg13g2_decap_8 FILLER_74_1018 ();
 sg13g2_decap_8 FILLER_74_1025 ();
 sg13g2_decap_8 FILLER_74_1032 ();
 sg13g2_decap_8 FILLER_74_1039 ();
 sg13g2_decap_8 FILLER_74_1046 ();
 sg13g2_decap_8 FILLER_74_1053 ();
 sg13g2_decap_8 FILLER_74_1060 ();
 sg13g2_decap_8 FILLER_74_1067 ();
 sg13g2_decap_8 FILLER_74_1074 ();
 sg13g2_decap_8 FILLER_74_1081 ();
 sg13g2_decap_8 FILLER_74_1088 ();
 sg13g2_decap_8 FILLER_74_1095 ();
 sg13g2_decap_8 FILLER_74_1102 ();
 sg13g2_decap_8 FILLER_74_1109 ();
 sg13g2_decap_8 FILLER_74_1116 ();
 sg13g2_decap_8 FILLER_74_1123 ();
 sg13g2_decap_8 FILLER_74_1130 ();
 sg13g2_decap_8 FILLER_74_1137 ();
 sg13g2_decap_8 FILLER_74_1144 ();
 sg13g2_decap_8 FILLER_74_1151 ();
 sg13g2_decap_8 FILLER_74_1158 ();
 sg13g2_decap_8 FILLER_74_1165 ();
 sg13g2_decap_8 FILLER_74_1172 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_decap_8 FILLER_74_1186 ();
 sg13g2_decap_8 FILLER_74_1193 ();
 sg13g2_decap_8 FILLER_74_1200 ();
 sg13g2_decap_8 FILLER_74_1207 ();
 sg13g2_decap_8 FILLER_74_1214 ();
 sg13g2_decap_8 FILLER_74_1221 ();
 sg13g2_decap_8 FILLER_74_1228 ();
 sg13g2_decap_8 FILLER_74_1235 ();
 sg13g2_decap_8 FILLER_74_1242 ();
 sg13g2_decap_8 FILLER_74_1249 ();
 sg13g2_decap_8 FILLER_74_1256 ();
 sg13g2_decap_8 FILLER_74_1263 ();
 sg13g2_decap_8 FILLER_74_1270 ();
 sg13g2_decap_8 FILLER_74_1277 ();
 sg13g2_decap_8 FILLER_74_1284 ();
 sg13g2_decap_8 FILLER_74_1291 ();
 sg13g2_decap_8 FILLER_74_1298 ();
 sg13g2_decap_8 FILLER_74_1305 ();
 sg13g2_decap_8 FILLER_74_1312 ();
 sg13g2_decap_8 FILLER_74_1319 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_4 ();
 sg13g2_decap_8 FILLER_75_10 ();
 sg13g2_decap_8 FILLER_75_17 ();
 sg13g2_decap_4 FILLER_75_24 ();
 sg13g2_fill_2 FILLER_75_69 ();
 sg13g2_fill_2 FILLER_75_80 ();
 sg13g2_fill_1 FILLER_75_91 ();
 sg13g2_fill_1 FILLER_75_107 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_269 ();
 sg13g2_fill_2 FILLER_75_284 ();
 sg13g2_fill_2 FILLER_75_299 ();
 sg13g2_fill_2 FILLER_75_337 ();
 sg13g2_fill_1 FILLER_75_363 ();
 sg13g2_fill_1 FILLER_75_383 ();
 sg13g2_fill_1 FILLER_75_432 ();
 sg13g2_fill_1 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_454 ();
 sg13g2_fill_1 FILLER_75_465 ();
 sg13g2_fill_1 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_511 ();
 sg13g2_fill_1 FILLER_75_595 ();
 sg13g2_fill_1 FILLER_75_664 ();
 sg13g2_fill_2 FILLER_75_695 ();
 sg13g2_fill_1 FILLER_75_711 ();
 sg13g2_fill_2 FILLER_75_756 ();
 sg13g2_fill_2 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_decap_8 FILLER_75_859 ();
 sg13g2_decap_8 FILLER_75_866 ();
 sg13g2_decap_8 FILLER_75_873 ();
 sg13g2_decap_8 FILLER_75_880 ();
 sg13g2_decap_8 FILLER_75_887 ();
 sg13g2_decap_8 FILLER_75_894 ();
 sg13g2_decap_8 FILLER_75_901 ();
 sg13g2_decap_8 FILLER_75_908 ();
 sg13g2_decap_8 FILLER_75_915 ();
 sg13g2_decap_8 FILLER_75_922 ();
 sg13g2_decap_8 FILLER_75_929 ();
 sg13g2_decap_8 FILLER_75_936 ();
 sg13g2_decap_8 FILLER_75_943 ();
 sg13g2_decap_8 FILLER_75_950 ();
 sg13g2_decap_8 FILLER_75_957 ();
 sg13g2_decap_8 FILLER_75_964 ();
 sg13g2_decap_8 FILLER_75_971 ();
 sg13g2_decap_8 FILLER_75_978 ();
 sg13g2_decap_8 FILLER_75_985 ();
 sg13g2_decap_8 FILLER_75_992 ();
 sg13g2_decap_8 FILLER_75_999 ();
 sg13g2_decap_8 FILLER_75_1006 ();
 sg13g2_decap_8 FILLER_75_1013 ();
 sg13g2_decap_8 FILLER_75_1020 ();
 sg13g2_decap_8 FILLER_75_1027 ();
 sg13g2_decap_8 FILLER_75_1034 ();
 sg13g2_decap_8 FILLER_75_1041 ();
 sg13g2_decap_8 FILLER_75_1048 ();
 sg13g2_decap_8 FILLER_75_1055 ();
 sg13g2_decap_8 FILLER_75_1062 ();
 sg13g2_decap_8 FILLER_75_1069 ();
 sg13g2_decap_8 FILLER_75_1076 ();
 sg13g2_decap_8 FILLER_75_1083 ();
 sg13g2_decap_8 FILLER_75_1090 ();
 sg13g2_decap_8 FILLER_75_1097 ();
 sg13g2_decap_8 FILLER_75_1104 ();
 sg13g2_decap_8 FILLER_75_1111 ();
 sg13g2_decap_8 FILLER_75_1118 ();
 sg13g2_decap_8 FILLER_75_1125 ();
 sg13g2_decap_8 FILLER_75_1132 ();
 sg13g2_decap_8 FILLER_75_1139 ();
 sg13g2_decap_8 FILLER_75_1146 ();
 sg13g2_decap_8 FILLER_75_1153 ();
 sg13g2_decap_8 FILLER_75_1160 ();
 sg13g2_decap_8 FILLER_75_1167 ();
 sg13g2_decap_8 FILLER_75_1174 ();
 sg13g2_decap_8 FILLER_75_1181 ();
 sg13g2_decap_8 FILLER_75_1188 ();
 sg13g2_decap_8 FILLER_75_1195 ();
 sg13g2_decap_8 FILLER_75_1202 ();
 sg13g2_decap_8 FILLER_75_1209 ();
 sg13g2_decap_8 FILLER_75_1216 ();
 sg13g2_decap_8 FILLER_75_1223 ();
 sg13g2_decap_8 FILLER_75_1230 ();
 sg13g2_decap_8 FILLER_75_1237 ();
 sg13g2_decap_8 FILLER_75_1244 ();
 sg13g2_decap_8 FILLER_75_1251 ();
 sg13g2_decap_8 FILLER_75_1258 ();
 sg13g2_decap_8 FILLER_75_1265 ();
 sg13g2_decap_8 FILLER_75_1272 ();
 sg13g2_decap_8 FILLER_75_1279 ();
 sg13g2_decap_8 FILLER_75_1286 ();
 sg13g2_decap_8 FILLER_75_1293 ();
 sg13g2_decap_8 FILLER_75_1300 ();
 sg13g2_decap_8 FILLER_75_1307 ();
 sg13g2_decap_8 FILLER_75_1314 ();
 sg13g2_decap_4 FILLER_75_1321 ();
 sg13g2_fill_1 FILLER_75_1325 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_4 FILLER_76_35 ();
 sg13g2_fill_1 FILLER_76_39 ();
 sg13g2_fill_2 FILLER_76_52 ();
 sg13g2_fill_2 FILLER_76_101 ();
 sg13g2_fill_2 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_125 ();
 sg13g2_fill_2 FILLER_76_225 ();
 sg13g2_fill_1 FILLER_76_255 ();
 sg13g2_fill_2 FILLER_76_376 ();
 sg13g2_fill_1 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_76_466 ();
 sg13g2_fill_2 FILLER_76_498 ();
 sg13g2_fill_1 FILLER_76_514 ();
 sg13g2_fill_2 FILLER_76_597 ();
 sg13g2_fill_1 FILLER_76_609 ();
 sg13g2_fill_2 FILLER_76_641 ();
 sg13g2_fill_1 FILLER_76_653 ();
 sg13g2_fill_1 FILLER_76_684 ();
 sg13g2_fill_1 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_761 ();
 sg13g2_fill_1 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_782 ();
 sg13g2_decap_8 FILLER_76_815 ();
 sg13g2_decap_8 FILLER_76_822 ();
 sg13g2_decap_8 FILLER_76_829 ();
 sg13g2_decap_8 FILLER_76_836 ();
 sg13g2_decap_8 FILLER_76_843 ();
 sg13g2_decap_8 FILLER_76_850 ();
 sg13g2_decap_8 FILLER_76_857 ();
 sg13g2_decap_8 FILLER_76_864 ();
 sg13g2_decap_8 FILLER_76_871 ();
 sg13g2_decap_8 FILLER_76_878 ();
 sg13g2_decap_8 FILLER_76_885 ();
 sg13g2_decap_8 FILLER_76_892 ();
 sg13g2_decap_8 FILLER_76_899 ();
 sg13g2_decap_8 FILLER_76_906 ();
 sg13g2_decap_8 FILLER_76_913 ();
 sg13g2_decap_8 FILLER_76_920 ();
 sg13g2_decap_8 FILLER_76_927 ();
 sg13g2_decap_8 FILLER_76_934 ();
 sg13g2_decap_8 FILLER_76_941 ();
 sg13g2_decap_8 FILLER_76_948 ();
 sg13g2_decap_8 FILLER_76_955 ();
 sg13g2_decap_8 FILLER_76_962 ();
 sg13g2_decap_8 FILLER_76_969 ();
 sg13g2_decap_8 FILLER_76_976 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_decap_8 FILLER_76_990 ();
 sg13g2_decap_8 FILLER_76_997 ();
 sg13g2_decap_8 FILLER_76_1004 ();
 sg13g2_decap_8 FILLER_76_1011 ();
 sg13g2_decap_8 FILLER_76_1018 ();
 sg13g2_decap_8 FILLER_76_1025 ();
 sg13g2_decap_8 FILLER_76_1032 ();
 sg13g2_decap_8 FILLER_76_1039 ();
 sg13g2_decap_8 FILLER_76_1046 ();
 sg13g2_decap_8 FILLER_76_1053 ();
 sg13g2_decap_8 FILLER_76_1060 ();
 sg13g2_decap_8 FILLER_76_1067 ();
 sg13g2_decap_8 FILLER_76_1074 ();
 sg13g2_decap_8 FILLER_76_1081 ();
 sg13g2_decap_8 FILLER_76_1088 ();
 sg13g2_decap_8 FILLER_76_1095 ();
 sg13g2_decap_8 FILLER_76_1102 ();
 sg13g2_decap_8 FILLER_76_1109 ();
 sg13g2_decap_8 FILLER_76_1116 ();
 sg13g2_decap_8 FILLER_76_1123 ();
 sg13g2_decap_8 FILLER_76_1130 ();
 sg13g2_decap_8 FILLER_76_1137 ();
 sg13g2_decap_8 FILLER_76_1144 ();
 sg13g2_decap_8 FILLER_76_1151 ();
 sg13g2_decap_8 FILLER_76_1158 ();
 sg13g2_decap_8 FILLER_76_1165 ();
 sg13g2_decap_8 FILLER_76_1172 ();
 sg13g2_decap_8 FILLER_76_1179 ();
 sg13g2_decap_8 FILLER_76_1186 ();
 sg13g2_decap_8 FILLER_76_1193 ();
 sg13g2_decap_8 FILLER_76_1200 ();
 sg13g2_decap_8 FILLER_76_1207 ();
 sg13g2_decap_8 FILLER_76_1214 ();
 sg13g2_decap_8 FILLER_76_1221 ();
 sg13g2_decap_8 FILLER_76_1228 ();
 sg13g2_decap_8 FILLER_76_1235 ();
 sg13g2_decap_8 FILLER_76_1242 ();
 sg13g2_decap_8 FILLER_76_1249 ();
 sg13g2_decap_8 FILLER_76_1256 ();
 sg13g2_decap_8 FILLER_76_1263 ();
 sg13g2_decap_8 FILLER_76_1270 ();
 sg13g2_decap_8 FILLER_76_1277 ();
 sg13g2_decap_8 FILLER_76_1284 ();
 sg13g2_decap_8 FILLER_76_1291 ();
 sg13g2_decap_8 FILLER_76_1298 ();
 sg13g2_decap_8 FILLER_76_1305 ();
 sg13g2_decap_8 FILLER_76_1312 ();
 sg13g2_decap_8 FILLER_76_1319 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_fill_2 FILLER_77_42 ();
 sg13g2_fill_1 FILLER_77_143 ();
 sg13g2_fill_2 FILLER_77_178 ();
 sg13g2_fill_1 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_207 ();
 sg13g2_fill_2 FILLER_77_217 ();
 sg13g2_fill_1 FILLER_77_265 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_308 ();
 sg13g2_fill_2 FILLER_77_314 ();
 sg13g2_fill_1 FILLER_77_352 ();
 sg13g2_fill_2 FILLER_77_439 ();
 sg13g2_fill_2 FILLER_77_631 ();
 sg13g2_fill_2 FILLER_77_643 ();
 sg13g2_fill_1 FILLER_77_645 ();
 sg13g2_fill_2 FILLER_77_660 ();
 sg13g2_fill_1 FILLER_77_662 ();
 sg13g2_fill_2 FILLER_77_671 ();
 sg13g2_fill_1 FILLER_77_673 ();
 sg13g2_fill_1 FILLER_77_704 ();
 sg13g2_fill_1 FILLER_77_715 ();
 sg13g2_fill_1 FILLER_77_726 ();
 sg13g2_fill_1 FILLER_77_737 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_fill_2 FILLER_77_791 ();
 sg13g2_fill_1 FILLER_77_793 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_decap_8 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_77_868 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_decap_8 FILLER_77_882 ();
 sg13g2_decap_8 FILLER_77_889 ();
 sg13g2_decap_8 FILLER_77_896 ();
 sg13g2_decap_8 FILLER_77_903 ();
 sg13g2_decap_8 FILLER_77_910 ();
 sg13g2_decap_8 FILLER_77_917 ();
 sg13g2_decap_8 FILLER_77_924 ();
 sg13g2_decap_8 FILLER_77_931 ();
 sg13g2_decap_8 FILLER_77_938 ();
 sg13g2_decap_8 FILLER_77_945 ();
 sg13g2_decap_8 FILLER_77_952 ();
 sg13g2_decap_8 FILLER_77_959 ();
 sg13g2_decap_8 FILLER_77_966 ();
 sg13g2_decap_8 FILLER_77_973 ();
 sg13g2_decap_8 FILLER_77_980 ();
 sg13g2_decap_8 FILLER_77_987 ();
 sg13g2_decap_8 FILLER_77_994 ();
 sg13g2_decap_8 FILLER_77_1001 ();
 sg13g2_decap_8 FILLER_77_1008 ();
 sg13g2_decap_8 FILLER_77_1015 ();
 sg13g2_decap_8 FILLER_77_1022 ();
 sg13g2_decap_8 FILLER_77_1029 ();
 sg13g2_decap_8 FILLER_77_1036 ();
 sg13g2_decap_8 FILLER_77_1043 ();
 sg13g2_decap_8 FILLER_77_1050 ();
 sg13g2_decap_8 FILLER_77_1057 ();
 sg13g2_decap_8 FILLER_77_1064 ();
 sg13g2_decap_8 FILLER_77_1071 ();
 sg13g2_decap_8 FILLER_77_1078 ();
 sg13g2_decap_8 FILLER_77_1085 ();
 sg13g2_decap_8 FILLER_77_1092 ();
 sg13g2_decap_8 FILLER_77_1099 ();
 sg13g2_decap_8 FILLER_77_1106 ();
 sg13g2_decap_8 FILLER_77_1113 ();
 sg13g2_decap_8 FILLER_77_1120 ();
 sg13g2_decap_8 FILLER_77_1127 ();
 sg13g2_decap_8 FILLER_77_1134 ();
 sg13g2_decap_8 FILLER_77_1141 ();
 sg13g2_decap_8 FILLER_77_1148 ();
 sg13g2_decap_8 FILLER_77_1155 ();
 sg13g2_decap_8 FILLER_77_1162 ();
 sg13g2_decap_8 FILLER_77_1169 ();
 sg13g2_decap_8 FILLER_77_1176 ();
 sg13g2_decap_8 FILLER_77_1183 ();
 sg13g2_decap_8 FILLER_77_1190 ();
 sg13g2_decap_8 FILLER_77_1197 ();
 sg13g2_decap_8 FILLER_77_1204 ();
 sg13g2_decap_8 FILLER_77_1211 ();
 sg13g2_decap_8 FILLER_77_1218 ();
 sg13g2_decap_8 FILLER_77_1225 ();
 sg13g2_decap_8 FILLER_77_1232 ();
 sg13g2_decap_8 FILLER_77_1239 ();
 sg13g2_decap_8 FILLER_77_1246 ();
 sg13g2_decap_8 FILLER_77_1253 ();
 sg13g2_decap_8 FILLER_77_1260 ();
 sg13g2_decap_8 FILLER_77_1267 ();
 sg13g2_decap_8 FILLER_77_1274 ();
 sg13g2_decap_8 FILLER_77_1281 ();
 sg13g2_decap_8 FILLER_77_1288 ();
 sg13g2_decap_8 FILLER_77_1295 ();
 sg13g2_decap_8 FILLER_77_1302 ();
 sg13g2_decap_8 FILLER_77_1309 ();
 sg13g2_decap_8 FILLER_77_1316 ();
 sg13g2_fill_2 FILLER_77_1323 ();
 sg13g2_fill_1 FILLER_77_1325 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_35 ();
 sg13g2_fill_2 FILLER_78_103 ();
 sg13g2_fill_1 FILLER_78_131 ();
 sg13g2_fill_2 FILLER_78_166 ();
 sg13g2_fill_1 FILLER_78_168 ();
 sg13g2_fill_2 FILLER_78_293 ();
 sg13g2_fill_2 FILLER_78_398 ();
 sg13g2_fill_2 FILLER_78_450 ();
 sg13g2_fill_1 FILLER_78_452 ();
 sg13g2_fill_2 FILLER_78_497 ();
 sg13g2_fill_2 FILLER_78_583 ();
 sg13g2_fill_1 FILLER_78_615 ();
 sg13g2_fill_2 FILLER_78_620 ();
 sg13g2_fill_2 FILLER_78_648 ();
 sg13g2_fill_2 FILLER_78_762 ();
 sg13g2_fill_1 FILLER_78_764 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_decap_8 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_78_847 ();
 sg13g2_decap_8 FILLER_78_854 ();
 sg13g2_decap_8 FILLER_78_861 ();
 sg13g2_decap_8 FILLER_78_868 ();
 sg13g2_decap_8 FILLER_78_875 ();
 sg13g2_decap_8 FILLER_78_882 ();
 sg13g2_decap_8 FILLER_78_889 ();
 sg13g2_decap_8 FILLER_78_896 ();
 sg13g2_decap_8 FILLER_78_903 ();
 sg13g2_decap_8 FILLER_78_910 ();
 sg13g2_decap_8 FILLER_78_917 ();
 sg13g2_decap_8 FILLER_78_924 ();
 sg13g2_decap_8 FILLER_78_931 ();
 sg13g2_decap_8 FILLER_78_938 ();
 sg13g2_decap_8 FILLER_78_945 ();
 sg13g2_decap_8 FILLER_78_952 ();
 sg13g2_decap_8 FILLER_78_959 ();
 sg13g2_decap_8 FILLER_78_966 ();
 sg13g2_decap_8 FILLER_78_973 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_decap_8 FILLER_78_987 ();
 sg13g2_decap_8 FILLER_78_994 ();
 sg13g2_decap_8 FILLER_78_1001 ();
 sg13g2_decap_8 FILLER_78_1008 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_decap_8 FILLER_78_1022 ();
 sg13g2_decap_8 FILLER_78_1029 ();
 sg13g2_decap_8 FILLER_78_1036 ();
 sg13g2_decap_8 FILLER_78_1043 ();
 sg13g2_decap_8 FILLER_78_1050 ();
 sg13g2_decap_8 FILLER_78_1057 ();
 sg13g2_decap_8 FILLER_78_1064 ();
 sg13g2_decap_8 FILLER_78_1071 ();
 sg13g2_decap_8 FILLER_78_1078 ();
 sg13g2_decap_8 FILLER_78_1085 ();
 sg13g2_decap_8 FILLER_78_1092 ();
 sg13g2_decap_8 FILLER_78_1099 ();
 sg13g2_decap_8 FILLER_78_1106 ();
 sg13g2_decap_8 FILLER_78_1113 ();
 sg13g2_decap_8 FILLER_78_1120 ();
 sg13g2_decap_8 FILLER_78_1127 ();
 sg13g2_decap_8 FILLER_78_1134 ();
 sg13g2_decap_8 FILLER_78_1141 ();
 sg13g2_decap_8 FILLER_78_1148 ();
 sg13g2_decap_8 FILLER_78_1155 ();
 sg13g2_decap_8 FILLER_78_1162 ();
 sg13g2_decap_8 FILLER_78_1169 ();
 sg13g2_decap_8 FILLER_78_1176 ();
 sg13g2_decap_8 FILLER_78_1183 ();
 sg13g2_decap_8 FILLER_78_1190 ();
 sg13g2_decap_8 FILLER_78_1197 ();
 sg13g2_decap_8 FILLER_78_1204 ();
 sg13g2_decap_8 FILLER_78_1211 ();
 sg13g2_decap_8 FILLER_78_1218 ();
 sg13g2_decap_8 FILLER_78_1225 ();
 sg13g2_decap_8 FILLER_78_1232 ();
 sg13g2_decap_8 FILLER_78_1239 ();
 sg13g2_decap_8 FILLER_78_1246 ();
 sg13g2_decap_8 FILLER_78_1253 ();
 sg13g2_decap_8 FILLER_78_1260 ();
 sg13g2_decap_8 FILLER_78_1267 ();
 sg13g2_decap_8 FILLER_78_1274 ();
 sg13g2_decap_8 FILLER_78_1281 ();
 sg13g2_decap_8 FILLER_78_1288 ();
 sg13g2_decap_8 FILLER_78_1295 ();
 sg13g2_decap_8 FILLER_78_1302 ();
 sg13g2_decap_8 FILLER_78_1309 ();
 sg13g2_decap_8 FILLER_78_1316 ();
 sg13g2_fill_2 FILLER_78_1323 ();
 sg13g2_fill_1 FILLER_78_1325 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_28 ();
 sg13g2_fill_1 FILLER_79_30 ();
 sg13g2_fill_2 FILLER_79_276 ();
 sg13g2_fill_2 FILLER_79_326 ();
 sg13g2_fill_1 FILLER_79_328 ();
 sg13g2_fill_1 FILLER_79_365 ();
 sg13g2_fill_1 FILLER_79_376 ();
 sg13g2_fill_2 FILLER_79_435 ();
 sg13g2_fill_1 FILLER_79_523 ();
 sg13g2_fill_1 FILLER_79_560 ();
 sg13g2_fill_2 FILLER_79_575 ();
 sg13g2_fill_1 FILLER_79_591 ();
 sg13g2_fill_1 FILLER_79_606 ();
 sg13g2_fill_1 FILLER_79_621 ();
 sg13g2_fill_1 FILLER_79_632 ();
 sg13g2_fill_1 FILLER_79_637 ();
 sg13g2_fill_1 FILLER_79_656 ();
 sg13g2_fill_1 FILLER_79_661 ();
 sg13g2_fill_2 FILLER_79_672 ();
 sg13g2_fill_2 FILLER_79_678 ();
 sg13g2_fill_2 FILLER_79_706 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_79_865 ();
 sg13g2_decap_8 FILLER_79_872 ();
 sg13g2_decap_8 FILLER_79_879 ();
 sg13g2_decap_8 FILLER_79_886 ();
 sg13g2_decap_8 FILLER_79_893 ();
 sg13g2_decap_8 FILLER_79_900 ();
 sg13g2_decap_8 FILLER_79_907 ();
 sg13g2_decap_8 FILLER_79_914 ();
 sg13g2_decap_8 FILLER_79_921 ();
 sg13g2_decap_8 FILLER_79_928 ();
 sg13g2_decap_8 FILLER_79_935 ();
 sg13g2_decap_8 FILLER_79_942 ();
 sg13g2_decap_8 FILLER_79_949 ();
 sg13g2_decap_8 FILLER_79_956 ();
 sg13g2_decap_8 FILLER_79_963 ();
 sg13g2_decap_8 FILLER_79_970 ();
 sg13g2_decap_8 FILLER_79_977 ();
 sg13g2_decap_8 FILLER_79_984 ();
 sg13g2_decap_8 FILLER_79_991 ();
 sg13g2_decap_8 FILLER_79_998 ();
 sg13g2_decap_8 FILLER_79_1005 ();
 sg13g2_decap_8 FILLER_79_1012 ();
 sg13g2_decap_8 FILLER_79_1019 ();
 sg13g2_decap_8 FILLER_79_1026 ();
 sg13g2_decap_8 FILLER_79_1033 ();
 sg13g2_decap_8 FILLER_79_1040 ();
 sg13g2_decap_8 FILLER_79_1047 ();
 sg13g2_decap_8 FILLER_79_1054 ();
 sg13g2_decap_8 FILLER_79_1061 ();
 sg13g2_decap_8 FILLER_79_1068 ();
 sg13g2_decap_8 FILLER_79_1075 ();
 sg13g2_decap_8 FILLER_79_1082 ();
 sg13g2_decap_8 FILLER_79_1089 ();
 sg13g2_decap_8 FILLER_79_1096 ();
 sg13g2_decap_8 FILLER_79_1103 ();
 sg13g2_decap_8 FILLER_79_1110 ();
 sg13g2_decap_8 FILLER_79_1117 ();
 sg13g2_decap_8 FILLER_79_1124 ();
 sg13g2_decap_8 FILLER_79_1131 ();
 sg13g2_decap_8 FILLER_79_1138 ();
 sg13g2_decap_8 FILLER_79_1145 ();
 sg13g2_decap_8 FILLER_79_1152 ();
 sg13g2_decap_8 FILLER_79_1159 ();
 sg13g2_decap_8 FILLER_79_1166 ();
 sg13g2_decap_8 FILLER_79_1173 ();
 sg13g2_decap_8 FILLER_79_1180 ();
 sg13g2_decap_8 FILLER_79_1187 ();
 sg13g2_decap_8 FILLER_79_1194 ();
 sg13g2_decap_8 FILLER_79_1201 ();
 sg13g2_decap_8 FILLER_79_1208 ();
 sg13g2_decap_8 FILLER_79_1215 ();
 sg13g2_decap_8 FILLER_79_1222 ();
 sg13g2_decap_8 FILLER_79_1229 ();
 sg13g2_decap_8 FILLER_79_1236 ();
 sg13g2_decap_8 FILLER_79_1243 ();
 sg13g2_decap_8 FILLER_79_1250 ();
 sg13g2_decap_8 FILLER_79_1257 ();
 sg13g2_decap_8 FILLER_79_1264 ();
 sg13g2_decap_8 FILLER_79_1271 ();
 sg13g2_decap_8 FILLER_79_1278 ();
 sg13g2_decap_8 FILLER_79_1285 ();
 sg13g2_decap_8 FILLER_79_1292 ();
 sg13g2_decap_8 FILLER_79_1299 ();
 sg13g2_decap_8 FILLER_79_1306 ();
 sg13g2_decap_8 FILLER_79_1313 ();
 sg13g2_decap_4 FILLER_79_1320 ();
 sg13g2_fill_2 FILLER_79_1324 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_21 ();
 sg13g2_fill_2 FILLER_80_197 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_fill_1 FILLER_80_288 ();
 sg13g2_fill_1 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_367 ();
 sg13g2_fill_1 FILLER_80_369 ();
 sg13g2_fill_2 FILLER_80_544 ();
 sg13g2_fill_2 FILLER_80_612 ();
 sg13g2_fill_2 FILLER_80_732 ();
 sg13g2_fill_1 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_799 ();
 sg13g2_decap_8 FILLER_80_806 ();
 sg13g2_decap_8 FILLER_80_813 ();
 sg13g2_decap_8 FILLER_80_820 ();
 sg13g2_decap_8 FILLER_80_827 ();
 sg13g2_decap_8 FILLER_80_834 ();
 sg13g2_decap_8 FILLER_80_841 ();
 sg13g2_decap_8 FILLER_80_848 ();
 sg13g2_decap_8 FILLER_80_855 ();
 sg13g2_decap_8 FILLER_80_862 ();
 sg13g2_decap_8 FILLER_80_869 ();
 sg13g2_decap_8 FILLER_80_876 ();
 sg13g2_decap_8 FILLER_80_883 ();
 sg13g2_decap_8 FILLER_80_890 ();
 sg13g2_decap_8 FILLER_80_897 ();
 sg13g2_decap_8 FILLER_80_904 ();
 sg13g2_decap_8 FILLER_80_911 ();
 sg13g2_decap_8 FILLER_80_918 ();
 sg13g2_decap_8 FILLER_80_925 ();
 sg13g2_decap_8 FILLER_80_932 ();
 sg13g2_decap_8 FILLER_80_939 ();
 sg13g2_decap_8 FILLER_80_946 ();
 sg13g2_decap_8 FILLER_80_953 ();
 sg13g2_decap_8 FILLER_80_960 ();
 sg13g2_decap_8 FILLER_80_967 ();
 sg13g2_decap_8 FILLER_80_974 ();
 sg13g2_decap_8 FILLER_80_981 ();
 sg13g2_decap_8 FILLER_80_988 ();
 sg13g2_decap_8 FILLER_80_995 ();
 sg13g2_decap_8 FILLER_80_1002 ();
 sg13g2_decap_8 FILLER_80_1009 ();
 sg13g2_decap_8 FILLER_80_1016 ();
 sg13g2_decap_8 FILLER_80_1023 ();
 sg13g2_decap_8 FILLER_80_1030 ();
 sg13g2_decap_8 FILLER_80_1037 ();
 sg13g2_decap_8 FILLER_80_1044 ();
 sg13g2_decap_8 FILLER_80_1051 ();
 sg13g2_decap_8 FILLER_80_1058 ();
 sg13g2_decap_8 FILLER_80_1065 ();
 sg13g2_decap_8 FILLER_80_1072 ();
 sg13g2_decap_8 FILLER_80_1079 ();
 sg13g2_decap_8 FILLER_80_1086 ();
 sg13g2_decap_8 FILLER_80_1093 ();
 sg13g2_decap_8 FILLER_80_1100 ();
 sg13g2_decap_8 FILLER_80_1107 ();
 sg13g2_decap_8 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1121 ();
 sg13g2_decap_8 FILLER_80_1128 ();
 sg13g2_decap_8 FILLER_80_1135 ();
 sg13g2_decap_8 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1149 ();
 sg13g2_decap_8 FILLER_80_1156 ();
 sg13g2_decap_8 FILLER_80_1163 ();
 sg13g2_decap_8 FILLER_80_1170 ();
 sg13g2_decap_8 FILLER_80_1177 ();
 sg13g2_decap_8 FILLER_80_1184 ();
 sg13g2_decap_8 FILLER_80_1191 ();
 sg13g2_decap_8 FILLER_80_1198 ();
 sg13g2_decap_8 FILLER_80_1205 ();
 sg13g2_decap_8 FILLER_80_1212 ();
 sg13g2_decap_8 FILLER_80_1219 ();
 sg13g2_decap_8 FILLER_80_1226 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_8 FILLER_80_1247 ();
 sg13g2_decap_8 FILLER_80_1254 ();
 sg13g2_decap_8 FILLER_80_1261 ();
 sg13g2_decap_8 FILLER_80_1268 ();
 sg13g2_decap_8 FILLER_80_1275 ();
 sg13g2_decap_8 FILLER_80_1282 ();
 sg13g2_decap_8 FILLER_80_1289 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_8 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1317 ();
 sg13g2_fill_2 FILLER_80_1324 ();
endmodule
