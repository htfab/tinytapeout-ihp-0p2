module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_1 _15001_ (.A(\cpu.dec.r_op[6] ),
    .X(_08279_));
 sg13g2_buf_1 _15002_ (.A(_08279_),
    .X(_08280_));
 sg13g2_buf_1 _15003_ (.A(_08280_),
    .X(_08281_));
 sg13g2_buf_1 _15004_ (.A(_00171_),
    .X(_08282_));
 sg13g2_buf_8 _15005_ (.A(\cpu.ex.ifetch ),
    .X(_08283_));
 sg13g2_inv_2 _15006_ (.Y(_08284_),
    .A(net1137));
 sg13g2_buf_1 _15007_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08285_));
 sg13g2_buf_2 _15008_ (.A(_00175_),
    .X(_08286_));
 sg13g2_a21o_1 _15009_ (.A2(_08285_),
    .A1(_08284_),
    .B1(_08286_),
    .X(_08287_));
 sg13g2_buf_4 _15010_ (.X(_08288_),
    .A(_08287_));
 sg13g2_buf_1 _15011_ (.A(\cpu.addr[13] ),
    .X(_08289_));
 sg13g2_buf_2 _15012_ (.A(\cpu.addr[15] ),
    .X(_08290_));
 sg13g2_buf_8 _15013_ (.A(_08290_),
    .X(_08291_));
 sg13g2_nor2b_1 _15014_ (.A(net1136),
    .B_N(net1076),
    .Y(_08292_));
 sg13g2_buf_8 _15015_ (.A(\cpu.addr[12] ),
    .X(_08293_));
 sg13g2_buf_8 _15016_ (.A(_08293_),
    .X(_08294_));
 sg13g2_buf_2 _15017_ (.A(\cpu.addr[14] ),
    .X(_08295_));
 sg13g2_buf_1 _15018_ (.A(_08295_),
    .X(_08296_));
 sg13g2_mux4_1 _15019_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S1(net1074),
    .X(_08297_));
 sg13g2_nand2_1 _15020_ (.Y(_08298_),
    .A(_08292_),
    .B(_08297_));
 sg13g2_buf_1 _15021_ (.A(_08295_),
    .X(_08299_));
 sg13g2_mux4_1 _15022_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S1(net1073),
    .X(_08300_));
 sg13g2_nor2_1 _15023_ (.A(net1136),
    .B(net1076),
    .Y(_08301_));
 sg13g2_nand2_1 _15024_ (.Y(_08302_),
    .A(_08300_),
    .B(_08301_));
 sg13g2_and2_1 _15025_ (.A(net1136),
    .B(_08290_),
    .X(_08303_));
 sg13g2_buf_1 _15026_ (.A(_08303_),
    .X(_08304_));
 sg13g2_mux4_1 _15027_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S1(net1074),
    .X(_08305_));
 sg13g2_mux4_1 _15028_ (.S0(_08294_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(_08296_),
    .X(_08306_));
 sg13g2_nor2b_1 _15029_ (.A(net1076),
    .B_N(net1136),
    .Y(_08307_));
 sg13g2_a22oi_1 _15030_ (.Y(_08308_),
    .B1(_08306_),
    .B2(_08307_),
    .A2(_08305_),
    .A1(_08304_));
 sg13g2_nand4_1 _15031_ (.B(_08298_),
    .C(_08302_),
    .A(_08288_),
    .Y(_08309_),
    .D(_08308_));
 sg13g2_a21oi_1 _15032_ (.A1(_08284_),
    .A2(_08285_),
    .Y(_08310_),
    .B1(_08286_));
 sg13g2_buf_1 _15033_ (.A(_08310_),
    .X(_08311_));
 sg13g2_mux4_1 _15034_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S1(net1074),
    .X(_08312_));
 sg13g2_nand2_1 _15035_ (.Y(_08313_),
    .A(_08292_),
    .B(_08312_));
 sg13g2_mux4_1 _15036_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S1(net1074),
    .X(_08314_));
 sg13g2_nand2_1 _15037_ (.Y(_08315_),
    .A(_08301_),
    .B(_08314_));
 sg13g2_mux4_1 _15038_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S1(_08295_),
    .X(_08316_));
 sg13g2_mux4_1 _15039_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net1074),
    .X(_08317_));
 sg13g2_a22oi_1 _15040_ (.Y(_08318_),
    .B1(_08317_),
    .B2(_08307_),
    .A2(_08316_),
    .A1(_08304_));
 sg13g2_nand4_1 _15041_ (.B(_08313_),
    .C(_08315_),
    .A(net826),
    .Y(_08319_),
    .D(_08318_));
 sg13g2_buf_1 _15042_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08320_));
 sg13g2_buf_2 _15043_ (.A(\cpu.ex.io_access ),
    .X(_08321_));
 sg13g2_inv_1 _15044_ (.Y(_08322_),
    .A(_08321_));
 sg13g2_buf_1 _15045_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08323_));
 sg13g2_inv_1 _15046_ (.Y(_08324_),
    .A(_08323_));
 sg13g2_buf_2 _15047_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08325_));
 sg13g2_inv_1 _15048_ (.Y(_08326_),
    .A(_08325_));
 sg13g2_nand2_1 _15049_ (.Y(_08327_),
    .A(_08324_),
    .B(_08326_));
 sg13g2_nand3_1 _15050_ (.B(_08322_),
    .C(_08327_),
    .A(net1135),
    .Y(_08328_));
 sg13g2_a21oi_1 _15051_ (.A1(_08309_),
    .A2(_08319_),
    .Y(_08329_),
    .B1(_08328_));
 sg13g2_buf_2 _15052_ (.A(_08329_),
    .X(_08330_));
 sg13g2_buf_2 _15053_ (.A(_00180_),
    .X(_08331_));
 sg13g2_buf_1 _15054_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08332_));
 sg13g2_nor2b_1 _15055_ (.A(net1134),
    .B_N(\cpu.cond[0] ),
    .Y(_08333_));
 sg13g2_nand2_1 _15056_ (.Y(_08334_),
    .A(_08331_),
    .B(_08333_));
 sg13g2_nand3_1 _15057_ (.B(_00179_),
    .C(_08334_),
    .A(net1135),
    .Y(_08335_));
 sg13g2_buf_1 _15058_ (.A(\cpu.cond[0] ),
    .X(_08336_));
 sg13g2_a21oi_2 _15059_ (.B1(_08331_),
    .Y(_08337_),
    .A2(net1133),
    .A1(net1134));
 sg13g2_nor2_1 _15060_ (.A(_08323_),
    .B(_08325_),
    .Y(_08338_));
 sg13g2_buf_2 _15061_ (.A(_08338_),
    .X(_08339_));
 sg13g2_nand2_1 _15062_ (.Y(_08340_),
    .A(_08282_),
    .B(_08339_));
 sg13g2_buf_1 _15063_ (.A(\cpu.ex.r_read_stall ),
    .X(_08341_));
 sg13g2_a21oi_1 _15064_ (.A1(_08337_),
    .A2(_08340_),
    .Y(_08342_),
    .B1(net1132));
 sg13g2_o21ai_1 _15065_ (.B1(_08328_),
    .Y(_08343_),
    .A1(_08335_),
    .A2(_08342_));
 sg13g2_mux4_1 _15066_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(net1136),
    .X(_08344_));
 sg13g2_nand3_1 _15067_ (.B(net1076),
    .C(_08344_),
    .A(net1073),
    .Y(_08345_));
 sg13g2_inv_2 _15068_ (.Y(_08346_),
    .A(net1076));
 sg13g2_mux4_1 _15069_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(net1136),
    .X(_08347_));
 sg13g2_nand3_1 _15070_ (.B(_08346_),
    .C(_08347_),
    .A(net1073),
    .Y(_08348_));
 sg13g2_mux4_1 _15071_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[11] ),
    .S1(_08289_),
    .X(_08349_));
 sg13g2_nor2b_1 _15072_ (.A(_08296_),
    .B_N(_08290_),
    .Y(_08350_));
 sg13g2_mux4_1 _15073_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[2] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[3] ),
    .S1(net1136),
    .X(_08351_));
 sg13g2_nor2_1 _15074_ (.A(net1073),
    .B(net1076),
    .Y(_08352_));
 sg13g2_a22oi_1 _15075_ (.Y(_08353_),
    .B1(_08351_),
    .B2(_08352_),
    .A2(_08350_),
    .A1(_08349_));
 sg13g2_nand3_1 _15076_ (.B(_08348_),
    .C(_08353_),
    .A(_08345_),
    .Y(_08354_));
 sg13g2_mux4_1 _15077_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[21] ),
    .S1(net1074),
    .X(_08355_));
 sg13g2_mux4_1 _15078_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[29] ),
    .S1(net1074),
    .X(_08356_));
 sg13g2_a22oi_1 _15079_ (.Y(_08357_),
    .B1(_08356_),
    .B2(_08292_),
    .A2(_08355_),
    .A1(_08301_));
 sg13g2_mux4_1 _15080_ (.S0(_08293_),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(_08295_),
    .X(_08358_));
 sg13g2_mux4_1 _15081_ (.S0(net1075),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1074),
    .X(_08359_));
 sg13g2_a22oi_1 _15082_ (.Y(_08360_),
    .B1(_08359_),
    .B2(_08304_),
    .A2(_08358_),
    .A1(_08307_));
 sg13g2_nand3_1 _15083_ (.B(_08357_),
    .C(_08360_),
    .A(_08310_),
    .Y(_08361_));
 sg13g2_o21ai_1 _15084_ (.B1(_08361_),
    .Y(_08362_),
    .A1(net826),
    .A2(_08354_));
 sg13g2_buf_4 _15085_ (.X(_08363_),
    .A(\cpu.ex.pc[15] ));
 sg13g2_buf_1 _15086_ (.A(\cpu.dec.supmode ),
    .X(_08364_));
 sg13g2_buf_8 _15087_ (.A(\cpu.ex.pc[14] ),
    .X(_08365_));
 sg13g2_mux2_1 _15088_ (.A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[4] ),
    .S(_08365_),
    .X(_08366_));
 sg13g2_mux2_1 _15089_ (.A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[5] ),
    .S(_08365_),
    .X(_08367_));
 sg13g2_mux2_1 _15090_ (.A0(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S(_08365_),
    .X(_08368_));
 sg13g2_mux2_1 _15091_ (.A0(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S(_08365_),
    .X(_08369_));
 sg13g2_buf_2 _15092_ (.A(\cpu.ex.pc[12] ),
    .X(_08370_));
 sg13g2_buf_4 _15093_ (.X(_08371_),
    .A(\cpu.ex.pc[13] ));
 sg13g2_mux4_1 _15094_ (.S0(_08370_),
    .A0(_08366_),
    .A1(_08367_),
    .A2(_08368_),
    .A3(_08369_),
    .S1(_08371_),
    .X(_08372_));
 sg13g2_nand2_1 _15095_ (.Y(_08373_),
    .A(_08320_),
    .B(_08283_));
 sg13g2_nor4_1 _15096_ (.A(_08363_),
    .B(net1131),
    .C(_08372_),
    .D(_08373_),
    .Y(_08374_));
 sg13g2_inv_4 _15097_ (.A(_08363_),
    .Y(_08375_));
 sg13g2_mux2_1 _15098_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(_08365_),
    .X(_08376_));
 sg13g2_buf_8 _15099_ (.A(_08365_),
    .X(_08377_));
 sg13g2_mux2_1 _15100_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(_08377_),
    .X(_08378_));
 sg13g2_mux2_1 _15101_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(_08365_),
    .X(_08379_));
 sg13g2_mux2_1 _15102_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(_08365_),
    .X(_08380_));
 sg13g2_mux4_1 _15103_ (.S0(_08370_),
    .A0(_08376_),
    .A1(_08378_),
    .A2(_08379_),
    .A3(_08380_),
    .S1(_08371_),
    .X(_08381_));
 sg13g2_nor4_1 _15104_ (.A(_08375_),
    .B(net1131),
    .C(_08373_),
    .D(_08381_),
    .Y(_08382_));
 sg13g2_inv_1 _15105_ (.Y(_08383_),
    .A(net1131));
 sg13g2_mux2_1 _15106_ (.A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .S(net1072),
    .X(_08384_));
 sg13g2_mux2_1 _15107_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(net1072),
    .X(_08385_));
 sg13g2_mux2_1 _15108_ (.A0(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S(net1072),
    .X(_08386_));
 sg13g2_mux2_1 _15109_ (.A0(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S(net1072),
    .X(_08387_));
 sg13g2_buf_8 _15110_ (.A(_08370_),
    .X(_08388_));
 sg13g2_mux4_1 _15111_ (.S0(_08388_),
    .A0(_08384_),
    .A1(_08385_),
    .A2(_08386_),
    .A3(_08387_),
    .S1(_08371_),
    .X(_08389_));
 sg13g2_nor4_1 _15112_ (.A(_08375_),
    .B(_08383_),
    .C(_08373_),
    .D(_08389_),
    .Y(_08390_));
 sg13g2_mux2_1 _15113_ (.A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .S(net1072),
    .X(_08391_));
 sg13g2_mux2_1 _15114_ (.A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[21] ),
    .S(net1072),
    .X(_08392_));
 sg13g2_mux2_1 _15115_ (.A0(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S(net1072),
    .X(_08393_));
 sg13g2_mux2_1 _15116_ (.A0(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S(net1072),
    .X(_08394_));
 sg13g2_mux4_1 _15117_ (.S0(_08388_),
    .A0(_08391_),
    .A1(_08392_),
    .A2(_08393_),
    .A3(_08394_),
    .S1(_08371_),
    .X(_08395_));
 sg13g2_nor4_1 _15118_ (.A(_08363_),
    .B(_08383_),
    .C(_08373_),
    .D(_08395_),
    .Y(_08396_));
 sg13g2_or4_1 _15119_ (.A(_08374_),
    .B(_08382_),
    .C(_08390_),
    .D(_08396_),
    .X(_08397_));
 sg13g2_buf_8 _15120_ (.A(_08397_),
    .X(_08398_));
 sg13g2_inv_1 _15121_ (.Y(_08399_),
    .A(net1132));
 sg13g2_nand3_1 _15122_ (.B(_08399_),
    .C(_08339_),
    .A(_08282_),
    .Y(_08400_));
 sg13g2_a22oi_1 _15123_ (.Y(_08401_),
    .B1(_08398_),
    .B2(_08400_),
    .A2(_08362_),
    .A1(_08343_));
 sg13g2_buf_8 _15124_ (.A(_08401_),
    .X(_08402_));
 sg13g2_nand2b_1 _15125_ (.Y(_08403_),
    .B(net459),
    .A_N(_08330_));
 sg13g2_buf_1 _15126_ (.A(_08403_),
    .X(_08404_));
 sg13g2_buf_1 _15127_ (.A(_08404_),
    .X(_08405_));
 sg13g2_buf_4 _15128_ (.X(_08406_),
    .A(net1071));
 sg13g2_buf_2 _15129_ (.A(_08406_),
    .X(_08407_));
 sg13g2_buf_2 _15130_ (.A(net825),
    .X(_08408_));
 sg13g2_buf_1 _15131_ (.A(net1135),
    .X(_08409_));
 sg13g2_buf_1 _15132_ (.A(_08406_),
    .X(_08410_));
 sg13g2_buf_2 _15133_ (.A(net824),
    .X(_08411_));
 sg13g2_buf_1 _15134_ (.A(_08371_),
    .X(_08412_));
 sg13g2_buf_1 _15135_ (.A(net1069),
    .X(_08413_));
 sg13g2_buf_2 _15136_ (.A(net934),
    .X(_08414_));
 sg13g2_mux4_1 _15137_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net823),
    .X(_08415_));
 sg13g2_buf_1 _15138_ (.A(_08413_),
    .X(_08416_));
 sg13g2_mux4_1 _15139_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net822),
    .X(_08417_));
 sg13g2_buf_2 _15140_ (.A(_08410_),
    .X(_08418_));
 sg13g2_mux4_1 _15141_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net823),
    .X(_08419_));
 sg13g2_mux4_1 _15142_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net823),
    .X(_08420_));
 sg13g2_buf_2 _15143_ (.A(_08375_),
    .X(_08421_));
 sg13g2_buf_2 _15144_ (.A(net933),
    .X(_08422_));
 sg13g2_buf_1 _15145_ (.A(_08377_),
    .X(_08423_));
 sg13g2_buf_2 _15146_ (.A(net932),
    .X(_08424_));
 sg13g2_mux4_1 _15147_ (.S0(net821),
    .A0(_08415_),
    .A1(_08417_),
    .A2(_08419_),
    .A3(_08420_),
    .S1(net820),
    .X(_08425_));
 sg13g2_nand2_1 _15148_ (.Y(_08426_),
    .A(net1131),
    .B(_08425_));
 sg13g2_buf_1 _15149_ (.A(_08383_),
    .X(_08427_));
 sg13g2_buf_1 _15150_ (.A(net931),
    .X(_08428_));
 sg13g2_mux4_1 _15151_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(net823),
    .X(_08429_));
 sg13g2_mux4_1 _15152_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net823),
    .X(_08430_));
 sg13g2_buf_1 _15153_ (.A(net1069),
    .X(_08431_));
 sg13g2_buf_1 _15154_ (.A(net930),
    .X(_08432_));
 sg13g2_mux4_1 _15155_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(net818),
    .X(_08433_));
 sg13g2_mux4_1 _15156_ (.S0(_08418_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(_08432_),
    .X(_08434_));
 sg13g2_mux4_1 _15157_ (.S0(net821),
    .A0(_08429_),
    .A1(_08430_),
    .A2(_08433_),
    .A3(_08434_),
    .S1(net820),
    .X(_08435_));
 sg13g2_nand2_1 _15158_ (.Y(_08436_),
    .A(net819),
    .B(_08435_));
 sg13g2_nand3_1 _15159_ (.B(_08426_),
    .C(_08436_),
    .A(net1070),
    .Y(_08437_));
 sg13g2_o21ai_1 _15160_ (.B1(_08437_),
    .Y(_08438_),
    .A1(net727),
    .A2(net1070));
 sg13g2_buf_2 _15161_ (.A(_08438_),
    .X(_08439_));
 sg13g2_buf_1 _15162_ (.A(\cpu.ex.pc[3] ),
    .X(_08440_));
 sg13g2_inv_2 _15163_ (.Y(_08441_),
    .A(_08440_));
 sg13g2_buf_2 _15164_ (.A(\cpu.ex.pc[4] ),
    .X(_08442_));
 sg13g2_buf_1 _15165_ (.A(_08440_),
    .X(_08443_));
 sg13g2_inv_2 _15166_ (.Y(_08444_),
    .A(_08442_));
 sg13g2_buf_1 _15167_ (.A(\cpu.ex.pc[2] ),
    .X(_08445_));
 sg13g2_buf_1 _15168_ (.A(_08445_),
    .X(_08446_));
 sg13g2_a21oi_1 _15169_ (.A1(net1068),
    .A2(_08444_),
    .Y(_08447_),
    .B1(net1067));
 sg13g2_a21oi_1 _15170_ (.A1(_08441_),
    .A2(_08442_),
    .Y(_08448_),
    .B1(_08447_));
 sg13g2_buf_2 _15171_ (.A(_00172_),
    .X(_08449_));
 sg13g2_buf_1 _15172_ (.A(_08449_),
    .X(_08450_));
 sg13g2_nand2b_1 _15173_ (.Y(_08451_),
    .B(net1066),
    .A_N(_08448_));
 sg13g2_buf_1 _15174_ (.A(_08451_),
    .X(_08452_));
 sg13g2_buf_1 _15175_ (.A(_08452_),
    .X(_08453_));
 sg13g2_buf_1 _15176_ (.A(net582),
    .X(_08454_));
 sg13g2_buf_1 _15177_ (.A(net517),
    .X(_08455_));
 sg13g2_inv_1 _15178_ (.Y(_08456_),
    .A(_08449_));
 sg13g2_buf_1 _15179_ (.A(_08456_),
    .X(_08457_));
 sg13g2_buf_1 _15180_ (.A(_08457_),
    .X(_08458_));
 sg13g2_buf_1 _15181_ (.A(net1067),
    .X(_08459_));
 sg13g2_buf_1 _15182_ (.A(net928),
    .X(_08460_));
 sg13g2_buf_2 _15183_ (.A(net816),
    .X(_08461_));
 sg13g2_buf_2 _15184_ (.A(net1068),
    .X(_08462_));
 sg13g2_buf_1 _15185_ (.A(net927),
    .X(_08463_));
 sg13g2_buf_2 _15186_ (.A(net815),
    .X(_08464_));
 sg13g2_buf_1 _15187_ (.A(net723),
    .X(_08465_));
 sg13g2_mux4_1 _15188_ (.S0(net724),
    .A0(\cpu.icache.r_tag[4][12] ),
    .A1(\cpu.icache.r_tag[5][12] ),
    .A2(\cpu.icache.r_tag[6][12] ),
    .A3(\cpu.icache.r_tag[7][12] ),
    .S1(net642),
    .X(_08466_));
 sg13g2_nand2_1 _15189_ (.Y(_08467_),
    .A(net817),
    .B(_08466_));
 sg13g2_inv_1 _15190_ (.Y(_08468_),
    .A(_08446_));
 sg13g2_nor3_1 _15191_ (.A(_08468_),
    .B(net1068),
    .C(_08442_),
    .Y(_08469_));
 sg13g2_buf_2 _15192_ (.A(_08469_),
    .X(_08470_));
 sg13g2_buf_1 _15193_ (.A(_08470_),
    .X(_08471_));
 sg13g2_buf_1 _15194_ (.A(net641),
    .X(_08472_));
 sg13g2_buf_1 _15195_ (.A(net581),
    .X(_08473_));
 sg13g2_buf_1 _15196_ (.A(net516),
    .X(_08474_));
 sg13g2_nand2_1 _15197_ (.Y(_08475_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(net457));
 sg13g2_and2_1 _15198_ (.A(_08445_),
    .B(_08440_),
    .X(_08476_));
 sg13g2_buf_1 _15199_ (.A(_08476_),
    .X(_08477_));
 sg13g2_and2_1 _15200_ (.A(_08449_),
    .B(net926),
    .X(_08478_));
 sg13g2_buf_2 _15201_ (.A(_08478_),
    .X(_08479_));
 sg13g2_buf_1 _15202_ (.A(_08479_),
    .X(_08480_));
 sg13g2_buf_1 _15203_ (.A(net640),
    .X(_08481_));
 sg13g2_buf_1 _15204_ (.A(net580),
    .X(_08482_));
 sg13g2_nor2_1 _15205_ (.A(_08445_),
    .B(_08441_),
    .Y(_08483_));
 sg13g2_and2_1 _15206_ (.A(_08444_),
    .B(_08483_),
    .X(_08484_));
 sg13g2_buf_2 _15207_ (.A(_08484_),
    .X(_08485_));
 sg13g2_buf_1 _15208_ (.A(_08485_),
    .X(_08486_));
 sg13g2_buf_1 _15209_ (.A(net639),
    .X(_08487_));
 sg13g2_buf_1 _15210_ (.A(net579),
    .X(_08488_));
 sg13g2_a22oi_1 _15211_ (.Y(_08489_),
    .B1(net514),
    .B2(\cpu.icache.r_tag[2][12] ),
    .A2(net515),
    .A1(\cpu.icache.r_tag[3][12] ));
 sg13g2_nand4_1 _15212_ (.B(_08467_),
    .C(_08475_),
    .A(net458),
    .Y(_08490_),
    .D(_08489_));
 sg13g2_o21ai_1 _15213_ (.B1(_08490_),
    .Y(_08491_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net458));
 sg13g2_xor2_1 _15214_ (.B(_08491_),
    .A(net362),
    .X(_08492_));
 sg13g2_mux4_1 _15215_ (.S0(net727),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net822),
    .X(_08493_));
 sg13g2_mux4_1 _15216_ (.S0(net727),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net822),
    .X(_08494_));
 sg13g2_mux4_1 _15217_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net823),
    .X(_08495_));
 sg13g2_mux4_1 _15218_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net823),
    .X(_08496_));
 sg13g2_mux4_1 _15219_ (.S0(net821),
    .A0(_08493_),
    .A1(_08494_),
    .A2(_08495_),
    .A3(_08496_),
    .S1(net820),
    .X(_08497_));
 sg13g2_nand2_1 _15220_ (.Y(_08498_),
    .A(net1131),
    .B(_08497_));
 sg13g2_mux4_1 _15221_ (.S0(_08411_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(_08414_),
    .X(_08499_));
 sg13g2_mux4_1 _15222_ (.S0(net727),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net822),
    .X(_08500_));
 sg13g2_mux4_1 _15223_ (.S0(_08411_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(_08414_),
    .X(_08501_));
 sg13g2_mux4_1 _15224_ (.S0(net726),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net823),
    .X(_08502_));
 sg13g2_mux4_1 _15225_ (.S0(net821),
    .A0(_08499_),
    .A1(_08500_),
    .A2(_08501_),
    .A3(_08502_),
    .S1(net820),
    .X(_08503_));
 sg13g2_nand2_1 _15226_ (.Y(_08504_),
    .A(net819),
    .B(_08503_));
 sg13g2_nand3_1 _15227_ (.B(_08498_),
    .C(_08504_),
    .A(net1070),
    .Y(_08505_));
 sg13g2_o21ai_1 _15228_ (.B1(_08505_),
    .Y(_08506_),
    .A1(net822),
    .A2(net1070));
 sg13g2_buf_2 _15229_ (.A(_08506_),
    .X(_08507_));
 sg13g2_nor3_2 _15230_ (.A(_08446_),
    .B(_08443_),
    .C(net1066),
    .Y(_08508_));
 sg13g2_buf_1 _15231_ (.A(_08508_),
    .X(_08509_));
 sg13g2_buf_1 _15232_ (.A(net814),
    .X(_08510_));
 sg13g2_buf_1 _15233_ (.A(net722),
    .X(_08511_));
 sg13g2_a22oi_1 _15234_ (.Y(_08512_),
    .B1(net638),
    .B2(\cpu.icache.r_tag[4][13] ),
    .A2(net457),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_a22oi_1 _15235_ (.Y(_08513_),
    .B1(net514),
    .B2(\cpu.icache.r_tag[2][13] ),
    .A2(net515),
    .A1(\cpu.icache.r_tag[3][13] ));
 sg13g2_buf_1 _15236_ (.A(net1066),
    .X(_08514_));
 sg13g2_buf_1 _15237_ (.A(net925),
    .X(_08515_));
 sg13g2_buf_1 _15238_ (.A(net813),
    .X(_08516_));
 sg13g2_buf_1 _15239_ (.A(_08483_),
    .X(_08517_));
 sg13g2_mux2_1 _15240_ (.A0(\cpu.icache.r_tag[5][13] ),
    .A1(\cpu.icache.r_tag[7][13] ),
    .S(net723),
    .X(_08518_));
 sg13g2_a22oi_1 _15241_ (.Y(_08519_),
    .B1(_08518_),
    .B2(net724),
    .A2(net812),
    .A1(\cpu.icache.r_tag[6][13] ));
 sg13g2_or2_1 _15242_ (.X(_08520_),
    .B(_08519_),
    .A(net721));
 sg13g2_nand4_1 _15243_ (.B(_08512_),
    .C(_08513_),
    .A(net458),
    .Y(_08521_),
    .D(_08520_));
 sg13g2_o21ai_1 _15244_ (.B1(_08521_),
    .Y(_08522_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net458));
 sg13g2_xor2_1 _15245_ (.B(_08522_),
    .A(net361),
    .X(_08523_));
 sg13g2_buf_4 _15246_ (.X(_08524_),
    .A(_00174_));
 sg13g2_buf_1 _15247_ (.A(_08524_),
    .X(_08525_));
 sg13g2_mux4_1 _15248_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net818),
    .X(_08526_));
 sg13g2_mux4_1 _15249_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net818),
    .X(_08527_));
 sg13g2_buf_2 _15250_ (.A(_08406_),
    .X(_08528_));
 sg13g2_buf_2 _15251_ (.A(net811),
    .X(_08529_));
 sg13g2_buf_2 _15252_ (.A(net1069),
    .X(_08530_));
 sg13g2_buf_1 _15253_ (.A(net924),
    .X(_08531_));
 sg13g2_mux4_1 _15254_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net810),
    .X(_08532_));
 sg13g2_mux4_1 _15255_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net810),
    .X(_08533_));
 sg13g2_buf_1 _15256_ (.A(net932),
    .X(_08534_));
 sg13g2_mux4_1 _15257_ (.S0(net821),
    .A0(_08526_),
    .A1(_08527_),
    .A2(_08532_),
    .A3(_08533_),
    .S1(net809),
    .X(_08535_));
 sg13g2_buf_2 _15258_ (.A(net811),
    .X(_08536_));
 sg13g2_buf_1 _15259_ (.A(net930),
    .X(_08537_));
 sg13g2_mux4_1 _15260_ (.S0(_08536_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(_08537_),
    .X(_08538_));
 sg13g2_mux4_1 _15261_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net808),
    .X(_08539_));
 sg13g2_buf_2 _15262_ (.A(net811),
    .X(_08540_));
 sg13g2_buf_1 _15263_ (.A(net924),
    .X(_08541_));
 sg13g2_mux4_1 _15264_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(net807),
    .X(_08542_));
 sg13g2_mux4_1 _15265_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net807),
    .X(_08543_));
 sg13g2_mux4_1 _15266_ (.S0(net933),
    .A0(_08538_),
    .A1(_08539_),
    .A2(_08542_),
    .A3(_08543_),
    .S1(_08534_),
    .X(_08544_));
 sg13g2_mux2_1 _15267_ (.A0(_08535_),
    .A1(_08544_),
    .S(net819),
    .X(_08545_));
 sg13g2_nand2b_1 _15268_ (.Y(_08546_),
    .B(_08545_),
    .A_N(net1065));
 sg13g2_buf_2 _15269_ (.A(_08546_),
    .X(_08547_));
 sg13g2_buf_1 _15270_ (.A(_08453_),
    .X(_08548_));
 sg13g2_buf_1 _15271_ (.A(net513),
    .X(_08549_));
 sg13g2_buf_1 _15272_ (.A(net639),
    .X(_08550_));
 sg13g2_buf_1 _15273_ (.A(net578),
    .X(_08551_));
 sg13g2_and2_1 _15274_ (.A(_08456_),
    .B(net926),
    .X(_08552_));
 sg13g2_buf_2 _15275_ (.A(_08552_),
    .X(_08553_));
 sg13g2_and2_1 _15276_ (.A(\cpu.icache.r_tag[4][18] ),
    .B(net814),
    .X(_08554_));
 sg13g2_a221oi_1 _15277_ (.B2(\cpu.icache.r_tag[7][18] ),
    .C1(_08554_),
    .B1(_08553_),
    .A1(\cpu.icache.r_tag[2][18] ),
    .Y(_08555_),
    .A2(net512));
 sg13g2_buf_1 _15278_ (.A(net581),
    .X(_08556_));
 sg13g2_and2_1 _15279_ (.A(_08457_),
    .B(_08483_),
    .X(_08557_));
 sg13g2_buf_1 _15280_ (.A(_08557_),
    .X(_08558_));
 sg13g2_buf_1 _15281_ (.A(_08558_),
    .X(_08559_));
 sg13g2_a22oi_1 _15282_ (.Y(_08560_),
    .B1(net637),
    .B2(\cpu.icache.r_tag[6][18] ),
    .A2(net511),
    .A1(\cpu.icache.r_tag[1][18] ));
 sg13g2_nor3_1 _15283_ (.A(_08468_),
    .B(net1068),
    .C(_08449_),
    .Y(_08561_));
 sg13g2_buf_2 _15284_ (.A(_08561_),
    .X(_08562_));
 sg13g2_buf_1 _15285_ (.A(_08562_),
    .X(_08563_));
 sg13g2_buf_1 _15286_ (.A(net636),
    .X(_08564_));
 sg13g2_a22oi_1 _15287_ (.Y(_08565_),
    .B1(net577),
    .B2(\cpu.icache.r_tag[5][18] ),
    .A2(net515),
    .A1(\cpu.icache.r_tag[3][18] ));
 sg13g2_nand4_1 _15288_ (.B(_08555_),
    .C(_08560_),
    .A(net456),
    .Y(_08566_),
    .D(_08565_));
 sg13g2_o21ai_1 _15289_ (.B1(_08566_),
    .Y(_08567_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net458));
 sg13g2_xnor2_1 _15290_ (.Y(_08568_),
    .A(net415),
    .B(_08567_));
 sg13g2_mux4_1 _15291_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net810),
    .X(_08569_));
 sg13g2_mux4_1 _15292_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net810),
    .X(_08570_));
 sg13g2_mux4_1 _15293_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net934),
    .X(_08571_));
 sg13g2_mux4_1 _15294_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(net934),
    .X(_08572_));
 sg13g2_mux4_1 _15295_ (.S0(_08421_),
    .A0(_08569_),
    .A1(_08570_),
    .A2(_08571_),
    .A3(_08572_),
    .S1(net809),
    .X(_08573_));
 sg13g2_mux4_1 _15296_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net807),
    .X(_08574_));
 sg13g2_mux4_1 _15297_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net807),
    .X(_08575_));
 sg13g2_mux4_1 _15298_ (.S0(_08407_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net934),
    .X(_08576_));
 sg13g2_mux4_1 _15299_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(net934),
    .X(_08577_));
 sg13g2_mux4_1 _15300_ (.S0(net933),
    .A0(_08574_),
    .A1(_08575_),
    .A2(_08576_),
    .A3(_08577_),
    .S1(net809),
    .X(_08578_));
 sg13g2_mux2_1 _15301_ (.A0(_08573_),
    .A1(_08578_),
    .S(net931),
    .X(_08579_));
 sg13g2_nand2b_1 _15302_ (.Y(_08580_),
    .B(_08579_),
    .A_N(_08525_));
 sg13g2_buf_1 _15303_ (.A(_08580_),
    .X(_08581_));
 sg13g2_and2_1 _15304_ (.A(\cpu.icache.r_tag[4][21] ),
    .B(net814),
    .X(_08582_));
 sg13g2_a221oi_1 _15305_ (.B2(\cpu.icache.r_tag[7][21] ),
    .C1(_08582_),
    .B1(_08553_),
    .A1(\cpu.icache.r_tag[2][21] ),
    .Y(_08583_),
    .A2(net512));
 sg13g2_a22oi_1 _15306_ (.Y(_08584_),
    .B1(net577),
    .B2(\cpu.icache.r_tag[5][21] ),
    .A2(net511),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_a22oi_1 _15307_ (.Y(_08585_),
    .B1(net637),
    .B2(\cpu.icache.r_tag[6][21] ),
    .A2(net515),
    .A1(\cpu.icache.r_tag[3][21] ));
 sg13g2_nand4_1 _15308_ (.B(_08583_),
    .C(_08584_),
    .A(net456),
    .Y(_08586_),
    .D(_08585_));
 sg13g2_o21ai_1 _15309_ (.B1(_08586_),
    .Y(_08587_),
    .A1(\cpu.icache.r_tag[0][21] ),
    .A2(net456));
 sg13g2_xnor2_1 _15310_ (.Y(_08588_),
    .A(net414),
    .B(_08587_));
 sg13g2_mux4_1 _15311_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1069),
    .X(_08589_));
 sg13g2_mux4_1 _15312_ (.S0(_08406_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net1069),
    .X(_08590_));
 sg13g2_mux4_1 _15313_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(_08371_),
    .X(_08591_));
 sg13g2_mux4_1 _15314_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net1069),
    .X(_08592_));
 sg13g2_mux4_1 _15315_ (.S0(_08375_),
    .A0(_08589_),
    .A1(_08590_),
    .A2(_08591_),
    .A3(_08592_),
    .S1(_08423_),
    .X(_08593_));
 sg13g2_mux4_1 _15316_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(_08412_),
    .X(_08594_));
 sg13g2_mux4_1 _15317_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net1069),
    .X(_08595_));
 sg13g2_mux4_1 _15318_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(_08371_),
    .X(_08596_));
 sg13g2_mux4_1 _15319_ (.S0(net1071),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(_08371_),
    .X(_08597_));
 sg13g2_mux4_1 _15320_ (.S0(_08375_),
    .A0(_08594_),
    .A1(_08595_),
    .A2(_08596_),
    .A3(_08597_),
    .S1(_08423_),
    .X(_08598_));
 sg13g2_mux2_1 _15321_ (.A0(_08593_),
    .A1(_08598_),
    .S(_08427_),
    .X(_08599_));
 sg13g2_nand2b_1 _15322_ (.Y(_08600_),
    .B(_08599_),
    .A_N(net1065));
 sg13g2_buf_2 _15323_ (.A(_08600_),
    .X(_08601_));
 sg13g2_nand2_1 _15324_ (.Y(_08602_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net722));
 sg13g2_a22oi_1 _15325_ (.Y(_08603_),
    .B1(_08553_),
    .B2(\cpu.icache.r_tag[7][23] ),
    .A2(net511),
    .A1(\cpu.icache.r_tag[1][23] ));
 sg13g2_nand3_1 _15326_ (.B(net925),
    .C(\cpu.icache.r_tag[3][23] ),
    .A(net723),
    .Y(_08604_));
 sg13g2_nor2_1 _15327_ (.A(net815),
    .B(net1066),
    .Y(_08605_));
 sg13g2_nand2_1 _15328_ (.Y(_08606_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(_08605_));
 sg13g2_buf_1 _15329_ (.A(_08468_),
    .X(_08607_));
 sg13g2_buf_1 _15330_ (.A(net806),
    .X(_08608_));
 sg13g2_a21oi_1 _15331_ (.A1(_08604_),
    .A2(_08606_),
    .Y(_08609_),
    .B1(net717));
 sg13g2_a221oi_1 _15332_ (.B2(\cpu.icache.r_tag[6][23] ),
    .C1(_08609_),
    .B1(net637),
    .A1(\cpu.icache.r_tag[2][23] ),
    .Y(_08610_),
    .A2(net512));
 sg13g2_nand4_1 _15333_ (.B(_08602_),
    .C(_08603_),
    .A(net517),
    .Y(_08611_),
    .D(_08610_));
 sg13g2_o21ai_1 _15334_ (.B1(_08611_),
    .Y(_08612_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net456));
 sg13g2_xnor2_1 _15335_ (.Y(_08613_),
    .A(_08601_),
    .B(_08612_));
 sg13g2_inv_1 _15336_ (.Y(_08614_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_buf_1 _15337_ (.A(_08614_),
    .X(_08615_));
 sg13g2_a22oi_1 _15338_ (.Y(_08616_),
    .B1(net814),
    .B2(\cpu.icache.r_tag[4][8] ),
    .A2(net641),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_a22oi_1 _15339_ (.Y(_08617_),
    .B1(net578),
    .B2(\cpu.icache.r_tag[2][8] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[3][8] ));
 sg13g2_mux2_1 _15340_ (.A0(\cpu.icache.r_tag[5][8] ),
    .A1(\cpu.icache.r_tag[7][8] ),
    .S(net927),
    .X(_08618_));
 sg13g2_a22oi_1 _15341_ (.Y(_08619_),
    .B1(_08618_),
    .B2(net928),
    .A2(net812),
    .A1(\cpu.icache.r_tag[6][8] ));
 sg13g2_or2_1 _15342_ (.X(_08620_),
    .B(_08619_),
    .A(_08514_));
 sg13g2_nand4_1 _15343_ (.B(_08616_),
    .C(_08617_),
    .A(_08453_),
    .Y(_08621_),
    .D(_08620_));
 sg13g2_o21ai_1 _15344_ (.B1(_08621_),
    .Y(_08622_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net582));
 sg13g2_xnor2_1 _15345_ (.Y(_08623_),
    .A(net1064),
    .B(_08622_));
 sg13g2_buf_1 _15346_ (.A(\cpu.ex.pc[6] ),
    .X(_08624_));
 sg13g2_buf_1 _15347_ (.A(net643),
    .X(_08625_));
 sg13g2_and2_1 _15348_ (.A(\cpu.icache.r_tag[7][6] ),
    .B(_08553_),
    .X(_08626_));
 sg13g2_a221oi_1 _15349_ (.B2(\cpu.icache.r_tag[6][6] ),
    .C1(_08626_),
    .B1(_08558_),
    .A1(\cpu.icache.r_tag[2][6] ),
    .Y(_08627_),
    .A2(net639));
 sg13g2_a22oi_1 _15350_ (.Y(_08628_),
    .B1(_08509_),
    .B2(\cpu.icache.r_tag[4][6] ),
    .A2(net641),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_a22oi_1 _15351_ (.Y(_08629_),
    .B1(_08562_),
    .B2(\cpu.icache.r_tag[5][6] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[3][6] ));
 sg13g2_nand4_1 _15352_ (.B(_08627_),
    .C(_08628_),
    .A(net576),
    .Y(_08630_),
    .D(_08629_));
 sg13g2_o21ai_1 _15353_ (.B1(_08630_),
    .Y(_08631_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net582));
 sg13g2_xor2_1 _15354_ (.B(_08631_),
    .A(_08624_),
    .X(_08632_));
 sg13g2_buf_1 _15355_ (.A(\cpu.ex.pc[7] ),
    .X(_08633_));
 sg13g2_a22oi_1 _15356_ (.Y(_08634_),
    .B1(_08562_),
    .B2(\cpu.icache.r_tag[5][7] ),
    .A2(_08486_),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_a22oi_1 _15357_ (.Y(_08635_),
    .B1(_08480_),
    .B2(\cpu.icache.r_tag[3][7] ),
    .A2(_08471_),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_mux2_1 _15358_ (.A0(\cpu.icache.r_tag[4][7] ),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(_08462_),
    .X(_08636_));
 sg13g2_a22oi_1 _15359_ (.Y(_08637_),
    .B1(_08636_),
    .B2(net806),
    .A2(_08477_),
    .A1(\cpu.icache.r_tag[7][7] ));
 sg13g2_or2_1 _15360_ (.X(_08638_),
    .B(_08637_),
    .A(net1066));
 sg13g2_nand4_1 _15361_ (.B(_08634_),
    .C(_08635_),
    .A(_08625_),
    .Y(_08639_),
    .D(_08638_));
 sg13g2_o21ai_1 _15362_ (.B1(_08639_),
    .Y(_08640_),
    .A1(\cpu.icache.r_tag[0][7] ),
    .A2(net582));
 sg13g2_xor2_1 _15363_ (.B(_08640_),
    .A(_08633_),
    .X(_08641_));
 sg13g2_inv_1 _15364_ (.Y(_08642_),
    .A(\cpu.ex.pc[11] ));
 sg13g2_buf_1 _15365_ (.A(_08642_),
    .X(_08643_));
 sg13g2_and2_1 _15366_ (.A(\cpu.icache.r_tag[4][11] ),
    .B(_08508_),
    .X(_08644_));
 sg13g2_a221oi_1 _15367_ (.B2(\cpu.icache.r_tag[7][11] ),
    .C1(_08644_),
    .B1(_08553_),
    .A1(\cpu.icache.r_tag[1][11] ),
    .Y(_08645_),
    .A2(_08471_));
 sg13g2_a22oi_1 _15368_ (.Y(_08646_),
    .B1(net637),
    .B2(\cpu.icache.r_tag[6][11] ),
    .A2(_08486_),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_a22oi_1 _15369_ (.Y(_08647_),
    .B1(_08562_),
    .B2(\cpu.icache.r_tag[5][11] ),
    .A2(net640),
    .A1(\cpu.icache.r_tag[3][11] ));
 sg13g2_nand4_1 _15370_ (.B(_08645_),
    .C(_08646_),
    .A(_08625_),
    .Y(_08648_),
    .D(_08647_));
 sg13g2_o21ai_1 _15371_ (.B1(_08648_),
    .Y(_08649_),
    .A1(\cpu.icache.r_tag[0][11] ),
    .A2(net582));
 sg13g2_xnor2_1 _15372_ (.Y(_08650_),
    .A(_08643_),
    .B(_08649_));
 sg13g2_nand4_1 _15373_ (.B(_08632_),
    .C(_08641_),
    .A(_08623_),
    .Y(_08651_),
    .D(_08650_));
 sg13g2_buf_1 _15374_ (.A(\cpu.ex.pc[10] ),
    .X(_08652_));
 sg13g2_buf_1 _15375_ (.A(net576),
    .X(_08653_));
 sg13g2_buf_1 _15376_ (.A(net1068),
    .X(_08654_));
 sg13g2_and2_1 _15377_ (.A(net923),
    .B(\cpu.icache.r_tag[6][10] ),
    .X(_08655_));
 sg13g2_a21oi_1 _15378_ (.A1(_08441_),
    .A2(\cpu.icache.r_tag[4][10] ),
    .Y(_08656_),
    .B1(_08655_));
 sg13g2_nor2_1 _15379_ (.A(net806),
    .B(_08443_),
    .Y(_08657_));
 sg13g2_buf_2 _15380_ (.A(_08657_),
    .X(_08658_));
 sg13g2_a22oi_1 _15381_ (.Y(_08659_),
    .B1(net926),
    .B2(\cpu.icache.r_tag[7][10] ),
    .A2(_08658_),
    .A1(\cpu.icache.r_tag[5][10] ));
 sg13g2_o21ai_1 _15382_ (.B1(_08659_),
    .Y(_08660_),
    .A1(net928),
    .A2(_08656_));
 sg13g2_nand2_1 _15383_ (.Y(_08661_),
    .A(_08458_),
    .B(_08660_));
 sg13g2_nand2_1 _15384_ (.Y(_08662_),
    .A(\cpu.icache.r_tag[1][10] ),
    .B(net516));
 sg13g2_a22oi_1 _15385_ (.Y(_08663_),
    .B1(net578),
    .B2(\cpu.icache.r_tag[2][10] ),
    .A2(net580),
    .A1(\cpu.icache.r_tag[3][10] ));
 sg13g2_nand4_1 _15386_ (.B(_08661_),
    .C(_08662_),
    .A(net509),
    .Y(_08664_),
    .D(_08663_));
 sg13g2_o21ai_1 _15387_ (.B1(_08664_),
    .Y(_08665_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(_08548_));
 sg13g2_xnor2_1 _15388_ (.Y(_08666_),
    .A(_08652_),
    .B(_08665_));
 sg13g2_buf_2 _15389_ (.A(\cpu.ex.pc[5] ),
    .X(_08667_));
 sg13g2_a22oi_1 _15390_ (.Y(_08668_),
    .B1(net636),
    .B2(\cpu.icache.r_tag[5][5] ),
    .A2(_08550_),
    .A1(\cpu.icache.r_tag[2][5] ));
 sg13g2_a22oi_1 _15391_ (.Y(_08669_),
    .B1(_08481_),
    .B2(\cpu.icache.r_tag[3][5] ),
    .A2(net581),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_buf_1 _15392_ (.A(net926),
    .X(_08670_));
 sg13g2_mux2_1 _15393_ (.A0(\cpu.icache.r_tag[4][5] ),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net923),
    .X(_08671_));
 sg13g2_a22oi_1 _15394_ (.Y(_08672_),
    .B1(_08671_),
    .B2(net806),
    .A2(net805),
    .A1(\cpu.icache.r_tag[7][5] ));
 sg13g2_or2_1 _15395_ (.X(_08673_),
    .B(_08672_),
    .A(net925));
 sg13g2_nand4_1 _15396_ (.B(_08668_),
    .C(_08669_),
    .A(net509),
    .Y(_08674_),
    .D(_08673_));
 sg13g2_o21ai_1 _15397_ (.B1(_08674_),
    .Y(_08675_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net517));
 sg13g2_xnor2_1 _15398_ (.Y(_08676_),
    .A(_08667_),
    .B(_08675_));
 sg13g2_mux4_1 _15399_ (.S0(net816),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net642),
    .X(_08677_));
 sg13g2_mux4_1 _15400_ (.S0(net816),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net642),
    .X(_08678_));
 sg13g2_mux2_1 _15401_ (.A0(_08677_),
    .A1(_08678_),
    .S(_08444_),
    .X(_08679_));
 sg13g2_buf_1 _15402_ (.A(\cpu.ex.pc[9] ),
    .X(_08680_));
 sg13g2_a22oi_1 _15403_ (.Y(_08681_),
    .B1(_08562_),
    .B2(\cpu.icache.r_tag[5][9] ),
    .A2(net578),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_a22oi_1 _15404_ (.Y(_08682_),
    .B1(_08481_),
    .B2(\cpu.icache.r_tag[3][9] ),
    .A2(_08472_),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_mux2_1 _15405_ (.A0(\cpu.icache.r_tag[4][9] ),
    .A1(\cpu.icache.r_tag[6][9] ),
    .S(net927),
    .X(_08683_));
 sg13g2_a22oi_1 _15406_ (.Y(_08684_),
    .B1(_08683_),
    .B2(net806),
    .A2(net926),
    .A1(\cpu.icache.r_tag[7][9] ));
 sg13g2_or2_1 _15407_ (.X(_08685_),
    .B(_08684_),
    .A(net925));
 sg13g2_nand4_1 _15408_ (.B(_08681_),
    .C(_08682_),
    .A(net582),
    .Y(_08686_),
    .D(_08685_));
 sg13g2_o21ai_1 _15409_ (.B1(_08686_),
    .Y(_08687_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(_08653_));
 sg13g2_xor2_1 _15410_ (.B(_08687_),
    .A(_08680_),
    .X(_08688_));
 sg13g2_nand2_1 _15411_ (.Y(_08689_),
    .A(_08679_),
    .B(_08688_));
 sg13g2_nor4_1 _15412_ (.A(_08651_),
    .B(_08666_),
    .C(_08676_),
    .D(_08689_),
    .Y(_08690_));
 sg13g2_nand4_1 _15413_ (.B(_08588_),
    .C(_08613_),
    .A(_08568_),
    .Y(_08691_),
    .D(_08690_));
 sg13g2_buf_2 _15414_ (.A(_08406_),
    .X(_08692_));
 sg13g2_mux4_1 _15415_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net924),
    .X(_08693_));
 sg13g2_mux4_1 _15416_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net924),
    .X(_08694_));
 sg13g2_buf_1 _15417_ (.A(net1069),
    .X(_08695_));
 sg13g2_mux4_1 _15418_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net922),
    .X(_08696_));
 sg13g2_mux4_1 _15419_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net922),
    .X(_08697_));
 sg13g2_mux4_1 _15420_ (.S0(net933),
    .A0(_08693_),
    .A1(_08694_),
    .A2(_08696_),
    .A3(_08697_),
    .S1(net932),
    .X(_08698_));
 sg13g2_mux4_1 _15421_ (.S0(_08692_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(net922),
    .X(_08699_));
 sg13g2_mux4_1 _15422_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net922),
    .X(_08700_));
 sg13g2_mux4_1 _15423_ (.S0(_08406_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(net922),
    .X(_08701_));
 sg13g2_mux4_1 _15424_ (.S0(_08406_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net922),
    .X(_08702_));
 sg13g2_mux4_1 _15425_ (.S0(_08375_),
    .A0(_08699_),
    .A1(_08700_),
    .A2(_08701_),
    .A3(_08702_),
    .S1(net932),
    .X(_08703_));
 sg13g2_mux2_1 _15426_ (.A0(_08698_),
    .A1(_08703_),
    .S(net931),
    .X(_08704_));
 sg13g2_nand2b_1 _15427_ (.Y(_08705_),
    .B(_08704_),
    .A_N(net1065));
 sg13g2_buf_2 _15428_ (.A(_08705_),
    .X(_08706_));
 sg13g2_a22oi_1 _15429_ (.Y(_08707_),
    .B1(_08509_),
    .B2(\cpu.icache.r_tag[4][19] ),
    .A2(_08473_),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_a22oi_1 _15430_ (.Y(_08708_),
    .B1(net636),
    .B2(\cpu.icache.r_tag[5][19] ),
    .A2(net579),
    .A1(\cpu.icache.r_tag[2][19] ));
 sg13g2_mux2_1 _15431_ (.A0(\cpu.icache.r_tag[7][19] ),
    .A1(\cpu.icache.r_tag[3][19] ),
    .S(_08450_),
    .X(_08709_));
 sg13g2_nor2_1 _15432_ (.A(net928),
    .B(_08450_),
    .Y(_08710_));
 sg13g2_a22oi_1 _15433_ (.Y(_08711_),
    .B1(_08710_),
    .B2(\cpu.icache.r_tag[6][19] ),
    .A2(_08709_),
    .A1(_08459_));
 sg13g2_nand2b_1 _15434_ (.Y(_08712_),
    .B(_08464_),
    .A_N(_08711_));
 sg13g2_nand4_1 _15435_ (.B(_08707_),
    .C(_08708_),
    .A(net509),
    .Y(_08713_),
    .D(_08712_));
 sg13g2_o21ai_1 _15436_ (.B1(_08713_),
    .Y(_08714_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(net517));
 sg13g2_xor2_1 _15437_ (.B(_08714_),
    .A(net455),
    .X(_08715_));
 sg13g2_mux4_1 _15438_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net924),
    .X(_08716_));
 sg13g2_mux4_1 _15439_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net924),
    .X(_08717_));
 sg13g2_mux4_1 _15440_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net922),
    .X(_08718_));
 sg13g2_mux4_1 _15441_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net922),
    .X(_08719_));
 sg13g2_mux4_1 _15442_ (.S0(net933),
    .A0(_08716_),
    .A1(_08717_),
    .A2(_08718_),
    .A3(_08719_),
    .S1(net932),
    .X(_08720_));
 sg13g2_mux4_1 _15443_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(_08530_),
    .X(_08721_));
 sg13g2_mux4_1 _15444_ (.S0(net804),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net924),
    .X(_08722_));
 sg13g2_mux4_1 _15445_ (.S0(_08406_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(_08695_),
    .X(_08723_));
 sg13g2_mux4_1 _15446_ (.S0(_08692_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(_08695_),
    .X(_08724_));
 sg13g2_mux4_1 _15447_ (.S0(net933),
    .A0(_08721_),
    .A1(_08722_),
    .A2(_08723_),
    .A3(_08724_),
    .S1(net932),
    .X(_08725_));
 sg13g2_mux2_1 _15448_ (.A0(_08720_),
    .A1(_08725_),
    .S(net931),
    .X(_08726_));
 sg13g2_nand2b_1 _15449_ (.Y(_08727_),
    .B(_08726_),
    .A_N(net1065));
 sg13g2_buf_2 _15450_ (.A(_08727_),
    .X(_08728_));
 sg13g2_a22oi_1 _15451_ (.Y(_08729_),
    .B1(_08563_),
    .B2(\cpu.icache.r_tag[5][16] ),
    .A2(net579),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_buf_1 _15452_ (.A(net580),
    .X(_08730_));
 sg13g2_a22oi_1 _15453_ (.Y(_08731_),
    .B1(_08730_),
    .B2(\cpu.icache.r_tag[3][16] ),
    .A2(_08472_),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_mux2_1 _15454_ (.A0(\cpu.icache.r_tag[4][16] ),
    .A1(\cpu.icache.r_tag[6][16] ),
    .S(_08654_),
    .X(_08732_));
 sg13g2_a22oi_1 _15455_ (.Y(_08733_),
    .B1(_08732_),
    .B2(_08607_),
    .A2(net805),
    .A1(\cpu.icache.r_tag[7][16] ));
 sg13g2_or2_1 _15456_ (.X(_08734_),
    .B(_08733_),
    .A(_08515_));
 sg13g2_nand4_1 _15457_ (.B(_08729_),
    .C(_08731_),
    .A(net509),
    .Y(_08735_),
    .D(_08734_));
 sg13g2_o21ai_1 _15458_ (.B1(_08735_),
    .Y(_08736_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net517));
 sg13g2_xor2_1 _15459_ (.B(_08736_),
    .A(_08728_),
    .X(_08737_));
 sg13g2_mux4_1 _15460_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net930),
    .X(_08738_));
 sg13g2_mux4_1 _15461_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(_08431_),
    .X(_08739_));
 sg13g2_mux4_1 _15462_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net930),
    .X(_08740_));
 sg13g2_mux4_1 _15463_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net930),
    .X(_08741_));
 sg13g2_mux4_1 _15464_ (.S0(net931),
    .A0(_08738_),
    .A1(_08739_),
    .A2(_08740_),
    .A3(_08741_),
    .S1(net932),
    .X(_08742_));
 sg13g2_a21oi_1 _15465_ (.A1(net1070),
    .A2(_08742_),
    .Y(_08743_),
    .B1(_08363_));
 sg13g2_inv_1 _15466_ (.Y(_08744_),
    .A(net1135));
 sg13g2_mux4_1 _15467_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(net934),
    .X(_08745_));
 sg13g2_mux4_1 _15468_ (.S0(_08407_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(_08413_),
    .X(_08746_));
 sg13g2_mux4_1 _15469_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(net930),
    .X(_08747_));
 sg13g2_mux4_1 _15470_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(_08431_),
    .X(_08748_));
 sg13g2_mux4_1 _15471_ (.S0(_08427_),
    .A0(_08745_),
    .A1(_08746_),
    .A2(_08747_),
    .A3(_08748_),
    .S1(net932),
    .X(_08749_));
 sg13g2_nor3_1 _15472_ (.A(net821),
    .B(_08744_),
    .C(_08749_),
    .Y(_08750_));
 sg13g2_or2_1 _15473_ (.X(_08751_),
    .B(_08750_),
    .A(_08743_));
 sg13g2_buf_2 _15474_ (.A(_08751_),
    .X(_08752_));
 sg13g2_and2_1 _15475_ (.A(_08654_),
    .B(\cpu.icache.r_tag[6][15] ),
    .X(_08753_));
 sg13g2_a21oi_1 _15476_ (.A1(_08441_),
    .A2(\cpu.icache.r_tag[4][15] ),
    .Y(_08754_),
    .B1(_08753_));
 sg13g2_a22oi_1 _15477_ (.Y(_08755_),
    .B1(_08670_),
    .B2(\cpu.icache.r_tag[7][15] ),
    .A2(_08658_),
    .A1(\cpu.icache.r_tag[5][15] ));
 sg13g2_o21ai_1 _15478_ (.B1(_08755_),
    .Y(_08756_),
    .A1(_08460_),
    .A2(_08754_));
 sg13g2_nand2_1 _15479_ (.Y(_08757_),
    .A(_08458_),
    .B(_08756_));
 sg13g2_nand2_1 _15480_ (.Y(_08758_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net511));
 sg13g2_a22oi_1 _15481_ (.Y(_08759_),
    .B1(_08487_),
    .B2(\cpu.icache.r_tag[2][15] ),
    .A2(_08730_),
    .A1(\cpu.icache.r_tag[3][15] ));
 sg13g2_nand4_1 _15482_ (.B(_08757_),
    .C(_08758_),
    .A(_08653_),
    .Y(_08760_),
    .D(_08759_));
 sg13g2_o21ai_1 _15483_ (.B1(_08760_),
    .Y(_08761_),
    .A1(\cpu.icache.r_tag[0][15] ),
    .A2(_08454_));
 sg13g2_xor2_1 _15484_ (.B(_08761_),
    .A(net453),
    .X(_08762_));
 sg13g2_mux4_1 _15485_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net930),
    .X(_08763_));
 sg13g2_mux4_1 _15486_ (.S0(net824),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net930),
    .X(_08764_));
 sg13g2_mux4_1 _15487_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net924),
    .X(_08765_));
 sg13g2_mux4_1 _15488_ (.S0(_08528_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(_08530_),
    .X(_08766_));
 sg13g2_mux4_1 _15489_ (.S0(net931),
    .A0(_08763_),
    .A1(_08764_),
    .A2(_08765_),
    .A3(_08766_),
    .S1(_08363_),
    .X(_08767_));
 sg13g2_nand2b_1 _15490_ (.Y(_08768_),
    .B(net1070),
    .A_N(_08767_));
 sg13g2_mux4_1 _15491_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net808),
    .X(_08769_));
 sg13g2_mux4_1 _15492_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net808),
    .X(_08770_));
 sg13g2_mux4_1 _15493_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net807),
    .X(_08771_));
 sg13g2_mux4_1 _15494_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net807),
    .X(_08772_));
 sg13g2_mux4_1 _15495_ (.S0(net931),
    .A0(_08769_),
    .A1(_08770_),
    .A2(_08771_),
    .A3(_08772_),
    .S1(_08363_),
    .X(_08773_));
 sg13g2_nor2_1 _15496_ (.A(net820),
    .B(_08744_),
    .Y(_08774_));
 sg13g2_a22oi_1 _15497_ (.Y(_08775_),
    .B1(_08773_),
    .B2(_08774_),
    .A2(_08768_),
    .A1(net820));
 sg13g2_buf_2 _15498_ (.A(_08775_),
    .X(_08776_));
 sg13g2_mux2_1 _15499_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net925),
    .X(_08777_));
 sg13g2_buf_1 _15500_ (.A(net805),
    .X(_08778_));
 sg13g2_a22oi_1 _15501_ (.Y(_08779_),
    .B1(_08777_),
    .B2(_08778_),
    .A2(_08510_),
    .A1(\cpu.icache.r_tag[4][14] ));
 sg13g2_a22oi_1 _15502_ (.Y(_08780_),
    .B1(net637),
    .B2(\cpu.icache.r_tag[6][14] ),
    .A2(_08473_),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_a22oi_1 _15503_ (.Y(_08781_),
    .B1(_08563_),
    .B2(\cpu.icache.r_tag[5][14] ),
    .A2(_08487_),
    .A1(\cpu.icache.r_tag[2][14] ));
 sg13g2_nand4_1 _15504_ (.B(_08779_),
    .C(_08780_),
    .A(_08548_),
    .Y(_08782_),
    .D(_08781_));
 sg13g2_o21ai_1 _15505_ (.B1(_08782_),
    .Y(_08783_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(_08454_));
 sg13g2_xor2_1 _15506_ (.B(_08783_),
    .A(_08776_),
    .X(_08784_));
 sg13g2_nor4_1 _15507_ (.A(_08715_),
    .B(_08737_),
    .C(_08762_),
    .D(_08784_),
    .Y(_08785_));
 sg13g2_mux4_1 _15508_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net818),
    .X(_08786_));
 sg13g2_mux4_1 _15509_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net818),
    .X(_08787_));
 sg13g2_mux4_1 _15510_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net808),
    .X(_08788_));
 sg13g2_mux4_1 _15511_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net808),
    .X(_08789_));
 sg13g2_mux4_1 _15512_ (.S0(net821),
    .A0(_08786_),
    .A1(_08787_),
    .A2(_08788_),
    .A3(_08789_),
    .S1(net809),
    .X(_08790_));
 sg13g2_mux4_1 _15513_ (.S0(_08418_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(_08432_),
    .X(_08791_));
 sg13g2_mux4_1 _15514_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net818),
    .X(_08792_));
 sg13g2_mux4_1 _15515_ (.S0(_08529_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(_08531_),
    .X(_08793_));
 sg13g2_mux4_1 _15516_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(net810),
    .X(_08794_));
 sg13g2_mux4_1 _15517_ (.S0(net821),
    .A0(_08791_),
    .A1(_08792_),
    .A2(_08793_),
    .A3(_08794_),
    .S1(_08534_),
    .X(_08795_));
 sg13g2_mux2_1 _15518_ (.A0(_08790_),
    .A1(_08795_),
    .S(net819),
    .X(_08796_));
 sg13g2_nand2b_1 _15519_ (.Y(_08797_),
    .B(_08796_),
    .A_N(net1065));
 sg13g2_buf_2 _15520_ (.A(_08797_),
    .X(_08798_));
 sg13g2_a22oi_1 _15521_ (.Y(_08799_),
    .B1(_08564_),
    .B2(\cpu.icache.r_tag[5][17] ),
    .A2(_08551_),
    .A1(\cpu.icache.r_tag[2][17] ));
 sg13g2_a22oi_1 _15522_ (.Y(_08800_),
    .B1(_08482_),
    .B2(\cpu.icache.r_tag[3][17] ),
    .A2(net457),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_mux2_1 _15523_ (.A0(\cpu.icache.r_tag[4][17] ),
    .A1(\cpu.icache.r_tag[6][17] ),
    .S(net815),
    .X(_08801_));
 sg13g2_a22oi_1 _15524_ (.Y(_08802_),
    .B1(_08801_),
    .B2(net717),
    .A2(_08670_),
    .A1(\cpu.icache.r_tag[7][17] ));
 sg13g2_or2_1 _15525_ (.X(_08803_),
    .B(_08802_),
    .A(_08516_));
 sg13g2_nand4_1 _15526_ (.B(_08799_),
    .C(_08800_),
    .A(net456),
    .Y(_08804_),
    .D(_08803_));
 sg13g2_o21ai_1 _15527_ (.B1(_08804_),
    .Y(_08805_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(_08455_));
 sg13g2_xnor2_1 _15528_ (.Y(_08806_),
    .A(net413),
    .B(_08805_));
 sg13g2_mux4_1 _15529_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net818),
    .X(_08807_));
 sg13g2_mux4_1 _15530_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net818),
    .X(_08808_));
 sg13g2_mux4_1 _15531_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net810),
    .X(_08809_));
 sg13g2_mux4_1 _15532_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net810),
    .X(_08810_));
 sg13g2_mux4_1 _15533_ (.S0(_08422_),
    .A0(_08807_),
    .A1(_08808_),
    .A2(_08809_),
    .A3(_08810_),
    .S1(net809),
    .X(_08811_));
 sg13g2_mux4_1 _15534_ (.S0(_08536_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(_08537_),
    .X(_08812_));
 sg13g2_mux4_1 _15535_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net808),
    .X(_08813_));
 sg13g2_mux4_1 _15536_ (.S0(_08540_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(_08541_),
    .X(_08814_));
 sg13g2_mux4_1 _15537_ (.S0(_08540_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(_08541_),
    .X(_08815_));
 sg13g2_mux4_1 _15538_ (.S0(net933),
    .A0(_08812_),
    .A1(_08813_),
    .A2(_08814_),
    .A3(_08815_),
    .S1(net809),
    .X(_08816_));
 sg13g2_mux2_1 _15539_ (.A0(_08811_),
    .A1(_08816_),
    .S(net819),
    .X(_08817_));
 sg13g2_nand2b_1 _15540_ (.Y(_08818_),
    .B(_08817_),
    .A_N(net1065));
 sg13g2_buf_1 _15541_ (.A(_08818_),
    .X(_08819_));
 sg13g2_a22oi_1 _15542_ (.Y(_08820_),
    .B1(net637),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(_08556_),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_a22oi_1 _15543_ (.Y(_08821_),
    .B1(_08488_),
    .B2(\cpu.icache.r_tag[2][22] ),
    .A2(_08482_),
    .A1(\cpu.icache.r_tag[3][22] ));
 sg13g2_nor2_1 _15544_ (.A(_08459_),
    .B(_08463_),
    .Y(_08822_));
 sg13g2_mux2_1 _15545_ (.A0(\cpu.icache.r_tag[5][22] ),
    .A1(\cpu.icache.r_tag[7][22] ),
    .S(_08463_),
    .X(_08823_));
 sg13g2_a22oi_1 _15546_ (.Y(_08824_),
    .B1(_08823_),
    .B2(_08460_),
    .A2(_08822_),
    .A1(\cpu.icache.r_tag[4][22] ));
 sg13g2_or2_1 _15547_ (.X(_08825_),
    .B(_08824_),
    .A(_08516_));
 sg13g2_nand4_1 _15548_ (.B(_08820_),
    .C(_08821_),
    .A(_08549_),
    .Y(_08826_),
    .D(_08825_));
 sg13g2_o21ai_1 _15549_ (.B1(_08826_),
    .Y(_08827_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(_08455_));
 sg13g2_xnor2_1 _15550_ (.Y(_08828_),
    .A(net412),
    .B(_08827_));
 sg13g2_mux4_1 _15551_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net808),
    .X(_08829_));
 sg13g2_mux4_1 _15552_ (.S0(net719),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(net808),
    .X(_08830_));
 sg13g2_mux4_1 _15553_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net807),
    .X(_08831_));
 sg13g2_mux4_1 _15554_ (.S0(net718),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(net807),
    .X(_08832_));
 sg13g2_mux4_1 _15555_ (.S0(_08421_),
    .A0(_08829_),
    .A1(_08830_),
    .A2(_08831_),
    .A3(_08832_),
    .S1(net809),
    .X(_08833_));
 sg13g2_mux4_1 _15556_ (.S0(_08529_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(_08531_),
    .X(_08834_));
 sg13g2_mux4_1 _15557_ (.S0(net720),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net810),
    .X(_08835_));
 sg13g2_mux4_1 _15558_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(net934),
    .X(_08836_));
 sg13g2_mux4_1 _15559_ (.S0(net825),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net934),
    .X(_08837_));
 sg13g2_mux4_1 _15560_ (.S0(net933),
    .A0(_08834_),
    .A1(_08835_),
    .A2(_08836_),
    .A3(_08837_),
    .S1(net809),
    .X(_08838_));
 sg13g2_mux2_1 _15561_ (.A0(_08833_),
    .A1(_08838_),
    .S(net931),
    .X(_08839_));
 sg13g2_nand2b_1 _15562_ (.Y(_08840_),
    .B(_08839_),
    .A_N(net1065));
 sg13g2_buf_1 _15563_ (.A(_08840_),
    .X(_08841_));
 sg13g2_a22oi_1 _15564_ (.Y(_08842_),
    .B1(_08559_),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(_08551_),
    .A1(\cpu.icache.r_tag[2][20] ));
 sg13g2_a22oi_1 _15565_ (.Y(_08843_),
    .B1(_08510_),
    .B2(\cpu.icache.r_tag[4][20] ),
    .A2(_08556_),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_mux2_1 _15566_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(_08514_),
    .X(_08844_));
 sg13g2_a22oi_1 _15567_ (.Y(_08845_),
    .B1(_08844_),
    .B2(_08464_),
    .A2(_08605_),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_nand2b_1 _15568_ (.Y(_08846_),
    .B(net724),
    .A_N(_08845_));
 sg13g2_nand4_1 _15569_ (.B(_08842_),
    .C(_08843_),
    .A(_08549_),
    .Y(_08847_),
    .D(_08846_));
 sg13g2_o21ai_1 _15570_ (.B1(_08847_),
    .Y(_08848_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net456));
 sg13g2_xnor2_1 _15571_ (.Y(_08849_),
    .A(net411),
    .B(_08848_));
 sg13g2_nand4_1 _15572_ (.B(_08806_),
    .C(_08828_),
    .A(_08785_),
    .Y(_08850_),
    .D(_08849_));
 sg13g2_or4_2 _15573_ (.A(_08492_),
    .B(_08523_),
    .C(_08691_),
    .D(_08850_),
    .X(_08851_));
 sg13g2_or3_1 _15574_ (.A(_08282_),
    .B(_08405_),
    .C(_08851_),
    .X(_08852_));
 sg13g2_buf_1 _15575_ (.A(_08852_),
    .X(_08853_));
 sg13g2_buf_1 _15576_ (.A(_08853_),
    .X(_08854_));
 sg13g2_buf_1 _15577_ (.A(net123),
    .X(_08855_));
 sg13g2_buf_1 _15578_ (.A(_08853_),
    .X(_08856_));
 sg13g2_buf_2 _15579_ (.A(\cpu.ex.pc[1] ),
    .X(_08857_));
 sg13g2_buf_1 _15580_ (.A(_08857_),
    .X(_08858_));
 sg13g2_nor2_1 _15581_ (.A(net929),
    .B(_08448_),
    .Y(_08859_));
 sg13g2_a22oi_1 _15582_ (.Y(_08860_),
    .B1(_08508_),
    .B2(\cpu.icache.r_data[4][5] ),
    .A2(_08470_),
    .A1(\cpu.icache.r_data[1][5] ));
 sg13g2_a22oi_1 _15583_ (.Y(_08861_),
    .B1(_08485_),
    .B2(\cpu.icache.r_data[2][5] ),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[3][5] ));
 sg13g2_mux2_1 _15584_ (.A0(\cpu.icache.r_data[5][5] ),
    .A1(\cpu.icache.r_data[7][5] ),
    .S(net1068),
    .X(_08862_));
 sg13g2_a22oi_1 _15585_ (.Y(_08863_),
    .B1(_08862_),
    .B2(net1067),
    .A2(_08483_),
    .A1(\cpu.icache.r_data[6][5] ));
 sg13g2_or2_1 _15586_ (.X(_08864_),
    .B(_08863_),
    .A(net1066));
 sg13g2_and4_1 _15587_ (.A(net643),
    .B(_08860_),
    .C(_08861_),
    .D(_08864_),
    .X(_08865_));
 sg13g2_a21oi_1 _15588_ (.A1(_00183_),
    .A2(_08859_),
    .Y(_08866_),
    .B1(_08865_));
 sg13g2_inv_1 _15589_ (.Y(_08867_),
    .A(_08857_));
 sg13g2_buf_1 _15590_ (.A(_08867_),
    .X(_08868_));
 sg13g2_nor2_1 _15591_ (.A(_00184_),
    .B(net643),
    .Y(_08869_));
 sg13g2_mux2_1 _15592_ (.A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(net927),
    .X(_08870_));
 sg13g2_a22oi_1 _15593_ (.Y(_08871_),
    .B1(_08870_),
    .B2(net806),
    .A2(net926),
    .A1(\cpu.icache.r_data[7][21] ));
 sg13g2_nor2_1 _15594_ (.A(net925),
    .B(_08871_),
    .Y(_08872_));
 sg13g2_a22oi_1 _15595_ (.Y(_08873_),
    .B1(net639),
    .B2(\cpu.icache.r_data[2][21] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][21] ));
 sg13g2_a22oi_1 _15596_ (.Y(_08874_),
    .B1(_08562_),
    .B2(\cpu.icache.r_data[5][21] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[3][21] ));
 sg13g2_nand2_1 _15597_ (.Y(_08875_),
    .A(_08873_),
    .B(_08874_));
 sg13g2_or4_1 _15598_ (.A(net921),
    .B(_08869_),
    .C(_08872_),
    .D(_08875_),
    .X(_08876_));
 sg13g2_o21ai_1 _15599_ (.B1(_08876_),
    .Y(_08877_),
    .A1(net1062),
    .A2(_08866_));
 sg13g2_buf_2 _15600_ (.A(_08877_),
    .X(_08878_));
 sg13g2_inv_1 _15601_ (.Y(_08879_),
    .A(_00185_));
 sg13g2_mux4_1 _15602_ (.S0(net1067),
    .A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[5][6] ),
    .A2(\cpu.icache.r_data[6][6] ),
    .A3(\cpu.icache.r_data[7][6] ),
    .S1(net1068),
    .X(_08880_));
 sg13g2_nand2_1 _15603_ (.Y(_08881_),
    .A(net929),
    .B(_08880_));
 sg13g2_nand2_1 _15604_ (.Y(_08882_),
    .A(\cpu.icache.r_data[1][6] ),
    .B(_08470_));
 sg13g2_a22oi_1 _15605_ (.Y(_08883_),
    .B1(_08485_),
    .B2(\cpu.icache.r_data[2][6] ),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[3][6] ));
 sg13g2_nand4_1 _15606_ (.B(_08881_),
    .C(_08882_),
    .A(net643),
    .Y(_08884_),
    .D(_08883_));
 sg13g2_o21ai_1 _15607_ (.B1(_08884_),
    .Y(_08885_),
    .A1(_08879_),
    .A2(net643));
 sg13g2_mux4_1 _15608_ (.S0(net1067),
    .A0(\cpu.icache.r_data[4][22] ),
    .A1(\cpu.icache.r_data[5][22] ),
    .A2(\cpu.icache.r_data[6][22] ),
    .A3(\cpu.icache.r_data[7][22] ),
    .S1(net927),
    .X(_08886_));
 sg13g2_and2_1 _15609_ (.A(net929),
    .B(_08886_),
    .X(_08887_));
 sg13g2_and2_1 _15610_ (.A(\cpu.icache.r_data[3][22] ),
    .B(_08479_),
    .X(_08888_));
 sg13g2_a221oi_1 _15611_ (.B2(\cpu.icache.r_data[2][22] ),
    .C1(_08888_),
    .B1(_08485_),
    .A1(\cpu.icache.r_data[1][22] ),
    .Y(_08889_),
    .A2(_08470_));
 sg13g2_o21ai_1 _15612_ (.B1(_08889_),
    .Y(_08890_),
    .A1(_00186_),
    .A2(net643));
 sg13g2_o21ai_1 _15613_ (.B1(_08857_),
    .Y(_08891_),
    .A1(_08887_),
    .A2(_08890_));
 sg13g2_o21ai_1 _15614_ (.B1(_08891_),
    .Y(_08892_),
    .A1(_08857_),
    .A2(_08885_));
 sg13g2_buf_2 _15615_ (.A(_08892_),
    .X(_08893_));
 sg13g2_inv_1 _15616_ (.Y(_08894_),
    .A(_08893_));
 sg13g2_nand2_1 _15617_ (.Y(_08895_),
    .A(_08878_),
    .B(_08894_));
 sg13g2_buf_1 _15618_ (.A(_08895_),
    .X(_08896_));
 sg13g2_buf_1 _15619_ (.A(net1062),
    .X(_08897_));
 sg13g2_a22oi_1 _15620_ (.Y(_08898_),
    .B1(net637),
    .B2(\cpu.icache.r_data[6][16] ),
    .A2(net457),
    .A1(\cpu.icache.r_data[1][16] ));
 sg13g2_a22oi_1 _15621_ (.Y(_08899_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][16] ),
    .A2(net514),
    .A1(\cpu.icache.r_data[2][16] ));
 sg13g2_mux2_1 _15622_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(net813),
    .X(_08900_));
 sg13g2_a22oi_1 _15623_ (.Y(_08901_),
    .B1(_08900_),
    .B2(net716),
    .A2(net577),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_buf_1 _15624_ (.A(_08859_),
    .X(_08902_));
 sg13g2_nand2_1 _15625_ (.Y(_08903_),
    .A(\cpu.icache.r_data[0][16] ),
    .B(net635));
 sg13g2_nand4_1 _15626_ (.B(_08899_),
    .C(_08901_),
    .A(_08898_),
    .Y(_08904_),
    .D(_08903_));
 sg13g2_a22oi_1 _15627_ (.Y(_08905_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][0] ),
    .A2(net516),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_a22oi_1 _15628_ (.Y(_08906_),
    .B1(net579),
    .B2(\cpu.icache.r_data[2][0] ),
    .A2(net580),
    .A1(\cpu.icache.r_data[3][0] ));
 sg13g2_mux2_1 _15629_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(\cpu.icache.r_data[7][0] ),
    .S(net923),
    .X(_08907_));
 sg13g2_a22oi_1 _15630_ (.Y(_08908_),
    .B1(_08907_),
    .B2(net928),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][0] ));
 sg13g2_or2_1 _15631_ (.X(_08909_),
    .B(_08908_),
    .A(net813));
 sg13g2_nand4_1 _15632_ (.B(_08905_),
    .C(_08906_),
    .A(net509),
    .Y(_08910_),
    .D(_08909_));
 sg13g2_o21ai_1 _15633_ (.B1(_08910_),
    .Y(_08911_),
    .A1(\cpu.icache.r_data[0][0] ),
    .A2(net517));
 sg13g2_nor2_1 _15634_ (.A(net920),
    .B(_08911_),
    .Y(_08912_));
 sg13g2_a21o_1 _15635_ (.A2(_08904_),
    .A1(net920),
    .B1(_08912_),
    .X(_08913_));
 sg13g2_buf_1 _15636_ (.A(_08913_),
    .X(_08914_));
 sg13g2_nor2_1 _15637_ (.A(_00200_),
    .B(net513),
    .Y(_08915_));
 sg13g2_mux2_1 _15638_ (.A0(\cpu.icache.r_data[4][17] ),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(net723),
    .X(_08916_));
 sg13g2_a22oi_1 _15639_ (.Y(_08917_),
    .B1(_08916_),
    .B2(net717),
    .A2(net716),
    .A1(\cpu.icache.r_data[7][17] ));
 sg13g2_nor2_1 _15640_ (.A(net721),
    .B(_08917_),
    .Y(_08918_));
 sg13g2_a22oi_1 _15641_ (.Y(_08919_),
    .B1(net512),
    .B2(\cpu.icache.r_data[2][17] ),
    .A2(net511),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_a22oi_1 _15642_ (.Y(_08920_),
    .B1(net636),
    .B2(\cpu.icache.r_data[5][17] ),
    .A2(net508),
    .A1(\cpu.icache.r_data[3][17] ));
 sg13g2_nand2_1 _15643_ (.Y(_08921_),
    .A(_08919_),
    .B(_08920_));
 sg13g2_nor3_1 _15644_ (.A(_08915_),
    .B(_08918_),
    .C(_08921_),
    .Y(_08922_));
 sg13g2_nand2_1 _15645_ (.Y(_08923_),
    .A(_00199_),
    .B(net635));
 sg13g2_a22oi_1 _15646_ (.Y(_08924_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][1] ),
    .A2(net511),
    .A1(\cpu.icache.r_data[1][1] ));
 sg13g2_a22oi_1 _15647_ (.Y(_08925_),
    .B1(net512),
    .B2(\cpu.icache.r_data[2][1] ),
    .A2(net508),
    .A1(\cpu.icache.r_data[3][1] ));
 sg13g2_mux2_1 _15648_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(\cpu.icache.r_data[7][1] ),
    .S(net815),
    .X(_08926_));
 sg13g2_a22oi_1 _15649_ (.Y(_08927_),
    .B1(_08926_),
    .B2(net816),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][1] ));
 sg13g2_or2_1 _15650_ (.X(_08928_),
    .B(_08927_),
    .A(net813));
 sg13g2_nand4_1 _15651_ (.B(_08924_),
    .C(_08925_),
    .A(net513),
    .Y(_08929_),
    .D(_08928_));
 sg13g2_a21oi_1 _15652_ (.A1(_08923_),
    .A2(_08929_),
    .Y(_08930_),
    .B1(net1062));
 sg13g2_a21o_1 _15653_ (.A2(_08922_),
    .A1(net920),
    .B1(_08930_),
    .X(_08931_));
 sg13g2_buf_1 _15654_ (.A(_08931_),
    .X(_08932_));
 sg13g2_buf_1 _15655_ (.A(_08932_),
    .X(_08933_));
 sg13g2_nand2_1 _15656_ (.Y(_08934_),
    .A(_08914_),
    .B(net221));
 sg13g2_buf_1 _15657_ (.A(_08934_),
    .X(_08935_));
 sg13g2_nor2_1 _15658_ (.A(_00198_),
    .B(net509),
    .Y(_08936_));
 sg13g2_mux2_1 _15659_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(\cpu.icache.r_data[7][31] ),
    .S(net815),
    .X(_08937_));
 sg13g2_a22oi_1 _15660_ (.Y(_08938_),
    .B1(_08937_),
    .B2(net724),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][31] ));
 sg13g2_nor2_1 _15661_ (.A(net721),
    .B(_08938_),
    .Y(_08939_));
 sg13g2_a22oi_1 _15662_ (.Y(_08940_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][31] ),
    .A2(net516),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_a22oi_1 _15663_ (.Y(_08941_),
    .B1(net512),
    .B2(\cpu.icache.r_data[2][31] ),
    .A2(net508),
    .A1(\cpu.icache.r_data[3][31] ));
 sg13g2_nand2_1 _15664_ (.Y(_08942_),
    .A(_08940_),
    .B(_08941_));
 sg13g2_nor3_1 _15665_ (.A(_08936_),
    .B(_08939_),
    .C(_08942_),
    .Y(_08943_));
 sg13g2_nand2_1 _15666_ (.Y(_08944_),
    .A(_00197_),
    .B(net635));
 sg13g2_a22oi_1 _15667_ (.Y(_08945_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][15] ),
    .A2(net516),
    .A1(\cpu.icache.r_data[1][15] ));
 sg13g2_a22oi_1 _15668_ (.Y(_08946_),
    .B1(net579),
    .B2(\cpu.icache.r_data[2][15] ),
    .A2(net508),
    .A1(\cpu.icache.r_data[3][15] ));
 sg13g2_mux2_1 _15669_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(\cpu.icache.r_data[7][15] ),
    .S(net923),
    .X(_08947_));
 sg13g2_a22oi_1 _15670_ (.Y(_08948_),
    .B1(_08947_),
    .B2(net816),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][15] ));
 sg13g2_or2_1 _15671_ (.X(_08949_),
    .B(_08948_),
    .A(net813));
 sg13g2_nand4_1 _15672_ (.B(_08945_),
    .C(_08946_),
    .A(net513),
    .Y(_08950_),
    .D(_08949_));
 sg13g2_a21oi_1 _15673_ (.A1(_08944_),
    .A2(_08950_),
    .Y(_08951_),
    .B1(net1062));
 sg13g2_a21oi_1 _15674_ (.A1(net920),
    .A2(_08943_),
    .Y(_08952_),
    .B1(_08951_));
 sg13g2_buf_1 _15675_ (.A(_08952_),
    .X(_08953_));
 sg13g2_a22oi_1 _15676_ (.Y(_08954_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][14] ),
    .A2(_08470_),
    .A1(\cpu.icache.r_data[1][14] ));
 sg13g2_a22oi_1 _15677_ (.Y(_08955_),
    .B1(net639),
    .B2(\cpu.icache.r_data[2][14] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[3][14] ));
 sg13g2_mux2_1 _15678_ (.A0(\cpu.icache.r_data[5][14] ),
    .A1(\cpu.icache.r_data[7][14] ),
    .S(net1068),
    .X(_08956_));
 sg13g2_a22oi_1 _15679_ (.Y(_08957_),
    .B1(_08956_),
    .B2(net928),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][14] ));
 sg13g2_or2_1 _15680_ (.X(_08958_),
    .B(_08957_),
    .A(net1066));
 sg13g2_and4_1 _15681_ (.A(net643),
    .B(_08954_),
    .C(_08955_),
    .D(_08958_),
    .X(_08959_));
 sg13g2_a21oi_1 _15682_ (.A1(_00195_),
    .A2(net635),
    .Y(_08960_),
    .B1(_08959_));
 sg13g2_nor2_1 _15683_ (.A(_00196_),
    .B(net576),
    .Y(_08961_));
 sg13g2_a22oi_1 _15684_ (.Y(_08962_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][30] ),
    .A2(net639),
    .A1(\cpu.icache.r_data[2][30] ));
 sg13g2_mux2_1 _15685_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net1066),
    .X(_08963_));
 sg13g2_a22oi_1 _15686_ (.Y(_08964_),
    .B1(_08963_),
    .B2(net805),
    .A2(_08558_),
    .A1(\cpu.icache.r_data[6][30] ));
 sg13g2_a22oi_1 _15687_ (.Y(_08965_),
    .B1(_08562_),
    .B2(\cpu.icache.r_data[5][30] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_nand3_1 _15688_ (.B(_08964_),
    .C(_08965_),
    .A(_08962_),
    .Y(_08966_));
 sg13g2_or3_1 _15689_ (.A(net921),
    .B(_08961_),
    .C(_08966_),
    .X(_08967_));
 sg13g2_o21ai_1 _15690_ (.B1(_08967_),
    .Y(_08968_),
    .A1(net1062),
    .A2(_08960_));
 sg13g2_buf_2 _15691_ (.A(_08968_),
    .X(_08969_));
 sg13g2_nand2b_1 _15692_ (.Y(_08970_),
    .B(_08859_),
    .A_N(_00194_));
 sg13g2_mux2_1 _15693_ (.A0(\cpu.icache.r_data[4][29] ),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(net927),
    .X(_08971_));
 sg13g2_a22oi_1 _15694_ (.Y(_08972_),
    .B1(_08971_),
    .B2(net806),
    .A2(net926),
    .A1(\cpu.icache.r_data[7][29] ));
 sg13g2_or2_1 _15695_ (.X(_08973_),
    .B(_08972_),
    .A(net925));
 sg13g2_a22oi_1 _15696_ (.Y(_08974_),
    .B1(net578),
    .B2(\cpu.icache.r_data[2][29] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[1][29] ));
 sg13g2_a22oi_1 _15697_ (.Y(_08975_),
    .B1(net636),
    .B2(\cpu.icache.r_data[5][29] ),
    .A2(net580),
    .A1(\cpu.icache.r_data[3][29] ));
 sg13g2_nand4_1 _15698_ (.B(_08973_),
    .C(_08974_),
    .A(_08970_),
    .Y(_08976_),
    .D(_08975_));
 sg13g2_nand2_1 _15699_ (.Y(_08977_),
    .A(_00193_),
    .B(_08859_));
 sg13g2_mux4_1 _15700_ (.S0(net928),
    .A0(\cpu.icache.r_data[4][13] ),
    .A1(\cpu.icache.r_data[5][13] ),
    .A2(\cpu.icache.r_data[6][13] ),
    .A3(\cpu.icache.r_data[7][13] ),
    .S1(net923),
    .X(_08978_));
 sg13g2_nand2_1 _15701_ (.Y(_08979_),
    .A(net929),
    .B(_08978_));
 sg13g2_nand2_1 _15702_ (.Y(_08980_),
    .A(\cpu.icache.r_data[1][13] ),
    .B(net641));
 sg13g2_a22oi_1 _15703_ (.Y(_08981_),
    .B1(net639),
    .B2(\cpu.icache.r_data[2][13] ),
    .A2(net640),
    .A1(\cpu.icache.r_data[3][13] ));
 sg13g2_nand4_1 _15704_ (.B(_08979_),
    .C(_08980_),
    .A(net576),
    .Y(_08982_),
    .D(_08981_));
 sg13g2_and3_1 _15705_ (.X(_08983_),
    .A(net921),
    .B(_08977_),
    .C(_08982_));
 sg13g2_a21oi_1 _15706_ (.A1(net1062),
    .A2(_08976_),
    .Y(_08984_),
    .B1(_08983_));
 sg13g2_buf_1 _15707_ (.A(_08984_),
    .X(_08985_));
 sg13g2_and2_1 _15708_ (.A(_08969_),
    .B(_08985_),
    .X(_08986_));
 sg13g2_buf_1 _15709_ (.A(_08986_),
    .X(_08987_));
 sg13g2_nand2_1 _15710_ (.Y(_08988_),
    .A(_08953_),
    .B(_08987_));
 sg13g2_buf_1 _15711_ (.A(_08988_),
    .X(_08989_));
 sg13g2_nor2_1 _15712_ (.A(_08935_),
    .B(net199),
    .Y(_08990_));
 sg13g2_buf_1 _15713_ (.A(net920),
    .X(_08991_));
 sg13g2_nand2b_1 _15714_ (.Y(_08992_),
    .B(net635),
    .A_N(_00192_));
 sg13g2_mux2_1 _15715_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(net642),
    .X(_08993_));
 sg13g2_a22oi_1 _15716_ (.Y(_08994_),
    .B1(_08993_),
    .B2(net717),
    .A2(net716),
    .A1(\cpu.icache.r_data[7][27] ));
 sg13g2_or2_1 _15717_ (.X(_08995_),
    .B(_08994_),
    .A(net721));
 sg13g2_buf_1 _15718_ (.A(net515),
    .X(_08996_));
 sg13g2_a22oi_1 _15719_ (.Y(_08997_),
    .B1(_08996_),
    .B2(\cpu.icache.r_data[3][27] ),
    .A2(net457),
    .A1(\cpu.icache.r_data[1][27] ));
 sg13g2_a22oi_1 _15720_ (.Y(_08998_),
    .B1(net577),
    .B2(\cpu.icache.r_data[5][27] ),
    .A2(net514),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_nand4_1 _15721_ (.B(_08995_),
    .C(_08997_),
    .A(_08992_),
    .Y(_08999_),
    .D(_08998_));
 sg13g2_nand2_1 _15722_ (.Y(_09000_),
    .A(_00191_),
    .B(_08902_));
 sg13g2_and2_1 _15723_ (.A(net723),
    .B(\cpu.icache.r_data[6][11] ),
    .X(_09001_));
 sg13g2_a21oi_1 _15724_ (.A1(_08441_),
    .A2(\cpu.icache.r_data[4][11] ),
    .Y(_09002_),
    .B1(_09001_));
 sg13g2_a22oi_1 _15725_ (.Y(_09003_),
    .B1(net716),
    .B2(\cpu.icache.r_data[7][11] ),
    .A2(_08658_),
    .A1(\cpu.icache.r_data[5][11] ));
 sg13g2_o21ai_1 _15726_ (.B1(_09003_),
    .Y(_09004_),
    .A1(_08461_),
    .A2(_09002_));
 sg13g2_nand2_1 _15727_ (.Y(_09005_),
    .A(net817),
    .B(_09004_));
 sg13g2_nand2_1 _15728_ (.Y(_09006_),
    .A(\cpu.icache.r_data[1][11] ),
    .B(net457));
 sg13g2_a22oi_1 _15729_ (.Y(_09007_),
    .B1(net514),
    .B2(\cpu.icache.r_data[2][11] ),
    .A2(net515),
    .A1(\cpu.icache.r_data[3][11] ));
 sg13g2_nand4_1 _15730_ (.B(_09005_),
    .C(_09006_),
    .A(net458),
    .Y(_09008_),
    .D(_09007_));
 sg13g2_and3_1 _15731_ (.X(_09009_),
    .A(net921),
    .B(_09000_),
    .C(_09008_));
 sg13g2_a21oi_1 _15732_ (.A1(net803),
    .A2(_08999_),
    .Y(_09010_),
    .B1(_09009_));
 sg13g2_buf_2 _15733_ (.A(_09010_),
    .X(_09011_));
 sg13g2_mux4_1 _15734_ (.S0(net816),
    .A0(\cpu.icache.r_data[4][26] ),
    .A1(\cpu.icache.r_data[5][26] ),
    .A2(\cpu.icache.r_data[6][26] ),
    .A3(\cpu.icache.r_data[7][26] ),
    .S1(_08465_),
    .X(_09012_));
 sg13g2_and2_1 _15735_ (.A(\cpu.icache.r_data[3][26] ),
    .B(net580),
    .X(_09013_));
 sg13g2_a221oi_1 _15736_ (.B2(\cpu.icache.r_data[2][26] ),
    .C1(_09013_),
    .B1(net579),
    .A1(\cpu.icache.r_data[1][26] ),
    .Y(_09014_),
    .A2(net516));
 sg13g2_o21ai_1 _15737_ (.B1(_09014_),
    .Y(_09015_),
    .A1(_00190_),
    .A2(net513));
 sg13g2_a21oi_1 _15738_ (.A1(net817),
    .A2(_09012_),
    .Y(_09016_),
    .B1(_09015_));
 sg13g2_nand2_1 _15739_ (.Y(_09017_),
    .A(_00189_),
    .B(_08902_));
 sg13g2_a22oi_1 _15740_ (.Y(_09018_),
    .B1(net636),
    .B2(\cpu.icache.r_data[5][10] ),
    .A2(net579),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_a22oi_1 _15741_ (.Y(_09019_),
    .B1(net508),
    .B2(\cpu.icache.r_data[3][10] ),
    .A2(net516),
    .A1(\cpu.icache.r_data[1][10] ));
 sg13g2_mux2_1 _15742_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(net923),
    .X(_09020_));
 sg13g2_a22oi_1 _15743_ (.Y(_09021_),
    .B1(_09020_),
    .B2(net806),
    .A2(net805),
    .A1(\cpu.icache.r_data[7][10] ));
 sg13g2_or2_1 _15744_ (.X(_09022_),
    .B(_09021_),
    .A(_08515_));
 sg13g2_nand4_1 _15745_ (.B(_09018_),
    .C(_09019_),
    .A(net513),
    .Y(_09023_),
    .D(_09022_));
 sg13g2_a21oi_1 _15746_ (.A1(_09017_),
    .A2(_09023_),
    .Y(_09024_),
    .B1(_08858_));
 sg13g2_a21oi_1 _15747_ (.A1(_08897_),
    .A2(_09016_),
    .Y(_09025_),
    .B1(_09024_));
 sg13g2_buf_1 _15748_ (.A(_09025_),
    .X(_09026_));
 sg13g2_inv_2 _15749_ (.Y(_09027_),
    .A(_09026_));
 sg13g2_nor2_2 _15750_ (.A(_09011_),
    .B(_09027_),
    .Y(_09028_));
 sg13g2_mux4_1 _15751_ (.S0(_08461_),
    .A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[5][28] ),
    .A2(\cpu.icache.r_data[6][28] ),
    .A3(\cpu.icache.r_data[7][28] ),
    .S1(_08465_),
    .X(_09029_));
 sg13g2_and2_1 _15752_ (.A(\cpu.icache.r_data[3][28] ),
    .B(net515),
    .X(_09030_));
 sg13g2_a221oi_1 _15753_ (.B2(\cpu.icache.r_data[2][28] ),
    .C1(_09030_),
    .B1(net514),
    .A1(\cpu.icache.r_data[1][28] ),
    .Y(_09031_),
    .A2(_08474_));
 sg13g2_o21ai_1 _15754_ (.B1(_09031_),
    .Y(_09032_),
    .A1(_00188_),
    .A2(net458));
 sg13g2_a21oi_1 _15755_ (.A1(net817),
    .A2(_09029_),
    .Y(_09033_),
    .B1(_09032_));
 sg13g2_nand2_1 _15756_ (.Y(_09034_),
    .A(_00187_),
    .B(net635));
 sg13g2_a22oi_1 _15757_ (.Y(_09035_),
    .B1(net577),
    .B2(\cpu.icache.r_data[5][12] ),
    .A2(net514),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15758_ (.Y(_09036_),
    .B1(net451),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(net457),
    .A1(\cpu.icache.r_data[1][12] ));
 sg13g2_mux2_1 _15759_ (.A0(\cpu.icache.r_data[4][12] ),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(net723),
    .X(_09037_));
 sg13g2_a22oi_1 _15760_ (.Y(_09038_),
    .B1(_09037_),
    .B2(net717),
    .A2(net716),
    .A1(\cpu.icache.r_data[7][12] ));
 sg13g2_or2_1 _15761_ (.X(_09039_),
    .B(_09038_),
    .A(net721));
 sg13g2_nand4_1 _15762_ (.B(_09035_),
    .C(_09036_),
    .A(net458),
    .Y(_09040_),
    .D(_09039_));
 sg13g2_a21oi_1 _15763_ (.A1(_09034_),
    .A2(_09040_),
    .Y(_09041_),
    .B1(net920));
 sg13g2_a21o_1 _15764_ (.A2(_09033_),
    .A1(net803),
    .B1(_09041_),
    .X(_09042_));
 sg13g2_buf_1 _15765_ (.A(_09042_),
    .X(_09043_));
 sg13g2_buf_1 _15766_ (.A(_09043_),
    .X(_09044_));
 sg13g2_nand3_1 _15767_ (.B(_09028_),
    .C(net198),
    .A(_08990_),
    .Y(_09045_));
 sg13g2_buf_1 _15768_ (.A(_09045_),
    .X(_09046_));
 sg13g2_nor3_1 _15769_ (.A(net122),
    .B(_08896_),
    .C(_09046_),
    .Y(_09047_));
 sg13g2_a21o_1 _15770_ (.A2(net108),
    .A1(net935),
    .B1(_09047_),
    .X(_00017_));
 sg13g2_buf_2 _15771_ (.A(\cpu.dec.r_op[4] ),
    .X(_09048_));
 sg13g2_buf_1 _15772_ (.A(_09048_),
    .X(_09049_));
 sg13g2_a21o_1 _15773_ (.A2(_08943_),
    .A1(net920),
    .B1(_08951_),
    .X(_09050_));
 sg13g2_buf_2 _15774_ (.A(_09050_),
    .X(_09051_));
 sg13g2_nand2_2 _15775_ (.Y(_09052_),
    .A(_08969_),
    .B(_08985_));
 sg13g2_nor2_1 _15776_ (.A(_09051_),
    .B(_09052_),
    .Y(_09053_));
 sg13g2_buf_1 _15777_ (.A(_09053_),
    .X(_09054_));
 sg13g2_a21oi_1 _15778_ (.A1(_08991_),
    .A2(_08904_),
    .Y(_09055_),
    .B1(_08912_));
 sg13g2_buf_1 _15779_ (.A(_09055_),
    .X(_09056_));
 sg13g2_nor2_1 _15780_ (.A(net220),
    .B(net221),
    .Y(_09057_));
 sg13g2_buf_2 _15781_ (.A(_09057_),
    .X(_09058_));
 sg13g2_nand3_1 _15782_ (.B(_09028_),
    .C(_09058_),
    .A(net197),
    .Y(_09059_));
 sg13g2_buf_1 _15783_ (.A(_09059_),
    .X(_09060_));
 sg13g2_nor4_1 _15784_ (.A(_08854_),
    .B(_08896_),
    .C(net198),
    .D(_09060_),
    .Y(_09061_));
 sg13g2_a21o_1 _15785_ (.A2(_08855_),
    .A1(net1061),
    .B1(_09061_),
    .X(_00015_));
 sg13g2_buf_1 _15786_ (.A(_08856_),
    .X(_09062_));
 sg13g2_buf_1 _15787_ (.A(_09011_),
    .X(_09063_));
 sg13g2_buf_1 _15788_ (.A(_09026_),
    .X(_09064_));
 sg13g2_nand3_1 _15789_ (.B(net196),
    .C(net219),
    .A(_08990_),
    .Y(_09065_));
 sg13g2_buf_1 _15790_ (.A(\cpu.dec.r_op[5] ),
    .X(_09066_));
 sg13g2_buf_1 _15791_ (.A(_08853_),
    .X(_09067_));
 sg13g2_nand2_1 _15792_ (.Y(_09068_),
    .A(net1130),
    .B(net121));
 sg13g2_o21ai_1 _15793_ (.B1(_09068_),
    .Y(_00016_),
    .A1(_09062_),
    .A2(_09065_));
 sg13g2_buf_2 _15794_ (.A(\cpu.dec.r_op[1] ),
    .X(_09069_));
 sg13g2_buf_1 _15795_ (.A(_08878_),
    .X(_09070_));
 sg13g2_nand2_1 _15796_ (.Y(_09071_),
    .A(_09070_),
    .B(_08893_));
 sg13g2_nor3_1 _15797_ (.A(net122),
    .B(_09060_),
    .C(_09071_),
    .Y(_09072_));
 sg13g2_a21o_1 _15798_ (.A2(net108),
    .A1(_09069_),
    .B1(_09072_),
    .X(_00012_));
 sg13g2_buf_2 _15799_ (.A(\cpu.dec.r_op[3] ),
    .X(_09073_));
 sg13g2_buf_1 _15800_ (.A(_09073_),
    .X(_09074_));
 sg13g2_or2_1 _15801_ (.X(_09075_),
    .B(_08893_),
    .A(_08878_));
 sg13g2_buf_1 _15802_ (.A(_09075_),
    .X(_09076_));
 sg13g2_nor3_1 _15803_ (.A(net122),
    .B(_09046_),
    .C(_09076_),
    .Y(_09077_));
 sg13g2_a21o_1 _15804_ (.A2(net108),
    .A1(net1060),
    .B1(_09077_),
    .X(_00014_));
 sg13g2_buf_1 _15805_ (.A(\cpu.dec.r_op[7] ),
    .X(_09078_));
 sg13g2_nor4_1 _15806_ (.A(net123),
    .B(_09070_),
    .C(_08894_),
    .D(_09060_),
    .Y(_09079_));
 sg13g2_a21o_1 _15807_ (.A2(net108),
    .A1(_09078_),
    .B1(_09079_),
    .X(_00018_));
 sg13g2_nor2b_1 _15808_ (.A(r_reset),
    .B_N(net1),
    .Y(_09080_));
 sg13g2_buf_2 _15809_ (.A(_09080_),
    .X(_09081_));
 sg13g2_buf_1 _15810_ (.A(_09081_),
    .X(_09082_));
 sg13g2_buf_1 _15811_ (.A(net919),
    .X(_09083_));
 sg13g2_buf_1 _15812_ (.A(_09083_),
    .X(_09084_));
 sg13g2_buf_1 _15813_ (.A(_00203_),
    .X(_09085_));
 sg13g2_inv_2 _15814_ (.Y(_09086_),
    .A(_09085_));
 sg13g2_buf_2 _15815_ (.A(\cpu.dec.r_trap ),
    .X(_09087_));
 sg13g2_buf_1 _15816_ (.A(\cpu.gpio.r_enable_in[2] ),
    .X(_09088_));
 sg13g2_buf_1 _15817_ (.A(ui_in[2]),
    .X(_09089_));
 sg13g2_buf_1 _15818_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_09090_));
 sg13g2_buf_1 _15819_ (.A(ui_in[4]),
    .X(_09091_));
 sg13g2_a22oi_1 _15820_ (.Y(_09092_),
    .B1(_09090_),
    .B2(_09091_),
    .A2(_09089_),
    .A1(_09088_));
 sg13g2_buf_1 _15821_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09093_));
 sg13g2_buf_1 _15822_ (.A(ui_in[1]),
    .X(_09094_));
 sg13g2_buf_1 _15823_ (.A(\cpu.gpio.r_enable_io[7] ),
    .X(_09095_));
 sg13g2_buf_1 _15824_ (.A(uio_in[7]),
    .X(_09096_));
 sg13g2_a22oi_1 _15825_ (.Y(_09097_),
    .B1(_09095_),
    .B2(_09096_),
    .A2(_09094_),
    .A1(_09093_));
 sg13g2_nand2_1 _15826_ (.Y(_09098_),
    .A(_09092_),
    .B(_09097_));
 sg13g2_buf_1 _15827_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_09099_));
 sg13g2_buf_2 _15828_ (.A(ui_in[6]),
    .X(_09100_));
 sg13g2_buf_1 _15829_ (.A(uio_in[6]),
    .X(_09101_));
 sg13g2_a22oi_1 _15830_ (.Y(_09102_),
    .B1(\cpu.gpio.r_enable_io[6] ),
    .B2(_09101_),
    .A2(_09100_),
    .A1(_09099_));
 sg13g2_buf_1 _15831_ (.A(\cpu.gpio.r_enable_io[4] ),
    .X(_09103_));
 sg13g2_buf_1 _15832_ (.A(uio_in[4]),
    .X(_09104_));
 sg13g2_buf_1 _15833_ (.A(\cpu.gpio.r_enable_io[5] ),
    .X(_09105_));
 sg13g2_a22oi_1 _15834_ (.Y(_09106_),
    .B1(_09105_),
    .B2(net3),
    .A2(_09104_),
    .A1(_09103_));
 sg13g2_buf_2 _15835_ (.A(ui_in[0]),
    .X(_09107_));
 sg13g2_buf_1 _15836_ (.A(\cpu.gpio.r_enable_in[7] ),
    .X(_09108_));
 sg13g2_buf_2 _15837_ (.A(ui_in[7]),
    .X(_09109_));
 sg13g2_a22oi_1 _15838_ (.Y(_09110_),
    .B1(_09108_),
    .B2(_09109_),
    .A2(_09107_),
    .A1(\cpu.gpio.r_enable_in[0] ));
 sg13g2_buf_1 _15839_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09111_));
 sg13g2_buf_2 _15840_ (.A(ui_in[3]),
    .X(_09112_));
 sg13g2_buf_1 _15841_ (.A(\cpu.gpio.r_enable_in[5] ),
    .X(_09113_));
 sg13g2_buf_2 _15842_ (.A(ui_in[5]),
    .X(_09114_));
 sg13g2_a22oi_1 _15843_ (.Y(_09115_),
    .B1(_09113_),
    .B2(_09114_),
    .A2(_09112_),
    .A1(_09111_));
 sg13g2_nand4_1 _15844_ (.B(_09106_),
    .C(_09110_),
    .A(_09102_),
    .Y(_09116_),
    .D(_09115_));
 sg13g2_buf_1 _15845_ (.A(_09116_),
    .X(_09117_));
 sg13g2_buf_1 _15846_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09118_));
 sg13g2_o21ai_1 _15847_ (.B1(_09118_),
    .Y(_09119_),
    .A1(_09098_),
    .A2(_09117_));
 sg13g2_buf_1 _15848_ (.A(\cpu.intr.r_swi ),
    .X(_09120_));
 sg13g2_buf_1 _15849_ (.A(\cpu.intr.spi_intr ),
    .X(_09121_));
 sg13g2_buf_1 _15850_ (.A(\cpu.intr.r_enable[5] ),
    .X(_09122_));
 sg13g2_a22oi_1 _15851_ (.Y(_09123_),
    .B1(_09121_),
    .B2(_09122_),
    .A2(_09120_),
    .A1(\cpu.intr.r_enable[3] ));
 sg13g2_buf_1 _15852_ (.A(\cpu.intr.r_enable[1] ),
    .X(_09124_));
 sg13g2_buf_1 _15853_ (.A(\cpu.intr.r_enable[2] ),
    .X(_09125_));
 sg13g2_a22oi_1 _15854_ (.Y(_09126_),
    .B1(\cpu.intr.r_timer ),
    .B2(_09125_),
    .A2(_09124_),
    .A1(\cpu.intr.r_clock ));
 sg13g2_buf_1 _15855_ (.A(\cpu.uart.r_x_int ),
    .X(_09127_));
 sg13g2_buf_1 _15856_ (.A(\cpu.uart.r_r_int ),
    .X(_09128_));
 sg13g2_buf_1 _15857_ (.A(\cpu.intr.r_enable[0] ),
    .X(_09129_));
 sg13g2_o21ai_1 _15858_ (.B1(_09129_),
    .Y(_09130_),
    .A1(_09127_),
    .A2(_09128_));
 sg13g2_nand3_1 _15859_ (.B(_09126_),
    .C(_09130_),
    .A(_09123_),
    .Y(_09131_));
 sg13g2_inv_1 _15860_ (.Y(_09132_),
    .A(_09131_));
 sg13g2_buf_1 _15861_ (.A(\cpu.ex.r_ie ),
    .X(_09133_));
 sg13g2_inv_2 _15862_ (.Y(_09134_),
    .A(_09133_));
 sg13g2_a21oi_2 _15863_ (.B1(_09134_),
    .Y(_09135_),
    .A2(_09132_),
    .A1(_09119_));
 sg13g2_and2_1 _15864_ (.A(net1131),
    .B(_09135_),
    .X(_09136_));
 sg13g2_nor3_2 _15865_ (.A(_09087_),
    .B(_08404_),
    .C(_09136_),
    .Y(_09137_));
 sg13g2_buf_1 _15866_ (.A(\cpu.addr[2] ),
    .X(_09138_));
 sg13g2_buf_1 _15867_ (.A(net1129),
    .X(_09139_));
 sg13g2_buf_1 _15868_ (.A(_09139_),
    .X(_09140_));
 sg13g2_buf_1 _15869_ (.A(_09140_),
    .X(_09141_));
 sg13g2_buf_2 _15870_ (.A(net801),
    .X(_09142_));
 sg13g2_buf_2 _15871_ (.A(\cpu.addr[1] ),
    .X(_09143_));
 sg13g2_nor2_2 _15872_ (.A(net714),
    .B(net1128),
    .Y(_09144_));
 sg13g2_nand3b_1 _15873_ (.B(_09137_),
    .C(_09144_),
    .Y(_09145_),
    .A_N(_00179_));
 sg13g2_inv_1 _15874_ (.Y(_09146_),
    .A(_08331_));
 sg13g2_mux2_1 _15875_ (.A0(_08331_),
    .A1(_08399_),
    .S(net1134),
    .X(_09147_));
 sg13g2_nand2_1 _15876_ (.Y(_09148_),
    .A(net1133),
    .B(_09147_));
 sg13g2_o21ai_1 _15877_ (.B1(_09148_),
    .Y(_09149_),
    .A1(_09146_),
    .A2(net1132));
 sg13g2_buf_1 _15878_ (.A(\cpu.addr[6] ),
    .X(_09150_));
 sg13g2_buf_1 _15879_ (.A(_09150_),
    .X(_09151_));
 sg13g2_buf_2 _15880_ (.A(\cpu.addr[8] ),
    .X(_09152_));
 sg13g2_inv_1 _15881_ (.Y(_09153_),
    .A(_09152_));
 sg13g2_buf_1 _15882_ (.A(\cpu.addr[7] ),
    .X(_09154_));
 sg13g2_buf_1 _15883_ (.A(_09154_),
    .X(_09155_));
 sg13g2_nand3_1 _15884_ (.B(_09153_),
    .C(net1057),
    .A(net1058),
    .Y(_09156_));
 sg13g2_buf_1 _15885_ (.A(_09156_),
    .X(_09157_));
 sg13g2_nor4_2 _15886_ (.A(_09086_),
    .B(_09145_),
    .C(_09149_),
    .Y(_09158_),
    .D(_09157_));
 sg13g2_buf_1 _15887_ (.A(\cpu.addr[3] ),
    .X(_09159_));
 sg13g2_buf_1 _15888_ (.A(_09159_),
    .X(_09160_));
 sg13g2_buf_1 _15889_ (.A(net1056),
    .X(_09161_));
 sg13g2_buf_1 _15890_ (.A(net917),
    .X(_09162_));
 sg13g2_buf_2 _15891_ (.A(_09162_),
    .X(_09163_));
 sg13g2_buf_1 _15892_ (.A(net713),
    .X(_09164_));
 sg13g2_buf_1 _15893_ (.A(net634),
    .X(_09165_));
 sg13g2_buf_1 _15894_ (.A(net575),
    .X(_09166_));
 sg13g2_nand3_1 _15895_ (.B(_08327_),
    .C(_09137_),
    .A(_08321_),
    .Y(_09167_));
 sg13g2_buf_2 _15896_ (.A(_09167_),
    .X(_09168_));
 sg13g2_or2_1 _15897_ (.X(_09169_),
    .B(_09168_),
    .A(net800));
 sg13g2_buf_2 _15898_ (.A(_09169_),
    .X(_09170_));
 sg13g2_buf_1 _15899_ (.A(\cpu.spi.r_state[1] ),
    .X(_09171_));
 sg13g2_o21ai_1 _15900_ (.B1(net1127),
    .Y(_09172_),
    .A1(net507),
    .A2(_09170_));
 sg13g2_buf_1 _15901_ (.A(\cpu.spi.r_state[6] ),
    .X(_09173_));
 sg13g2_buf_1 _15902_ (.A(_09173_),
    .X(_09174_));
 sg13g2_buf_1 _15903_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09175_));
 sg13g2_buf_1 _15904_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09176_));
 sg13g2_nor3_1 _15905_ (.A(_09175_),
    .B(_09176_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09177_));
 sg13g2_nor3_2 _15906_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .C(\cpu.spi.r_timeout_count[2] ),
    .Y(_09178_));
 sg13g2_nor2b_1 _15907_ (.A(\cpu.spi.r_timeout_count[3] ),
    .B_N(_09178_),
    .Y(_09179_));
 sg13g2_nand2b_1 _15908_ (.Y(_09180_),
    .B(_09179_),
    .A_N(\cpu.spi.r_timeout_count[4] ));
 sg13g2_nor2_1 _15909_ (.A(\cpu.spi.r_timeout_count[5] ),
    .B(_09180_),
    .Y(_09181_));
 sg13g2_nand2b_1 _15910_ (.Y(_09182_),
    .B(_09181_),
    .A_N(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _15911_ (.A(_09182_),
    .X(_09183_));
 sg13g2_o21ai_1 _15912_ (.B1(\cpu.spi.r_searching ),
    .Y(_09184_),
    .A1(\cpu.spi.r_timeout_count[7] ),
    .A2(_09183_));
 sg13g2_nand2_1 _15913_ (.Y(_09185_),
    .A(_09177_),
    .B(_09184_));
 sg13g2_buf_1 _15914_ (.A(\cpu.spi.r_in[3] ),
    .X(_09186_));
 sg13g2_buf_1 _15915_ (.A(\cpu.spi.r_in[6] ),
    .X(_09187_));
 sg13g2_buf_1 _15916_ (.A(\cpu.spi.r_in[1] ),
    .X(_09188_));
 sg13g2_buf_1 _15917_ (.A(\cpu.spi.r_in[0] ),
    .X(_09189_));
 sg13g2_nand2_1 _15918_ (.Y(_09190_),
    .A(_09188_),
    .B(_09189_));
 sg13g2_nand3_1 _15919_ (.B(_09187_),
    .C(_09190_),
    .A(_09186_),
    .Y(_09191_));
 sg13g2_buf_1 _15920_ (.A(\cpu.spi.r_in[2] ),
    .X(_09192_));
 sg13g2_buf_1 _15921_ (.A(\cpu.spi.r_in[5] ),
    .X(_09193_));
 sg13g2_buf_1 _15922_ (.A(\cpu.spi.r_in[4] ),
    .X(_09194_));
 sg13g2_nand4_1 _15923_ (.B(_09193_),
    .C(_09194_),
    .A(_09192_),
    .Y(_09195_),
    .D(\cpu.spi.r_in[7] ));
 sg13g2_nor2_1 _15924_ (.A(_09191_),
    .B(_09195_),
    .Y(_09196_));
 sg13g2_o21ai_1 _15925_ (.B1(\cpu.spi.r_searching ),
    .Y(_09197_),
    .A1(_00202_),
    .A2(_09196_));
 sg13g2_nand2_1 _15926_ (.Y(_09198_),
    .A(_09185_),
    .B(_09197_));
 sg13g2_buf_1 _15927_ (.A(\cpu.spi.r_count[7] ),
    .X(_09199_));
 sg13g2_buf_1 _15928_ (.A(\cpu.spi.r_count[3] ),
    .X(_09200_));
 sg13g2_buf_1 _15929_ (.A(\cpu.spi.r_count[0] ),
    .X(_09201_));
 sg13g2_nor2_1 _15930_ (.A(_09201_),
    .B(\cpu.spi.r_count[1] ),
    .Y(_09202_));
 sg13g2_nand2b_1 _15931_ (.Y(_09203_),
    .B(_09202_),
    .A_N(\cpu.spi.r_count[2] ));
 sg13g2_nor3_1 _15932_ (.A(_09200_),
    .B(\cpu.spi.r_count[4] ),
    .C(_09203_),
    .Y(_09204_));
 sg13g2_nor2b_1 _15933_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09204_),
    .Y(_09205_));
 sg13g2_nor2b_1 _15934_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09205_),
    .Y(_09206_));
 sg13g2_buf_1 _15935_ (.A(_09206_),
    .X(_09207_));
 sg13g2_nor2b_1 _15936_ (.A(_09199_),
    .B_N(_09207_),
    .Y(_09208_));
 sg13g2_buf_1 _15937_ (.A(_09208_),
    .X(_09209_));
 sg13g2_buf_1 _15938_ (.A(_09209_),
    .X(_09210_));
 sg13g2_buf_1 _15939_ (.A(net410),
    .X(_09211_));
 sg13g2_nand3_1 _15940_ (.B(_09198_),
    .C(net360),
    .A(net1055),
    .Y(_09212_));
 sg13g2_o21ai_1 _15941_ (.B1(_09212_),
    .Y(_09213_),
    .A1(_09158_),
    .A2(_09172_));
 sg13g2_and2_1 _15942_ (.A(net715),
    .B(_09213_),
    .X(_00030_));
 sg13g2_nand4_1 _15943_ (.B(_09185_),
    .C(_09197_),
    .A(net1055),
    .Y(_09214_),
    .D(net410));
 sg13g2_buf_1 _15944_ (.A(_09214_),
    .X(_09215_));
 sg13g2_buf_1 _15945_ (.A(\cpu.spi.r_state[2] ),
    .X(_09216_));
 sg13g2_buf_1 _15946_ (.A(_09171_),
    .X(_09217_));
 sg13g2_nor2_1 _15947_ (.A(net507),
    .B(_09170_),
    .Y(_09218_));
 sg13g2_buf_1 _15948_ (.A(_09218_),
    .X(_09219_));
 sg13g2_buf_1 _15949_ (.A(_09219_),
    .X(_09220_));
 sg13g2_buf_1 _15950_ (.A(net106),
    .X(_09221_));
 sg13g2_nand2_1 _15951_ (.Y(_09222_),
    .A(net1054),
    .B(net88));
 sg13g2_buf_1 _15952_ (.A(\cpu.spi.r_state[4] ),
    .X(_09223_));
 sg13g2_nand2b_1 _15953_ (.Y(_09224_),
    .B(_09207_),
    .A_N(_09199_));
 sg13g2_buf_2 _15954_ (.A(_09224_),
    .X(_09225_));
 sg13g2_nor3_1 _15955_ (.A(\cpu.spi.r_state[5] ),
    .B(net1125),
    .C(_09225_),
    .Y(_09226_));
 sg13g2_nand2_1 _15956_ (.Y(_09227_),
    .A(_09222_),
    .B(_09226_));
 sg13g2_o21ai_1 _15957_ (.B1(_09227_),
    .Y(_09228_),
    .A1(net1126),
    .A2(net360));
 sg13g2_nand2b_1 _15958_ (.Y(_09229_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_2 _15959_ (.A(_09229_),
    .X(_09230_));
 sg13g2_buf_2 _15960_ (.A(net1053),
    .X(_09231_));
 sg13g2_buf_1 _15961_ (.A(net916),
    .X(_09232_));
 sg13g2_buf_1 _15962_ (.A(net798),
    .X(_09233_));
 sg13g2_a21oi_1 _15963_ (.A1(_09215_),
    .A2(_09228_),
    .Y(_00031_),
    .B1(_09233_));
 sg13g2_inv_1 _15964_ (.Y(_09234_),
    .A(net1127));
 sg13g2_nor2_2 _15965_ (.A(_09234_),
    .B(_09219_),
    .Y(_09235_));
 sg13g2_buf_1 _15966_ (.A(\cpu.spi.r_state[3] ),
    .X(_09236_));
 sg13g2_a21oi_1 _15967_ (.A1(_09158_),
    .A2(_09235_),
    .Y(_09237_),
    .B1(_09236_));
 sg13g2_nor2_1 _15968_ (.A(net916),
    .B(_09211_),
    .Y(_09238_));
 sg13g2_nor2b_1 _15969_ (.A(_09237_),
    .B_N(_09238_),
    .Y(_00032_));
 sg13g2_buf_2 _15970_ (.A(\cpu.spi.r_state[0] ),
    .X(_09239_));
 sg13g2_inv_1 _15971_ (.Y(_09240_),
    .A(_09239_));
 sg13g2_buf_1 _15972_ (.A(net714),
    .X(_09241_));
 sg13g2_buf_1 _15973_ (.A(_09241_),
    .X(_09242_));
 sg13g2_buf_2 _15974_ (.A(_09242_),
    .X(_09243_));
 sg13g2_buf_1 _15975_ (.A(net1128),
    .X(_09244_));
 sg13g2_buf_1 _15976_ (.A(net1052),
    .X(_09245_));
 sg13g2_buf_1 _15977_ (.A(net915),
    .X(_09246_));
 sg13g2_nor3_1 _15978_ (.A(net506),
    .B(net797),
    .C(_09170_),
    .Y(_09247_));
 sg13g2_nand2_1 _15979_ (.Y(_09248_),
    .A(_09085_),
    .B(_09247_));
 sg13g2_nor3_2 _15980_ (.A(_09240_),
    .B(net916),
    .C(_09248_),
    .Y(_09249_));
 sg13g2_a21o_1 _15981_ (.A2(_09238_),
    .A1(_09223_),
    .B1(_09249_),
    .X(_00033_));
 sg13g2_buf_1 _15982_ (.A(net1127),
    .X(_09250_));
 sg13g2_buf_1 _15983_ (.A(net1051),
    .X(_09251_));
 sg13g2_a21oi_1 _15984_ (.A1(net914),
    .A2(_09221_),
    .Y(_09252_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_nor2b_1 _15985_ (.A(_09252_),
    .B_N(_09238_),
    .Y(_00034_));
 sg13g2_buf_1 _15986_ (.A(net916),
    .X(_09253_));
 sg13g2_buf_1 _15987_ (.A(net796),
    .X(_09254_));
 sg13g2_and2_1 _15988_ (.A(_09173_),
    .B(_09225_),
    .X(_09255_));
 sg13g2_a21oi_1 _15989_ (.A1(net1126),
    .A2(net360),
    .Y(_09256_),
    .B1(_09255_));
 sg13g2_nor2_1 _15990_ (.A(net711),
    .B(_09256_),
    .Y(_00035_));
 sg13g2_buf_1 _15991_ (.A(\cpu.ex.r_div_running ),
    .X(_09257_));
 sg13g2_buf_2 _15992_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09258_));
 sg13g2_buf_1 _15993_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09259_));
 sg13g2_buf_1 _15994_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09260_));
 sg13g2_nand2_1 _15995_ (.Y(_09261_),
    .A(\cpu.dec.iready ),
    .B(_00181_));
 sg13g2_or2_1 _15996_ (.X(_09262_),
    .B(_09261_),
    .A(\cpu.ex.r_branch_stall ));
 sg13g2_buf_1 _15997_ (.A(_09262_),
    .X(_09263_));
 sg13g2_nor2_1 _15998_ (.A(_09230_),
    .B(_09263_),
    .Y(_09264_));
 sg13g2_buf_1 _15999_ (.A(_09264_),
    .X(_09265_));
 sg13g2_and2_1 _16000_ (.A(\cpu.dec.div ),
    .B(net710),
    .X(_09266_));
 sg13g2_buf_1 _16001_ (.A(_09266_),
    .X(_09267_));
 sg13g2_and2_1 _16002_ (.A(\cpu.dec.mult ),
    .B(net710),
    .X(_09268_));
 sg13g2_buf_1 _16003_ (.A(_09268_),
    .X(_09269_));
 sg13g2_nor2_1 _16004_ (.A(_09267_),
    .B(_09269_),
    .Y(_09270_));
 sg13g2_buf_2 _16005_ (.A(_09270_),
    .X(_09271_));
 sg13g2_nand2_1 _16006_ (.Y(_09272_),
    .A(_09260_),
    .B(_09271_));
 sg13g2_buf_2 _16007_ (.A(_09272_),
    .X(\cpu.ex.c_mult_off[0] ));
 sg13g2_nor4_2 _16008_ (.A(_09258_),
    .B(_09259_),
    .C(\cpu.ex.r_mult_off[3] ),
    .Y(_09273_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16009_ (.A(net573),
    .X(_09274_));
 sg13g2_buf_1 _16010_ (.A(_09274_),
    .X(_09275_));
 sg13g2_o21ai_1 _16011_ (.B1(_09081_),
    .Y(_09276_),
    .A1(_09257_),
    .A2(net450));
 sg13g2_a21oi_1 _16012_ (.A1(_09257_),
    .A2(_09273_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09276_));
 sg13g2_buf_1 _16013_ (.A(\cpu.ex.r_mult_running ),
    .X(_09277_));
 sg13g2_buf_1 _16014_ (.A(_09269_),
    .X(_09278_));
 sg13g2_o21ai_1 _16015_ (.B1(_09081_),
    .Y(_09279_),
    .A1(net1124),
    .A2(net504));
 sg13g2_a21oi_1 _16016_ (.A1(net1124),
    .A2(_09273_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09279_));
 sg13g2_a21oi_1 _16017_ (.A1(_09239_),
    .A2(_09248_),
    .Y(_09280_),
    .B1(net1053));
 sg13g2_o21ai_1 _16018_ (.B1(_09280_),
    .Y(_00029_),
    .A1(_09225_),
    .A2(_09237_));
 sg13g2_buf_1 _16019_ (.A(\cpu.dcache.flush_write ),
    .X(_09281_));
 sg13g2_buf_8 _16020_ (.A(_08294_),
    .X(_09282_));
 sg13g2_buf_8 _16021_ (.A(_09282_),
    .X(_09283_));
 sg13g2_buf_2 _16022_ (.A(net795),
    .X(_09284_));
 sg13g2_buf_2 _16023_ (.A(net1136),
    .X(_09285_));
 sg13g2_buf_2 _16024_ (.A(_09285_),
    .X(_09286_));
 sg13g2_buf_1 _16025_ (.A(net913),
    .X(_09287_));
 sg13g2_mux4_1 _16026_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net794),
    .X(_09288_));
 sg13g2_mux4_1 _16027_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net794),
    .X(_09289_));
 sg13g2_buf_2 _16028_ (.A(_09285_),
    .X(_09290_));
 sg13g2_mux4_1 _16029_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net912),
    .X(_09291_));
 sg13g2_mux4_1 _16030_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net912),
    .X(_09292_));
 sg13g2_buf_2 _16031_ (.A(_08346_),
    .X(_09293_));
 sg13g2_buf_2 _16032_ (.A(net793),
    .X(_09294_));
 sg13g2_buf_1 _16033_ (.A(net1073),
    .X(_09295_));
 sg13g2_mux4_1 _16034_ (.S0(net708),
    .A0(_09288_),
    .A1(_09289_),
    .A2(_09291_),
    .A3(_09292_),
    .S1(net911),
    .X(_09296_));
 sg13g2_nand2_1 _16035_ (.Y(_09297_),
    .A(net826),
    .B(_09296_));
 sg13g2_buf_1 _16036_ (.A(_08288_),
    .X(_09298_));
 sg13g2_mux4_1 _16037_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(net794),
    .X(_09299_));
 sg13g2_mux4_1 _16038_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(net794),
    .X(_09300_));
 sg13g2_buf_2 _16039_ (.A(_09282_),
    .X(_09301_));
 sg13g2_mux4_1 _16040_ (.S0(_09301_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(_09290_),
    .X(_09302_));
 sg13g2_mux4_1 _16041_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net912),
    .X(_09303_));
 sg13g2_mux4_1 _16042_ (.S0(net708),
    .A0(_09299_),
    .A1(_09300_),
    .A2(_09302_),
    .A3(_09303_),
    .S1(net911),
    .X(_09304_));
 sg13g2_nand2_1 _16043_ (.Y(_09305_),
    .A(_09298_),
    .B(_09304_));
 sg13g2_a21oi_2 _16044_ (.B1(_08524_),
    .Y(_09306_),
    .A2(_09305_),
    .A1(_09297_));
 sg13g2_buf_1 _16045_ (.A(_09306_),
    .X(_09307_));
 sg13g2_buf_1 _16046_ (.A(_00208_),
    .X(_09308_));
 sg13g2_buf_1 _16047_ (.A(_09308_),
    .X(_09309_));
 sg13g2_inv_2 _16048_ (.Y(_09310_),
    .A(net1050));
 sg13g2_mux2_1 _16049_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(\cpu.dcache.r_tag[3][19] ),
    .S(_09163_),
    .X(_09311_));
 sg13g2_nor2b_1 _16050_ (.A(net1059),
    .B_N(net1056),
    .Y(_09312_));
 sg13g2_buf_1 _16051_ (.A(_09312_),
    .X(_09313_));
 sg13g2_buf_1 _16052_ (.A(_09313_),
    .X(_09314_));
 sg13g2_a22oi_1 _16053_ (.Y(_09315_),
    .B1(net706),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(_09311_),
    .A1(net801));
 sg13g2_nor2_1 _16054_ (.A(_09310_),
    .B(_09315_),
    .Y(_09316_));
 sg13g2_buf_1 _16055_ (.A(\cpu.addr[4] ),
    .X(_09317_));
 sg13g2_inv_1 _16056_ (.Y(_09318_),
    .A(_09317_));
 sg13g2_buf_1 _16057_ (.A(_09318_),
    .X(_09319_));
 sg13g2_mux2_1 _16058_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(\cpu.dcache.r_tag[7][19] ),
    .S(net799),
    .X(_09320_));
 sg13g2_nor2_1 _16059_ (.A(net1059),
    .B(net917),
    .Y(_09321_));
 sg13g2_buf_1 _16060_ (.A(_09321_),
    .X(_09322_));
 sg13g2_a22oi_1 _16061_ (.Y(_09323_),
    .B1(_09322_),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(_09320_),
    .A1(net801));
 sg13g2_inv_1 _16062_ (.Y(_09324_),
    .A(_00230_));
 sg13g2_and2_1 _16063_ (.A(net1129),
    .B(_09308_),
    .X(_09325_));
 sg13g2_buf_2 _16064_ (.A(_09325_),
    .X(_09326_));
 sg13g2_or2_1 _16065_ (.X(_09327_),
    .B(_09159_),
    .A(net1123));
 sg13g2_buf_2 _16066_ (.A(_09327_),
    .X(_09328_));
 sg13g2_nor2_1 _16067_ (.A(_09326_),
    .B(_09328_),
    .Y(_09329_));
 sg13g2_buf_1 _16068_ (.A(_09329_),
    .X(_09330_));
 sg13g2_buf_1 _16069_ (.A(_09330_),
    .X(_09331_));
 sg13g2_nor2b_1 _16070_ (.A(net1129),
    .B_N(net1123),
    .Y(_09332_));
 sg13g2_buf_1 _16071_ (.A(_09332_),
    .X(_09333_));
 sg13g2_and2_1 _16072_ (.A(net1056),
    .B(_09333_),
    .X(_09334_));
 sg13g2_buf_1 _16073_ (.A(_09334_),
    .X(_09335_));
 sg13g2_buf_1 _16074_ (.A(_09335_),
    .X(_09336_));
 sg13g2_a22oi_1 _16075_ (.Y(_09337_),
    .B1(net631),
    .B2(\cpu.dcache.r_tag[6][19] ),
    .A2(net632),
    .A1(_09324_));
 sg13g2_o21ai_1 _16076_ (.B1(_09337_),
    .Y(_09338_),
    .A1(net910),
    .A2(_09323_));
 sg13g2_nor2_1 _16077_ (.A(_09316_),
    .B(_09338_),
    .Y(_09339_));
 sg13g2_xnor2_1 _16078_ (.Y(_09340_),
    .A(net409),
    .B(_09339_));
 sg13g2_mux4_1 _16079_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net912),
    .X(_09341_));
 sg13g2_mux4_1 _16080_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net912),
    .X(_09342_));
 sg13g2_buf_2 _16081_ (.A(_09282_),
    .X(_09343_));
 sg13g2_buf_1 _16082_ (.A(_09285_),
    .X(_09344_));
 sg13g2_mux4_1 _16083_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net909),
    .X(_09345_));
 sg13g2_mux4_1 _16084_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net909),
    .X(_09346_));
 sg13g2_mux4_1 _16085_ (.S0(net793),
    .A0(_09341_),
    .A1(_09342_),
    .A2(_09345_),
    .A3(_09346_),
    .S1(net911),
    .X(_09347_));
 sg13g2_nand2_1 _16086_ (.Y(_09348_),
    .A(_08311_),
    .B(_09347_));
 sg13g2_mux4_1 _16087_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(_09344_),
    .X(_09349_));
 sg13g2_mux4_1 _16088_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net909),
    .X(_09350_));
 sg13g2_buf_8 _16089_ (.A(_09282_),
    .X(_09351_));
 sg13g2_buf_1 _16090_ (.A(_09285_),
    .X(_09352_));
 sg13g2_mux4_1 _16091_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net908),
    .X(_09353_));
 sg13g2_mux4_1 _16092_ (.S0(_09351_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(_09352_),
    .X(_09354_));
 sg13g2_mux4_1 _16093_ (.S0(_09293_),
    .A0(_09349_),
    .A1(_09350_),
    .A2(_09353_),
    .A3(_09354_),
    .S1(_09295_),
    .X(_09355_));
 sg13g2_nand2_1 _16094_ (.Y(_09356_),
    .A(net707),
    .B(_09355_));
 sg13g2_a21oi_2 _16095_ (.B1(_08524_),
    .Y(_09357_),
    .A2(_09356_),
    .A1(_09348_));
 sg13g2_nand2_1 _16096_ (.Y(_09358_),
    .A(_00228_),
    .B(_09331_));
 sg13g2_inv_1 _16097_ (.Y(_09359_),
    .A(_09358_));
 sg13g2_nand2_1 _16098_ (.Y(_09360_),
    .A(_09139_),
    .B(_09308_));
 sg13g2_nor2_1 _16099_ (.A(net1123),
    .B(_09160_),
    .Y(_09361_));
 sg13g2_buf_2 _16100_ (.A(_09361_),
    .X(_09362_));
 sg13g2_nand2_1 _16101_ (.Y(_09363_),
    .A(_09360_),
    .B(_09362_));
 sg13g2_buf_2 _16102_ (.A(_09363_),
    .X(_09364_));
 sg13g2_nor2b_1 _16103_ (.A(net1129),
    .B_N(_09308_),
    .Y(_09365_));
 sg13g2_and2_1 _16104_ (.A(net917),
    .B(_09365_),
    .X(_09366_));
 sg13g2_buf_1 _16105_ (.A(_09366_),
    .X(_09367_));
 sg13g2_a22oi_1 _16106_ (.Y(_09368_),
    .B1(_09367_),
    .B2(\cpu.dcache.r_tag[2][17] ),
    .A2(_09335_),
    .A1(\cpu.dcache.r_tag[6][17] ));
 sg13g2_nand2_1 _16107_ (.Y(_09369_),
    .A(net1129),
    .B(net1123));
 sg13g2_nor2_1 _16108_ (.A(net917),
    .B(_09369_),
    .Y(_09370_));
 sg13g2_buf_1 _16109_ (.A(net1056),
    .X(_09371_));
 sg13g2_nor2_1 _16110_ (.A(net907),
    .B(_09360_),
    .Y(_09372_));
 sg13g2_a22oi_1 _16111_ (.Y(_09373_),
    .B1(_09372_),
    .B2(\cpu.dcache.r_tag[1][17] ),
    .A2(_09370_),
    .A1(\cpu.dcache.r_tag[5][17] ));
 sg13g2_inv_1 _16112_ (.Y(_09374_),
    .A(net1056));
 sg13g2_and2_1 _16113_ (.A(_09374_),
    .B(_09333_),
    .X(_09375_));
 sg13g2_buf_1 _16114_ (.A(_09375_),
    .X(_09376_));
 sg13g2_nor2_1 _16115_ (.A(_09374_),
    .B(_09369_),
    .Y(_09377_));
 sg13g2_and3_1 _16116_ (.X(_09378_),
    .A(_09138_),
    .B(_09160_),
    .C(_09308_));
 sg13g2_buf_1 _16117_ (.A(_09378_),
    .X(_09379_));
 sg13g2_and2_1 _16118_ (.A(\cpu.dcache.r_tag[3][17] ),
    .B(_09379_),
    .X(_09380_));
 sg13g2_a221oi_1 _16119_ (.B2(\cpu.dcache.r_tag[7][17] ),
    .C1(_09380_),
    .B1(_09377_),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .Y(_09381_),
    .A2(_09376_));
 sg13g2_and4_1 _16120_ (.A(_09364_),
    .B(_09368_),
    .C(_09373_),
    .D(_09381_),
    .X(_09382_));
 sg13g2_buf_1 _16121_ (.A(_09382_),
    .X(_09383_));
 sg13g2_or3_1 _16122_ (.A(_09357_),
    .B(_09359_),
    .C(_09383_),
    .X(_09384_));
 sg13g2_buf_1 _16123_ (.A(_09357_),
    .X(_09385_));
 sg13g2_o21ai_1 _16124_ (.B1(net449),
    .Y(_09386_),
    .A1(_09359_),
    .A2(_09383_));
 sg13g2_buf_1 _16125_ (.A(_09374_),
    .X(_09387_));
 sg13g2_inv_1 _16126_ (.Y(_09388_),
    .A(\cpu.dcache.r_tag[2][22] ));
 sg13g2_nand3b_1 _16127_ (.B(net1056),
    .C(_09308_),
    .Y(_09389_),
    .A_N(net1129));
 sg13g2_buf_2 _16128_ (.A(_09389_),
    .X(_09390_));
 sg13g2_nand4_1 _16129_ (.B(net917),
    .C(net1050),
    .A(net1059),
    .Y(_09391_),
    .D(\cpu.dcache.r_tag[3][22] ));
 sg13g2_o21ai_1 _16130_ (.B1(_09391_),
    .Y(_09392_),
    .A1(_09388_),
    .A2(_09390_));
 sg13g2_inv_1 _16131_ (.Y(_09393_),
    .A(\cpu.dcache.r_tag[5][22] ));
 sg13g2_nand3b_1 _16132_ (.B(net1123),
    .C(net1129),
    .Y(_09394_),
    .A_N(_09159_));
 sg13g2_buf_2 _16133_ (.A(_09394_),
    .X(_09395_));
 sg13g2_nand4_1 _16134_ (.B(net1123),
    .C(net917),
    .A(net1059),
    .Y(_09396_),
    .D(\cpu.dcache.r_tag[7][22] ));
 sg13g2_o21ai_1 _16135_ (.B1(_09396_),
    .Y(_09397_),
    .A1(_09393_),
    .A2(_09395_));
 sg13g2_inv_1 _16136_ (.Y(_09398_),
    .A(\cpu.dcache.r_tag[6][22] ));
 sg13g2_nand3b_1 _16137_ (.B(net1123),
    .C(net1056),
    .Y(_09399_),
    .A_N(net1129));
 sg13g2_buf_2 _16138_ (.A(_09399_),
    .X(_09400_));
 sg13g2_nor2_1 _16139_ (.A(_09398_),
    .B(_09400_),
    .Y(_09401_));
 sg13g2_and3_1 _16140_ (.X(_09402_),
    .A(_09374_),
    .B(\cpu.dcache.r_tag[4][22] ),
    .C(_09333_));
 sg13g2_nor4_1 _16141_ (.A(_09392_),
    .B(_09397_),
    .C(_09401_),
    .D(_09402_),
    .Y(_09403_));
 sg13g2_nor2_1 _16142_ (.A(\cpu.dcache.r_tag[0][22] ),
    .B(_09328_),
    .Y(_09404_));
 sg13g2_a221oi_1 _16143_ (.B2(_09403_),
    .C1(_09404_),
    .B1(_09328_),
    .A1(net789),
    .Y(_09405_),
    .A2(_09326_));
 sg13g2_inv_1 _16144_ (.Y(_09406_),
    .A(\cpu.dcache.r_tag[1][22] ));
 sg13g2_nand2_1 _16145_ (.Y(_09407_),
    .A(net789),
    .B(_09326_));
 sg13g2_buf_1 _16146_ (.A(_09407_),
    .X(_09408_));
 sg13g2_a21oi_1 _16147_ (.A1(_09406_),
    .A2(_09403_),
    .Y(_09409_),
    .B1(_09408_));
 sg13g2_mux4_1 _16148_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net913),
    .X(_09410_));
 sg13g2_mux4_1 _16149_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(net913),
    .X(_09411_));
 sg13g2_mux4_1 _16150_ (.S0(_09282_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(_09285_),
    .X(_09412_));
 sg13g2_mux4_1 _16151_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net913),
    .X(_09413_));
 sg13g2_mux4_1 _16152_ (.S0(_08346_),
    .A0(_09410_),
    .A1(_09411_),
    .A2(_09412_),
    .A3(_09413_),
    .S1(net1073),
    .X(_09414_));
 sg13g2_mux4_1 _16153_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net913),
    .X(_09415_));
 sg13g2_mux4_1 _16154_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(net913),
    .X(_09416_));
 sg13g2_mux4_1 _16155_ (.S0(_09282_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(_09285_),
    .X(_09417_));
 sg13g2_mux4_1 _16156_ (.S0(_09282_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(_09285_),
    .X(_09418_));
 sg13g2_mux4_1 _16157_ (.S0(_08346_),
    .A0(_09415_),
    .A1(_09416_),
    .A2(_09417_),
    .A3(_09418_),
    .S1(net1073),
    .X(_09419_));
 sg13g2_mux2_1 _16158_ (.A0(_09414_),
    .A1(_09419_),
    .S(_08288_),
    .X(_09420_));
 sg13g2_nand2b_1 _16159_ (.Y(_09421_),
    .B(_09420_),
    .A_N(_08524_));
 sg13g2_buf_1 _16160_ (.A(_09421_),
    .X(_09422_));
 sg13g2_o21ai_1 _16161_ (.B1(_09422_),
    .Y(_09423_),
    .A1(_09405_),
    .A2(_09409_));
 sg13g2_or3_1 _16162_ (.A(_09422_),
    .B(_09405_),
    .C(_09409_),
    .X(_09424_));
 sg13g2_nand4_1 _16163_ (.B(_09386_),
    .C(_09423_),
    .A(_09384_),
    .Y(_09425_),
    .D(_09424_));
 sg13g2_buf_2 _16164_ (.A(net708),
    .X(_09426_));
 sg13g2_buf_2 _16165_ (.A(net790),
    .X(_09427_));
 sg13g2_buf_2 _16166_ (.A(net908),
    .X(_09428_));
 sg13g2_mux4_1 _16167_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net788),
    .X(_09429_));
 sg13g2_mux4_1 _16168_ (.S0(_09427_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(net788),
    .X(_09430_));
 sg13g2_buf_2 _16169_ (.A(_09285_),
    .X(_09431_));
 sg13g2_buf_1 _16170_ (.A(net906),
    .X(_09432_));
 sg13g2_mux4_1 _16171_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net787),
    .X(_09433_));
 sg13g2_mux4_1 _16172_ (.S0(_09427_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(net788),
    .X(_09434_));
 sg13g2_buf_1 _16173_ (.A(_08299_),
    .X(_09435_));
 sg13g2_mux4_1 _16174_ (.S0(_08288_),
    .A0(_09429_),
    .A1(_09430_),
    .A2(_09433_),
    .A3(_09434_),
    .S1(net905),
    .X(_09436_));
 sg13g2_nand3_1 _16175_ (.B(net630),
    .C(_09436_),
    .A(net1135),
    .Y(_09437_));
 sg13g2_buf_1 _16176_ (.A(_09437_),
    .X(_09438_));
 sg13g2_buf_2 _16177_ (.A(_09343_),
    .X(_09439_));
 sg13g2_buf_2 _16178_ (.A(_09290_),
    .X(_09440_));
 sg13g2_mux4_1 _16179_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net786),
    .X(_09441_));
 sg13g2_mux4_1 _16180_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(_09440_),
    .X(_09442_));
 sg13g2_mux4_1 _16181_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net788),
    .X(_09443_));
 sg13g2_mux4_1 _16182_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net788),
    .X(_09444_));
 sg13g2_mux4_1 _16183_ (.S0(_08288_),
    .A0(_09441_),
    .A1(_09442_),
    .A2(_09443_),
    .A3(_09444_),
    .S1(net905),
    .X(_09445_));
 sg13g2_buf_1 _16184_ (.A(net1076),
    .X(_09446_));
 sg13g2_o21ai_1 _16185_ (.B1(net904),
    .Y(_09447_),
    .A1(_08744_),
    .A2(_09445_));
 sg13g2_mux2_1 _16186_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(\cpu.dcache.r_tag[3][15] ),
    .S(net799),
    .X(_09448_));
 sg13g2_a22oi_1 _16187_ (.Y(_09449_),
    .B1(_09448_),
    .B2(net801),
    .A2(_09313_),
    .A1(\cpu.dcache.r_tag[2][15] ));
 sg13g2_nand2b_1 _16188_ (.Y(_09450_),
    .B(net1050),
    .A_N(_09449_));
 sg13g2_mux2_1 _16189_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(\cpu.dcache.r_tag[7][15] ),
    .S(net799),
    .X(_09451_));
 sg13g2_a22oi_1 _16190_ (.Y(_09452_),
    .B1(_09451_),
    .B2(net801),
    .A2(net705),
    .A1(\cpu.dcache.r_tag[4][15] ));
 sg13g2_buf_1 _16191_ (.A(net1123),
    .X(_09453_));
 sg13g2_buf_1 _16192_ (.A(net1049),
    .X(_09454_));
 sg13g2_nand2b_1 _16193_ (.Y(_09455_),
    .B(net903),
    .A_N(_09452_));
 sg13g2_inv_1 _16194_ (.Y(_09456_),
    .A(_00226_));
 sg13g2_a22oi_1 _16195_ (.Y(_09457_),
    .B1(net631),
    .B2(\cpu.dcache.r_tag[6][15] ),
    .A2(_09330_),
    .A1(_09456_));
 sg13g2_nand3_1 _16196_ (.B(_09455_),
    .C(_09457_),
    .A(_09450_),
    .Y(_09458_));
 sg13g2_a21oi_1 _16197_ (.A1(_09438_),
    .A2(_09447_),
    .Y(_09459_),
    .B1(_09458_));
 sg13g2_nand3_1 _16198_ (.B(_09438_),
    .C(_09447_),
    .A(_09458_),
    .Y(_09460_));
 sg13g2_buf_2 _16199_ (.A(_09282_),
    .X(_09461_));
 sg13g2_buf_8 _16200_ (.A(net785),
    .X(_09462_));
 sg13g2_mux4_1 _16201_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net787),
    .X(_09463_));
 sg13g2_mux4_1 _16202_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net787),
    .X(_09464_));
 sg13g2_buf_2 _16203_ (.A(net795),
    .X(_09465_));
 sg13g2_buf_1 _16204_ (.A(net913),
    .X(_09466_));
 sg13g2_mux4_1 _16205_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net784),
    .X(_09467_));
 sg13g2_mux4_1 _16206_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net784),
    .X(_09468_));
 sg13g2_mux4_1 _16207_ (.S0(net708),
    .A0(_09463_),
    .A1(_09464_),
    .A2(_09467_),
    .A3(_09468_),
    .S1(net905),
    .X(_09469_));
 sg13g2_nand2_1 _16208_ (.Y(_09470_),
    .A(net826),
    .B(_09469_));
 sg13g2_mux4_1 _16209_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(net784),
    .X(_09471_));
 sg13g2_mux4_1 _16210_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(net784),
    .X(_09472_));
 sg13g2_mux4_1 _16211_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net794),
    .X(_09473_));
 sg13g2_mux4_1 _16212_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net784),
    .X(_09474_));
 sg13g2_mux4_1 _16213_ (.S0(net708),
    .A0(_09471_),
    .A1(_09472_),
    .A2(_09473_),
    .A3(_09474_),
    .S1(net905),
    .X(_09475_));
 sg13g2_nand2_1 _16214_ (.Y(_09476_),
    .A(_09298_),
    .B(_09475_));
 sg13g2_a21oi_2 _16215_ (.B1(_08524_),
    .Y(_09477_),
    .A2(_09476_),
    .A1(_09470_));
 sg13g2_buf_1 _16216_ (.A(_09367_),
    .X(_09478_));
 sg13g2_buf_1 _16217_ (.A(_09370_),
    .X(_09479_));
 sg13g2_a22oi_1 _16218_ (.Y(_09480_),
    .B1(net700),
    .B2(\cpu.dcache.r_tag[5][23] ),
    .A2(net629),
    .A1(\cpu.dcache.r_tag[2][23] ));
 sg13g2_buf_1 _16219_ (.A(_09372_),
    .X(_09481_));
 sg13g2_a22oi_1 _16220_ (.Y(_09482_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[1][23] ),
    .A2(net631),
    .A1(\cpu.dcache.r_tag[6][23] ));
 sg13g2_buf_1 _16221_ (.A(_09379_),
    .X(_09483_));
 sg13g2_buf_1 _16222_ (.A(_09377_),
    .X(_09484_));
 sg13g2_a22oi_1 _16223_ (.Y(_09485_),
    .B1(net697),
    .B2(\cpu.dcache.r_tag[7][23] ),
    .A2(net698),
    .A1(\cpu.dcache.r_tag[3][23] ));
 sg13g2_inv_1 _16224_ (.Y(_09486_),
    .A(_00231_));
 sg13g2_buf_1 _16225_ (.A(_09376_),
    .X(_09487_));
 sg13g2_a22oi_1 _16226_ (.Y(_09488_),
    .B1(net628),
    .B2(\cpu.dcache.r_tag[4][23] ),
    .A2(_09330_),
    .A1(_09486_));
 sg13g2_nand4_1 _16227_ (.B(_09482_),
    .C(_09485_),
    .A(_09480_),
    .Y(_09489_),
    .D(_09488_));
 sg13g2_xnor2_1 _16228_ (.Y(_09490_),
    .A(_09477_),
    .B(_09489_));
 sg13g2_nand3b_1 _16229_ (.B(_09460_),
    .C(_09490_),
    .Y(_09491_),
    .A_N(_09459_));
 sg13g2_buf_1 _16230_ (.A(_09435_),
    .X(_09492_));
 sg13g2_inv_1 _16231_ (.Y(_09493_),
    .A(net783));
 sg13g2_mux4_1 _16232_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(net786),
    .X(_09494_));
 sg13g2_mux4_1 _16233_ (.S0(_09439_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(net786),
    .X(_09495_));
 sg13g2_mux4_1 _16234_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(_09428_),
    .X(_09496_));
 sg13g2_mux4_1 _16235_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(_09428_),
    .X(_09497_));
 sg13g2_mux4_1 _16236_ (.S0(_08288_),
    .A0(_09494_),
    .A1(_09495_),
    .A2(_09496_),
    .A3(_09497_),
    .S1(net1076),
    .X(_09498_));
 sg13g2_nand3_1 _16237_ (.B(_09493_),
    .C(_09498_),
    .A(net1070),
    .Y(_09499_));
 sg13g2_buf_1 _16238_ (.A(_09499_),
    .X(_09500_));
 sg13g2_mux4_1 _16239_ (.S0(_09439_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net786),
    .X(_09501_));
 sg13g2_mux4_1 _16240_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net786),
    .X(_09502_));
 sg13g2_mux4_1 _16241_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net786),
    .X(_09503_));
 sg13g2_mux4_1 _16242_ (.S0(net703),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(net786),
    .X(_09504_));
 sg13g2_mux4_1 _16243_ (.S0(_08288_),
    .A0(_09501_),
    .A1(_09502_),
    .A2(_09503_),
    .A3(_09504_),
    .S1(_08291_),
    .X(_09505_));
 sg13g2_o21ai_1 _16244_ (.B1(net783),
    .Y(_09506_),
    .A1(_08744_),
    .A2(_09505_));
 sg13g2_nand2b_1 _16245_ (.Y(_09507_),
    .B(net632),
    .A_N(_00225_));
 sg13g2_a22oi_1 _16246_ (.Y(_09508_),
    .B1(_09481_),
    .B2(\cpu.dcache.r_tag[1][14] ),
    .A2(net698),
    .A1(\cpu.dcache.r_tag[3][14] ));
 sg13g2_a22oi_1 _16247_ (.Y(_09509_),
    .B1(net700),
    .B2(\cpu.dcache.r_tag[5][14] ),
    .A2(net629),
    .A1(\cpu.dcache.r_tag[2][14] ));
 sg13g2_and2_1 _16248_ (.A(net1059),
    .B(net1056),
    .X(_09510_));
 sg13g2_buf_1 _16249_ (.A(_09510_),
    .X(_09511_));
 sg13g2_mux2_1 _16250_ (.A0(\cpu.dcache.r_tag[4][14] ),
    .A1(\cpu.dcache.r_tag[6][14] ),
    .S(net907),
    .X(_09512_));
 sg13g2_inv_2 _16251_ (.Y(_09513_),
    .A(net1059));
 sg13g2_a22oi_1 _16252_ (.Y(_09514_),
    .B1(_09512_),
    .B2(_09513_),
    .A2(_09511_),
    .A1(\cpu.dcache.r_tag[7][14] ));
 sg13g2_nand2b_1 _16253_ (.Y(_09515_),
    .B(_09454_),
    .A_N(_09514_));
 sg13g2_nand4_1 _16254_ (.B(_09508_),
    .C(_09509_),
    .A(_09507_),
    .Y(_09516_),
    .D(_09515_));
 sg13g2_a21oi_1 _16255_ (.A1(_09500_),
    .A2(_09506_),
    .Y(_09517_),
    .B1(_09516_));
 sg13g2_nand3_1 _16256_ (.B(_09500_),
    .C(_09506_),
    .A(_09516_),
    .Y(_09518_));
 sg13g2_mux4_1 _16257_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net906),
    .X(_09519_));
 sg13g2_mux4_1 _16258_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net906),
    .X(_09520_));
 sg13g2_mux4_1 _16259_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(net906),
    .X(_09521_));
 sg13g2_mux4_1 _16260_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net906),
    .X(_09522_));
 sg13g2_mux4_1 _16261_ (.S0(net793),
    .A0(_09519_),
    .A1(_09520_),
    .A2(_09521_),
    .A3(_09522_),
    .S1(net911),
    .X(_09523_));
 sg13g2_nand2_1 _16262_ (.Y(_09524_),
    .A(net826),
    .B(_09523_));
 sg13g2_mux4_1 _16263_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net906),
    .X(_09525_));
 sg13g2_mux4_1 _16264_ (.S0(_09461_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(_09431_),
    .X(_09526_));
 sg13g2_mux4_1 _16265_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(_09286_),
    .X(_09527_));
 sg13g2_mux4_1 _16266_ (.S0(_09461_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(_09431_),
    .X(_09528_));
 sg13g2_mux4_1 _16267_ (.S0(net793),
    .A0(_09525_),
    .A1(_09526_),
    .A2(_09527_),
    .A3(_09528_),
    .S1(net911),
    .X(_09529_));
 sg13g2_nand2_1 _16268_ (.Y(_09530_),
    .A(net707),
    .B(_09529_));
 sg13g2_a21oi_2 _16269_ (.B1(_08524_),
    .Y(_09531_),
    .A2(_09530_),
    .A1(_09524_));
 sg13g2_buf_2 _16270_ (.A(_09531_),
    .X(_09532_));
 sg13g2_nand2b_1 _16271_ (.Y(_09533_),
    .B(net632),
    .A_N(_00229_));
 sg13g2_a22oi_1 _16272_ (.Y(_09534_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[1][18] ),
    .A2(net698),
    .A1(\cpu.dcache.r_tag[3][18] ));
 sg13g2_a22oi_1 _16273_ (.Y(_09535_),
    .B1(net700),
    .B2(\cpu.dcache.r_tag[5][18] ),
    .A2(net629),
    .A1(\cpu.dcache.r_tag[2][18] ));
 sg13g2_mux2_1 _16274_ (.A0(\cpu.dcache.r_tag[4][18] ),
    .A1(\cpu.dcache.r_tag[6][18] ),
    .S(net799),
    .X(_09536_));
 sg13g2_buf_1 _16275_ (.A(_09513_),
    .X(_09537_));
 sg13g2_a22oi_1 _16276_ (.Y(_09538_),
    .B1(_09536_),
    .B2(net782),
    .A2(_09511_),
    .A1(\cpu.dcache.r_tag[7][18] ));
 sg13g2_nand2b_1 _16277_ (.Y(_09539_),
    .B(_09454_),
    .A_N(_09538_));
 sg13g2_nand4_1 _16278_ (.B(_09534_),
    .C(_09535_),
    .A(_09533_),
    .Y(_09540_),
    .D(_09539_));
 sg13g2_xnor2_1 _16279_ (.Y(_09541_),
    .A(_09532_),
    .B(_09540_));
 sg13g2_nand3b_1 _16280_ (.B(_09518_),
    .C(_09541_),
    .Y(_09542_),
    .A_N(_09517_));
 sg13g2_nor4_1 _16281_ (.A(_09340_),
    .B(_09425_),
    .C(_09491_),
    .D(_09542_),
    .Y(_09543_));
 sg13g2_nand2b_1 _16282_ (.Y(_09544_),
    .B(net632),
    .A_N(_00224_));
 sg13g2_a22oi_1 _16283_ (.Y(_09545_),
    .B1(net628),
    .B2(\cpu.dcache.r_tag[4][13] ),
    .A2(net699),
    .A1(\cpu.dcache.r_tag[1][13] ));
 sg13g2_a22oi_1 _16284_ (.Y(_09546_),
    .B1(_09478_),
    .B2(\cpu.dcache.r_tag[2][13] ),
    .A2(_09483_),
    .A1(\cpu.dcache.r_tag[3][13] ));
 sg13g2_mux2_1 _16285_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(\cpu.dcache.r_tag[7][13] ),
    .S(net713),
    .X(_09547_));
 sg13g2_a22oi_1 _16286_ (.Y(_09548_),
    .B1(_09547_),
    .B2(net801),
    .A2(_09313_),
    .A1(\cpu.dcache.r_tag[6][13] ));
 sg13g2_nand2b_1 _16287_ (.Y(_09549_),
    .B(net903),
    .A_N(_09548_));
 sg13g2_nand4_1 _16288_ (.B(_09545_),
    .C(_09546_),
    .A(_09544_),
    .Y(_09550_),
    .D(_09549_));
 sg13g2_mux4_1 _16289_ (.S0(_09284_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net794),
    .X(_09551_));
 sg13g2_mux4_1 _16290_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(net794),
    .X(_09552_));
 sg13g2_mux4_1 _16291_ (.S0(_09284_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(_09287_),
    .X(_09553_));
 sg13g2_mux4_1 _16292_ (.S0(net709),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net794),
    .X(_09554_));
 sg13g2_mux4_1 _16293_ (.S0(_09294_),
    .A0(_09551_),
    .A1(_09552_),
    .A2(_09553_),
    .A3(_09554_),
    .S1(net905),
    .X(_09555_));
 sg13g2_mux4_1 _16294_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net906),
    .X(_09556_));
 sg13g2_mux4_1 _16295_ (.S0(net785),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net906),
    .X(_09557_));
 sg13g2_mux4_1 _16296_ (.S0(net795),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net913),
    .X(_09558_));
 sg13g2_mux4_1 _16297_ (.S0(_09283_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(_09286_),
    .X(_09559_));
 sg13g2_mux4_1 _16298_ (.S0(net793),
    .A0(_09556_),
    .A1(_09557_),
    .A2(_09558_),
    .A3(_09559_),
    .S1(_08299_),
    .X(_09560_));
 sg13g2_and2_1 _16299_ (.A(_08311_),
    .B(_09560_),
    .X(_09561_));
 sg13g2_a21oi_1 _16300_ (.A1(net707),
    .A2(_09555_),
    .Y(_09562_),
    .B1(_09561_));
 sg13g2_buf_1 _16301_ (.A(net786),
    .X(_09563_));
 sg13g2_nor2_1 _16302_ (.A(net1135),
    .B(net696),
    .Y(_09564_));
 sg13g2_a21oi_1 _16303_ (.A1(_08409_),
    .A2(_09562_),
    .Y(_09565_),
    .B1(_09564_));
 sg13g2_buf_2 _16304_ (.A(_09565_),
    .X(_09566_));
 sg13g2_xor2_1 _16305_ (.B(_09566_),
    .A(_09550_),
    .X(_09567_));
 sg13g2_nand2b_1 _16306_ (.Y(_09568_),
    .B(net632),
    .A_N(_00223_));
 sg13g2_a22oi_1 _16307_ (.Y(_09569_),
    .B1(_09487_),
    .B2(\cpu.dcache.r_tag[4][12] ),
    .A2(net699),
    .A1(\cpu.dcache.r_tag[1][12] ));
 sg13g2_a22oi_1 _16308_ (.Y(_09570_),
    .B1(_09478_),
    .B2(\cpu.dcache.r_tag[2][12] ),
    .A2(_09483_),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_mux2_1 _16309_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(\cpu.dcache.r_tag[7][12] ),
    .S(net713),
    .X(_09571_));
 sg13g2_a22oi_1 _16310_ (.Y(_09572_),
    .B1(_09571_),
    .B2(net714),
    .A2(_09313_),
    .A1(\cpu.dcache.r_tag[6][12] ));
 sg13g2_nand2b_1 _16311_ (.Y(_09573_),
    .B(net903),
    .A_N(_09572_));
 sg13g2_nand4_1 _16312_ (.B(_09569_),
    .C(_09570_),
    .A(_09568_),
    .Y(_09574_),
    .D(_09573_));
 sg13g2_buf_1 _16313_ (.A(net792),
    .X(_09575_));
 sg13g2_inv_1 _16314_ (.Y(_09576_),
    .A(net695));
 sg13g2_mux4_1 _16315_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(net909),
    .X(_09577_));
 sg13g2_mux4_1 _16316_ (.S0(_09343_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(_09344_),
    .X(_09578_));
 sg13g2_mux4_1 _16317_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(net908),
    .X(_09579_));
 sg13g2_mux4_1 _16318_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net908),
    .X(_09580_));
 sg13g2_mux4_1 _16319_ (.S0(_09293_),
    .A0(_09577_),
    .A1(_09578_),
    .A2(_09579_),
    .A3(_09580_),
    .S1(_09295_),
    .X(_09581_));
 sg13g2_mux4_1 _16320_ (.S0(_09351_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(_09352_),
    .X(_09582_));
 sg13g2_mux4_1 _16321_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net908),
    .X(_09583_));
 sg13g2_mux4_1 _16322_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(net908),
    .X(_09584_));
 sg13g2_mux4_1 _16323_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net908),
    .X(_09585_));
 sg13g2_mux4_1 _16324_ (.S0(net793),
    .A0(_09582_),
    .A1(_09583_),
    .A2(_09584_),
    .A3(_09585_),
    .S1(net911),
    .X(_09586_));
 sg13g2_mux2_1 _16325_ (.A0(_09581_),
    .A1(_09586_),
    .S(net707),
    .X(_09587_));
 sg13g2_nand2_1 _16326_ (.Y(_09588_),
    .A(_08320_),
    .B(_09587_));
 sg13g2_o21ai_1 _16327_ (.B1(_09588_),
    .Y(_09589_),
    .A1(_08409_),
    .A2(_09576_));
 sg13g2_buf_1 _16328_ (.A(_09589_),
    .X(_09590_));
 sg13g2_xor2_1 _16329_ (.B(_09590_),
    .A(_09574_),
    .X(_09591_));
 sg13g2_nor2_1 _16330_ (.A(_09567_),
    .B(_09591_),
    .Y(_09592_));
 sg13g2_buf_1 _16331_ (.A(_09408_),
    .X(_09593_));
 sg13g2_buf_1 _16332_ (.A(_09328_),
    .X(_09594_));
 sg13g2_a22oi_1 _16333_ (.Y(_09595_),
    .B1(_09367_),
    .B2(\cpu.dcache.r_tag[2][21] ),
    .A2(_09379_),
    .A1(\cpu.dcache.r_tag[3][21] ));
 sg13g2_a22oi_1 _16334_ (.Y(_09596_),
    .B1(_09479_),
    .B2(\cpu.dcache.r_tag[5][21] ),
    .A2(net631),
    .A1(\cpu.dcache.r_tag[6][21] ));
 sg13g2_a22oi_1 _16335_ (.Y(_09597_),
    .B1(net697),
    .B2(\cpu.dcache.r_tag[7][21] ),
    .A2(_09376_),
    .A1(\cpu.dcache.r_tag[4][21] ));
 sg13g2_and3_1 _16336_ (.X(_09598_),
    .A(_09595_),
    .B(_09596_),
    .C(_09597_));
 sg13g2_buf_1 _16337_ (.A(_09598_),
    .X(_09599_));
 sg13g2_nor2_1 _16338_ (.A(\cpu.dcache.r_tag[0][21] ),
    .B(_09594_),
    .Y(_09600_));
 sg13g2_a21o_1 _16339_ (.A2(_09599_),
    .A1(_09594_),
    .B1(_09600_),
    .X(_09601_));
 sg13g2_nor2_1 _16340_ (.A(\cpu.dcache.r_tag[1][21] ),
    .B(_09408_),
    .Y(_09602_));
 sg13g2_mux4_1 _16341_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net912),
    .X(_09603_));
 sg13g2_mux4_1 _16342_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net912),
    .X(_09604_));
 sg13g2_mux4_1 _16343_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net909),
    .X(_09605_));
 sg13g2_mux4_1 _16344_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net909),
    .X(_09606_));
 sg13g2_mux4_1 _16345_ (.S0(net793),
    .A0(_09603_),
    .A1(_09604_),
    .A2(_09605_),
    .A3(_09606_),
    .S1(net911),
    .X(_09607_));
 sg13g2_nand2_1 _16346_ (.Y(_09608_),
    .A(net826),
    .B(_09607_));
 sg13g2_mux4_1 _16347_ (.S0(_09301_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(net909),
    .X(_09609_));
 sg13g2_mux4_1 _16348_ (.S0(net792),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net912),
    .X(_09610_));
 sg13g2_mux4_1 _16349_ (.S0(net790),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(net908),
    .X(_09611_));
 sg13g2_mux4_1 _16350_ (.S0(net791),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net909),
    .X(_09612_));
 sg13g2_mux4_1 _16351_ (.S0(net793),
    .A0(_09609_),
    .A1(_09610_),
    .A2(_09611_),
    .A3(_09612_),
    .S1(net911),
    .X(_09613_));
 sg13g2_nand2_1 _16352_ (.Y(_09614_),
    .A(net707),
    .B(_09613_));
 sg13g2_a21oi_2 _16353_ (.B1(_08524_),
    .Y(_09615_),
    .A2(_09614_),
    .A1(_09608_));
 sg13g2_buf_2 _16354_ (.A(_09615_),
    .X(_09616_));
 sg13g2_a221oi_1 _16355_ (.B2(_09599_),
    .C1(_09616_),
    .B1(_09602_),
    .A1(_09593_),
    .Y(_09617_),
    .A2(_09601_));
 sg13g2_inv_1 _16356_ (.Y(_09618_),
    .A(_09616_));
 sg13g2_a221oi_1 _16357_ (.B2(_09599_),
    .C1(_09600_),
    .B1(net781),
    .A1(net789),
    .Y(_09619_),
    .A2(_09326_));
 sg13g2_inv_1 _16358_ (.Y(_09620_),
    .A(\cpu.dcache.r_tag[1][21] ));
 sg13g2_a21oi_1 _16359_ (.A1(_09620_),
    .A2(_09599_),
    .Y(_09621_),
    .B1(_09408_));
 sg13g2_nor3_1 _16360_ (.A(_09618_),
    .B(_09619_),
    .C(_09621_),
    .Y(_09622_));
 sg13g2_mux4_1 _16361_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net787),
    .X(_09623_));
 sg13g2_mux4_1 _16362_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net787),
    .X(_09624_));
 sg13g2_mux4_1 _16363_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net784),
    .X(_09625_));
 sg13g2_mux4_1 _16364_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net784),
    .X(_09626_));
 sg13g2_mux4_1 _16365_ (.S0(net708),
    .A0(_09623_),
    .A1(_09624_),
    .A2(_09625_),
    .A3(_09626_),
    .S1(net905),
    .X(_09627_));
 sg13g2_nand2_1 _16366_ (.Y(_09628_),
    .A(net826),
    .B(_09627_));
 sg13g2_mux4_1 _16367_ (.S0(_09465_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(_09466_),
    .X(_09629_));
 sg13g2_mux4_1 _16368_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net784),
    .X(_09630_));
 sg13g2_mux4_1 _16369_ (.S0(_09465_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(_09287_),
    .X(_09631_));
 sg13g2_mux4_1 _16370_ (.S0(net701),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(_09466_),
    .X(_09632_));
 sg13g2_mux4_1 _16371_ (.S0(net708),
    .A0(_09629_),
    .A1(_09630_),
    .A2(_09631_),
    .A3(_09632_),
    .S1(net905),
    .X(_09633_));
 sg13g2_nand2_1 _16372_ (.Y(_09634_),
    .A(net707),
    .B(_09633_));
 sg13g2_a21oi_2 _16373_ (.B1(_08524_),
    .Y(_09635_),
    .A2(_09634_),
    .A1(_09628_));
 sg13g2_buf_1 _16374_ (.A(_09635_),
    .X(_09636_));
 sg13g2_a22oi_1 _16375_ (.Y(_09637_),
    .B1(net629),
    .B2(\cpu.dcache.r_tag[2][20] ),
    .A2(net698),
    .A1(\cpu.dcache.r_tag[3][20] ));
 sg13g2_a22oi_1 _16376_ (.Y(_09638_),
    .B1(net697),
    .B2(\cpu.dcache.r_tag[7][20] ),
    .A2(net699),
    .A1(\cpu.dcache.r_tag[1][20] ));
 sg13g2_mux2_1 _16377_ (.A0(\cpu.dcache.r_tag[4][20] ),
    .A1(\cpu.dcache.r_tag[6][20] ),
    .S(net799),
    .X(_09639_));
 sg13g2_nor2b_1 _16378_ (.A(net917),
    .B_N(net1059),
    .Y(_09640_));
 sg13g2_buf_2 _16379_ (.A(_09640_),
    .X(_09641_));
 sg13g2_a22oi_1 _16380_ (.Y(_09642_),
    .B1(_09641_),
    .B2(\cpu.dcache.r_tag[5][20] ),
    .A2(_09639_),
    .A1(net782));
 sg13g2_nand2b_1 _16381_ (.Y(_09643_),
    .B(net903),
    .A_N(_09642_));
 sg13g2_nand4_1 _16382_ (.B(_09637_),
    .C(_09638_),
    .A(_09364_),
    .Y(_09644_),
    .D(_09643_));
 sg13g2_o21ai_1 _16383_ (.B1(_09644_),
    .Y(_09645_),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .A2(_09364_));
 sg13g2_xnor2_1 _16384_ (.Y(_09646_),
    .A(net406),
    .B(_09645_));
 sg13g2_nor3_1 _16385_ (.A(_09617_),
    .B(_09622_),
    .C(_09646_),
    .Y(_09647_));
 sg13g2_mux4_1 _16386_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(net788),
    .X(_09648_));
 sg13g2_mux4_1 _16387_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net788),
    .X(_09649_));
 sg13g2_mux4_1 _16388_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net787),
    .X(_09650_));
 sg13g2_mux4_1 _16389_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net787),
    .X(_09651_));
 sg13g2_mux4_1 _16390_ (.S0(_09294_),
    .A0(_09648_),
    .A1(_09649_),
    .A2(_09650_),
    .A3(_09651_),
    .S1(net905),
    .X(_09652_));
 sg13g2_nand2_1 _16391_ (.Y(_09653_),
    .A(net826),
    .B(_09652_));
 sg13g2_mux4_1 _16392_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(_09432_),
    .X(_09654_));
 sg13g2_mux4_1 _16393_ (.S0(net704),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net788),
    .X(_09655_));
 sg13g2_mux4_1 _16394_ (.S0(_09462_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(net787),
    .X(_09656_));
 sg13g2_mux4_1 _16395_ (.S0(_09462_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09432_),
    .X(_09657_));
 sg13g2_mux4_1 _16396_ (.S0(net708),
    .A0(_09654_),
    .A1(_09655_),
    .A2(_09656_),
    .A3(_09657_),
    .S1(_09435_),
    .X(_09658_));
 sg13g2_nand2_1 _16397_ (.Y(_09659_),
    .A(net707),
    .B(_09658_));
 sg13g2_a21oi_2 _16398_ (.B1(_08525_),
    .Y(_09660_),
    .A2(_09659_),
    .A1(_09653_));
 sg13g2_buf_1 _16399_ (.A(_09660_),
    .X(_09661_));
 sg13g2_a22oi_1 _16400_ (.Y(_09662_),
    .B1(_09367_),
    .B2(\cpu.dcache.r_tag[2][16] ),
    .A2(net631),
    .A1(\cpu.dcache.r_tag[6][16] ));
 sg13g2_a22oi_1 _16401_ (.Y(_09663_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[1][16] ),
    .A2(_09479_),
    .A1(\cpu.dcache.r_tag[5][16] ));
 sg13g2_and2_1 _16402_ (.A(\cpu.dcache.r_tag[3][16] ),
    .B(_09379_),
    .X(_09664_));
 sg13g2_a221oi_1 _16403_ (.B2(\cpu.dcache.r_tag[7][16] ),
    .C1(_09664_),
    .B1(net697),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .Y(_09665_),
    .A2(_09487_));
 sg13g2_and4_1 _16404_ (.A(_09364_),
    .B(_09662_),
    .C(_09663_),
    .D(_09665_),
    .X(_09666_));
 sg13g2_a21oi_1 _16405_ (.A1(_00227_),
    .A2(net632),
    .Y(_09667_),
    .B1(_09666_));
 sg13g2_nand2_1 _16406_ (.Y(_09668_),
    .A(_09661_),
    .B(_09667_));
 sg13g2_or2_1 _16407_ (.X(_09669_),
    .B(_09667_),
    .A(_09660_));
 sg13g2_nand2_1 _16408_ (.Y(_09670_),
    .A(_00218_),
    .B(_09362_));
 sg13g2_a22oi_1 _16409_ (.Y(_09671_),
    .B1(_09370_),
    .B2(\cpu.dcache.r_tag[5][9] ),
    .A2(net631),
    .A1(\cpu.dcache.r_tag[6][9] ));
 sg13g2_a22oi_1 _16410_ (.Y(_09672_),
    .B1(_09484_),
    .B2(\cpu.dcache.r_tag[7][9] ),
    .A2(_09367_),
    .A1(\cpu.dcache.r_tag[2][9] ));
 sg13g2_a22oi_1 _16411_ (.Y(_09673_),
    .B1(_09376_),
    .B2(\cpu.dcache.r_tag[4][9] ),
    .A2(_09379_),
    .A1(\cpu.dcache.r_tag[3][9] ));
 sg13g2_nand4_1 _16412_ (.B(_09671_),
    .C(_09672_),
    .A(_09328_),
    .Y(_09674_),
    .D(_09673_));
 sg13g2_nand3_1 _16413_ (.B(_09670_),
    .C(_09674_),
    .A(_09408_),
    .Y(_09675_));
 sg13g2_buf_1 _16414_ (.A(_09675_),
    .X(_09676_));
 sg13g2_nand3_1 _16415_ (.B(_09672_),
    .C(_09673_),
    .A(_09671_),
    .Y(_09677_));
 sg13g2_buf_1 _16416_ (.A(net699),
    .X(_09678_));
 sg13g2_o21ai_1 _16417_ (.B1(net627),
    .Y(_09679_),
    .A1(\cpu.dcache.r_tag[1][9] ),
    .A2(_09677_));
 sg13g2_nand3_1 _16418_ (.B(_09676_),
    .C(_09679_),
    .A(_00217_),
    .Y(_09680_));
 sg13g2_a21o_1 _16419_ (.A2(_09679_),
    .A1(_09676_),
    .B1(_00217_),
    .X(_09681_));
 sg13g2_nand3_1 _16420_ (.B(net1050),
    .C(\cpu.dcache.r_tag[1][10] ),
    .A(net918),
    .Y(_09682_));
 sg13g2_nand3b_1 _16421_ (.B(net1049),
    .C(\cpu.dcache.r_tag[4][10] ),
    .Y(_09683_),
    .A_N(net918));
 sg13g2_nand3_1 _16422_ (.B(_09682_),
    .C(_09683_),
    .A(net789),
    .Y(_09684_));
 sg13g2_mux2_1 _16423_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(\cpu.dcache.r_tag[3][10] ),
    .S(net918),
    .X(_09685_));
 sg13g2_a21o_1 _16424_ (.A2(_09685_),
    .A1(net1050),
    .B1(_09387_),
    .X(_09686_));
 sg13g2_mux2_1 _16425_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(\cpu.dcache.r_tag[7][10] ),
    .S(net907),
    .X(_09687_));
 sg13g2_and2_1 _16426_ (.A(net799),
    .B(\cpu.dcache.r_tag[6][10] ),
    .X(_09688_));
 sg13g2_mux2_1 _16427_ (.A0(_09687_),
    .A1(_09688_),
    .S(_09513_),
    .X(_09689_));
 sg13g2_a221oi_1 _16428_ (.B2(net1049),
    .C1(_09331_),
    .B1(_09689_),
    .A1(_09684_),
    .Y(_09690_),
    .A2(_09686_));
 sg13g2_a21o_1 _16429_ (.A2(net632),
    .A1(_00220_),
    .B1(_09690_),
    .X(_09691_));
 sg13g2_xnor2_1 _16430_ (.Y(_09692_),
    .A(_00219_),
    .B(_09691_));
 sg13g2_nand2_1 _16431_ (.Y(_09693_),
    .A(\cpu.dcache.r_tag[7][7] ),
    .B(net697));
 sg13g2_inv_1 _16432_ (.Y(_09694_),
    .A(_00214_));
 sg13g2_a22oi_1 _16433_ (.Y(_09695_),
    .B1(net698),
    .B2(\cpu.dcache.r_tag[3][7] ),
    .A2(_09330_),
    .A1(_09694_));
 sg13g2_a22oi_1 _16434_ (.Y(_09696_),
    .B1(net699),
    .B2(\cpu.dcache.r_tag[1][7] ),
    .A2(net629),
    .A1(\cpu.dcache.r_tag[2][7] ));
 sg13g2_mux2_1 _16435_ (.A0(\cpu.dcache.r_tag[4][7] ),
    .A1(\cpu.dcache.r_tag[6][7] ),
    .S(net907),
    .X(_09697_));
 sg13g2_a22oi_1 _16436_ (.Y(_09698_),
    .B1(_09697_),
    .B2(_09513_),
    .A2(_09641_),
    .A1(\cpu.dcache.r_tag[5][7] ));
 sg13g2_nand2b_1 _16437_ (.Y(_09699_),
    .B(net1049),
    .A_N(_09698_));
 sg13g2_and4_1 _16438_ (.A(_09693_),
    .B(_09695_),
    .C(_09696_),
    .D(_09699_),
    .X(_09700_));
 sg13g2_xnor2_1 _16439_ (.Y(_09701_),
    .A(_00213_),
    .B(_09700_));
 sg13g2_inv_1 _16440_ (.Y(_09702_),
    .A(_00216_));
 sg13g2_a22oi_1 _16441_ (.Y(_09703_),
    .B1(net698),
    .B2(\cpu.dcache.r_tag[3][8] ),
    .A2(_09330_),
    .A1(_09702_));
 sg13g2_nand2_1 _16442_ (.Y(_09704_),
    .A(\cpu.dcache.r_tag[2][8] ),
    .B(net629));
 sg13g2_a22oi_1 _16443_ (.Y(_09705_),
    .B1(_09481_),
    .B2(\cpu.dcache.r_tag[1][8] ),
    .A2(_09336_),
    .A1(\cpu.dcache.r_tag[6][8] ));
 sg13g2_mux2_1 _16444_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(\cpu.dcache.r_tag[7][8] ),
    .S(net907),
    .X(_09706_));
 sg13g2_a22oi_1 _16445_ (.Y(_09707_),
    .B1(_09706_),
    .B2(net801),
    .A2(net705),
    .A1(\cpu.dcache.r_tag[4][8] ));
 sg13g2_nand2b_1 _16446_ (.Y(_09708_),
    .B(net1049),
    .A_N(_09707_));
 sg13g2_and4_1 _16447_ (.A(_09703_),
    .B(_09704_),
    .C(_09705_),
    .D(_09708_),
    .X(_09709_));
 sg13g2_xnor2_1 _16448_ (.Y(_09710_),
    .A(_00215_),
    .B(_09709_));
 sg13g2_mux2_1 _16449_ (.A0(\cpu.dcache.r_tag[4][6] ),
    .A1(\cpu.dcache.r_tag[6][6] ),
    .S(_09161_),
    .X(_09711_));
 sg13g2_a22oi_1 _16450_ (.Y(_09712_),
    .B1(_09711_),
    .B2(_09513_),
    .A2(_09641_),
    .A1(\cpu.dcache.r_tag[5][6] ));
 sg13g2_nor2_1 _16451_ (.A(net910),
    .B(_09712_),
    .Y(_09713_));
 sg13g2_nand3b_1 _16452_ (.B(net907),
    .C(\cpu.dcache.r_tag[2][6] ),
    .Y(_09714_),
    .A_N(net918));
 sg13g2_nand3b_1 _16453_ (.B(\cpu.dcache.r_tag[1][6] ),
    .C(net918),
    .Y(_09715_),
    .A_N(_09161_));
 sg13g2_a21oi_1 _16454_ (.A1(_09714_),
    .A2(_09715_),
    .Y(_09716_),
    .B1(_09310_));
 sg13g2_a22oi_1 _16455_ (.Y(_09717_),
    .B1(\cpu.dcache.r_tag[3][6] ),
    .B2(net1050),
    .A2(\cpu.dcache.r_tag[7][6] ),
    .A1(net1049));
 sg13g2_nor2b_1 _16456_ (.A(_09717_),
    .B_N(_09511_),
    .Y(_09718_));
 sg13g2_nor3_1 _16457_ (.A(_00212_),
    .B(_09326_),
    .C(_09328_),
    .Y(_09719_));
 sg13g2_nor3_1 _16458_ (.A(_09716_),
    .B(_09718_),
    .C(_09719_),
    .Y(_09720_));
 sg13g2_nand3b_1 _16459_ (.B(_09720_),
    .C(_00211_),
    .Y(_09721_),
    .A_N(_09713_));
 sg13g2_or3_1 _16460_ (.A(_09716_),
    .B(_09718_),
    .C(_09719_),
    .X(_09722_));
 sg13g2_inv_1 _16461_ (.Y(_09723_),
    .A(_00211_));
 sg13g2_o21ai_1 _16462_ (.B1(_09723_),
    .Y(_09724_),
    .A1(_09713_),
    .A2(_09722_));
 sg13g2_mux2_1 _16463_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(\cpu.dcache.r_tag[7][11] ),
    .S(net907),
    .X(_09725_));
 sg13g2_a22oi_1 _16464_ (.Y(_09726_),
    .B1(_09725_),
    .B2(net801),
    .A2(_09313_),
    .A1(\cpu.dcache.r_tag[6][11] ));
 sg13g2_nor2_1 _16465_ (.A(_09319_),
    .B(_09726_),
    .Y(_09727_));
 sg13g2_nand3_1 _16466_ (.B(_09309_),
    .C(\cpu.dcache.r_tag[2][11] ),
    .A(net799),
    .Y(_09728_));
 sg13g2_nand3b_1 _16467_ (.B(\cpu.dcache.r_tag[4][11] ),
    .C(net1049),
    .Y(_09729_),
    .A_N(_09371_));
 sg13g2_a21oi_1 _16468_ (.A1(_09728_),
    .A2(_09729_),
    .Y(_09730_),
    .B1(net918));
 sg13g2_nor3_1 _16469_ (.A(_00222_),
    .B(_09326_),
    .C(_09328_),
    .Y(_09731_));
 sg13g2_nand2_1 _16470_ (.Y(_09732_),
    .A(net799),
    .B(\cpu.dcache.r_tag[3][11] ));
 sg13g2_nand2b_1 _16471_ (.Y(_09733_),
    .B(\cpu.dcache.r_tag[1][11] ),
    .A_N(_09371_));
 sg13g2_a21oi_1 _16472_ (.A1(_09732_),
    .A2(_09733_),
    .Y(_09734_),
    .B1(_09360_));
 sg13g2_nor3_1 _16473_ (.A(_09730_),
    .B(_09731_),
    .C(_09734_),
    .Y(_09735_));
 sg13g2_nand3b_1 _16474_ (.B(_09735_),
    .C(_00221_),
    .Y(_09736_),
    .A_N(_09727_));
 sg13g2_or3_1 _16475_ (.A(_09730_),
    .B(_09731_),
    .C(_09734_),
    .X(_09737_));
 sg13g2_inv_1 _16476_ (.Y(_09738_),
    .A(_00221_));
 sg13g2_o21ai_1 _16477_ (.B1(_09738_),
    .Y(_09739_),
    .A1(_09727_),
    .A2(_09737_));
 sg13g2_buf_2 _16478_ (.A(_00209_),
    .X(_09740_));
 sg13g2_inv_2 _16479_ (.Y(_09741_),
    .A(_09740_));
 sg13g2_nand3_1 _16480_ (.B(net1050),
    .C(\cpu.dcache.r_tag[1][5] ),
    .A(net918),
    .Y(_09742_));
 sg13g2_nand3b_1 _16481_ (.B(_09453_),
    .C(\cpu.dcache.r_tag[4][5] ),
    .Y(_09743_),
    .A_N(net918));
 sg13g2_nand3_1 _16482_ (.B(_09742_),
    .C(_09743_),
    .A(_09387_),
    .Y(_09744_));
 sg13g2_mux2_1 _16483_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(\cpu.dcache.r_tag[3][5] ),
    .S(net1059),
    .X(_09745_));
 sg13g2_a21o_1 _16484_ (.A2(_09745_),
    .A1(_09309_),
    .B1(_09374_),
    .X(_09746_));
 sg13g2_mux2_1 _16485_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(\cpu.dcache.r_tag[7][5] ),
    .S(net917),
    .X(_09747_));
 sg13g2_and2_1 _16486_ (.A(net907),
    .B(\cpu.dcache.r_tag[6][5] ),
    .X(_09748_));
 sg13g2_mux2_1 _16487_ (.A0(_09747_),
    .A1(_09748_),
    .S(_09513_),
    .X(_09749_));
 sg13g2_nor3_1 _16488_ (.A(_00210_),
    .B(_09326_),
    .C(_09328_),
    .Y(_09750_));
 sg13g2_a221oi_1 _16489_ (.B2(net1049),
    .C1(_09750_),
    .B1(_09749_),
    .A1(_09744_),
    .Y(_09751_),
    .A2(_09746_));
 sg13g2_xnor2_1 _16490_ (.Y(_09752_),
    .A(_09741_),
    .B(_09751_));
 sg13g2_a221oi_1 _16491_ (.B2(_09739_),
    .C1(_09752_),
    .B1(_09736_),
    .A1(_09721_),
    .Y(_09753_),
    .A2(_09724_));
 sg13g2_nand4_1 _16492_ (.B(_09701_),
    .C(_09710_),
    .A(_09692_),
    .Y(_09754_),
    .D(_09753_));
 sg13g2_a221oi_1 _16493_ (.B2(_09681_),
    .C1(_09754_),
    .B1(_09680_),
    .A1(_09668_),
    .Y(_09755_),
    .A2(_09669_));
 sg13g2_nand4_1 _16494_ (.B(_09592_),
    .C(_09647_),
    .A(_09543_),
    .Y(_09756_),
    .D(_09755_));
 sg13g2_mux4_1 _16495_ (.S0(net714),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net713),
    .X(_09757_));
 sg13g2_mux4_1 _16496_ (.S0(net714),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net713),
    .X(_09758_));
 sg13g2_mux2_1 _16497_ (.A0(_09757_),
    .A1(_09758_),
    .S(net910),
    .X(_09759_));
 sg13g2_mux4_1 _16498_ (.S0(net714),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(net634),
    .X(_09760_));
 sg13g2_mux4_1 _16499_ (.S0(net714),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net713),
    .X(_09761_));
 sg13g2_mux2_1 _16500_ (.A0(_09760_),
    .A1(_09761_),
    .S(net910),
    .X(_09762_));
 sg13g2_and3_1 _16501_ (.X(_09763_),
    .A(_09137_),
    .B(_09759_),
    .C(_09762_));
 sg13g2_o21ai_1 _16502_ (.B1(_09763_),
    .Y(_09764_),
    .A1(_09281_),
    .A2(_09756_));
 sg13g2_buf_2 _16503_ (.A(_09764_),
    .X(_09765_));
 sg13g2_nand2b_1 _16504_ (.Y(_09766_),
    .B(_09759_),
    .A_N(_09756_));
 sg13g2_buf_1 _16505_ (.A(_09766_),
    .X(_09767_));
 sg13g2_nand2b_1 _16506_ (.Y(_09768_),
    .B(_09767_),
    .A_N(_09281_));
 sg13g2_buf_1 _16507_ (.A(_08322_),
    .X(_09769_));
 sg13g2_and2_1 _16508_ (.A(net902),
    .B(_09137_),
    .X(_09770_));
 sg13g2_buf_1 _16509_ (.A(_09770_),
    .X(_09771_));
 sg13g2_inv_1 _16510_ (.Y(_09772_),
    .A(_09771_));
 sg13g2_a21oi_1 _16511_ (.A1(_09765_),
    .A2(_09768_),
    .Y(_09773_),
    .B1(_09772_));
 sg13g2_nand2_1 _16512_ (.Y(_09774_),
    .A(_08339_),
    .B(_09149_));
 sg13g2_a22oi_1 _16513_ (.Y(_09775_),
    .B1(_09773_),
    .B2(_09774_),
    .A2(_08851_),
    .A1(net1137));
 sg13g2_buf_1 _16514_ (.A(_09775_),
    .X(_09776_));
 sg13g2_nand2_1 _16515_ (.Y(_09777_),
    .A(\cpu.qspi.r_state[17] ),
    .B(_09776_));
 sg13g2_buf_1 _16516_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09778_));
 sg13g2_buf_2 _16517_ (.A(\cpu.qspi.r_ind ),
    .X(_09779_));
 sg13g2_buf_1 _16518_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09780_));
 sg13g2_buf_2 _16519_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09781_));
 sg13g2_nor3_1 _16520_ (.A(_09780_),
    .B(_09781_),
    .C(\cpu.qspi.r_count[2] ),
    .Y(_09782_));
 sg13g2_nor2b_1 _16521_ (.A(\cpu.qspi.r_count[3] ),
    .B_N(_09782_),
    .Y(_09783_));
 sg13g2_buf_1 _16522_ (.A(_09783_),
    .X(_09784_));
 sg13g2_and2_1 _16523_ (.A(_00232_),
    .B(_09784_),
    .X(_09785_));
 sg13g2_buf_1 _16524_ (.A(_09785_),
    .X(_09786_));
 sg13g2_buf_1 _16525_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09787_));
 sg13g2_buf_1 _16526_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09788_));
 sg13g2_a221oi_1 _16527_ (.B2(_09787_),
    .C1(_09788_),
    .B1(_09786_),
    .A1(_09778_),
    .Y(_09789_),
    .A2(_09779_));
 sg13g2_a21oi_1 _16528_ (.A1(_09777_),
    .A2(_09789_),
    .Y(_00026_),
    .B1(net712));
 sg13g2_buf_2 _16529_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09790_));
 sg13g2_nand2_1 _16530_ (.Y(_09791_),
    .A(_00232_),
    .B(_09784_));
 sg13g2_buf_1 _16531_ (.A(_09791_),
    .X(_09792_));
 sg13g2_nor2_1 _16532_ (.A(net1137),
    .B(_09765_),
    .Y(_09793_));
 sg13g2_buf_2 _16533_ (.A(_09793_),
    .X(_09794_));
 sg13g2_buf_2 _16534_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09795_));
 sg13g2_a22oi_1 _16535_ (.Y(_09796_),
    .B1(_09794_),
    .B2(_09795_),
    .A2(net626),
    .A1(_09790_));
 sg13g2_nor2_1 _16536_ (.A(net711),
    .B(_09796_),
    .Y(_00025_));
 sg13g2_buf_1 _16537_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09797_));
 sg13g2_buf_1 _16538_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09798_));
 sg13g2_a21oi_1 _16539_ (.A1(_09797_),
    .A2(_09786_),
    .Y(_09799_),
    .B1(_09798_));
 sg13g2_nor2_1 _16540_ (.A(net711),
    .B(_09799_),
    .Y(_00022_));
 sg13g2_buf_1 _16541_ (.A(_00258_),
    .X(_09800_));
 sg13g2_buf_1 _16542_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09801_));
 sg13g2_nand2_1 _16543_ (.Y(_09802_),
    .A(net1122),
    .B(net626));
 sg13g2_a21oi_1 _16544_ (.A1(_09800_),
    .A2(_09802_),
    .Y(_00023_),
    .B1(net712));
 sg13g2_buf_1 _16545_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09803_));
 sg13g2_buf_1 _16546_ (.A(_09477_),
    .X(_09804_));
 sg13g2_nor2_1 _16547_ (.A(_08284_),
    .B(_08601_),
    .Y(_09805_));
 sg13g2_a21oi_1 _16548_ (.A1(_08284_),
    .A2(_09804_),
    .Y(_09806_),
    .B1(_09805_));
 sg13g2_nor3_1 _16549_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .B(_09803_),
    .C(_09806_),
    .Y(_09807_));
 sg13g2_buf_2 _16550_ (.A(_09807_),
    .X(_09808_));
 sg13g2_inv_1 _16551_ (.Y(_09809_),
    .A(_09803_));
 sg13g2_inv_1 _16552_ (.Y(_09810_),
    .A(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_nor3_1 _16553_ (.A(net1137),
    .B(_09810_),
    .C(_09765_),
    .Y(_09811_));
 sg13g2_and2_1 _16554_ (.A(_09810_),
    .B(_09806_),
    .X(_09812_));
 sg13g2_nor3_1 _16555_ (.A(_09809_),
    .B(_09811_),
    .C(_09812_),
    .Y(_09813_));
 sg13g2_buf_2 _16556_ (.A(_09813_),
    .X(_09814_));
 sg13g2_a22oi_1 _16557_ (.Y(_09815_),
    .B1(_09814_),
    .B2(\cpu.qspi.r_quad[1] ),
    .A2(_09808_),
    .A1(\cpu.qspi.r_quad[2] ));
 sg13g2_inv_1 _16558_ (.Y(_09816_),
    .A(\cpu.qspi.r_quad[0] ));
 sg13g2_or2_1 _16559_ (.X(_09817_),
    .B(_09814_),
    .A(_09808_));
 sg13g2_buf_1 _16560_ (.A(_09817_),
    .X(_09818_));
 sg13g2_or2_1 _16561_ (.X(_09819_),
    .B(_09818_),
    .A(_09816_));
 sg13g2_and2_1 _16562_ (.A(_09815_),
    .B(_09819_),
    .X(_09820_));
 sg13g2_buf_1 _16563_ (.A(_09820_),
    .X(_09821_));
 sg13g2_inv_1 _16564_ (.Y(_09822_),
    .A(\cpu.qspi.r_state[17] ));
 sg13g2_nor3_1 _16565_ (.A(_09822_),
    .B(net916),
    .C(_09776_),
    .Y(_09823_));
 sg13g2_nand2_1 _16566_ (.Y(_09824_),
    .A(_09821_),
    .B(_09823_));
 sg13g2_nand3_1 _16567_ (.B(net802),
    .C(net626),
    .A(_09797_),
    .Y(_09825_));
 sg13g2_nand2_1 _16568_ (.Y(_00028_),
    .A(_09824_),
    .B(_09825_));
 sg13g2_nand2_1 _16569_ (.Y(_09826_),
    .A(_09787_),
    .B(_09791_));
 sg13g2_buf_2 _16570_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09827_));
 sg13g2_nand2_1 _16571_ (.Y(_09828_),
    .A(_09827_),
    .B(_09786_));
 sg13g2_a21oi_1 _16572_ (.A1(_09826_),
    .A2(_09828_),
    .Y(_00027_),
    .B1(net712));
 sg13g2_inv_1 _16573_ (.Y(_09829_),
    .A(_09778_));
 sg13g2_buf_1 _16574_ (.A(net802),
    .X(_09830_));
 sg13g2_o21ai_1 _16575_ (.B1(_09830_),
    .Y(_00021_),
    .A1(_09829_),
    .A2(_09779_));
 sg13g2_buf_2 _16576_ (.A(\cpu.dec.r_op[10] ),
    .X(_09831_));
 sg13g2_nand2_1 _16577_ (.Y(_09832_),
    .A(_09011_),
    .B(_09027_));
 sg13g2_nor4_1 _16578_ (.A(_08854_),
    .B(_08935_),
    .C(_08989_),
    .D(_09832_),
    .Y(_09833_));
 sg13g2_a21o_1 _16579_ (.A2(net108),
    .A1(_09831_),
    .B1(_09833_),
    .X(_00011_));
 sg13g2_buf_2 _16580_ (.A(\cpu.dec.r_op[9] ),
    .X(_09834_));
 sg13g2_inv_1 _16581_ (.Y(_09835_),
    .A(_09834_));
 sg13g2_buf_1 _16582_ (.A(_08856_),
    .X(_09836_));
 sg13g2_buf_1 _16583_ (.A(_08853_),
    .X(_09837_));
 sg13g2_nor2_1 _16584_ (.A(net196),
    .B(net219),
    .Y(_09838_));
 sg13g2_nand3_1 _16585_ (.B(_09058_),
    .C(_09838_),
    .A(net197),
    .Y(_09839_));
 sg13g2_o21ai_1 _16586_ (.B1(_09839_),
    .Y(_09840_),
    .A1(_09046_),
    .A2(_09071_));
 sg13g2_nor2_1 _16587_ (.A(net120),
    .B(_09840_),
    .Y(_09841_));
 sg13g2_a21oi_1 _16588_ (.A1(_09835_),
    .A2(net105),
    .Y(_00020_),
    .B1(_09841_));
 sg13g2_buf_2 _16589_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09842_));
 sg13g2_a21oi_1 _16590_ (.A1(_09827_),
    .A2(net626),
    .Y(_09843_),
    .B1(_09842_));
 sg13g2_nor2_1 _16591_ (.A(net711),
    .B(_09843_),
    .Y(_00024_));
 sg13g2_nand3b_1 _16592_ (.B(_08893_),
    .C(net198),
    .Y(_09844_),
    .A_N(net287));
 sg13g2_a21oi_1 _16593_ (.A1(net219),
    .A2(_09844_),
    .Y(_09845_),
    .B1(net196));
 sg13g2_nand2_1 _16594_ (.Y(_09846_),
    .A(_08990_),
    .B(_09845_));
 sg13g2_buf_1 _16595_ (.A(\cpu.dec.r_op[2] ),
    .X(_09847_));
 sg13g2_buf_1 _16596_ (.A(net1121),
    .X(_09848_));
 sg13g2_nand2_1 _16597_ (.Y(_09849_),
    .A(net1048),
    .B(_09067_));
 sg13g2_o21ai_1 _16598_ (.B1(_09849_),
    .Y(_00013_),
    .A1(_09062_),
    .A2(_09846_));
 sg13g2_buf_2 _16599_ (.A(\cpu.dec.r_op[8] ),
    .X(_09850_));
 sg13g2_nand2_1 _16600_ (.Y(_09851_),
    .A(_09051_),
    .B(_08987_));
 sg13g2_buf_1 _16601_ (.A(_09851_),
    .X(_09852_));
 sg13g2_a21oi_1 _16602_ (.A1(net920),
    .A2(_08922_),
    .Y(_09853_),
    .B1(_08930_));
 sg13g2_buf_2 _16603_ (.A(_09853_),
    .X(_09854_));
 sg13g2_nand2_1 _16604_ (.Y(_09855_),
    .A(net220),
    .B(_09854_));
 sg13g2_buf_1 _16605_ (.A(_09855_),
    .X(_09856_));
 sg13g2_nor3_1 _16606_ (.A(net122),
    .B(net195),
    .C(_09856_),
    .Y(_09857_));
 sg13g2_a21o_1 _16607_ (.A2(_08855_),
    .A1(_09850_),
    .B1(_09857_),
    .X(_00019_));
 sg13g2_buf_1 _16608_ (.A(\cpu.uart.r_div[11] ),
    .X(_09858_));
 sg13g2_nor3_1 _16609_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09859_));
 sg13g2_nor2b_1 _16610_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09859_),
    .Y(_09860_));
 sg13g2_nor2b_1 _16611_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09860_),
    .Y(_09861_));
 sg13g2_nor2b_1 _16612_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09861_),
    .Y(_09862_));
 sg13g2_nor2b_1 _16613_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09862_),
    .Y(_09863_));
 sg13g2_nand2b_1 _16614_ (.Y(_09864_),
    .B(_09863_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16615_ (.A(\cpu.uart.r_div[8] ),
    .B(_09864_),
    .Y(_09865_));
 sg13g2_nand2b_1 _16616_ (.Y(_09866_),
    .B(_09865_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16617_ (.A(_09866_),
    .X(_09867_));
 sg13g2_nor3_1 _16618_ (.A(_09858_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09867_),
    .Y(_09868_));
 sg13g2_buf_2 _16619_ (.A(_09868_),
    .X(_09869_));
 sg13g2_nor2_1 _16620_ (.A(net1053),
    .B(_09869_),
    .Y(_09870_));
 sg13g2_buf_1 _16621_ (.A(_09870_),
    .X(_09871_));
 sg13g2_buf_1 _16622_ (.A(net244),
    .X(_09872_));
 sg13g2_mux2_1 _16623_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00260_),
    .S(net218),
    .X(_00079_));
 sg13g2_xnor2_1 _16624_ (.Y(_09873_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16625_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09873_),
    .S(net218),
    .X(_00082_));
 sg13g2_o21ai_1 _16626_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09874_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16627_ (.A(_09859_),
    .B_N(_09874_),
    .Y(_09875_));
 sg13g2_nor2_1 _16628_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net244),
    .Y(_09876_));
 sg13g2_a21oi_1 _16629_ (.A1(net218),
    .A2(_09875_),
    .Y(_00083_),
    .B1(_09876_));
 sg13g2_xnor2_1 _16630_ (.Y(_09877_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09859_));
 sg13g2_nor2_1 _16631_ (.A(\cpu.uart.r_div_value[3] ),
    .B(net244),
    .Y(_09878_));
 sg13g2_a21oi_1 _16632_ (.A1(_09872_),
    .A2(_09877_),
    .Y(_00084_),
    .B1(_09878_));
 sg13g2_xnor2_1 _16633_ (.Y(_09879_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09860_));
 sg13g2_nor2_1 _16634_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net244),
    .Y(_09880_));
 sg13g2_a21oi_1 _16635_ (.A1(net218),
    .A2(_09879_),
    .Y(_00085_),
    .B1(_09880_));
 sg13g2_xnor2_1 _16636_ (.Y(_09881_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09861_));
 sg13g2_nor2_1 _16637_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net244),
    .Y(_09882_));
 sg13g2_a21oi_1 _16638_ (.A1(net218),
    .A2(_09881_),
    .Y(_00086_),
    .B1(_09882_));
 sg13g2_xnor2_1 _16639_ (.Y(_09883_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09862_));
 sg13g2_nor2_1 _16640_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net244),
    .Y(_09884_));
 sg13g2_a21oi_1 _16641_ (.A1(net218),
    .A2(_09883_),
    .Y(_00087_),
    .B1(_09884_));
 sg13g2_xnor2_1 _16642_ (.Y(_09885_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09863_));
 sg13g2_nor2_1 _16643_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net244),
    .Y(_09886_));
 sg13g2_a21oi_1 _16644_ (.A1(net218),
    .A2(_09885_),
    .Y(_00088_),
    .B1(_09886_));
 sg13g2_xor2_1 _16645_ (.B(_09864_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09887_));
 sg13g2_nor2_1 _16646_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net244),
    .Y(_09888_));
 sg13g2_a21oi_1 _16647_ (.A1(net218),
    .A2(_09887_),
    .Y(_00089_),
    .B1(_09888_));
 sg13g2_xnor2_1 _16648_ (.Y(_09889_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09865_));
 sg13g2_nor2_1 _16649_ (.A(\cpu.uart.r_div_value[9] ),
    .B(_09871_),
    .Y(_09890_));
 sg13g2_a21oi_1 _16650_ (.A1(_09872_),
    .A2(_09889_),
    .Y(_00090_),
    .B1(_09890_));
 sg13g2_buf_1 _16651_ (.A(\cpu.uart.r_div_value[10] ),
    .X(_09891_));
 sg13g2_inv_1 _16652_ (.Y(_09892_),
    .A(_09891_));
 sg13g2_nand2_1 _16653_ (.Y(_09893_),
    .A(net919),
    .B(_09867_));
 sg13g2_o21ai_1 _16654_ (.B1(_09893_),
    .Y(_09894_),
    .A1(_09858_),
    .A2(_09891_));
 sg13g2_inv_1 _16655_ (.Y(_09895_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16656_ (.A(_09895_),
    .B(net798),
    .C(_09867_),
    .Y(_09896_));
 sg13g2_a221oi_1 _16657_ (.B2(_09895_),
    .C1(_09896_),
    .B1(_09894_),
    .A1(_09892_),
    .Y(_00080_),
    .A2(net796));
 sg13g2_nor2_1 _16658_ (.A(\cpu.uart.r_div[10] ),
    .B(_09867_),
    .Y(_09897_));
 sg13g2_nand2_1 _16659_ (.Y(_09898_),
    .A(_09858_),
    .B(net802));
 sg13g2_o21ai_1 _16660_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09899_),
    .A1(net798),
    .A2(_09869_));
 sg13g2_o21ai_1 _16661_ (.B1(_09899_),
    .Y(_00081_),
    .A1(_09897_),
    .A2(_09898_));
 sg13g2_inv_2 _16662_ (.Y(_09900_),
    .A(net1128));
 sg13g2_buf_1 _16663_ (.A(_09900_),
    .X(_09901_));
 sg13g2_buf_1 _16664_ (.A(_09901_),
    .X(_09902_));
 sg13g2_buf_1 _16665_ (.A(net903),
    .X(_09903_));
 sg13g2_buf_1 _16666_ (.A(_09511_),
    .X(_09904_));
 sg13g2_nand2_1 _16667_ (.Y(_09905_),
    .A(_09903_),
    .B(net693));
 sg13g2_buf_2 _16668_ (.A(_09905_),
    .X(_09906_));
 sg13g2_buf_1 _16669_ (.A(\cpu.addr[5] ),
    .X(_09907_));
 sg13g2_nor3_2 _16670_ (.A(net1120),
    .B(_09152_),
    .C(net1057),
    .Y(_09908_));
 sg13g2_nand2_1 _16671_ (.Y(_09909_),
    .A(_09150_),
    .B(_09908_));
 sg13g2_buf_1 _16672_ (.A(_09909_),
    .X(_09910_));
 sg13g2_nor4_1 _16673_ (.A(net780),
    .B(_09168_),
    .C(_09906_),
    .D(net692),
    .Y(_09911_));
 sg13g2_buf_1 _16674_ (.A(_09911_),
    .X(_09912_));
 sg13g2_buf_1 _16675_ (.A(\cpu.intr.r_timer_count[15] ),
    .X(_09913_));
 sg13g2_buf_1 _16676_ (.A(\cpu.intr.r_timer_count[14] ),
    .X(_09914_));
 sg13g2_buf_1 _16677_ (.A(\cpu.intr.r_timer_count[11] ),
    .X(_09915_));
 sg13g2_buf_1 _16678_ (.A(\cpu.intr.r_timer_count[8] ),
    .X(_09916_));
 sg13g2_buf_2 _16679_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09917_));
 sg13g2_nor3_2 _16680_ (.A(_09917_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09918_));
 sg13g2_nor2b_1 _16681_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09918_),
    .Y(_09919_));
 sg13g2_nor2b_1 _16682_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09919_),
    .Y(_09920_));
 sg13g2_nor2b_1 _16683_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09920_),
    .Y(_09921_));
 sg13g2_nor2b_1 _16684_ (.A(\cpu.intr.r_timer_count[6] ),
    .B_N(_09921_),
    .Y(_09922_));
 sg13g2_nand2b_1 _16685_ (.Y(_09923_),
    .B(_09922_),
    .A_N(\cpu.intr.r_timer_count[7] ));
 sg13g2_nor3_2 _16686_ (.A(\cpu.intr.r_timer_count[9] ),
    .B(_09916_),
    .C(_09923_),
    .Y(_09924_));
 sg13g2_nand2b_1 _16687_ (.Y(_09925_),
    .B(_09924_),
    .A_N(\cpu.intr.r_timer_count[10] ));
 sg13g2_nor3_2 _16688_ (.A(_09915_),
    .B(\cpu.intr.r_timer_count[12] ),
    .C(_09925_),
    .Y(_09926_));
 sg13g2_nand2b_1 _16689_ (.Y(_09927_),
    .B(_09926_),
    .A_N(\cpu.intr.r_timer_count[13] ));
 sg13g2_nor3_1 _16690_ (.A(_09913_),
    .B(_09914_),
    .C(_09927_),
    .Y(_09928_));
 sg13g2_buf_1 _16691_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09929_));
 sg13g2_buf_1 _16692_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09930_));
 sg13g2_buf_2 _16693_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09931_));
 sg13g2_buf_1 _16694_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09932_));
 sg13g2_buf_1 _16695_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09933_));
 sg13g2_buf_1 _16696_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09934_));
 sg13g2_buf_1 _16697_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09935_));
 sg13g2_nor4_1 _16698_ (.A(_09932_),
    .B(_09933_),
    .C(_09934_),
    .D(_09935_),
    .Y(_09936_));
 sg13g2_nand2b_1 _16699_ (.Y(_09937_),
    .B(_09936_),
    .A_N(\cpu.intr.r_timer_count[20] ));
 sg13g2_nor4_2 _16700_ (.A(_09929_),
    .B(_09930_),
    .C(_09931_),
    .Y(_09938_),
    .D(_09937_));
 sg13g2_nand2_1 _16701_ (.Y(_09939_),
    .A(_09928_),
    .B(_09938_));
 sg13g2_buf_2 _16702_ (.A(_09939_),
    .X(_09940_));
 sg13g2_nand2b_1 _16703_ (.Y(_09941_),
    .B(_09940_),
    .A_N(_09912_));
 sg13g2_buf_1 _16704_ (.A(_09941_),
    .X(_09942_));
 sg13g2_buf_1 _16705_ (.A(_09942_),
    .X(_09943_));
 sg13g2_mux2_1 _16706_ (.A0(_00266_),
    .A1(\cpu.intr.r_timer_reload[0] ),
    .S(_09943_),
    .X(_00055_));
 sg13g2_buf_1 _16707_ (.A(_09942_),
    .X(_09944_));
 sg13g2_xor2_1 _16708_ (.B(\cpu.intr.r_timer_count[0] ),
    .A(_09917_),
    .X(_09945_));
 sg13g2_nand2_1 _16709_ (.Y(_09946_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net104));
 sg13g2_o21ai_1 _16710_ (.B1(_09946_),
    .Y(_00066_),
    .A1(net103),
    .A2(_09945_));
 sg13g2_o21ai_1 _16711_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_09947_),
    .A1(_09917_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16712_ (.A(_09918_),
    .B_N(_09947_),
    .Y(_09948_));
 sg13g2_nand2_1 _16713_ (.Y(_09949_),
    .A(\cpu.intr.r_timer_reload[2] ),
    .B(net104));
 sg13g2_o21ai_1 _16714_ (.B1(_09949_),
    .Y(_00071_),
    .A1(net103),
    .A2(_09948_));
 sg13g2_xnor2_1 _16715_ (.Y(_09950_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09918_));
 sg13g2_nand2_1 _16716_ (.Y(_09951_),
    .A(\cpu.intr.r_timer_reload[3] ),
    .B(net104));
 sg13g2_o21ai_1 _16717_ (.B1(_09951_),
    .Y(_00072_),
    .A1(net103),
    .A2(_09950_));
 sg13g2_xnor2_1 _16718_ (.Y(_09952_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09919_));
 sg13g2_nand2_1 _16719_ (.Y(_09953_),
    .A(\cpu.intr.r_timer_reload[4] ),
    .B(net104));
 sg13g2_o21ai_1 _16720_ (.B1(_09953_),
    .Y(_00073_),
    .A1(_09944_),
    .A2(_09952_));
 sg13g2_xnor2_1 _16721_ (.Y(_09954_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09920_));
 sg13g2_buf_1 _16722_ (.A(_09942_),
    .X(_09955_));
 sg13g2_nand2_1 _16723_ (.Y(_09956_),
    .A(\cpu.intr.r_timer_reload[5] ),
    .B(_09955_));
 sg13g2_o21ai_1 _16724_ (.B1(_09956_),
    .Y(_00074_),
    .A1(_09944_),
    .A2(_09954_));
 sg13g2_xnor2_1 _16725_ (.Y(_09957_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09921_));
 sg13g2_nand2_1 _16726_ (.Y(_09958_),
    .A(\cpu.intr.r_timer_reload[6] ),
    .B(net102));
 sg13g2_o21ai_1 _16727_ (.B1(_09958_),
    .Y(_00075_),
    .A1(net103),
    .A2(_09957_));
 sg13g2_xnor2_1 _16728_ (.Y(_09959_),
    .A(\cpu.intr.r_timer_count[7] ),
    .B(_09922_));
 sg13g2_nand2_1 _16729_ (.Y(_09960_),
    .A(\cpu.intr.r_timer_reload[7] ),
    .B(net102));
 sg13g2_o21ai_1 _16730_ (.B1(_09960_),
    .Y(_00076_),
    .A1(net103),
    .A2(_09959_));
 sg13g2_xor2_1 _16731_ (.B(_09923_),
    .A(_09916_),
    .X(_09961_));
 sg13g2_nand2_1 _16732_ (.Y(_09962_),
    .A(\cpu.intr.r_timer_reload[8] ),
    .B(net102));
 sg13g2_o21ai_1 _16733_ (.B1(_09962_),
    .Y(_00077_),
    .A1(net103),
    .A2(_09961_));
 sg13g2_o21ai_1 _16734_ (.B1(\cpu.intr.r_timer_count[9] ),
    .Y(_09963_),
    .A1(_09916_),
    .A2(_09923_));
 sg13g2_nor2b_1 _16735_ (.A(_09924_),
    .B_N(_09963_),
    .Y(_09964_));
 sg13g2_nand2_1 _16736_ (.Y(_09965_),
    .A(\cpu.intr.r_timer_reload[9] ),
    .B(net102));
 sg13g2_o21ai_1 _16737_ (.B1(_09965_),
    .Y(_00078_),
    .A1(net103),
    .A2(_09964_));
 sg13g2_xnor2_1 _16738_ (.Y(_09966_),
    .A(\cpu.intr.r_timer_count[10] ),
    .B(_09924_));
 sg13g2_nand2_1 _16739_ (.Y(_09967_),
    .A(\cpu.intr.r_timer_reload[10] ),
    .B(net102));
 sg13g2_o21ai_1 _16740_ (.B1(_09967_),
    .Y(_00056_),
    .A1(net103),
    .A2(_09966_));
 sg13g2_xor2_1 _16741_ (.B(_09925_),
    .A(_09915_),
    .X(_09968_));
 sg13g2_nand2_1 _16742_ (.Y(_09969_),
    .A(\cpu.intr.r_timer_reload[11] ),
    .B(net102));
 sg13g2_o21ai_1 _16743_ (.B1(_09969_),
    .Y(_00057_),
    .A1(net104),
    .A2(_09968_));
 sg13g2_o21ai_1 _16744_ (.B1(\cpu.intr.r_timer_count[12] ),
    .Y(_09970_),
    .A1(_09915_),
    .A2(_09925_));
 sg13g2_nor2b_1 _16745_ (.A(_09926_),
    .B_N(_09970_),
    .Y(_09971_));
 sg13g2_nand2_1 _16746_ (.Y(_09972_),
    .A(\cpu.intr.r_timer_reload[12] ),
    .B(net102));
 sg13g2_o21ai_1 _16747_ (.B1(_09972_),
    .Y(_00058_),
    .A1(net104),
    .A2(_09971_));
 sg13g2_xnor2_1 _16748_ (.Y(_09973_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_09926_));
 sg13g2_nand2_1 _16749_ (.Y(_09974_),
    .A(\cpu.intr.r_timer_reload[13] ),
    .B(net102));
 sg13g2_o21ai_1 _16750_ (.B1(_09974_),
    .Y(_00059_),
    .A1(net104),
    .A2(_09973_));
 sg13g2_xor2_1 _16751_ (.B(_09927_),
    .A(_09914_),
    .X(_09975_));
 sg13g2_nand2_1 _16752_ (.Y(_09976_),
    .A(\cpu.intr.r_timer_reload[14] ),
    .B(_09955_));
 sg13g2_o21ai_1 _16753_ (.B1(_09976_),
    .Y(_00060_),
    .A1(net104),
    .A2(_09975_));
 sg13g2_nor2_1 _16754_ (.A(_09914_),
    .B(_09927_),
    .Y(_09977_));
 sg13g2_xnor2_1 _16755_ (.Y(_09978_),
    .A(_09913_),
    .B(_09977_));
 sg13g2_nand2_1 _16756_ (.Y(_09979_),
    .A(\cpu.intr.r_timer_reload[15] ),
    .B(_09942_));
 sg13g2_o21ai_1 _16757_ (.B1(_09979_),
    .Y(_00061_),
    .A1(_09943_),
    .A2(_09978_));
 sg13g2_buf_1 _16758_ (.A(_09912_),
    .X(_09980_));
 sg13g2_nand2b_1 _16759_ (.Y(_09981_),
    .B(_09977_),
    .A_N(_09913_));
 sg13g2_buf_1 _16760_ (.A(_09981_),
    .X(_09982_));
 sg13g2_inv_1 _16761_ (.Y(_09983_),
    .A(\cpu.intr.r_timer_reload[16] ));
 sg13g2_a21oi_1 _16762_ (.A1(_09983_),
    .A2(_09938_),
    .Y(_09984_),
    .B1(_09933_));
 sg13g2_and2_1 _16763_ (.A(_09928_),
    .B(_09984_),
    .X(_09985_));
 sg13g2_a21oi_1 _16764_ (.A1(_09933_),
    .A2(_09982_),
    .Y(_09986_),
    .B1(_09985_));
 sg13g2_buf_1 _16765_ (.A(\cpu.dcache.wdata[0] ),
    .X(_09987_));
 sg13g2_buf_1 _16766_ (.A(_09987_),
    .X(_09988_));
 sg13g2_buf_1 _16767_ (.A(_09912_),
    .X(_09989_));
 sg13g2_nand2_1 _16768_ (.Y(_09990_),
    .A(net1047),
    .B(net143));
 sg13g2_o21ai_1 _16769_ (.B1(_09990_),
    .Y(_00062_),
    .A1(net144),
    .A2(_09986_));
 sg13g2_inv_1 _16770_ (.Y(_09991_),
    .A(\cpu.intr.r_timer_reload[17] ));
 sg13g2_a21oi_1 _16771_ (.A1(_09991_),
    .A2(_09938_),
    .Y(_09992_),
    .B1(_09932_));
 sg13g2_nor2_1 _16772_ (.A(_09933_),
    .B(_09982_),
    .Y(_09993_));
 sg13g2_mux2_1 _16773_ (.A0(_09932_),
    .A1(_09992_),
    .S(_09993_),
    .X(_09994_));
 sg13g2_buf_1 _16774_ (.A(\cpu.dcache.wdata[1] ),
    .X(_09995_));
 sg13g2_buf_1 _16775_ (.A(_09995_),
    .X(_09996_));
 sg13g2_buf_1 _16776_ (.A(net1046),
    .X(_09997_));
 sg13g2_mux2_1 _16777_ (.A0(_09994_),
    .A1(net900),
    .S(_09989_),
    .X(_00063_));
 sg13g2_or3_1 _16778_ (.A(_09932_),
    .B(_09933_),
    .C(_09982_),
    .X(_09998_));
 sg13g2_xnor2_1 _16779_ (.Y(_09999_),
    .A(_09935_),
    .B(_09998_));
 sg13g2_o21ai_1 _16780_ (.B1(_09999_),
    .Y(_10000_),
    .A1(\cpu.intr.r_timer_reload[18] ),
    .A2(_09940_));
 sg13g2_buf_1 _16781_ (.A(\cpu.dcache.wdata[2] ),
    .X(_10001_));
 sg13g2_buf_1 _16782_ (.A(_10001_),
    .X(_10002_));
 sg13g2_nand2_1 _16783_ (.Y(_10003_),
    .A(net1045),
    .B(net143));
 sg13g2_o21ai_1 _16784_ (.B1(_10003_),
    .Y(_00064_),
    .A1(net144),
    .A2(_10000_));
 sg13g2_or2_1 _16785_ (.X(_10004_),
    .B(_09998_),
    .A(_09935_));
 sg13g2_xnor2_1 _16786_ (.Y(_10005_),
    .A(_09934_),
    .B(_10004_));
 sg13g2_o21ai_1 _16787_ (.B1(_10005_),
    .Y(_10006_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09940_));
 sg13g2_buf_1 _16788_ (.A(\cpu.dcache.wdata[3] ),
    .X(_10007_));
 sg13g2_buf_1 _16789_ (.A(_10007_),
    .X(_10008_));
 sg13g2_nand2_1 _16790_ (.Y(_10009_),
    .A(net1044),
    .B(_09989_));
 sg13g2_o21ai_1 _16791_ (.B1(_10009_),
    .Y(_00065_),
    .A1(_09980_),
    .A2(_10006_));
 sg13g2_nor2_1 _16792_ (.A(_09934_),
    .B(_10004_),
    .Y(_10010_));
 sg13g2_xor2_1 _16793_ (.B(_10010_),
    .A(\cpu.intr.r_timer_count[20] ),
    .X(_10011_));
 sg13g2_o21ai_1 _16794_ (.B1(_10011_),
    .Y(_10012_),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .A2(_09940_));
 sg13g2_buf_2 _16795_ (.A(\cpu.dcache.wdata[4] ),
    .X(_10013_));
 sg13g2_buf_1 _16796_ (.A(_10013_),
    .X(_10014_));
 sg13g2_nand2_1 _16797_ (.Y(_10015_),
    .A(net1043),
    .B(_09912_));
 sg13g2_o21ai_1 _16798_ (.B1(_10015_),
    .Y(_00067_),
    .A1(net143),
    .A2(_10012_));
 sg13g2_or2_1 _16799_ (.X(_10016_),
    .B(_09937_),
    .A(_09982_));
 sg13g2_xnor2_1 _16800_ (.Y(_10017_),
    .A(_09929_),
    .B(_10016_));
 sg13g2_o21ai_1 _16801_ (.B1(_10017_),
    .Y(_10018_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09940_));
 sg13g2_buf_2 _16802_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10019_));
 sg13g2_buf_1 _16803_ (.A(_10019_),
    .X(_10020_));
 sg13g2_nand2_1 _16804_ (.Y(_10021_),
    .A(net1042),
    .B(_09912_));
 sg13g2_o21ai_1 _16805_ (.B1(_10021_),
    .Y(_00068_),
    .A1(net143),
    .A2(_10018_));
 sg13g2_or2_1 _16806_ (.X(_10022_),
    .B(_10016_),
    .A(_09929_));
 sg13g2_buf_1 _16807_ (.A(_10022_),
    .X(_10023_));
 sg13g2_nor2_1 _16808_ (.A(_09930_),
    .B(\cpu.intr.r_timer_reload[22] ),
    .Y(_10024_));
 sg13g2_nor3_1 _16809_ (.A(_09931_),
    .B(_10023_),
    .C(_10024_),
    .Y(_10025_));
 sg13g2_a21oi_1 _16810_ (.A1(_09931_),
    .A2(_10023_),
    .Y(_10026_),
    .B1(_10025_));
 sg13g2_buf_1 _16811_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10027_));
 sg13g2_nand2_1 _16812_ (.Y(_10028_),
    .A(net1119),
    .B(_09912_));
 sg13g2_o21ai_1 _16813_ (.B1(_10028_),
    .Y(_00069_),
    .A1(net143),
    .A2(_10026_));
 sg13g2_nor2_1 _16814_ (.A(_09931_),
    .B(_10023_),
    .Y(_10029_));
 sg13g2_nand2_1 _16815_ (.Y(_10030_),
    .A(\cpu.intr.r_timer_reload[23] ),
    .B(_10029_));
 sg13g2_o21ai_1 _16816_ (.B1(_09930_),
    .Y(_10031_),
    .A1(_09931_),
    .A2(_10023_));
 sg13g2_o21ai_1 _16817_ (.B1(_10031_),
    .Y(_10032_),
    .A1(_09930_),
    .A2(_10030_));
 sg13g2_buf_1 _16818_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10033_));
 sg13g2_buf_1 _16819_ (.A(net1118),
    .X(_10034_));
 sg13g2_mux2_1 _16820_ (.A0(_10032_),
    .A1(net1041),
    .S(net143),
    .X(_00070_));
 sg13g2_buf_1 _16821_ (.A(net628),
    .X(_10035_));
 sg13g2_buf_1 _16822_ (.A(_10035_),
    .X(_10036_));
 sg13g2_nor2_1 _16823_ (.A(_09168_),
    .B(net692),
    .Y(_10037_));
 sg13g2_buf_1 _16824_ (.A(_10037_),
    .X(_10038_));
 sg13g2_nand2_1 _16825_ (.Y(_10039_),
    .A(net503),
    .B(_10038_));
 sg13g2_buf_1 _16826_ (.A(_10039_),
    .X(_10040_));
 sg13g2_nand2_1 _16827_ (.Y(_10041_),
    .A(net789),
    .B(_09333_));
 sg13g2_buf_2 _16828_ (.A(_10041_),
    .X(_10042_));
 sg13g2_nor2_1 _16829_ (.A(net1052),
    .B(_10042_),
    .Y(_10043_));
 sg13g2_buf_1 _16830_ (.A(_10043_),
    .X(_10044_));
 sg13g2_buf_1 _16831_ (.A(net502),
    .X(_10045_));
 sg13g2_and2_1 _16832_ (.A(_10038_),
    .B(net447),
    .X(_10046_));
 sg13g2_buf_1 _16833_ (.A(_10046_),
    .X(_10047_));
 sg13g2_buf_1 _16834_ (.A(_10047_),
    .X(_10048_));
 sg13g2_buf_1 _16835_ (.A(net1047),
    .X(_10049_));
 sg13g2_a22oi_1 _16836_ (.Y(_10050_),
    .B1(net101),
    .B2(net899),
    .A2(net119),
    .A1(_00267_));
 sg13g2_inv_1 _16837_ (.Y(_00036_),
    .A(_10050_));
 sg13g2_buf_1 _16838_ (.A(_09995_),
    .X(_10051_));
 sg13g2_buf_1 _16839_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10052_));
 sg13g2_buf_2 _16840_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10053_));
 sg13g2_xor2_1 _16841_ (.B(_10053_),
    .A(_10052_),
    .X(_10054_));
 sg13g2_buf_1 _16842_ (.A(net119),
    .X(_10055_));
 sg13g2_a22oi_1 _16843_ (.Y(_10056_),
    .B1(_10054_),
    .B2(net100),
    .A2(net101),
    .A1(net1040));
 sg13g2_inv_1 _16844_ (.Y(_00043_),
    .A(_10056_));
 sg13g2_buf_1 _16845_ (.A(net1045),
    .X(_10057_));
 sg13g2_buf_2 _16846_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10058_));
 sg13g2_nand2_1 _16847_ (.Y(_10059_),
    .A(_10052_),
    .B(_10053_));
 sg13g2_xnor2_1 _16848_ (.Y(_10060_),
    .A(_10058_),
    .B(_10059_));
 sg13g2_a22oi_1 _16849_ (.Y(_10061_),
    .B1(_10060_),
    .B2(net100),
    .A2(net101),
    .A1(net898));
 sg13g2_inv_1 _16850_ (.Y(_00044_),
    .A(_10061_));
 sg13g2_buf_1 _16851_ (.A(_10007_),
    .X(_10062_));
 sg13g2_buf_2 _16852_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10063_));
 sg13g2_nand2_1 _16853_ (.Y(_10064_),
    .A(_10053_),
    .B(_10058_));
 sg13g2_nor2_1 _16854_ (.A(_00267_),
    .B(_10064_),
    .Y(_10065_));
 sg13g2_xor2_1 _16855_ (.B(_10065_),
    .A(_10063_),
    .X(_10066_));
 sg13g2_a22oi_1 _16856_ (.Y(_10067_),
    .B1(_10066_),
    .B2(net100),
    .A2(net101),
    .A1(net1039));
 sg13g2_inv_1 _16857_ (.Y(_00045_),
    .A(_10067_));
 sg13g2_buf_2 _16858_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10068_));
 sg13g2_and4_1 _16859_ (.A(_10052_),
    .B(_10053_),
    .C(_10058_),
    .D(_10063_),
    .X(_10069_));
 sg13g2_buf_1 _16860_ (.A(_10069_),
    .X(_10070_));
 sg13g2_xor2_1 _16861_ (.B(_10070_),
    .A(_10068_),
    .X(_10071_));
 sg13g2_a22oi_1 _16862_ (.Y(_10072_),
    .B1(_10071_),
    .B2(net100),
    .A2(net101),
    .A1(net1043));
 sg13g2_inv_1 _16863_ (.Y(_00046_),
    .A(_10072_));
 sg13g2_buf_2 _16864_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10073_));
 sg13g2_and3_1 _16865_ (.X(_10074_),
    .A(_10063_),
    .B(_10068_),
    .C(_10065_));
 sg13g2_buf_1 _16866_ (.A(_10074_),
    .X(_10075_));
 sg13g2_xor2_1 _16867_ (.B(_10075_),
    .A(_10073_),
    .X(_10076_));
 sg13g2_a22oi_1 _16868_ (.Y(_10077_),
    .B1(_10076_),
    .B2(net100),
    .A2(net101),
    .A1(net1042));
 sg13g2_inv_1 _16869_ (.Y(_00047_),
    .A(_10077_));
 sg13g2_buf_1 _16870_ (.A(_10027_),
    .X(_10078_));
 sg13g2_buf_2 _16871_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10079_));
 sg13g2_nand3_1 _16872_ (.B(_10073_),
    .C(_10070_),
    .A(_10068_),
    .Y(_10080_));
 sg13g2_xnor2_1 _16873_ (.Y(_10081_),
    .A(_10079_),
    .B(_10080_));
 sg13g2_a22oi_1 _16874_ (.Y(_10082_),
    .B1(_10081_),
    .B2(net100),
    .A2(net101),
    .A1(net1038));
 sg13g2_inv_1 _16875_ (.Y(_00048_),
    .A(_10082_));
 sg13g2_buf_1 _16876_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10083_));
 sg13g2_nand3_1 _16877_ (.B(_10079_),
    .C(_10075_),
    .A(_10073_),
    .Y(_10084_));
 sg13g2_xnor2_1 _16878_ (.Y(_10085_),
    .A(_10083_),
    .B(_10084_));
 sg13g2_a22oi_1 _16879_ (.Y(_10086_),
    .B1(_10085_),
    .B2(net100),
    .A2(_10048_),
    .A1(net1041));
 sg13g2_inv_1 _16880_ (.Y(_00049_),
    .A(_10086_));
 sg13g2_buf_2 _16881_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10087_));
 sg13g2_buf_2 _16882_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10088_));
 sg13g2_nand2_1 _16883_ (.Y(_10089_),
    .A(_10068_),
    .B(_10070_));
 sg13g2_nand3_1 _16884_ (.B(_10079_),
    .C(_10083_),
    .A(_10073_),
    .Y(_10090_));
 sg13g2_nor2_1 _16885_ (.A(_10089_),
    .B(_10090_),
    .Y(_10091_));
 sg13g2_xor2_1 _16886_ (.B(_10091_),
    .A(_10088_),
    .X(_10092_));
 sg13g2_a22oi_1 _16887_ (.Y(_10093_),
    .B1(_10092_),
    .B2(_10055_),
    .A2(net101),
    .A1(_10087_));
 sg13g2_inv_1 _16888_ (.Y(_00050_),
    .A(_10093_));
 sg13g2_buf_2 _16889_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10094_));
 sg13g2_buf_1 _16890_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10095_));
 sg13g2_nand2_1 _16891_ (.Y(_10096_),
    .A(_10088_),
    .B(_10091_));
 sg13g2_xnor2_1 _16892_ (.Y(_10097_),
    .A(_10095_),
    .B(_10096_));
 sg13g2_a22oi_1 _16893_ (.Y(_10098_),
    .B1(_10097_),
    .B2(_10055_),
    .A2(_10048_),
    .A1(_10094_));
 sg13g2_inv_1 _16894_ (.Y(_00051_),
    .A(_10098_));
 sg13g2_buf_2 _16895_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10099_));
 sg13g2_buf_1 _16896_ (.A(_10047_),
    .X(_10100_));
 sg13g2_buf_1 _16897_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10101_));
 sg13g2_nand3_1 _16898_ (.B(_10095_),
    .C(_10091_),
    .A(_10088_),
    .Y(_10102_));
 sg13g2_xnor2_1 _16899_ (.Y(_10103_),
    .A(_10101_),
    .B(_10102_));
 sg13g2_a22oi_1 _16900_ (.Y(_10104_),
    .B1(_10103_),
    .B2(net100),
    .A2(net99),
    .A1(_10099_));
 sg13g2_inv_1 _16901_ (.Y(_00037_),
    .A(_10104_));
 sg13g2_buf_2 _16902_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10105_));
 sg13g2_buf_1 _16903_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10106_));
 sg13g2_nand3_1 _16904_ (.B(_10095_),
    .C(_10101_),
    .A(_10088_),
    .Y(_10107_));
 sg13g2_nor2_1 _16905_ (.A(_10090_),
    .B(_10107_),
    .Y(_10108_));
 sg13g2_nand2_1 _16906_ (.Y(_10109_),
    .A(_10075_),
    .B(_10108_));
 sg13g2_xnor2_1 _16907_ (.Y(_10110_),
    .A(_10106_),
    .B(_10109_));
 sg13g2_buf_1 _16908_ (.A(net119),
    .X(_10111_));
 sg13g2_a22oi_1 _16909_ (.Y(_10112_),
    .B1(_10110_),
    .B2(net98),
    .A2(net99),
    .A1(_10105_));
 sg13g2_inv_1 _16910_ (.Y(_00038_),
    .A(_10112_));
 sg13g2_buf_2 _16911_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10113_));
 sg13g2_buf_2 _16912_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10114_));
 sg13g2_and2_1 _16913_ (.A(_10106_),
    .B(_10108_),
    .X(_10115_));
 sg13g2_nor2b_1 _16914_ (.A(_10089_),
    .B_N(_10115_),
    .Y(_10116_));
 sg13g2_xor2_1 _16915_ (.B(_10116_),
    .A(_10114_),
    .X(_10117_));
 sg13g2_a22oi_1 _16916_ (.Y(_10118_),
    .B1(_10117_),
    .B2(net98),
    .A2(net99),
    .A1(_10113_));
 sg13g2_inv_1 _16917_ (.Y(_00039_),
    .A(_10118_));
 sg13g2_buf_2 _16918_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10119_));
 sg13g2_buf_2 _16919_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10120_));
 sg13g2_nand3_1 _16920_ (.B(_10075_),
    .C(_10115_),
    .A(_10114_),
    .Y(_10121_));
 sg13g2_buf_1 _16921_ (.A(_10121_),
    .X(_10122_));
 sg13g2_xnor2_1 _16922_ (.Y(_10123_),
    .A(_10120_),
    .B(_10122_));
 sg13g2_a22oi_1 _16923_ (.Y(_10124_),
    .B1(_10123_),
    .B2(net98),
    .A2(net99),
    .A1(_10119_));
 sg13g2_inv_1 _16924_ (.Y(_00040_),
    .A(_10124_));
 sg13g2_buf_2 _16925_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10125_));
 sg13g2_buf_1 _16926_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10126_));
 sg13g2_nand3_1 _16927_ (.B(_10120_),
    .C(_10116_),
    .A(_10114_),
    .Y(_10127_));
 sg13g2_xnor2_1 _16928_ (.Y(_10128_),
    .A(_10126_),
    .B(_10127_));
 sg13g2_a22oi_1 _16929_ (.Y(_10129_),
    .B1(_10128_),
    .B2(net98),
    .A2(net99),
    .A1(_10125_));
 sg13g2_inv_1 _16930_ (.Y(_00041_),
    .A(_10129_));
 sg13g2_buf_2 _16931_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10130_));
 sg13g2_buf_1 _16932_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10131_));
 sg13g2_nand2_1 _16933_ (.Y(_10132_),
    .A(_10120_),
    .B(_10126_));
 sg13g2_nor2_1 _16934_ (.A(_10122_),
    .B(_10132_),
    .Y(_10133_));
 sg13g2_xor2_1 _16935_ (.B(_10133_),
    .A(_10131_),
    .X(_10134_));
 sg13g2_a22oi_1 _16936_ (.Y(_10135_),
    .B1(_10134_),
    .B2(net98),
    .A2(net99),
    .A1(_10130_));
 sg13g2_inv_1 _16937_ (.Y(_00042_),
    .A(_10135_));
 sg13g2_buf_2 _16938_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10136_));
 sg13g2_inv_1 _16939_ (.Y(_10137_),
    .A(_10136_));
 sg13g2_buf_1 _16940_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10138_));
 sg13g2_inv_1 _16941_ (.Y(_10139_),
    .A(_10138_));
 sg13g2_buf_2 _16942_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10140_));
 sg13g2_nand2_1 _16943_ (.Y(_10141_),
    .A(_10139_),
    .B(_10140_));
 sg13g2_buf_1 _16944_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10142_));
 sg13g2_buf_1 _16945_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10143_));
 sg13g2_buf_8 _16946_ (.A(_10143_),
    .X(_10144_));
 sg13g2_nand2_1 _16947_ (.Y(_10145_),
    .A(net1116),
    .B(net1037));
 sg13g2_nor3_1 _16948_ (.A(_10137_),
    .B(_10141_),
    .C(_10145_),
    .Y(_10146_));
 sg13g2_buf_1 _16949_ (.A(_10146_),
    .X(_10147_));
 sg13g2_buf_1 _16950_ (.A(net691),
    .X(_10148_));
 sg13g2_buf_1 _16951_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10149_));
 sg13g2_inv_1 _16952_ (.Y(_10150_),
    .A(net1115));
 sg13g2_buf_1 _16953_ (.A(_10150_),
    .X(_10151_));
 sg13g2_buf_2 _16954_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10152_));
 sg13g2_xnor2_1 _16955_ (.Y(_10153_),
    .A(net1117),
    .B(_10152_));
 sg13g2_buf_2 _16956_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10154_));
 sg13g2_xnor2_1 _16957_ (.Y(_10155_),
    .A(net1037),
    .B(_10154_));
 sg13g2_nand2_1 _16958_ (.Y(_10156_),
    .A(_10153_),
    .B(_10155_));
 sg13g2_buf_1 _16959_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10157_));
 sg13g2_buf_1 _16960_ (.A(_10157_),
    .X(_10158_));
 sg13g2_xor2_1 _16961_ (.B(net1036),
    .A(_10140_),
    .X(_10159_));
 sg13g2_buf_8 _16962_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10160_));
 sg13g2_xor2_1 _16963_ (.B(net1114),
    .A(net1116),
    .X(_10161_));
 sg13g2_nor2_1 _16964_ (.A(net1116),
    .B(_10143_),
    .Y(_10162_));
 sg13g2_nor2_1 _16965_ (.A(net1117),
    .B(_10140_),
    .Y(_10163_));
 sg13g2_a21o_1 _16966_ (.A2(_10163_),
    .A1(_10162_),
    .B1(_10137_),
    .X(_10164_));
 sg13g2_nor4_2 _16967_ (.A(_10156_),
    .B(_10159_),
    .C(_10161_),
    .Y(_10165_),
    .D(_10164_));
 sg13g2_buf_8 _16968_ (.A(_10165_),
    .X(_10166_));
 sg13g2_inv_1 _16969_ (.Y(_10167_),
    .A(net1114));
 sg13g2_buf_8 _16970_ (.A(_10152_),
    .X(_10168_));
 sg13g2_nor3_1 _16971_ (.A(_10154_),
    .B(net1034),
    .C(net1036),
    .Y(_10169_));
 sg13g2_and2_1 _16972_ (.A(net1035),
    .B(_10169_),
    .X(_10170_));
 sg13g2_or2_1 _16973_ (.X(_10171_),
    .B(_10170_),
    .A(net624));
 sg13g2_buf_2 _16974_ (.A(_10171_),
    .X(_10172_));
 sg13g2_buf_1 _16975_ (.A(net1114),
    .X(_10173_));
 sg13g2_buf_8 _16976_ (.A(net1033),
    .X(_10174_));
 sg13g2_buf_1 _16977_ (.A(_10174_),
    .X(_10175_));
 sg13g2_buf_1 _16978_ (.A(_10175_),
    .X(_10176_));
 sg13g2_buf_8 _16979_ (.A(net1034),
    .X(_10177_));
 sg13g2_buf_8 _16980_ (.A(net895),
    .X(_10178_));
 sg13g2_buf_1 _16981_ (.A(_10178_),
    .X(_10179_));
 sg13g2_nand2_1 _16982_ (.Y(_10180_),
    .A(net690),
    .B(net689));
 sg13g2_buf_8 _16983_ (.A(_10154_),
    .X(_10181_));
 sg13g2_buf_1 _16984_ (.A(_10157_),
    .X(_10182_));
 sg13g2_nor2b_1 _16985_ (.A(net1032),
    .B_N(net1031),
    .Y(_10183_));
 sg13g2_buf_1 _16986_ (.A(_10183_),
    .X(_10184_));
 sg13g2_buf_8 _16987_ (.A(net1036),
    .X(_10185_));
 sg13g2_buf_8 _16988_ (.A(net1032),
    .X(_10186_));
 sg13g2_nor2b_2 _16989_ (.A(net894),
    .B_N(net893),
    .Y(_10187_));
 sg13g2_a22oi_1 _16990_ (.Y(_10188_),
    .B1(_10187_),
    .B2(\cpu.ex.r_11[15] ),
    .A2(_10184_),
    .A1(\cpu.ex.r_14[15] ));
 sg13g2_buf_1 _16991_ (.A(net894),
    .X(_10189_));
 sg13g2_buf_1 _16992_ (.A(_10189_),
    .X(_10190_));
 sg13g2_nand3b_1 _16993_ (.B(net690),
    .C(\cpu.ex.r_epc[15] ),
    .Y(_10191_),
    .A_N(net688));
 sg13g2_buf_1 _16994_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10192_));
 sg13g2_nand3b_1 _16995_ (.B(net688),
    .C(_10192_),
    .Y(_10193_),
    .A_N(_10175_));
 sg13g2_buf_8 _16996_ (.A(net1032),
    .X(_10194_));
 sg13g2_buf_1 _16997_ (.A(net892),
    .X(_10195_));
 sg13g2_buf_1 _16998_ (.A(net775),
    .X(_10196_));
 sg13g2_nand2b_1 _16999_ (.Y(_10197_),
    .B(net687),
    .A_N(net689));
 sg13g2_a21o_1 _17000_ (.A2(_10193_),
    .A1(_10191_),
    .B1(_10197_),
    .X(_10198_));
 sg13g2_o21ai_1 _17001_ (.B1(_10198_),
    .Y(_10199_),
    .A1(_10180_),
    .A2(_10188_));
 sg13g2_buf_1 _17002_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10200_));
 sg13g2_nor2_2 _17003_ (.A(net1034),
    .B(net1036),
    .Y(_10201_));
 sg13g2_buf_8 _17004_ (.A(_10201_),
    .X(_10202_));
 sg13g2_nor2b_1 _17005_ (.A(_10181_),
    .B_N(_10173_),
    .Y(_10203_));
 sg13g2_buf_2 _17006_ (.A(_10203_),
    .X(_10204_));
 sg13g2_nand3_1 _17007_ (.B(_10202_),
    .C(_10204_),
    .A(_10200_),
    .Y(_10205_));
 sg13g2_inv_2 _17008_ (.Y(_10206_),
    .A(net1031));
 sg13g2_buf_1 _17009_ (.A(_10206_),
    .X(_10207_));
 sg13g2_nor2b_1 _17010_ (.A(net1114),
    .B_N(_10152_),
    .Y(_10208_));
 sg13g2_buf_1 _17011_ (.A(_10208_),
    .X(_10209_));
 sg13g2_buf_1 _17012_ (.A(_10209_),
    .X(_10210_));
 sg13g2_mux2_1 _17013_ (.A0(\cpu.ex.r_8[15] ),
    .A1(\cpu.ex.r_9[15] ),
    .S(net687),
    .X(_10211_));
 sg13g2_nand3_1 _17014_ (.B(net772),
    .C(_10211_),
    .A(net773),
    .Y(_10212_));
 sg13g2_buf_1 _17015_ (.A(_10190_),
    .X(_10213_));
 sg13g2_mux2_1 _17016_ (.A0(\cpu.ex.r_12[15] ),
    .A1(\cpu.ex.r_13[15] ),
    .S(_10196_),
    .X(_10214_));
 sg13g2_nand3_1 _17017_ (.B(_10210_),
    .C(_10214_),
    .A(net623),
    .Y(_10215_));
 sg13g2_nand3_1 _17018_ (.B(_10212_),
    .C(_10215_),
    .A(_10205_),
    .Y(_10216_));
 sg13g2_inv_1 _17019_ (.Y(_10217_),
    .A(_10154_));
 sg13g2_buf_1 _17020_ (.A(_10217_),
    .X(_10218_));
 sg13g2_buf_1 _17021_ (.A(net891),
    .X(_10219_));
 sg13g2_buf_1 _17022_ (.A(net771),
    .X(_10220_));
 sg13g2_and2_1 _17023_ (.A(net1033),
    .B(net895),
    .X(_10221_));
 sg13g2_buf_2 _17024_ (.A(_10221_),
    .X(_10222_));
 sg13g2_nand3_1 _17025_ (.B(net686),
    .C(_10222_),
    .A(\cpu.ex.r_10[15] ),
    .Y(_10223_));
 sg13g2_buf_1 _17026_ (.A(net687),
    .X(_10224_));
 sg13g2_nor2_1 _17027_ (.A(net1033),
    .B(_10177_),
    .Y(_10225_));
 sg13g2_buf_1 _17028_ (.A(_10225_),
    .X(_10226_));
 sg13g2_nand3_1 _17029_ (.B(net622),
    .C(_10226_),
    .A(\cpu.ex.r_lr[15] ),
    .Y(_10227_));
 sg13g2_a21oi_1 _17030_ (.A1(_10223_),
    .A2(_10227_),
    .Y(_10228_),
    .B1(net623));
 sg13g2_buf_8 _17031_ (.A(_10177_),
    .X(_10229_));
 sg13g2_nor2_1 _17032_ (.A(net893),
    .B(net770),
    .Y(_10230_));
 sg13g2_nand2_1 _17033_ (.Y(_10231_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(_10230_));
 sg13g2_nor2b_1 _17034_ (.A(_00253_),
    .B_N(_10178_),
    .Y(_10232_));
 sg13g2_nor2b_1 _17035_ (.A(net689),
    .B_N(\cpu.ex.r_mult[31] ),
    .Y(_10233_));
 sg13g2_o21ai_1 _17036_ (.B1(net622),
    .Y(_10234_),
    .A1(_10232_),
    .A2(_10233_));
 sg13g2_nand2_1 _17037_ (.Y(_10235_),
    .A(net690),
    .B(_10213_));
 sg13g2_a21oi_1 _17038_ (.A1(_10231_),
    .A2(_10234_),
    .Y(_10236_),
    .B1(_10235_));
 sg13g2_nor4_1 _17039_ (.A(_10199_),
    .B(_10216_),
    .C(_10228_),
    .D(_10236_),
    .Y(_10237_));
 sg13g2_buf_1 _17040_ (.A(net624),
    .X(_10238_));
 sg13g2_nand2_1 _17041_ (.Y(_10239_),
    .A(net904),
    .B(net570));
 sg13g2_o21ai_1 _17042_ (.B1(_10239_),
    .Y(_10240_),
    .A1(_10172_),
    .A2(_10237_));
 sg13g2_buf_1 _17043_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10241_));
 sg13g2_buf_1 _17044_ (.A(_10241_),
    .X(_10242_));
 sg13g2_buf_1 _17045_ (.A(_10242_),
    .X(_10243_));
 sg13g2_mux2_1 _17046_ (.A0(\cpu.dec.imm[15] ),
    .A1(_10240_),
    .S(net890),
    .X(_10244_));
 sg13g2_nor2_1 _17047_ (.A(_10151_),
    .B(_00176_),
    .Y(_10245_));
 sg13g2_a21o_1 _17048_ (.A2(_10244_),
    .A1(net897),
    .B1(_10245_),
    .X(_10246_));
 sg13g2_buf_1 _17049_ (.A(_10246_),
    .X(_10247_));
 sg13g2_inv_1 _17050_ (.Y(_10248_),
    .A(_00177_));
 sg13g2_nor2_1 _17051_ (.A(_10165_),
    .B(_10170_),
    .Y(_10249_));
 sg13g2_buf_1 _17052_ (.A(_10249_),
    .X(_10250_));
 sg13g2_buf_1 _17053_ (.A(net569),
    .X(_10251_));
 sg13g2_nor2b_1 _17054_ (.A(net1033),
    .B_N(_10154_),
    .Y(_10252_));
 sg13g2_buf_1 _17055_ (.A(_10252_),
    .X(_10253_));
 sg13g2_mux2_1 _17056_ (.A0(\cpu.ex.r_8[14] ),
    .A1(\cpu.ex.r_10[14] ),
    .S(_10176_),
    .X(_10254_));
 sg13g2_a22oi_1 _17057_ (.Y(_10255_),
    .B1(_10254_),
    .B2(_10220_),
    .A2(_10253_),
    .A1(\cpu.ex.r_9[14] ));
 sg13g2_nor2b_1 _17058_ (.A(net896),
    .B_N(net894),
    .Y(_10256_));
 sg13g2_buf_2 _17059_ (.A(_10256_),
    .X(_10257_));
 sg13g2_mux2_1 _17060_ (.A0(\cpu.ex.r_12[14] ),
    .A1(\cpu.ex.r_13[14] ),
    .S(net687),
    .X(_10258_));
 sg13g2_nand2_1 _17061_ (.Y(_10259_),
    .A(_10257_),
    .B(_10258_));
 sg13g2_o21ai_1 _17062_ (.B1(_10259_),
    .Y(_10260_),
    .A1(net623),
    .A2(_10255_));
 sg13g2_nand2_1 _17063_ (.Y(_10261_),
    .A(net689),
    .B(_10260_));
 sg13g2_nor3_1 _17064_ (.A(_00252_),
    .B(net773),
    .C(_10180_),
    .Y(_10262_));
 sg13g2_and3_1 _17065_ (.X(_10263_),
    .A(\cpu.ex.r_lr[14] ),
    .B(net773),
    .C(_10226_));
 sg13g2_o21ai_1 _17066_ (.B1(net622),
    .Y(_10264_),
    .A1(_10262_),
    .A2(_10263_));
 sg13g2_nor2b_1 _17067_ (.A(_10168_),
    .B_N(_10158_),
    .Y(_10265_));
 sg13g2_buf_2 _17068_ (.A(_10265_),
    .X(_10266_));
 sg13g2_nand2_1 _17069_ (.Y(_10267_),
    .A(\cpu.ex.r_stmp[14] ),
    .B(_10266_));
 sg13g2_nor2b_1 _17070_ (.A(net1031),
    .B_N(net1034),
    .Y(_10268_));
 sg13g2_buf_2 _17071_ (.A(_10268_),
    .X(_10269_));
 sg13g2_nand3_1 _17072_ (.B(net622),
    .C(_10269_),
    .A(\cpu.ex.r_11[14] ),
    .Y(_10270_));
 sg13g2_o21ai_1 _17073_ (.B1(_10270_),
    .Y(_10271_),
    .A1(_10224_),
    .A2(_10267_));
 sg13g2_inv_1 _17074_ (.Y(_10272_),
    .A(\cpu.ex.r_14[14] ));
 sg13g2_nand3b_1 _17075_ (.B(net1033),
    .C(net1034),
    .Y(_10273_),
    .A_N(net1032));
 sg13g2_buf_1 _17076_ (.A(_10273_),
    .X(_10274_));
 sg13g2_buf_1 _17077_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_10275_));
 sg13g2_nand3_1 _17078_ (.B(net622),
    .C(net685),
    .A(_10275_),
    .Y(_10276_));
 sg13g2_o21ai_1 _17079_ (.B1(_10276_),
    .Y(_10277_),
    .A1(_10272_),
    .A2(_10274_));
 sg13g2_buf_1 _17080_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10278_));
 sg13g2_nand3_1 _17081_ (.B(net774),
    .C(_10204_),
    .A(_10278_),
    .Y(_10279_));
 sg13g2_nor2b_1 _17082_ (.A(_10152_),
    .B_N(\cpu.dec.r_rs2[1] ),
    .Y(_10280_));
 sg13g2_buf_1 _17083_ (.A(_10280_),
    .X(_10281_));
 sg13g2_mux2_1 _17084_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(\cpu.ex.r_mult[30] ),
    .S(net623),
    .X(_10282_));
 sg13g2_nand3_1 _17085_ (.B(net889),
    .C(_10282_),
    .A(net622),
    .Y(_10283_));
 sg13g2_nand2_1 _17086_ (.Y(_10284_),
    .A(_10279_),
    .B(_10283_));
 sg13g2_a221oi_1 _17087_ (.B2(net623),
    .C1(_10284_),
    .B1(_10277_),
    .A1(_10176_),
    .Y(_10285_),
    .A2(_10271_));
 sg13g2_nand3_1 _17088_ (.B(_10264_),
    .C(_10285_),
    .A(_10261_),
    .Y(_10286_));
 sg13g2_a22oi_1 _17089_ (.Y(_10287_),
    .B1(net501),
    .B2(_10286_),
    .A2(net570),
    .A1(net783));
 sg13g2_nor2_1 _17090_ (.A(net890),
    .B(\cpu.dec.imm[14] ),
    .Y(_10288_));
 sg13g2_a21oi_1 _17091_ (.A1(net890),
    .A2(_10287_),
    .Y(_10289_),
    .B1(_10288_));
 sg13g2_mux2_1 _17092_ (.A0(_10248_),
    .A1(_10289_),
    .S(net897),
    .X(_10290_));
 sg13g2_buf_2 _17093_ (.A(_10290_),
    .X(_10291_));
 sg13g2_buf_2 _17094_ (.A(_10291_),
    .X(_10292_));
 sg13g2_buf_1 _17095_ (.A(_00275_),
    .X(_10293_));
 sg13g2_nor2_1 _17096_ (.A(_10150_),
    .B(_10293_),
    .Y(_10294_));
 sg13g2_buf_1 _17097_ (.A(net1115),
    .X(_10295_));
 sg13g2_nor2_1 _17098_ (.A(net1030),
    .B(\cpu.dec.imm[9] ),
    .Y(_10296_));
 sg13g2_buf_2 _17099_ (.A(\cpu.addr[9] ),
    .X(_10297_));
 sg13g2_nand2_1 _17100_ (.Y(_10298_),
    .A(_10154_),
    .B(_10160_));
 sg13g2_buf_1 _17101_ (.A(_10298_),
    .X(_10299_));
 sg13g2_nor2_1 _17102_ (.A(_00247_),
    .B(net888),
    .Y(_10300_));
 sg13g2_buf_8 _17103_ (.A(net896),
    .X(_10301_));
 sg13g2_nand2_1 _17104_ (.Y(_10302_),
    .A(\cpu.ex.r_14[9] ),
    .B(net769));
 sg13g2_nand2b_1 _17105_ (.Y(_10303_),
    .B(\cpu.ex.r_12[9] ),
    .A_N(net896));
 sg13g2_a21oi_1 _17106_ (.A1(_10302_),
    .A2(_10303_),
    .Y(_10304_),
    .B1(net775));
 sg13g2_and2_1 _17107_ (.A(_10168_),
    .B(net1036),
    .X(_10305_));
 sg13g2_buf_1 _17108_ (.A(_10305_),
    .X(_10306_));
 sg13g2_o21ai_1 _17109_ (.B1(net768),
    .Y(_10307_),
    .A1(_10300_),
    .A2(_10304_));
 sg13g2_nand2b_1 _17110_ (.Y(_10308_),
    .B(net1114),
    .A_N(_10154_));
 sg13g2_nor2_1 _17111_ (.A(net895),
    .B(_10308_),
    .Y(_10309_));
 sg13g2_buf_1 _17112_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10310_));
 sg13g2_mux2_1 _17113_ (.A0(_10310_),
    .A1(\cpu.ex.r_stmp[9] ),
    .S(net776),
    .X(_10311_));
 sg13g2_nand2b_1 _17114_ (.Y(_10312_),
    .B(_10152_),
    .A_N(_10154_));
 sg13g2_buf_1 _17115_ (.A(_10312_),
    .X(_10313_));
 sg13g2_nor2_1 _17116_ (.A(net1031),
    .B(_10313_),
    .Y(_10314_));
 sg13g2_mux2_1 _17117_ (.A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_10[9] ),
    .S(net769),
    .X(_10315_));
 sg13g2_a22oi_1 _17118_ (.Y(_10316_),
    .B1(_10314_),
    .B2(_10315_),
    .A2(_10311_),
    .A1(_10309_));
 sg13g2_a22oi_1 _17119_ (.Y(_10317_),
    .B1(net685),
    .B2(\cpu.ex.r_lr[9] ),
    .A2(_10222_),
    .A1(\cpu.ex.r_11[9] ));
 sg13g2_nand2b_1 _17120_ (.Y(_10318_),
    .B(_10187_),
    .A_N(_10317_));
 sg13g2_mux2_1 _17121_ (.A0(\cpu.ex.r_9[9] ),
    .A1(\cpu.ex.r_13[9] ),
    .S(_10185_),
    .X(_10319_));
 sg13g2_mux2_1 _17122_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(\cpu.ex.r_mult[25] ),
    .S(net894),
    .X(_10320_));
 sg13g2_a22oi_1 _17123_ (.Y(_10321_),
    .B1(_10320_),
    .B2(net889),
    .A2(_10319_),
    .A1(_10209_));
 sg13g2_nand2b_1 _17124_ (.Y(_10322_),
    .B(net775),
    .A_N(_10321_));
 sg13g2_nand4_1 _17125_ (.B(_10316_),
    .C(_10318_),
    .A(_10307_),
    .Y(_10323_),
    .D(_10322_));
 sg13g2_inv_1 _17126_ (.Y(_10324_),
    .A(_10241_));
 sg13g2_a221oi_1 _17127_ (.B2(_10323_),
    .C1(net1028),
    .B1(net569),
    .A1(_10297_),
    .Y(_10325_),
    .A2(net624));
 sg13g2_nor3_2 _17128_ (.A(net1029),
    .B(_10296_),
    .C(_10325_),
    .Y(_10326_));
 sg13g2_nor2_1 _17129_ (.A(_10294_),
    .B(_10326_),
    .Y(_10327_));
 sg13g2_buf_1 _17130_ (.A(_10327_),
    .X(_10328_));
 sg13g2_buf_1 _17131_ (.A(_10328_),
    .X(_10329_));
 sg13g2_buf_2 _17132_ (.A(_00277_),
    .X(_10330_));
 sg13g2_nand2b_1 _17133_ (.Y(_10331_),
    .B(net1115),
    .A_N(_10330_));
 sg13g2_buf_1 _17134_ (.A(_10331_),
    .X(_10332_));
 sg13g2_nor2_1 _17135_ (.A(net1030),
    .B(\cpu.dec.imm[6] ),
    .Y(_10333_));
 sg13g2_inv_1 _17136_ (.Y(_10334_),
    .A(_00244_));
 sg13g2_a22oi_1 _17137_ (.Y(_10335_),
    .B1(net768),
    .B2(_10334_),
    .A2(_10201_),
    .A1(\cpu.ex.r_epc[6] ));
 sg13g2_or2_1 _17138_ (.X(_10336_),
    .B(_10335_),
    .A(net888));
 sg13g2_nor2_2 _17139_ (.A(net1114),
    .B(net1036),
    .Y(_10337_));
 sg13g2_and2_1 _17140_ (.A(_10160_),
    .B(_10158_),
    .X(_10338_));
 sg13g2_buf_2 _17141_ (.A(_10338_),
    .X(_10339_));
 sg13g2_a22oi_1 _17142_ (.Y(_10340_),
    .B1(_10339_),
    .B2(\cpu.ex.r_mult[22] ),
    .A2(_10337_),
    .A1(\cpu.ex.r_lr[6] ));
 sg13g2_nor2b_1 _17143_ (.A(net895),
    .B_N(net1032),
    .Y(_10341_));
 sg13g2_buf_1 _17144_ (.A(_10341_),
    .X(_10342_));
 sg13g2_nand2b_1 _17145_ (.Y(_10343_),
    .B(_10342_),
    .A_N(_10340_));
 sg13g2_mux2_1 _17146_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_10[6] ),
    .S(net1033),
    .X(_10344_));
 sg13g2_mux2_1 _17147_ (.A0(\cpu.ex.r_12[6] ),
    .A1(\cpu.ex.r_13[6] ),
    .S(_10181_),
    .X(_10345_));
 sg13g2_nand2b_1 _17148_ (.Y(_10346_),
    .B(net1034),
    .A_N(net1114));
 sg13g2_buf_1 _17149_ (.A(_10346_),
    .X(_10347_));
 sg13g2_nor2_1 _17150_ (.A(_10206_),
    .B(_10347_),
    .Y(_10348_));
 sg13g2_nand2_1 _17151_ (.Y(_10349_),
    .A(\cpu.ex.r_11[6] ),
    .B(net1033));
 sg13g2_nand2b_1 _17152_ (.Y(_10350_),
    .B(\cpu.ex.r_9[6] ),
    .A_N(_10173_));
 sg13g2_nand3b_1 _17153_ (.B(net1034),
    .C(net1032),
    .Y(_10351_),
    .A_N(_10182_));
 sg13g2_a21oi_1 _17154_ (.A1(_10349_),
    .A2(_10350_),
    .Y(_10352_),
    .B1(_10351_));
 sg13g2_a221oi_1 _17155_ (.B2(_10348_),
    .C1(_10352_),
    .B1(_10345_),
    .A1(_10314_),
    .Y(_10353_),
    .A2(_10344_));
 sg13g2_buf_1 _17156_ (.A(\cpu.ex.r_sp[6] ),
    .X(_10354_));
 sg13g2_mux2_1 _17157_ (.A0(_10354_),
    .A1(\cpu.ex.r_stmp[6] ),
    .S(_10182_),
    .X(_10355_));
 sg13g2_inv_2 _17158_ (.Y(_10356_),
    .A(net895));
 sg13g2_a22oi_1 _17159_ (.Y(_10357_),
    .B1(_10355_),
    .B2(_10356_),
    .A2(_10306_),
    .A1(\cpu.ex.r_14[6] ));
 sg13g2_nand2b_1 _17160_ (.Y(_10358_),
    .B(_10204_),
    .A_N(_10357_));
 sg13g2_nand4_1 _17161_ (.B(_10343_),
    .C(_10353_),
    .A(_10336_),
    .Y(_10359_),
    .D(_10358_));
 sg13g2_a221oi_1 _17162_ (.B2(_10359_),
    .C1(net1028),
    .B1(net569),
    .A1(_09150_),
    .Y(_10360_),
    .A2(net624));
 sg13g2_or3_1 _17163_ (.A(net1115),
    .B(_10333_),
    .C(_10360_),
    .X(_10361_));
 sg13g2_buf_2 _17164_ (.A(_10361_),
    .X(_10362_));
 sg13g2_and2_1 _17165_ (.A(_10332_),
    .B(_10362_),
    .X(_10363_));
 sg13g2_buf_1 _17166_ (.A(_10363_),
    .X(_10364_));
 sg13g2_buf_1 _17167_ (.A(_00274_),
    .X(_10365_));
 sg13g2_nor2_1 _17168_ (.A(net897),
    .B(_10365_),
    .Y(_10366_));
 sg13g2_nor2_1 _17169_ (.A(net1030),
    .B(\cpu.dec.imm[10] ),
    .Y(_10367_));
 sg13g2_buf_2 _17170_ (.A(\cpu.addr[10] ),
    .X(_10368_));
 sg13g2_nor2b_1 _17171_ (.A(_00248_),
    .B_N(net893),
    .Y(_10369_));
 sg13g2_mux2_1 _17172_ (.A0(\cpu.ex.r_8[10] ),
    .A1(\cpu.ex.r_9[10] ),
    .S(_10186_),
    .X(_10370_));
 sg13g2_a22oi_1 _17173_ (.Y(_10371_),
    .B1(_10370_),
    .B2(_10337_),
    .A2(_10369_),
    .A1(_10339_));
 sg13g2_mux2_1 _17174_ (.A0(\cpu.ex.r_12[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(_10174_),
    .X(_10372_));
 sg13g2_nand2_1 _17175_ (.Y(_10373_),
    .A(_10184_),
    .B(_10372_));
 sg13g2_a21oi_1 _17176_ (.A1(_10371_),
    .A2(_10373_),
    .Y(_10374_),
    .B1(_10356_));
 sg13g2_or2_1 _17177_ (.X(_10375_),
    .B(net894),
    .A(_10229_));
 sg13g2_buf_1 _17178_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10376_));
 sg13g2_a22oi_1 _17179_ (.Y(_10377_),
    .B1(_10253_),
    .B2(\cpu.ex.r_lr[10] ),
    .A2(_10204_),
    .A1(_10376_));
 sg13g2_nor2_1 _17180_ (.A(_10375_),
    .B(_10377_),
    .Y(_10378_));
 sg13g2_nand3_1 _17181_ (.B(net776),
    .C(_10209_),
    .A(\cpu.ex.r_13[10] ),
    .Y(_10379_));
 sg13g2_nand3_1 _17182_ (.B(_10301_),
    .C(_10202_),
    .A(\cpu.ex.r_epc[10] ),
    .Y(_10380_));
 sg13g2_a21oi_1 _17183_ (.A1(_10379_),
    .A2(_10380_),
    .Y(_10381_),
    .B1(net771));
 sg13g2_a221oi_1 _17184_ (.B2(\cpu.ex.r_10[10] ),
    .C1(net892),
    .B1(_10269_),
    .A1(\cpu.ex.r_stmp[10] ),
    .Y(_10382_),
    .A2(_10266_));
 sg13g2_a221oi_1 _17185_ (.B2(\cpu.ex.r_11[10] ),
    .C1(net891),
    .B1(_10269_),
    .A1(\cpu.ex.r_mult[26] ),
    .Y(_10383_),
    .A2(_10266_));
 sg13g2_nor3_1 _17186_ (.A(_10167_),
    .B(_10382_),
    .C(_10383_),
    .Y(_10384_));
 sg13g2_or4_1 _17187_ (.A(_10374_),
    .B(_10378_),
    .C(_10381_),
    .D(_10384_),
    .X(_10385_));
 sg13g2_a221oi_1 _17188_ (.B2(_10385_),
    .C1(net1028),
    .B1(net569),
    .A1(_10368_),
    .Y(_10386_),
    .A2(_10166_));
 sg13g2_nor3_1 _17189_ (.A(net1029),
    .B(_10367_),
    .C(_10386_),
    .Y(_10387_));
 sg13g2_nor2_1 _17190_ (.A(_10366_),
    .B(_10387_),
    .Y(_10388_));
 sg13g2_buf_2 _17191_ (.A(_10388_),
    .X(_10389_));
 sg13g2_buf_1 _17192_ (.A(_10389_),
    .X(_10390_));
 sg13g2_nand3_1 _17193_ (.B(net286),
    .C(net285),
    .A(net243),
    .Y(_10391_));
 sg13g2_buf_1 _17194_ (.A(_00178_),
    .X(_10392_));
 sg13g2_mux2_1 _17195_ (.A0(\cpu.ex.r_8[13] ),
    .A1(\cpu.ex.r_12[13] ),
    .S(net688),
    .X(_10393_));
 sg13g2_buf_1 _17196_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10394_));
 sg13g2_mux2_1 _17197_ (.A0(_10394_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net688),
    .X(_10395_));
 sg13g2_a22oi_1 _17198_ (.Y(_10396_),
    .B1(_10395_),
    .B2(net889),
    .A2(_10393_),
    .A1(_10210_));
 sg13g2_inv_1 _17199_ (.Y(_10397_),
    .A(_10396_));
 sg13g2_nand3_1 _17200_ (.B(net686),
    .C(_10222_),
    .A(\cpu.ex.r_10[13] ),
    .Y(_10398_));
 sg13g2_nand3_1 _17201_ (.B(net622),
    .C(net685),
    .A(\cpu.ex.r_lr[13] ),
    .Y(_10399_));
 sg13g2_nand3_1 _17202_ (.B(_10398_),
    .C(_10399_),
    .A(net773),
    .Y(_10400_));
 sg13g2_buf_1 _17203_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10401_));
 sg13g2_nand3_1 _17204_ (.B(net622),
    .C(net685),
    .A(_10401_),
    .Y(_10402_));
 sg13g2_nand3_1 _17205_ (.B(net686),
    .C(_10222_),
    .A(\cpu.ex.r_14[13] ),
    .Y(_10403_));
 sg13g2_nand3_1 _17206_ (.B(_10402_),
    .C(_10403_),
    .A(net623),
    .Y(_10404_));
 sg13g2_nand2b_1 _17207_ (.Y(_10405_),
    .B(net689),
    .A_N(_00251_));
 sg13g2_nand2b_1 _17208_ (.Y(_10406_),
    .B(\cpu.ex.r_mult[29] ),
    .A_N(_10179_));
 sg13g2_nand3_1 _17209_ (.B(net690),
    .C(net688),
    .A(net687),
    .Y(_10407_));
 sg13g2_a21oi_1 _17210_ (.A1(_10405_),
    .A2(_10406_),
    .Y(_10408_),
    .B1(_10407_));
 sg13g2_nand3b_1 _17211_ (.B(net690),
    .C(\cpu.ex.r_epc[13] ),
    .Y(_10409_),
    .A_N(net689));
 sg13g2_nand3b_1 _17212_ (.B(net689),
    .C(\cpu.ex.r_9[13] ),
    .Y(_10410_),
    .A_N(net690));
 sg13g2_nand2b_1 _17213_ (.Y(_10411_),
    .B(net687),
    .A_N(net688));
 sg13g2_a21oi_1 _17214_ (.A1(_10409_),
    .A2(_10410_),
    .Y(_10412_),
    .B1(_10411_));
 sg13g2_nand3b_1 _17215_ (.B(net688),
    .C(\cpu.ex.r_13[13] ),
    .Y(_10413_),
    .A_N(net690));
 sg13g2_nand3b_1 _17216_ (.B(net690),
    .C(\cpu.ex.r_11[13] ),
    .Y(_10414_),
    .A_N(net688));
 sg13g2_nand2_1 _17217_ (.Y(_10415_),
    .A(_10196_),
    .B(net689));
 sg13g2_a21oi_1 _17218_ (.A1(_10413_),
    .A2(_10414_),
    .Y(_10416_),
    .B1(_10415_));
 sg13g2_or3_1 _17219_ (.A(_10408_),
    .B(_10412_),
    .C(_10416_),
    .X(_10417_));
 sg13g2_a221oi_1 _17220_ (.B2(_10404_),
    .C1(_10417_),
    .B1(_10400_),
    .A1(_10220_),
    .Y(_10418_),
    .A2(_10397_));
 sg13g2_nand2_1 _17221_ (.Y(_10419_),
    .A(net696),
    .B(_10238_));
 sg13g2_o21ai_1 _17222_ (.B1(_10419_),
    .Y(_10420_),
    .A1(_10172_),
    .A2(_10418_));
 sg13g2_inv_1 _17223_ (.Y(_10421_),
    .A(\cpu.dec.imm[13] ));
 sg13g2_nor2_1 _17224_ (.A(net890),
    .B(_10421_),
    .Y(_10422_));
 sg13g2_a21oi_1 _17225_ (.A1(net890),
    .A2(_10420_),
    .Y(_10423_),
    .B1(_10422_));
 sg13g2_mux2_1 _17226_ (.A0(_10392_),
    .A1(_10423_),
    .S(net897),
    .X(_10424_));
 sg13g2_buf_1 _17227_ (.A(_10424_),
    .X(_10425_));
 sg13g2_buf_1 _17228_ (.A(_10425_),
    .X(_10426_));
 sg13g2_buf_2 _17229_ (.A(_00270_),
    .X(_10427_));
 sg13g2_nand2b_1 _17230_ (.Y(_10428_),
    .B(net1029),
    .A_N(_10427_));
 sg13g2_buf_1 _17231_ (.A(_10428_),
    .X(_10429_));
 sg13g2_nor2_1 _17232_ (.A(net890),
    .B(\cpu.dec.imm[8] ),
    .Y(_10430_));
 sg13g2_nand3_1 _17233_ (.B(net892),
    .C(net889),
    .A(\cpu.ex.r_epc[8] ),
    .Y(_10431_));
 sg13g2_nand3_1 _17234_ (.B(_10218_),
    .C(net772),
    .A(\cpu.ex.r_8[8] ),
    .Y(_10432_));
 sg13g2_a21oi_1 _17235_ (.A1(_10431_),
    .A2(_10432_),
    .Y(_10433_),
    .B1(net776));
 sg13g2_buf_1 _17236_ (.A(net894),
    .X(_10434_));
 sg13g2_nor2b_1 _17237_ (.A(_00246_),
    .B_N(_10434_),
    .Y(_10435_));
 sg13g2_nor2b_1 _17238_ (.A(_10434_),
    .B_N(\cpu.ex.r_11[8] ),
    .Y(_10436_));
 sg13g2_o21ai_1 _17239_ (.B1(_10222_),
    .Y(_10437_),
    .A1(_10435_),
    .A2(_10436_));
 sg13g2_nand3_1 _17240_ (.B(net1035),
    .C(net774),
    .A(\cpu.ex.r_lr[8] ),
    .Y(_10438_));
 sg13g2_a21oi_1 _17241_ (.A1(_10437_),
    .A2(_10438_),
    .Y(_10439_),
    .B1(net771));
 sg13g2_a22oi_1 _17242_ (.Y(_10440_),
    .B1(net772),
    .B2(\cpu.ex.r_13[8] ),
    .A2(net889),
    .A1(\cpu.ex.r_mult[24] ));
 sg13g2_nor3_1 _17243_ (.A(net771),
    .B(_10206_),
    .C(_10440_),
    .Y(_10441_));
 sg13g2_nor2b_1 _17244_ (.A(net776),
    .B_N(net896),
    .Y(_10442_));
 sg13g2_a22oi_1 _17245_ (.Y(_10443_),
    .B1(_10442_),
    .B2(\cpu.ex.r_10[8] ),
    .A2(_10257_),
    .A1(\cpu.ex.r_12[8] ));
 sg13g2_nor2_1 _17246_ (.A(_10313_),
    .B(_10443_),
    .Y(_10444_));
 sg13g2_nor4_1 _17247_ (.A(_10433_),
    .B(_10439_),
    .C(_10441_),
    .D(_10444_),
    .Y(_10445_));
 sg13g2_nand3_1 _17248_ (.B(_10218_),
    .C(_10339_),
    .A(\cpu.ex.r_14[8] ),
    .Y(_10446_));
 sg13g2_nand3_1 _17249_ (.B(_10195_),
    .C(_10337_),
    .A(\cpu.ex.r_9[8] ),
    .Y(_10447_));
 sg13g2_nand2_1 _17250_ (.Y(_10448_),
    .A(_10446_),
    .B(_10447_));
 sg13g2_buf_1 _17251_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10449_));
 sg13g2_mux2_1 _17252_ (.A0(_10449_),
    .A1(\cpu.ex.r_stmp[8] ),
    .S(net776),
    .X(_10450_));
 sg13g2_a22oi_1 _17253_ (.Y(_10451_),
    .B1(_10450_),
    .B2(_10309_),
    .A2(_10448_),
    .A1(net777));
 sg13g2_a21oi_1 _17254_ (.A1(_10445_),
    .A2(_10451_),
    .Y(_10452_),
    .B1(_10172_));
 sg13g2_and2_1 _17255_ (.A(_09152_),
    .B(net570),
    .X(_10453_));
 sg13g2_nor3_1 _17256_ (.A(net1028),
    .B(_10452_),
    .C(_10453_),
    .Y(_10454_));
 sg13g2_or3_1 _17257_ (.A(net1029),
    .B(_10430_),
    .C(_10454_),
    .X(_10455_));
 sg13g2_buf_1 _17258_ (.A(_10455_),
    .X(_10456_));
 sg13g2_buf_2 _17259_ (.A(_00276_),
    .X(_10457_));
 sg13g2_buf_1 _17260_ (.A(\cpu.dec.user_io ),
    .X(_10458_));
 sg13g2_a22oi_1 _17261_ (.Y(_10459_),
    .B1(_10269_),
    .B2(\cpu.ex.r_8[7] ),
    .A2(_10266_),
    .A1(_10458_));
 sg13g2_buf_1 _17262_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10460_));
 sg13g2_nand3_1 _17263_ (.B(net769),
    .C(net774),
    .A(_10460_),
    .Y(_10461_));
 sg13g2_o21ai_1 _17264_ (.B1(_10461_),
    .Y(_10462_),
    .A1(net778),
    .A2(_10459_));
 sg13g2_a22oi_1 _17265_ (.Y(_10463_),
    .B1(net768),
    .B2(\cpu.ex.r_13[7] ),
    .A2(net774),
    .A1(\cpu.ex.r_lr[7] ));
 sg13g2_o21ai_1 _17266_ (.B1(net1035),
    .Y(_10464_),
    .A1(net891),
    .A2(_10463_));
 sg13g2_mux2_1 _17267_ (.A0(\cpu.ex.r_stmp[7] ),
    .A1(\cpu.ex.r_14[7] ),
    .S(net895),
    .X(_10465_));
 sg13g2_a22oi_1 _17268_ (.Y(_10466_),
    .B1(_10465_),
    .B2(net891),
    .A2(_10342_),
    .A1(\cpu.ex.r_mult[23] ));
 sg13g2_mux2_1 _17269_ (.A0(\cpu.ex.r_10[7] ),
    .A1(\cpu.ex.r_11[7] ),
    .S(net893),
    .X(_10467_));
 sg13g2_a21oi_1 _17270_ (.A1(_10269_),
    .A2(_10467_),
    .Y(_10468_),
    .B1(net1035));
 sg13g2_o21ai_1 _17271_ (.B1(_10468_),
    .Y(_10469_),
    .A1(_10206_),
    .A2(_10466_));
 sg13g2_inv_1 _17272_ (.Y(_10470_),
    .A(_00245_));
 sg13g2_a22oi_1 _17273_ (.Y(_10471_),
    .B1(_10306_),
    .B2(_10470_),
    .A2(net774),
    .A1(\cpu.ex.r_epc[7] ));
 sg13g2_nand3b_1 _17274_ (.B(net766),
    .C(\cpu.ex.r_12[7] ),
    .Y(_10472_),
    .A_N(net893));
 sg13g2_nand3b_1 _17275_ (.B(net893),
    .C(\cpu.ex.r_9[7] ),
    .Y(_10473_),
    .A_N(_10185_));
 sg13g2_a21o_1 _17276_ (.A2(_10473_),
    .A1(_10472_),
    .B1(_10347_),
    .X(_10474_));
 sg13g2_o21ai_1 _17277_ (.B1(_10474_),
    .Y(_10475_),
    .A1(net888),
    .A2(_10471_));
 sg13g2_a221oi_1 _17278_ (.B2(_10469_),
    .C1(_10475_),
    .B1(_10464_),
    .A1(net771),
    .Y(_10476_),
    .A2(_10462_));
 sg13g2_nand2_1 _17279_ (.Y(_10477_),
    .A(_09154_),
    .B(net624));
 sg13g2_o21ai_1 _17280_ (.B1(_10477_),
    .Y(_10478_),
    .A1(_10172_),
    .A2(_10476_));
 sg13g2_nor2b_1 _17281_ (.A(_10242_),
    .B_N(\cpu.dec.imm[7] ),
    .Y(_10479_));
 sg13g2_a21oi_1 _17282_ (.A1(net1030),
    .A2(_10478_),
    .Y(_10480_),
    .B1(_10479_));
 sg13g2_mux2_1 _17283_ (.A0(_10457_),
    .A1(_10480_),
    .S(net897),
    .X(_10481_));
 sg13g2_buf_1 _17284_ (.A(_10481_),
    .X(_10482_));
 sg13g2_buf_1 _17285_ (.A(_10482_),
    .X(_10483_));
 sg13g2_nand4_1 _17286_ (.B(net767),
    .C(net284),
    .A(net217),
    .Y(_10484_),
    .D(net242));
 sg13g2_nor4_1 _17287_ (.A(_10247_),
    .B(net168),
    .C(_10391_),
    .D(_10484_),
    .Y(_10485_));
 sg13g2_buf_1 _17288_ (.A(_00173_),
    .X(_10486_));
 sg13g2_nor2_2 _17289_ (.A(_10151_),
    .B(_10486_),
    .Y(_10487_));
 sg13g2_buf_1 _17290_ (.A(\cpu.dec.imm[3] ),
    .X(_10488_));
 sg13g2_nor2_1 _17291_ (.A(_10488_),
    .B(_10243_),
    .Y(_10489_));
 sg13g2_nor2_1 _17292_ (.A(net775),
    .B(net776),
    .Y(_10490_));
 sg13g2_inv_1 _17293_ (.Y(_10491_),
    .A(\cpu.ex.r_8[3] ));
 sg13g2_buf_1 _17294_ (.A(\cpu.ex.r_sp[3] ),
    .X(_10492_));
 sg13g2_nand3b_1 _17295_ (.B(net769),
    .C(_10492_),
    .Y(_10493_),
    .A_N(net777));
 sg13g2_o21ai_1 _17296_ (.B1(_10493_),
    .Y(_10494_),
    .A1(_10491_),
    .A2(_10347_));
 sg13g2_nor2b_1 _17297_ (.A(net888),
    .B_N(net768),
    .Y(_10495_));
 sg13g2_inv_1 _17298_ (.Y(_10496_),
    .A(_00241_));
 sg13g2_nand2_1 _17299_ (.Y(_10497_),
    .A(\cpu.ex.r_11[3] ),
    .B(net778));
 sg13g2_nand2b_1 _17300_ (.Y(_10498_),
    .B(\cpu.ex.r_9[3] ),
    .A_N(net769));
 sg13g2_a21oi_1 _17301_ (.A1(_10497_),
    .A2(_10498_),
    .Y(_10499_),
    .B1(_10351_));
 sg13g2_a221oi_1 _17302_ (.B2(_10496_),
    .C1(_10499_),
    .B1(_10495_),
    .A1(_10490_),
    .Y(_10500_),
    .A2(_10494_));
 sg13g2_mux2_1 _17303_ (.A0(\cpu.ex.r_stmp[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net770),
    .X(_10501_));
 sg13g2_mux2_1 _17304_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(\cpu.ex.r_mult[19] ),
    .S(net766),
    .X(_10502_));
 sg13g2_a22oi_1 _17305_ (.Y(_10503_),
    .B1(_10502_),
    .B2(_10342_),
    .A2(_10184_),
    .A1(_10501_));
 sg13g2_nand2b_1 _17306_ (.Y(_10504_),
    .B(net778),
    .A_N(_10503_));
 sg13g2_buf_1 _17307_ (.A(\cpu.ex.mmu_read[3] ),
    .X(_10505_));
 sg13g2_mux4_1 _17308_ (.S0(net777),
    .A0(net1135),
    .A1(\cpu.ex.r_12[3] ),
    .A2(_10505_),
    .A3(\cpu.ex.r_13[3] ),
    .S1(net775),
    .X(_10506_));
 sg13g2_nand2_1 _17309_ (.Y(_10507_),
    .A(_10257_),
    .B(_10506_));
 sg13g2_inv_1 _17310_ (.Y(_10508_),
    .A(\cpu.ex.r_10[3] ));
 sg13g2_nor2_1 _17311_ (.A(_10508_),
    .B(_10274_),
    .Y(_10509_));
 sg13g2_and3_1 _17312_ (.X(_10510_),
    .A(\cpu.ex.r_lr[3] ),
    .B(net775),
    .C(net685));
 sg13g2_o21ai_1 _17313_ (.B1(net773),
    .Y(_10511_),
    .A1(_10509_),
    .A2(_10510_));
 sg13g2_nand4_1 _17314_ (.B(_10504_),
    .C(_10507_),
    .A(_10500_),
    .Y(_10512_),
    .D(_10511_));
 sg13g2_a221oi_1 _17315_ (.B2(_10512_),
    .C1(net1028),
    .B1(net569),
    .A1(_09162_),
    .Y(_10513_),
    .A2(net570));
 sg13g2_nor3_2 _17316_ (.A(_10295_),
    .B(_10489_),
    .C(_10513_),
    .Y(_10514_));
 sg13g2_mux2_1 _17317_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(\cpu.ex.r_11[2] ),
    .S(net777),
    .X(_10515_));
 sg13g2_buf_1 _17318_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10516_));
 sg13g2_mux2_1 _17319_ (.A0(net1113),
    .A1(\cpu.ex.r_13[2] ),
    .S(net777),
    .X(_10517_));
 sg13g2_a22oi_1 _17320_ (.Y(_10518_),
    .B1(_10517_),
    .B2(_10257_),
    .A2(_10515_),
    .A1(_10442_));
 sg13g2_nand2b_1 _17321_ (.Y(_10519_),
    .B(net687),
    .A_N(_10518_));
 sg13g2_and3_1 _17322_ (.X(_10520_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net775),
    .C(net685));
 sg13g2_inv_1 _17323_ (.Y(_10521_),
    .A(\cpu.ex.r_10[2] ));
 sg13g2_nor2_1 _17324_ (.A(_10521_),
    .B(_10274_),
    .Y(_10522_));
 sg13g2_o21ai_1 _17325_ (.B1(net773),
    .Y(_10523_),
    .A1(_10520_),
    .A2(_10522_));
 sg13g2_buf_1 _17326_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10524_));
 sg13g2_nor2b_1 _17327_ (.A(_00240_),
    .B_N(net892),
    .Y(_10525_));
 sg13g2_a22oi_1 _17328_ (.Y(_10526_),
    .B1(net768),
    .B2(_10525_),
    .A2(_10169_),
    .A1(_10524_));
 sg13g2_nand2b_1 _17329_ (.Y(_10527_),
    .B(net778),
    .A_N(_10526_));
 sg13g2_nor2_1 _17330_ (.A(net766),
    .B(_10347_),
    .Y(_10528_));
 sg13g2_mux2_1 _17331_ (.A0(\cpu.ex.r_8[2] ),
    .A1(\cpu.ex.r_9[2] ),
    .S(_10194_),
    .X(_10529_));
 sg13g2_mux2_1 _17332_ (.A0(net1131),
    .A1(\cpu.ex.r_stmp[2] ),
    .S(net896),
    .X(_10530_));
 sg13g2_and3_1 _17333_ (.X(_10531_),
    .A(\cpu.ex.r_mult[18] ),
    .B(net892),
    .C(net896));
 sg13g2_a21o_1 _17334_ (.A2(_10530_),
    .A1(net891),
    .B1(_10531_),
    .X(_10532_));
 sg13g2_mux2_1 _17335_ (.A0(\cpu.ex.r_12[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net896),
    .X(_10533_));
 sg13g2_nor2b_1 _17336_ (.A(_10186_),
    .B_N(net770),
    .Y(_10534_));
 sg13g2_and3_1 _17337_ (.X(_10535_),
    .A(net776),
    .B(_10533_),
    .C(_10534_));
 sg13g2_a221oi_1 _17338_ (.B2(_10532_),
    .C1(_10535_),
    .B1(_10266_),
    .A1(_10528_),
    .Y(_10536_),
    .A2(_10529_));
 sg13g2_nand4_1 _17339_ (.B(_10523_),
    .C(_10527_),
    .A(_10519_),
    .Y(_10537_),
    .D(_10536_));
 sg13g2_a22oi_1 _17340_ (.Y(_10538_),
    .B1(net569),
    .B2(_10537_),
    .A2(net570),
    .A1(_09141_));
 sg13g2_nand2_1 _17341_ (.Y(_10539_),
    .A(_10150_),
    .B(net1030));
 sg13g2_buf_1 _17342_ (.A(net1029),
    .X(_10540_));
 sg13g2_inv_1 _17343_ (.Y(_10541_),
    .A(_00271_));
 sg13g2_buf_1 _17344_ (.A(\cpu.dec.imm[2] ),
    .X(_10542_));
 sg13g2_and3_1 _17345_ (.X(_10543_),
    .A(_10542_),
    .B(_10150_),
    .C(net1028));
 sg13g2_a21oi_1 _17346_ (.A1(net887),
    .A2(_10541_),
    .Y(_10544_),
    .B1(_10543_));
 sg13g2_o21ai_1 _17347_ (.B1(_10544_),
    .Y(_10545_),
    .A1(_10538_),
    .A2(_10539_));
 sg13g2_buf_1 _17348_ (.A(_10545_),
    .X(_10546_));
 sg13g2_buf_1 _17349_ (.A(_10546_),
    .X(_10547_));
 sg13g2_nor3_1 _17350_ (.A(_10487_),
    .B(_10514_),
    .C(_10547_),
    .Y(_10548_));
 sg13g2_buf_2 _17351_ (.A(_10548_),
    .X(_10549_));
 sg13g2_buf_1 _17352_ (.A(\cpu.dec.imm[0] ),
    .X(_10550_));
 sg13g2_nor2_1 _17353_ (.A(_10550_),
    .B(_10243_),
    .Y(_10551_));
 sg13g2_a22oi_1 _17354_ (.Y(_10552_),
    .B1(_10339_),
    .B2(\cpu.ex.r_14[0] ),
    .A2(_10337_),
    .A1(\cpu.ex.r_8[0] ));
 sg13g2_mux2_1 _17355_ (.A0(_09133_),
    .A1(\cpu.ex.r_12[0] ),
    .S(net777),
    .X(_10553_));
 sg13g2_nand3_1 _17356_ (.B(_10257_),
    .C(_10553_),
    .A(_10219_),
    .Y(_10554_));
 sg13g2_o21ai_1 _17357_ (.B1(_10554_),
    .Y(_10555_),
    .A1(_10313_),
    .A2(_10552_));
 sg13g2_a22oi_1 _17358_ (.Y(_10556_),
    .B1(_10253_),
    .B2(\cpu.ex.r_9[0] ),
    .A2(_10204_),
    .A1(\cpu.ex.r_10[0] ));
 sg13g2_nor2b_1 _17359_ (.A(_10556_),
    .B_N(_10269_),
    .Y(_10557_));
 sg13g2_nand3_1 _17360_ (.B(_10195_),
    .C(net772),
    .A(\cpu.ex.r_13[0] ),
    .Y(_10558_));
 sg13g2_nand3_1 _17361_ (.B(_10219_),
    .C(net889),
    .A(\cpu.ex.r_stmp[0] ),
    .Y(_10559_));
 sg13g2_a21oi_1 _17362_ (.A1(_10558_),
    .A2(_10559_),
    .Y(_10560_),
    .B1(_10207_));
 sg13g2_buf_1 _17363_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10561_));
 sg13g2_mux4_1 _17364_ (.S0(net777),
    .A0(_10561_),
    .A1(\cpu.ex.r_11[0] ),
    .A2(\cpu.ex.r_mult[16] ),
    .A3(\cpu.ex.r_15[0] ),
    .S1(_10190_),
    .X(_10562_));
 sg13g2_nor2b_1 _17365_ (.A(_10299_),
    .B_N(_10562_),
    .Y(_10563_));
 sg13g2_or4_1 _17366_ (.A(_10555_),
    .B(_10557_),
    .C(_10560_),
    .D(_10563_),
    .X(_10564_));
 sg13g2_a221oi_1 _17367_ (.B2(_10564_),
    .C1(net1028),
    .B1(net569),
    .A1(net1134),
    .Y(_10565_),
    .A2(net570));
 sg13g2_nor3_2 _17368_ (.A(_10540_),
    .B(_10551_),
    .C(_10565_),
    .Y(_10566_));
 sg13g2_buf_1 _17369_ (.A(_10566_),
    .X(_10567_));
 sg13g2_a22oi_1 _17370_ (.Y(_10568_),
    .B1(net768),
    .B2(\cpu.ex.r_13[1] ),
    .A2(net774),
    .A1(\cpu.ex.r_lr[1] ));
 sg13g2_nand2b_1 _17371_ (.Y(_10569_),
    .B(_10253_),
    .A_N(_10568_));
 sg13g2_nor2_1 _17372_ (.A(_10229_),
    .B(net888),
    .Y(_10570_));
 sg13g2_mux2_1 _17373_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(\cpu.ex.r_mult[17] ),
    .S(net766),
    .X(_10571_));
 sg13g2_inv_1 _17374_ (.Y(_10572_),
    .A(\cpu.ex.r_9[1] ));
 sg13g2_nor2_1 _17375_ (.A(_10572_),
    .B(net891),
    .Y(_10573_));
 sg13g2_a22oi_1 _17376_ (.Y(_10574_),
    .B1(_10573_),
    .B2(_10528_),
    .A2(_10571_),
    .A1(_10570_));
 sg13g2_and3_1 _17377_ (.X(_10575_),
    .A(\cpu.ex.mmu_read[1] ),
    .B(net892),
    .C(_10225_));
 sg13g2_inv_1 _17378_ (.Y(_10576_),
    .A(\cpu.ex.r_14[1] ));
 sg13g2_nor2_1 _17379_ (.A(_10576_),
    .B(_10274_),
    .Y(_10577_));
 sg13g2_o21ai_1 _17380_ (.B1(net776),
    .Y(_10578_),
    .A1(_10575_),
    .A2(_10577_));
 sg13g2_and3_1 _17381_ (.X(_10579_),
    .A(_10569_),
    .B(_10574_),
    .C(_10578_));
 sg13g2_a22oi_1 _17382_ (.Y(_10580_),
    .B1(_10269_),
    .B2(\cpu.ex.r_10[1] ),
    .A2(_10266_),
    .A1(\cpu.ex.r_stmp[1] ));
 sg13g2_nor2b_1 _17383_ (.A(_00239_),
    .B_N(net894),
    .Y(_10581_));
 sg13g2_nor2b_1 _17384_ (.A(net766),
    .B_N(\cpu.ex.r_11[1] ),
    .Y(_10582_));
 sg13g2_and2_1 _17385_ (.A(net893),
    .B(net770),
    .X(_10583_));
 sg13g2_o21ai_1 _17386_ (.B1(_10583_),
    .Y(_10584_),
    .A1(_10581_),
    .A2(_10582_));
 sg13g2_o21ai_1 _17387_ (.B1(_10584_),
    .Y(_10585_),
    .A1(net892),
    .A2(_10580_));
 sg13g2_buf_1 _17388_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10586_));
 sg13g2_and3_1 _17389_ (.X(_10587_),
    .A(\cpu.ex.r_12[1] ),
    .B(net895),
    .C(net894));
 sg13g2_a221oi_1 _17390_ (.B2(\cpu.ex.r_8[1] ),
    .C1(_10587_),
    .B1(_10269_),
    .A1(_10586_),
    .Y(_10588_),
    .A2(_10266_));
 sg13g2_buf_1 _17391_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10589_));
 sg13g2_nand3_1 _17392_ (.B(net769),
    .C(net774),
    .A(_10589_),
    .Y(_10590_));
 sg13g2_o21ai_1 _17393_ (.B1(_10590_),
    .Y(_10591_),
    .A1(net778),
    .A2(_10588_));
 sg13g2_a22oi_1 _17394_ (.Y(_10592_),
    .B1(_10591_),
    .B2(net771),
    .A2(_10585_),
    .A1(net778));
 sg13g2_a21o_1 _17395_ (.A2(_10592_),
    .A1(_10579_),
    .B1(_10172_),
    .X(_10593_));
 sg13g2_buf_1 _17396_ (.A(_10593_),
    .X(_10594_));
 sg13g2_a21oi_1 _17397_ (.A1(\cpu.addr[1] ),
    .A2(net624),
    .Y(_10595_),
    .B1(_10539_));
 sg13g2_buf_1 _17398_ (.A(_00182_),
    .X(_10596_));
 sg13g2_buf_1 _17399_ (.A(\cpu.dec.imm[1] ),
    .X(_10597_));
 sg13g2_nor3_1 _17400_ (.A(_10597_),
    .B(_10149_),
    .C(net1030),
    .Y(_10598_));
 sg13g2_a21o_1 _17401_ (.A2(_10596_),
    .A1(net1115),
    .B1(_10598_),
    .X(_10599_));
 sg13g2_a21oi_1 _17402_ (.A1(_10594_),
    .A2(_10595_),
    .Y(_10600_),
    .B1(_10599_));
 sg13g2_buf_8 _17403_ (.A(_10600_),
    .X(_10601_));
 sg13g2_nor2_1 _17404_ (.A(net359),
    .B(net282),
    .Y(_10602_));
 sg13g2_nand2_1 _17405_ (.Y(_10603_),
    .A(_10549_),
    .B(_10602_));
 sg13g2_buf_2 _17406_ (.A(_10603_),
    .X(_10604_));
 sg13g2_nor2_1 _17407_ (.A(_10241_),
    .B(\cpu.dec.imm[5] ),
    .Y(_10605_));
 sg13g2_mux2_1 _17408_ (.A0(\cpu.ex.r_9[5] ),
    .A1(\cpu.ex.r_13[5] ),
    .S(net1036),
    .X(_10606_));
 sg13g2_a22oi_1 _17409_ (.Y(_10607_),
    .B1(_10606_),
    .B2(net895),
    .A2(_10201_),
    .A1(\cpu.ex.r_lr[5] ));
 sg13g2_nand2b_1 _17410_ (.Y(_10608_),
    .B(_10253_),
    .A_N(_10607_));
 sg13g2_nand2b_1 _17411_ (.Y(_10609_),
    .B(net1031),
    .A_N(_00243_));
 sg13g2_nand2b_1 _17412_ (.Y(_10610_),
    .B(\cpu.ex.r_11[5] ),
    .A_N(net1036));
 sg13g2_a21oi_1 _17413_ (.A1(_10609_),
    .A2(_10610_),
    .Y(_10611_),
    .B1(net888));
 sg13g2_nand3b_1 _17414_ (.B(net1033),
    .C(\cpu.ex.r_10[5] ),
    .Y(_10612_),
    .A_N(net1031));
 sg13g2_nand3b_1 _17415_ (.B(net1031),
    .C(\cpu.ex.r_12[5] ),
    .Y(_10613_),
    .A_N(net1114));
 sg13g2_a21oi_1 _17416_ (.A1(_10612_),
    .A2(_10613_),
    .Y(_10614_),
    .B1(net893));
 sg13g2_o21ai_1 _17417_ (.B1(net770),
    .Y(_10615_),
    .A1(_10611_),
    .A2(_10614_));
 sg13g2_nand3_1 _17418_ (.B(net1032),
    .C(net889),
    .A(\cpu.ex.r_epc[5] ),
    .Y(_10616_));
 sg13g2_nand3_1 _17419_ (.B(net891),
    .C(_10209_),
    .A(\cpu.ex.r_8[5] ),
    .Y(_10617_));
 sg13g2_a21o_1 _17420_ (.A2(_10617_),
    .A1(_10616_),
    .B1(net766),
    .X(_10618_));
 sg13g2_inv_1 _17421_ (.Y(_10619_),
    .A(\cpu.ex.r_14[5] ));
 sg13g2_nand3b_1 _17422_ (.B(net1032),
    .C(\cpu.ex.r_mult[21] ),
    .Y(_10620_),
    .A_N(net1034));
 sg13g2_o21ai_1 _17423_ (.B1(_10620_),
    .Y(_10621_),
    .A1(_10619_),
    .A2(_10313_));
 sg13g2_buf_1 _17424_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10622_));
 sg13g2_mux2_1 _17425_ (.A0(_10622_),
    .A1(\cpu.ex.r_stmp[5] ),
    .S(net1031),
    .X(_10623_));
 sg13g2_a22oi_1 _17426_ (.Y(_10624_),
    .B1(_10309_),
    .B2(_10623_),
    .A2(_10621_),
    .A1(_10339_));
 sg13g2_nand4_1 _17427_ (.B(_10615_),
    .C(_10618_),
    .A(_10608_),
    .Y(_10625_),
    .D(_10624_));
 sg13g2_a221oi_1 _17428_ (.B2(_10625_),
    .C1(net1028),
    .B1(net569),
    .A1(_09907_),
    .Y(_10626_),
    .A2(net624));
 sg13g2_or3_1 _17429_ (.A(net1115),
    .B(_10605_),
    .C(_10626_),
    .X(_10627_));
 sg13g2_buf_1 _17430_ (.A(_10627_),
    .X(_10628_));
 sg13g2_buf_1 _17431_ (.A(_00278_),
    .X(_10629_));
 sg13g2_nand2b_1 _17432_ (.Y(_10630_),
    .B(net1115),
    .A_N(_10629_));
 sg13g2_buf_1 _17433_ (.A(_10630_),
    .X(_10631_));
 sg13g2_and2_1 _17434_ (.A(_10628_),
    .B(_10631_),
    .X(_10632_));
 sg13g2_buf_1 _17435_ (.A(_10632_),
    .X(_10633_));
 sg13g2_buf_1 _17436_ (.A(_10633_),
    .X(_10634_));
 sg13g2_buf_1 _17437_ (.A(net241),
    .X(_10635_));
 sg13g2_mux2_1 _17438_ (.A0(\cpu.ex.r_lr[4] ),
    .A1(\cpu.ex.r_9[4] ),
    .S(net770),
    .X(_10636_));
 sg13g2_a22oi_1 _17439_ (.Y(_10637_),
    .B1(_10636_),
    .B2(net1035),
    .A2(_10222_),
    .A1(\cpu.ex.r_11[4] ));
 sg13g2_nand3_1 _17440_ (.B(net891),
    .C(net772),
    .A(\cpu.ex.r_8[4] ),
    .Y(_10638_));
 sg13g2_o21ai_1 _17441_ (.B1(_10638_),
    .Y(_10639_),
    .A1(net771),
    .A2(_10637_));
 sg13g2_a221oi_1 _17442_ (.B2(_08285_),
    .C1(net769),
    .B1(_10230_),
    .A1(\cpu.ex.r_13[4] ),
    .Y(_10640_),
    .A2(_10583_));
 sg13g2_a221oi_1 _17443_ (.B2(\cpu.ex.r_14[4] ),
    .C1(net1035),
    .B1(_10534_),
    .A1(\cpu.ex.r_mult[20] ),
    .Y(_10641_),
    .A2(_10342_));
 sg13g2_nor3_1 _17444_ (.A(_10206_),
    .B(_10640_),
    .C(_10641_),
    .Y(_10642_));
 sg13g2_a21oi_1 _17445_ (.A1(net773),
    .A2(_10639_),
    .Y(_10643_),
    .B1(_10642_));
 sg13g2_buf_1 _17446_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10644_));
 sg13g2_mux2_1 _17447_ (.A0(_10644_),
    .A1(\cpu.ex.r_10[4] ),
    .S(net770),
    .X(_10645_));
 sg13g2_a22oi_1 _17448_ (.Y(_10646_),
    .B1(_10645_),
    .B2(_10206_),
    .A2(_10266_),
    .A1(\cpu.ex.r_stmp[4] ));
 sg13g2_a21oi_1 _17449_ (.A1(\cpu.ex.r_12[4] ),
    .A2(net768),
    .Y(_10647_),
    .B1(net778));
 sg13g2_a21oi_1 _17450_ (.A1(net778),
    .A2(_10646_),
    .Y(_10648_),
    .B1(_10647_));
 sg13g2_inv_1 _17451_ (.Y(_10649_),
    .A(_00242_));
 sg13g2_a22oi_1 _17452_ (.Y(_10650_),
    .B1(net768),
    .B2(_10649_),
    .A2(net774),
    .A1(\cpu.ex.r_epc[4] ));
 sg13g2_nor2_1 _17453_ (.A(net888),
    .B(_10650_),
    .Y(_10651_));
 sg13g2_a21oi_1 _17454_ (.A1(net771),
    .A2(_10648_),
    .Y(_10652_),
    .B1(_10651_));
 sg13g2_a21oi_1 _17455_ (.A1(_10643_),
    .A2(_10652_),
    .Y(_10653_),
    .B1(_10172_));
 sg13g2_a21o_1 _17456_ (.A2(net624),
    .A1(_09453_),
    .B1(_10539_),
    .X(_10654_));
 sg13g2_nor3_1 _17457_ (.A(net1115),
    .B(net1030),
    .C(\cpu.dec.imm[4] ),
    .Y(_10655_));
 sg13g2_a21oi_1 _17458_ (.A1(_08449_),
    .A2(_10295_),
    .Y(_10656_),
    .B1(_10655_));
 sg13g2_o21ai_1 _17459_ (.B1(_10656_),
    .Y(_10657_),
    .A1(_10653_),
    .A2(_10654_));
 sg13g2_buf_1 _17460_ (.A(_10657_),
    .X(_10658_));
 sg13g2_buf_1 _17461_ (.A(net358),
    .X(_10659_));
 sg13g2_nand2_1 _17462_ (.Y(_10660_),
    .A(net216),
    .B(net281));
 sg13g2_buf_1 _17463_ (.A(_00272_),
    .X(_10661_));
 sg13g2_nand2b_1 _17464_ (.Y(_10662_),
    .B(net887),
    .A_N(_10661_));
 sg13g2_nor2_1 _17465_ (.A(net890),
    .B(\cpu.dec.imm[12] ),
    .Y(_10663_));
 sg13g2_buf_1 _17466_ (.A(\cpu.ex.r_sp[12] ),
    .X(_10664_));
 sg13g2_and2_1 _17467_ (.A(\cpu.ex.r_10[12] ),
    .B(net777),
    .X(_10665_));
 sg13g2_a21oi_1 _17468_ (.A1(_10664_),
    .A2(_10356_),
    .Y(_10666_),
    .B1(_10665_));
 sg13g2_nand3_1 _17469_ (.B(net687),
    .C(net772),
    .A(\cpu.ex.r_9[12] ),
    .Y(_10667_));
 sg13g2_o21ai_1 _17470_ (.B1(_10667_),
    .Y(_10668_),
    .A1(_10308_),
    .A2(_10666_));
 sg13g2_a22oi_1 _17471_ (.Y(_10669_),
    .B1(net685),
    .B2(\cpu.ex.r_lr[12] ),
    .A2(_10222_),
    .A1(\cpu.ex.r_11[12] ));
 sg13g2_nor2_1 _17472_ (.A(net686),
    .B(_10669_),
    .Y(_10670_));
 sg13g2_o21ai_1 _17473_ (.B1(net773),
    .Y(_10671_),
    .A1(_10668_),
    .A2(_10670_));
 sg13g2_a22oi_1 _17474_ (.Y(_10672_),
    .B1(net772),
    .B2(\cpu.ex.r_13[12] ),
    .A2(net889),
    .A1(\cpu.ex.r_mult[28] ));
 sg13g2_nor2_1 _17475_ (.A(net686),
    .B(_10672_),
    .Y(_10673_));
 sg13g2_and3_1 _17476_ (.X(_10674_),
    .A(\cpu.ex.r_12[12] ),
    .B(net686),
    .C(net772));
 sg13g2_o21ai_1 _17477_ (.B1(net623),
    .Y(_10675_),
    .A1(_10673_),
    .A2(_10674_));
 sg13g2_buf_2 _17478_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10676_));
 sg13g2_a22oi_1 _17479_ (.Y(_10677_),
    .B1(_10442_),
    .B2(\cpu.ex.r_epc[12] ),
    .A2(_10257_),
    .A1(_10676_));
 sg13g2_nand3_1 _17480_ (.B(net686),
    .C(_10339_),
    .A(\cpu.ex.r_stmp[12] ),
    .Y(_10678_));
 sg13g2_o21ai_1 _17481_ (.B1(_10678_),
    .Y(_10679_),
    .A1(net686),
    .A2(_10677_));
 sg13g2_nor3_1 _17482_ (.A(_00250_),
    .B(_10356_),
    .C(net888),
    .Y(_10680_));
 sg13g2_a22oi_1 _17483_ (.Y(_10681_),
    .B1(_10680_),
    .B2(net623),
    .A2(_10679_),
    .A1(_10356_));
 sg13g2_a22oi_1 _17484_ (.Y(_10682_),
    .B1(_10339_),
    .B2(\cpu.ex.r_14[12] ),
    .A2(_10337_),
    .A1(\cpu.ex.r_8[12] ));
 sg13g2_nand2b_1 _17485_ (.Y(_10683_),
    .B(_10534_),
    .A_N(_10682_));
 sg13g2_nand4_1 _17486_ (.B(_10675_),
    .C(_10681_),
    .A(_10671_),
    .Y(_10684_),
    .D(_10683_));
 sg13g2_a221oi_1 _17487_ (.B2(_10684_),
    .C1(_10324_),
    .B1(net501),
    .A1(net695),
    .Y(_10685_),
    .A2(net570));
 sg13g2_or3_1 _17488_ (.A(net887),
    .B(_10663_),
    .C(_10685_),
    .X(_10686_));
 sg13g2_buf_1 _17489_ (.A(_10686_),
    .X(_10687_));
 sg13g2_nand2_1 _17490_ (.Y(_10688_),
    .A(_10662_),
    .B(_10687_));
 sg13g2_buf_2 _17491_ (.A(_10688_),
    .X(_10689_));
 sg13g2_buf_1 _17492_ (.A(_10689_),
    .X(_10690_));
 sg13g2_nor2_1 _17493_ (.A(net897),
    .B(_00273_),
    .Y(_10691_));
 sg13g2_nor2_1 _17494_ (.A(net1030),
    .B(\cpu.dec.imm[11] ),
    .Y(_10692_));
 sg13g2_buf_2 _17495_ (.A(\cpu.addr[11] ),
    .X(_10693_));
 sg13g2_a221oi_1 _17496_ (.B2(\cpu.ex.r_9[11] ),
    .C1(net769),
    .B1(_10187_),
    .A1(\cpu.ex.r_12[11] ),
    .Y(_10694_),
    .A2(_10184_));
 sg13g2_a221oi_1 _17497_ (.B2(\cpu.ex.r_11[11] ),
    .C1(net1035),
    .B1(_10187_),
    .A1(\cpu.ex.r_14[11] ),
    .Y(_10695_),
    .A2(_10184_));
 sg13g2_or3_1 _17498_ (.A(_10356_),
    .B(_10694_),
    .C(_10695_),
    .X(_10696_));
 sg13g2_buf_1 _17499_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10697_));
 sg13g2_nor2_1 _17500_ (.A(_10375_),
    .B(_10308_),
    .Y(_10698_));
 sg13g2_mux2_1 _17501_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(\cpu.ex.r_mult[27] ),
    .S(net766),
    .X(_10699_));
 sg13g2_nand2b_1 _17502_ (.Y(_10700_),
    .B(_10301_),
    .A_N(_00249_));
 sg13g2_nand2b_1 _17503_ (.Y(_10701_),
    .B(\cpu.ex.r_13[11] ),
    .A_N(net896));
 sg13g2_nand3_1 _17504_ (.B(net770),
    .C(net766),
    .A(_10194_),
    .Y(_10702_));
 sg13g2_a21oi_1 _17505_ (.A1(_10700_),
    .A2(_10701_),
    .Y(_10703_),
    .B1(_10702_));
 sg13g2_a221oi_1 _17506_ (.B2(_10570_),
    .C1(_10703_),
    .B1(_10699_),
    .A1(_10697_),
    .Y(_10704_),
    .A2(_10698_));
 sg13g2_and3_1 _17507_ (.X(_10705_),
    .A(\cpu.ex.r_lr[11] ),
    .B(net892),
    .C(net685));
 sg13g2_inv_1 _17508_ (.Y(_10706_),
    .A(\cpu.ex.r_10[11] ));
 sg13g2_nor2_1 _17509_ (.A(_10706_),
    .B(_10274_),
    .Y(_10707_));
 sg13g2_o21ai_1 _17510_ (.B1(_10207_),
    .Y(_10708_),
    .A1(_10705_),
    .A2(_10707_));
 sg13g2_nand3_1 _17511_ (.B(_10206_),
    .C(_10209_),
    .A(\cpu.ex.r_8[11] ),
    .Y(_10709_));
 sg13g2_nand3_1 _17512_ (.B(_10189_),
    .C(_10281_),
    .A(\cpu.ex.r_stmp[11] ),
    .Y(_10710_));
 sg13g2_a21o_1 _17513_ (.A2(_10710_),
    .A1(_10709_),
    .B1(net775),
    .X(_10711_));
 sg13g2_nand4_1 _17514_ (.B(_10704_),
    .C(_10708_),
    .A(_10696_),
    .Y(_10712_),
    .D(_10711_));
 sg13g2_a221oi_1 _17515_ (.B2(_10712_),
    .C1(_10324_),
    .B1(_10250_),
    .A1(_10693_),
    .Y(_10713_),
    .A2(_10166_));
 sg13g2_nor3_2 _17516_ (.A(net1029),
    .B(_10692_),
    .C(_10713_),
    .Y(_10714_));
 sg13g2_or2_1 _17517_ (.X(_10715_),
    .B(_10714_),
    .A(_10691_));
 sg13g2_buf_1 _17518_ (.A(_10715_),
    .X(_10716_));
 sg13g2_buf_1 _17519_ (.A(_10716_),
    .X(_10717_));
 sg13g2_nor4_1 _17520_ (.A(_10604_),
    .B(_10660_),
    .C(net194),
    .D(net240),
    .Y(_10718_));
 sg13g2_nor2_1 _17521_ (.A(net1124),
    .B(net504),
    .Y(_10719_));
 sg13g2_o21ai_1 _17522_ (.B1(_10719_),
    .Y(_10720_),
    .A1(_09257_),
    .A2(_09275_));
 sg13g2_a21oi_1 _17523_ (.A1(_10485_),
    .A2(_10718_),
    .Y(_10721_),
    .B1(_10720_));
 sg13g2_buf_2 _17524_ (.A(_10721_),
    .X(_10722_));
 sg13g2_inv_1 _17525_ (.Y(_10723_),
    .A(_10722_));
 sg13g2_buf_1 _17526_ (.A(_10723_),
    .X(_10724_));
 sg13g2_buf_2 _17527_ (.A(_00285_),
    .X(_10725_));
 sg13g2_nor2_1 _17528_ (.A(_10725_),
    .B(net573),
    .Y(_10726_));
 sg13g2_buf_1 _17529_ (.A(_10726_),
    .X(_10727_));
 sg13g2_or2_1 _17530_ (.X(_10728_),
    .B(_10326_),
    .A(_10294_));
 sg13g2_buf_2 _17531_ (.A(_10728_),
    .X(_10729_));
 sg13g2_mux2_1 _17532_ (.A0(_10725_),
    .A1(net446),
    .S(_10729_),
    .X(_10730_));
 sg13g2_buf_2 _17533_ (.A(_00283_),
    .X(_10731_));
 sg13g2_a22oi_1 _17534_ (.Y(_10732_),
    .B1(_10730_),
    .B2(_10731_),
    .A2(net243),
    .A1(_09275_));
 sg13g2_nor2_2 _17535_ (.A(_10731_),
    .B(net573),
    .Y(_10733_));
 sg13g2_xnor2_1 _17536_ (.Y(_10734_),
    .A(_10725_),
    .B(_10328_));
 sg13g2_nand3_1 _17537_ (.B(_10733_),
    .C(_10734_),
    .A(_10716_),
    .Y(_10735_));
 sg13g2_o21ai_1 _17538_ (.B1(_10735_),
    .Y(_10736_),
    .A1(net240),
    .A2(_10732_));
 sg13g2_buf_2 _17539_ (.A(_00286_),
    .X(_10737_));
 sg13g2_and3_1 _17540_ (.X(_10738_),
    .A(_10737_),
    .B(net767),
    .C(net284));
 sg13g2_a21oi_1 _17541_ (.A1(net767),
    .A2(net284),
    .Y(_10739_),
    .B1(_10737_));
 sg13g2_buf_2 _17542_ (.A(_00284_),
    .X(_10740_));
 sg13g2_nand2_1 _17543_ (.Y(_10741_),
    .A(\cpu.dec.div ),
    .B(net710));
 sg13g2_buf_1 _17544_ (.A(_10741_),
    .X(_10742_));
 sg13g2_nand2b_1 _17545_ (.Y(_10743_),
    .B(_10742_),
    .A_N(_10740_));
 sg13g2_nor2_1 _17546_ (.A(_10389_),
    .B(_10743_),
    .Y(_10744_));
 sg13g2_o21ai_1 _17547_ (.B1(_10744_),
    .Y(_10745_),
    .A1(_10738_),
    .A2(_10739_));
 sg13g2_and2_1 _17548_ (.A(net767),
    .B(net284),
    .X(_10746_));
 sg13g2_buf_1 _17549_ (.A(_10746_),
    .X(_10747_));
 sg13g2_nand3_1 _17550_ (.B(_10747_),
    .C(net285),
    .A(net450),
    .Y(_10748_));
 sg13g2_inv_1 _17551_ (.Y(_10749_),
    .A(_10737_));
 sg13g2_nand2_2 _17552_ (.Y(_10750_),
    .A(_10749_),
    .B(_10742_));
 sg13g2_a21oi_1 _17553_ (.A1(net767),
    .A2(net284),
    .Y(_10751_),
    .B1(_10750_));
 sg13g2_and2_1 _17554_ (.A(_10740_),
    .B(_10389_),
    .X(_10752_));
 sg13g2_o21ai_1 _17555_ (.B1(_10752_),
    .Y(_10753_),
    .A1(_10738_),
    .A2(_10751_));
 sg13g2_nand3_1 _17556_ (.B(_10748_),
    .C(_10753_),
    .A(_10745_),
    .Y(_10754_));
 sg13g2_nor2_1 _17557_ (.A(_10737_),
    .B(net573),
    .Y(_10755_));
 sg13g2_buf_1 _17558_ (.A(_10755_),
    .X(_10756_));
 sg13g2_nand4_1 _17559_ (.B(net767),
    .C(net284),
    .A(_10328_),
    .Y(_10757_),
    .D(_10756_));
 sg13g2_and3_1 _17560_ (.X(_10758_),
    .A(net767),
    .B(net446),
    .C(_10756_));
 sg13g2_a22oi_1 _17561_ (.Y(_10759_),
    .B1(_10758_),
    .B2(net284),
    .A2(_10727_),
    .A1(_10328_));
 sg13g2_nor2_1 _17562_ (.A(_10691_),
    .B(_10714_),
    .Y(_10760_));
 sg13g2_buf_1 _17563_ (.A(_10760_),
    .X(_10761_));
 sg13g2_nor2_1 _17564_ (.A(_10740_),
    .B(net505),
    .Y(_10762_));
 sg13g2_nand2_1 _17565_ (.Y(_10763_),
    .A(net280),
    .B(_10762_));
 sg13g2_nand2_1 _17566_ (.Y(_10764_),
    .A(_10389_),
    .B(net280));
 sg13g2_a22oi_1 _17567_ (.Y(_10765_),
    .B1(_10763_),
    .B2(_10764_),
    .A2(_10759_),
    .A1(_10757_));
 sg13g2_nand2_1 _17568_ (.Y(_10766_),
    .A(_10389_),
    .B(_10733_));
 sg13g2_or3_1 _17569_ (.A(_10731_),
    .B(_10740_),
    .C(_09274_),
    .X(_10767_));
 sg13g2_a22oi_1 _17570_ (.Y(_10768_),
    .B1(_10766_),
    .B2(_10767_),
    .A2(_10759_),
    .A1(_10757_));
 sg13g2_nor3_1 _17571_ (.A(_10731_),
    .B(_10740_),
    .C(net505),
    .Y(_10769_));
 sg13g2_a22oi_1 _17572_ (.Y(_10770_),
    .B1(_10769_),
    .B2(_10389_),
    .A2(_10733_),
    .A1(net280));
 sg13g2_o21ai_1 _17573_ (.B1(_10770_),
    .Y(_10771_),
    .A1(_10764_),
    .A2(_10743_));
 sg13g2_or3_1 _17574_ (.A(_10765_),
    .B(_10768_),
    .C(_10771_),
    .X(_10772_));
 sg13g2_buf_1 _17575_ (.A(_10772_),
    .X(_10773_));
 sg13g2_a21oi_2 _17576_ (.B1(_10773_),
    .Y(_10774_),
    .A2(_10754_),
    .A1(_10736_));
 sg13g2_inv_1 _17577_ (.Y(_10775_),
    .A(_09259_));
 sg13g2_nor3_1 _17578_ (.A(_09258_),
    .B(_10775_),
    .C(\cpu.ex.c_mult_off[0] ),
    .Y(_10776_));
 sg13g2_inv_1 _17579_ (.Y(_10777_),
    .A(_09118_));
 sg13g2_nor2_1 _17580_ (.A(_10777_),
    .B(_09134_),
    .Y(_10778_));
 sg13g2_o21ai_1 _17581_ (.B1(_10778_),
    .Y(_10779_),
    .A1(_09098_),
    .A2(_09117_));
 sg13g2_a21oi_1 _17582_ (.A1(_09133_),
    .A2(_09131_),
    .Y(_10780_),
    .B1(_09087_));
 sg13g2_buf_1 _17583_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10781_));
 sg13g2_buf_8 _17584_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10782_));
 sg13g2_nor2_1 _17585_ (.A(_10781_),
    .B(_10782_),
    .Y(_10783_));
 sg13g2_buf_2 _17586_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10784_));
 sg13g2_buf_8 _17587_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10785_));
 sg13g2_nor2_1 _17588_ (.A(_10784_),
    .B(_10785_),
    .Y(_10786_));
 sg13g2_a21oi_1 _17589_ (.A1(_10783_),
    .A2(_10786_),
    .Y(_10787_),
    .B1(_00254_));
 sg13g2_nand3_1 _17590_ (.B(_10780_),
    .C(_10787_),
    .A(_10779_),
    .Y(_10788_));
 sg13g2_buf_1 _17591_ (.A(_10788_),
    .X(_10789_));
 sg13g2_nor2_2 _17592_ (.A(_08330_),
    .B(_10789_),
    .Y(_10790_));
 sg13g2_buf_2 _17593_ (.A(\cpu.br ),
    .X(_10791_));
 sg13g2_inv_1 _17594_ (.Y(_10792_),
    .A(_10791_));
 sg13g2_a21o_1 _17595_ (.A2(_10790_),
    .A1(net459),
    .B1(_10792_),
    .X(_10793_));
 sg13g2_buf_2 _17596_ (.A(_10793_),
    .X(_10794_));
 sg13g2_buf_8 _17597_ (.A(_10794_),
    .X(_10795_));
 sg13g2_buf_8 _17598_ (.A(net279),
    .X(_10796_));
 sg13g2_buf_8 _17599_ (.A(net1111),
    .X(_10797_));
 sg13g2_buf_8 _17600_ (.A(_10782_),
    .X(_10798_));
 sg13g2_and2_1 _17601_ (.A(net1027),
    .B(net1026),
    .X(_10799_));
 sg13g2_buf_1 _17602_ (.A(_10799_),
    .X(_10800_));
 sg13g2_buf_1 _17603_ (.A(net1027),
    .X(_10801_));
 sg13g2_buf_1 _17604_ (.A(_10798_),
    .X(_10802_));
 sg13g2_nor2_1 _17605_ (.A(net886),
    .B(net885),
    .Y(_10803_));
 sg13g2_a22oi_1 _17606_ (.Y(_10804_),
    .B1(_10803_),
    .B2(\cpu.ex.r_lr[12] ),
    .A2(_10800_),
    .A1(\cpu.ex.r_mult[28] ));
 sg13g2_buf_8 _17607_ (.A(_10784_),
    .X(_10805_));
 sg13g2_buf_8 _17608_ (.A(net1025),
    .X(_10806_));
 sg13g2_inv_2 _17609_ (.Y(_10807_),
    .A(net884));
 sg13g2_buf_8 _17610_ (.A(net1112),
    .X(_10808_));
 sg13g2_buf_8 _17611_ (.A(net1024),
    .X(_10809_));
 sg13g2_nor2_1 _17612_ (.A(_10807_),
    .B(net883),
    .Y(_10810_));
 sg13g2_nor2b_1 _17613_ (.A(_10804_),
    .B_N(_10810_),
    .Y(_10811_));
 sg13g2_buf_8 _17614_ (.A(net1026),
    .X(_10812_));
 sg13g2_buf_8 _17615_ (.A(net882),
    .X(_10813_));
 sg13g2_nor2b_1 _17616_ (.A(_10784_),
    .B_N(net1111),
    .Y(_10814_));
 sg13g2_buf_1 _17617_ (.A(_10814_),
    .X(_10815_));
 sg13g2_buf_1 _17618_ (.A(_10815_),
    .X(_10816_));
 sg13g2_nand3_1 _17619_ (.B(\cpu.ex.r_14[12] ),
    .C(net764),
    .A(net765),
    .Y(_10817_));
 sg13g2_inv_1 _17620_ (.Y(_10818_),
    .A(net1026));
 sg13g2_buf_1 _17621_ (.A(_10818_),
    .X(_10819_));
 sg13g2_nor2b_1 _17622_ (.A(net1027),
    .B_N(net1025),
    .Y(_10820_));
 sg13g2_buf_2 _17623_ (.A(_10820_),
    .X(_10821_));
 sg13g2_nand3_1 _17624_ (.B(\cpu.ex.r_9[12] ),
    .C(_10821_),
    .A(net763),
    .Y(_10822_));
 sg13g2_inv_2 _17625_ (.Y(_10823_),
    .A(net1024));
 sg13g2_a21oi_1 _17626_ (.A1(_10817_),
    .A2(_10822_),
    .Y(_10824_),
    .B1(_10823_));
 sg13g2_nand2_1 _17627_ (.Y(_10825_),
    .A(net1112),
    .B(net1026));
 sg13g2_nand2b_1 _17628_ (.Y(_10826_),
    .B(_10784_),
    .A_N(net1111));
 sg13g2_buf_1 _17629_ (.A(_10826_),
    .X(_10827_));
 sg13g2_nor2_1 _17630_ (.A(_10825_),
    .B(_10827_),
    .Y(_10828_));
 sg13g2_buf_2 _17631_ (.A(_10828_),
    .X(_10829_));
 sg13g2_nand4_1 _17632_ (.B(net1111),
    .C(net1112),
    .A(_10805_),
    .Y(_10830_),
    .D(_10782_));
 sg13g2_buf_2 _17633_ (.A(_10830_),
    .X(_10831_));
 sg13g2_nor2_1 _17634_ (.A(_00250_),
    .B(_10831_),
    .Y(_10832_));
 sg13g2_a21oi_1 _17635_ (.A1(\cpu.ex.r_13[12] ),
    .A2(_10829_),
    .Y(_10833_),
    .B1(_10832_));
 sg13g2_and2_1 _17636_ (.A(_10784_),
    .B(\cpu.dec.r_rs1[1] ),
    .X(_10834_));
 sg13g2_buf_1 _17637_ (.A(_10834_),
    .X(_10835_));
 sg13g2_and2_1 _17638_ (.A(_10783_),
    .B(net881),
    .X(_10836_));
 sg13g2_buf_1 _17639_ (.A(_10836_),
    .X(_10837_));
 sg13g2_buf_1 _17640_ (.A(_10837_),
    .X(_10838_));
 sg13g2_and2_1 _17641_ (.A(net1112),
    .B(_10782_),
    .X(_10839_));
 sg13g2_buf_8 _17642_ (.A(_10839_),
    .X(_10840_));
 sg13g2_and2_1 _17643_ (.A(_10786_),
    .B(_10840_),
    .X(_10841_));
 sg13g2_buf_1 _17644_ (.A(_10841_),
    .X(_10842_));
 sg13g2_a22oi_1 _17645_ (.Y(_10843_),
    .B1(net684),
    .B2(\cpu.ex.r_12[12] ),
    .A2(net621),
    .A1(\cpu.ex.r_epc[12] ));
 sg13g2_nand3b_1 _17646_ (.B(_10833_),
    .C(_10843_),
    .Y(_10844_),
    .A_N(_10824_));
 sg13g2_nor2b_2 _17647_ (.A(net1025),
    .B_N(net1112),
    .Y(_10845_));
 sg13g2_nand3_1 _17648_ (.B(\cpu.ex.r_8[12] ),
    .C(_10845_),
    .A(net763),
    .Y(_10846_));
 sg13g2_buf_8 _17649_ (.A(net884),
    .X(_10847_));
 sg13g2_nor2b_1 _17650_ (.A(net1112),
    .B_N(_10782_),
    .Y(_10848_));
 sg13g2_buf_1 _17651_ (.A(_10848_),
    .X(_10849_));
 sg13g2_buf_1 _17652_ (.A(_10849_),
    .X(_10850_));
 sg13g2_nand3_1 _17653_ (.B(_10676_),
    .C(net761),
    .A(_10847_),
    .Y(_10851_));
 sg13g2_buf_1 _17654_ (.A(net1027),
    .X(_10852_));
 sg13g2_a21o_1 _17655_ (.A2(_10851_),
    .A1(_10846_),
    .B1(net880),
    .X(_10853_));
 sg13g2_and2_1 _17656_ (.A(_10815_),
    .B(_10849_),
    .X(_10854_));
 sg13g2_buf_1 _17657_ (.A(_10854_),
    .X(_10855_));
 sg13g2_nor2b_1 _17658_ (.A(_10782_),
    .B_N(\cpu.dec.r_rs1[3] ),
    .Y(_10856_));
 sg13g2_buf_1 _17659_ (.A(_10856_),
    .X(_10857_));
 sg13g2_and2_1 _17660_ (.A(_10835_),
    .B(_10857_),
    .X(_10858_));
 sg13g2_buf_2 _17661_ (.A(_10858_),
    .X(_10859_));
 sg13g2_a22oi_1 _17662_ (.Y(_10860_),
    .B1(_10859_),
    .B2(\cpu.ex.r_11[12] ),
    .A2(_10855_),
    .A1(\cpu.ex.r_stmp[12] ));
 sg13g2_and2_1 _17663_ (.A(_10815_),
    .B(_10857_),
    .X(_10861_));
 sg13g2_buf_2 _17664_ (.A(_10861_),
    .X(_10862_));
 sg13g2_buf_1 _17665_ (.A(_10783_),
    .X(_10863_));
 sg13g2_and2_1 _17666_ (.A(net879),
    .B(net764),
    .X(_10864_));
 sg13g2_a22oi_1 _17667_ (.Y(_10865_),
    .B1(_10864_),
    .B2(_10664_),
    .A2(_10862_),
    .A1(\cpu.ex.r_10[12] ));
 sg13g2_nand3_1 _17668_ (.B(_10860_),
    .C(_10865_),
    .A(_10853_),
    .Y(_10866_));
 sg13g2_nor3_1 _17669_ (.A(_10811_),
    .B(_10844_),
    .C(_10866_),
    .Y(_10867_));
 sg13g2_xor2_1 _17670_ (.B(_10781_),
    .A(net1117),
    .X(_10868_));
 sg13g2_xor2_1 _17671_ (.B(_10784_),
    .A(_10143_),
    .X(_10869_));
 sg13g2_xor2_1 _17672_ (.B(_10782_),
    .A(_10140_),
    .X(_10870_));
 sg13g2_xor2_1 _17673_ (.B(_10785_),
    .A(_10142_),
    .X(_10871_));
 sg13g2_nor4_1 _17674_ (.A(_10868_),
    .B(_10869_),
    .C(_10870_),
    .D(_10871_),
    .Y(_10872_));
 sg13g2_nand2b_1 _17675_ (.Y(_10873_),
    .B(_10872_),
    .A_N(_10164_));
 sg13g2_buf_2 _17676_ (.A(_10873_),
    .X(_10874_));
 sg13g2_buf_8 _17677_ (.A(_10874_),
    .X(_10875_));
 sg13g2_mux2_1 _17678_ (.A0(_09576_),
    .A1(_10867_),
    .S(net620),
    .X(_10876_));
 sg13g2_nand2b_1 _17679_ (.Y(_10877_),
    .B(net279),
    .A_N(_10876_));
 sg13g2_o21ai_1 _17680_ (.B1(_10877_),
    .Y(_10878_),
    .A1(_10661_),
    .A2(net239));
 sg13g2_buf_1 _17681_ (.A(_10878_),
    .X(_10879_));
 sg13g2_xor2_1 _17682_ (.B(_09258_),
    .A(_09260_),
    .X(_10880_));
 sg13g2_nor3_1 _17683_ (.A(_09260_),
    .B(_09258_),
    .C(_09259_),
    .Y(_10881_));
 sg13g2_o21ai_1 _17684_ (.B1(_09259_),
    .Y(_10882_),
    .A1(_09260_),
    .A2(_09258_));
 sg13g2_nor2b_1 _17685_ (.A(_10881_),
    .B_N(_10882_),
    .Y(_10883_));
 sg13g2_o21ai_1 _17686_ (.B1(_09271_),
    .Y(_10884_),
    .A1(_10880_),
    .A2(_10883_));
 sg13g2_nor2_1 _17687_ (.A(net1073),
    .B(_10875_),
    .Y(_10885_));
 sg13g2_buf_1 _17688_ (.A(net762),
    .X(_10886_));
 sg13g2_buf_8 _17689_ (.A(_10857_),
    .X(_10887_));
 sg13g2_a22oi_1 _17690_ (.Y(_10888_),
    .B1(net760),
    .B2(\cpu.ex.r_11[14] ),
    .A2(_10850_),
    .A1(\cpu.ex.r_mult[30] ));
 sg13g2_a221oi_1 _17691_ (.B2(\cpu.ex.r_9[14] ),
    .C1(_10801_),
    .B1(net760),
    .A1(_10275_),
    .Y(_10889_),
    .A2(_10849_));
 sg13g2_a21oi_1 _17692_ (.A1(_10852_),
    .A2(_10888_),
    .Y(_10890_),
    .B1(_10889_));
 sg13g2_nand2_1 _17693_ (.Y(_10891_),
    .A(net683),
    .B(_10890_));
 sg13g2_buf_1 _17694_ (.A(net883),
    .X(_10892_));
 sg13g2_nand2b_1 _17695_ (.Y(_10893_),
    .B(net1111),
    .A_N(_10784_));
 sg13g2_buf_1 _17696_ (.A(_10893_),
    .X(_10894_));
 sg13g2_nor2_1 _17697_ (.A(_10818_),
    .B(net878),
    .Y(_10895_));
 sg13g2_nor2_1 _17698_ (.A(_10802_),
    .B(_10827_),
    .Y(_10896_));
 sg13g2_a22oi_1 _17699_ (.Y(_10897_),
    .B1(_10896_),
    .B2(\cpu.ex.r_lr[14] ),
    .A2(_10895_),
    .A1(\cpu.ex.r_stmp[14] ));
 sg13g2_or2_1 _17700_ (.X(_10898_),
    .B(_10897_),
    .A(_10892_));
 sg13g2_and2_1 _17701_ (.A(_10786_),
    .B(_10887_),
    .X(_10899_));
 sg13g2_buf_2 _17702_ (.A(_10899_),
    .X(_10900_));
 sg13g2_a22oi_1 _17703_ (.Y(_10901_),
    .B1(_10900_),
    .B2(\cpu.ex.r_8[14] ),
    .A2(_10829_),
    .A1(\cpu.ex.r_13[14] ));
 sg13g2_nor2b_1 _17704_ (.A(net1112),
    .B_N(net1111),
    .Y(_10902_));
 sg13g2_buf_1 _17705_ (.A(_10902_),
    .X(_10903_));
 sg13g2_mux2_1 _17706_ (.A0(_10278_),
    .A1(\cpu.ex.r_epc[14] ),
    .S(net884),
    .X(_10904_));
 sg13g2_nand3_1 _17707_ (.B(_10903_),
    .C(_10904_),
    .A(_10819_),
    .Y(_10905_));
 sg13g2_a22oi_1 _17708_ (.Y(_10906_),
    .B1(net684),
    .B2(\cpu.ex.r_12[14] ),
    .A2(_10862_),
    .A1(\cpu.ex.r_10[14] ));
 sg13g2_nor2_2 _17709_ (.A(_10825_),
    .B(_10894_),
    .Y(_10907_));
 sg13g2_nor2_1 _17710_ (.A(_00252_),
    .B(_10831_),
    .Y(_10908_));
 sg13g2_a21oi_1 _17711_ (.A1(\cpu.ex.r_14[14] ),
    .A2(_10907_),
    .Y(_10909_),
    .B1(_10908_));
 sg13g2_and4_1 _17712_ (.A(_10901_),
    .B(_10905_),
    .C(_10906_),
    .D(_10909_),
    .X(_10910_));
 sg13g2_nand4_1 _17713_ (.B(_10891_),
    .C(_10898_),
    .A(_10874_),
    .Y(_10911_),
    .D(_10910_));
 sg13g2_nor2b_1 _17714_ (.A(_10885_),
    .B_N(_10911_),
    .Y(_10912_));
 sg13g2_mux2_1 _17715_ (.A0(_10248_),
    .A1(_10912_),
    .S(_10794_),
    .X(_10913_));
 sg13g2_buf_8 _17716_ (.A(_10913_),
    .X(_10914_));
 sg13g2_inv_1 _17717_ (.Y(_10915_),
    .A(_00176_));
 sg13g2_nor2_1 _17718_ (.A(_08291_),
    .B(net620),
    .Y(_10916_));
 sg13g2_nor2b_1 _17719_ (.A(_10797_),
    .B_N(net1112),
    .Y(_10917_));
 sg13g2_buf_2 _17720_ (.A(_10917_),
    .X(_10918_));
 sg13g2_nand3_1 _17721_ (.B(\cpu.ex.r_9[15] ),
    .C(_10918_),
    .A(_10818_),
    .Y(_10919_));
 sg13g2_nand3_1 _17722_ (.B(\cpu.ex.r_mult[31] ),
    .C(_10849_),
    .A(_10801_),
    .Y(_10920_));
 sg13g2_a21oi_1 _17723_ (.A1(_10919_),
    .A2(_10920_),
    .Y(_10921_),
    .B1(_10807_));
 sg13g2_a221oi_1 _17724_ (.B2(\cpu.ex.r_8[15] ),
    .C1(_10921_),
    .B1(_10900_),
    .A1(\cpu.ex.r_epc[15] ),
    .Y(_10922_),
    .A2(net621));
 sg13g2_nor2_1 _17725_ (.A(_10847_),
    .B(_10825_),
    .Y(_10923_));
 sg13g2_mux2_1 _17726_ (.A0(\cpu.ex.r_lr[15] ),
    .A1(_10192_),
    .S(net882),
    .X(_10924_));
 sg13g2_a22oi_1 _17727_ (.Y(_10925_),
    .B1(_10924_),
    .B2(_10810_),
    .A2(_10923_),
    .A1(\cpu.ex.r_12[15] ));
 sg13g2_or2_1 _17728_ (.X(_10926_),
    .B(_10925_),
    .A(_10852_));
 sg13g2_a22oi_1 _17729_ (.Y(_10927_),
    .B1(_10907_),
    .B2(\cpu.ex.r_14[15] ),
    .A2(_10862_),
    .A1(\cpu.ex.r_10[15] ));
 sg13g2_nand2_1 _17730_ (.Y(_10928_),
    .A(\cpu.ex.r_13[15] ),
    .B(_10829_));
 sg13g2_or2_1 _17731_ (.X(_10929_),
    .B(_10831_),
    .A(_00253_));
 sg13g2_nor2_1 _17732_ (.A(_10808_),
    .B(net878),
    .Y(_10930_));
 sg13g2_mux2_1 _17733_ (.A0(_10200_),
    .A1(\cpu.ex.r_stmp[15] ),
    .S(net882),
    .X(_10931_));
 sg13g2_a22oi_1 _17734_ (.Y(_10932_),
    .B1(_10930_),
    .B2(_10931_),
    .A2(_10859_),
    .A1(\cpu.ex.r_11[15] ));
 sg13g2_and4_1 _17735_ (.A(_10927_),
    .B(_10928_),
    .C(_10929_),
    .D(_10932_),
    .X(_10933_));
 sg13g2_nand4_1 _17736_ (.B(_10922_),
    .C(_10926_),
    .A(_10874_),
    .Y(_10934_),
    .D(_10933_));
 sg13g2_nor2b_1 _17737_ (.A(_10916_),
    .B_N(_10934_),
    .Y(_10935_));
 sg13g2_mux2_1 _17738_ (.A0(_10915_),
    .A1(_10935_),
    .S(_10794_),
    .X(_10936_));
 sg13g2_buf_8 _17739_ (.A(_10936_),
    .X(_10937_));
 sg13g2_mux2_1 _17740_ (.A0(_10914_),
    .A1(net237),
    .S(\cpu.ex.c_mult_off[0] ),
    .X(_10938_));
 sg13g2_inv_1 _17741_ (.Y(_10939_),
    .A(_09260_));
 sg13g2_nand4_1 _17742_ (.B(_09258_),
    .C(_09259_),
    .A(_10939_),
    .Y(_10940_),
    .D(_09271_));
 sg13g2_buf_8 _17743_ (.A(_10874_),
    .X(_10941_));
 sg13g2_nand3_1 _17744_ (.B(\cpu.ex.r_8[13] ),
    .C(_10845_),
    .A(net763),
    .Y(_10942_));
 sg13g2_nand3_1 _17745_ (.B(_10401_),
    .C(_10850_),
    .A(_10886_),
    .Y(_10943_));
 sg13g2_a21o_1 _17746_ (.A2(_10943_),
    .A1(_10942_),
    .B1(net880),
    .X(_10944_));
 sg13g2_a22oi_1 _17747_ (.Y(_10945_),
    .B1(_10821_),
    .B2(\cpu.ex.r_lr[13] ),
    .A2(_10815_),
    .A1(_10394_));
 sg13g2_nand2b_1 _17748_ (.Y(_10946_),
    .B(net879),
    .A_N(_10945_));
 sg13g2_nor2_1 _17749_ (.A(_00251_),
    .B(_10831_),
    .Y(_10947_));
 sg13g2_a21oi_1 _17750_ (.A1(\cpu.ex.r_11[13] ),
    .A2(_10859_),
    .Y(_10948_),
    .B1(_10947_));
 sg13g2_a22oi_1 _17751_ (.Y(_10949_),
    .B1(_10862_),
    .B2(\cpu.ex.r_10[13] ),
    .A2(net621),
    .A1(\cpu.ex.r_epc[13] ));
 sg13g2_a22oi_1 _17752_ (.Y(_10950_),
    .B1(_10907_),
    .B2(\cpu.ex.r_14[13] ),
    .A2(net684),
    .A1(\cpu.ex.r_12[13] ));
 sg13g2_and4_1 _17753_ (.A(_10946_),
    .B(_10948_),
    .C(_10949_),
    .D(_10950_),
    .X(_10951_));
 sg13g2_and2_1 _17754_ (.A(_10835_),
    .B(_10849_),
    .X(_10952_));
 sg13g2_buf_1 _17755_ (.A(_10952_),
    .X(_10953_));
 sg13g2_nor2_1 _17756_ (.A(_10823_),
    .B(_10827_),
    .Y(_10954_));
 sg13g2_mux2_1 _17757_ (.A0(\cpu.ex.r_9[13] ),
    .A1(\cpu.ex.r_13[13] ),
    .S(_10802_),
    .X(_10955_));
 sg13g2_and2_1 _17758_ (.A(_10954_),
    .B(_10955_),
    .X(_10956_));
 sg13g2_a221oi_1 _17759_ (.B2(\cpu.ex.r_mult[29] ),
    .C1(_10956_),
    .B1(_10953_),
    .A1(\cpu.ex.r_stmp[13] ),
    .Y(_10957_),
    .A2(_10855_));
 sg13g2_nand4_1 _17760_ (.B(_10944_),
    .C(_10951_),
    .A(net620),
    .Y(_10958_),
    .D(_10957_));
 sg13g2_o21ai_1 _17761_ (.B1(_10958_),
    .Y(_10959_),
    .A1(_09440_),
    .A2(_10941_));
 sg13g2_mux2_1 _17762_ (.A0(_10392_),
    .A1(_10959_),
    .S(_10795_),
    .X(_10960_));
 sg13g2_buf_2 _17763_ (.A(_10960_),
    .X(_10961_));
 sg13g2_xnor2_1 _17764_ (.Y(_10962_),
    .A(\cpu.ex.r_mult_off[3] ),
    .B(_10881_));
 sg13g2_nand2_1 _17765_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(_09271_),
    .B(_10962_));
 sg13g2_o21ai_1 _17766_ (.B1(\cpu.ex.c_mult_off[3] ),
    .Y(_10963_),
    .A1(_10940_),
    .A2(_10961_));
 sg13g2_a221oi_1 _17767_ (.B2(_10938_),
    .C1(_10963_),
    .B1(_10884_),
    .A1(_10776_),
    .Y(_10964_),
    .A2(net193));
 sg13g2_nand2_1 _17768_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(_09271_),
    .B(_10883_));
 sg13g2_nor2_1 _17769_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(\cpu.ex.c_mult_off[2] ),
    .Y(_10965_));
 sg13g2_inv_1 _17770_ (.Y(_10966_),
    .A(_09258_));
 sg13g2_inv_2 _17771_ (.Y(_10967_),
    .A(_10874_));
 sg13g2_nor2_1 _17772_ (.A(_10823_),
    .B(net878),
    .Y(_10968_));
 sg13g2_nor2_1 _17773_ (.A(_10809_),
    .B(_10827_),
    .Y(_10969_));
 sg13g2_a22oi_1 _17774_ (.Y(_10970_),
    .B1(_10969_),
    .B2(\cpu.ex.r_lr[8] ),
    .A2(_10968_),
    .A1(\cpu.ex.r_10[8] ));
 sg13g2_and3_1 _17775_ (.X(_10971_),
    .A(\cpu.ex.r_stmp[8] ),
    .B(_10815_),
    .C(net761));
 sg13g2_a221oi_1 _17776_ (.B2(\cpu.ex.r_13[8] ),
    .C1(_10971_),
    .B1(_10829_),
    .A1(\cpu.ex.r_epc[8] ),
    .Y(_10972_),
    .A2(_10837_));
 sg13g2_o21ai_1 _17777_ (.B1(_10972_),
    .Y(_10973_),
    .A1(net765),
    .A2(_10970_));
 sg13g2_nor2b_1 _17778_ (.A(net884),
    .B_N(net1026),
    .Y(_10974_));
 sg13g2_nor2b_1 _17779_ (.A(net882),
    .B_N(net884),
    .Y(_10975_));
 sg13g2_a22oi_1 _17780_ (.Y(_10976_),
    .B1(_10975_),
    .B2(\cpu.ex.r_9[8] ),
    .A2(_10974_),
    .A1(\cpu.ex.r_12[8] ));
 sg13g2_nand2b_1 _17781_ (.Y(_10977_),
    .B(_10918_),
    .A_N(_10976_));
 sg13g2_and2_1 _17782_ (.A(net884),
    .B(net882),
    .X(_10978_));
 sg13g2_nor2_2 _17783_ (.A(_10806_),
    .B(_10812_),
    .Y(_10979_));
 sg13g2_a22oi_1 _17784_ (.Y(_10980_),
    .B1(_10979_),
    .B2(_10449_),
    .A2(_10978_),
    .A1(\cpu.ex.r_mult[24] ));
 sg13g2_nand2b_1 _17785_ (.Y(_10981_),
    .B(_10903_),
    .A_N(_10980_));
 sg13g2_a22oi_1 _17786_ (.Y(_10982_),
    .B1(_10900_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(_10859_),
    .A1(\cpu.ex.r_11[8] ));
 sg13g2_nor2_1 _17787_ (.A(_00246_),
    .B(_10831_),
    .Y(_10983_));
 sg13g2_a21oi_1 _17788_ (.A1(\cpu.ex.r_14[8] ),
    .A2(_10907_),
    .Y(_10984_),
    .B1(_10983_));
 sg13g2_nand4_1 _17789_ (.B(_10981_),
    .C(_10982_),
    .A(_10977_),
    .Y(_10985_),
    .D(_10984_));
 sg13g2_or3_1 _17790_ (.A(_10967_),
    .B(_10973_),
    .C(_10985_),
    .X(_10986_));
 sg13g2_o21ai_1 _17791_ (.B1(_10986_),
    .Y(_10987_),
    .A1(_09152_),
    .A2(net620));
 sg13g2_mux2_1 _17792_ (.A0(_10427_),
    .A1(_10987_),
    .S(_10795_),
    .X(_10988_));
 sg13g2_buf_2 _17793_ (.A(_10988_),
    .X(_10989_));
 sg13g2_nand3_1 _17794_ (.B(net1024),
    .C(net1026),
    .A(net1027),
    .Y(_10990_));
 sg13g2_buf_1 _17795_ (.A(_10990_),
    .X(_10991_));
 sg13g2_nor3_1 _17796_ (.A(net1027),
    .B(net1024),
    .C(net882),
    .Y(_10992_));
 sg13g2_nand2_1 _17797_ (.Y(_10993_),
    .A(\cpu.ex.r_lr[10] ),
    .B(_10992_));
 sg13g2_o21ai_1 _17798_ (.B1(_10993_),
    .Y(_10994_),
    .A1(_00248_),
    .A2(_10991_));
 sg13g2_nand2_1 _17799_ (.Y(_10995_),
    .A(net683),
    .B(_10994_));
 sg13g2_a22oi_1 _17800_ (.Y(_10996_),
    .B1(_10918_),
    .B2(\cpu.ex.r_8[10] ),
    .A2(_10903_),
    .A1(_10376_));
 sg13g2_nand2b_1 _17801_ (.Y(_10997_),
    .B(_10979_),
    .A_N(_10996_));
 sg13g2_a22oi_1 _17802_ (.Y(_10998_),
    .B1(_10842_),
    .B2(\cpu.ex.r_12[10] ),
    .A2(_10838_),
    .A1(\cpu.ex.r_epc[10] ));
 sg13g2_a22oi_1 _17803_ (.Y(_10999_),
    .B1(_10859_),
    .B2(\cpu.ex.r_11[10] ),
    .A2(_10855_),
    .A1(\cpu.ex.r_stmp[10] ));
 sg13g2_and2_1 _17804_ (.A(_10821_),
    .B(_10887_),
    .X(_11000_));
 sg13g2_a22oi_1 _17805_ (.Y(_11001_),
    .B1(_11000_),
    .B2(\cpu.ex.r_9[10] ),
    .A2(_10907_),
    .A1(\cpu.ex.r_14[10] ));
 sg13g2_and4_1 _17806_ (.A(_10997_),
    .B(_10998_),
    .C(_10999_),
    .D(_11001_),
    .X(_11002_));
 sg13g2_and2_1 _17807_ (.A(\cpu.ex.r_mult[26] ),
    .B(_10953_),
    .X(_11003_));
 sg13g2_a221oi_1 _17808_ (.B2(\cpu.ex.r_10[10] ),
    .C1(_11003_),
    .B1(_10862_),
    .A1(\cpu.ex.r_13[10] ),
    .Y(_11004_),
    .A2(_10829_));
 sg13g2_nand4_1 _17809_ (.B(_10995_),
    .C(_11002_),
    .A(net619),
    .Y(_11005_),
    .D(_11004_));
 sg13g2_o21ai_1 _17810_ (.B1(_11005_),
    .Y(_11006_),
    .A1(_10368_),
    .A2(net619));
 sg13g2_mux2_1 _17811_ (.A0(_10365_),
    .A1(_11006_),
    .S(net279),
    .X(_11007_));
 sg13g2_buf_1 _17812_ (.A(_11007_),
    .X(_11008_));
 sg13g2_nand2_2 _17813_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_09271_),
    .B(_10880_));
 sg13g2_a22oi_1 _17814_ (.Y(_11009_),
    .B1(_11008_),
    .B2(\cpu.ex.c_mult_off[1] ),
    .A2(_10989_),
    .A1(_10966_));
 sg13g2_nor2b_1 _17815_ (.A(\cpu.ex.c_mult_off[2] ),
    .B_N(\cpu.ex.c_mult_off[0] ),
    .Y(_11010_));
 sg13g2_inv_1 _17816_ (.Y(_11011_),
    .A(_10293_));
 sg13g2_inv_1 _17817_ (.Y(_11012_),
    .A(_10297_));
 sg13g2_mux4_1 _17818_ (.S0(net762),
    .A0(\cpu.ex.r_8[9] ),
    .A1(\cpu.ex.r_9[9] ),
    .A2(\cpu.ex.r_12[9] ),
    .A3(\cpu.ex.r_13[9] ),
    .S1(net885),
    .X(_11013_));
 sg13g2_and2_1 _17819_ (.A(_10918_),
    .B(_11013_),
    .X(_11014_));
 sg13g2_nand3_1 _17820_ (.B(net881),
    .C(net761),
    .A(\cpu.ex.r_mult[25] ),
    .Y(_11015_));
 sg13g2_nand3_1 _17821_ (.B(net879),
    .C(net881),
    .A(\cpu.ex.r_epc[9] ),
    .Y(_11016_));
 sg13g2_nand3_1 _17822_ (.B(net881),
    .C(net760),
    .A(\cpu.ex.r_11[9] ),
    .Y(_11017_));
 sg13g2_nand3_1 _17823_ (.B(net764),
    .C(net761),
    .A(\cpu.ex.r_stmp[9] ),
    .Y(_11018_));
 sg13g2_nand4_1 _17824_ (.B(_11016_),
    .C(_11017_),
    .A(_11015_),
    .Y(_11019_),
    .D(_11018_));
 sg13g2_or2_1 _17825_ (.X(_11020_),
    .B(_10991_),
    .A(_00247_));
 sg13g2_nand2_1 _17826_ (.Y(_11021_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_10992_));
 sg13g2_a21oi_1 _17827_ (.A1(_11020_),
    .A2(_11021_),
    .Y(_11022_),
    .B1(_10807_));
 sg13g2_mux2_1 _17828_ (.A0(\cpu.ex.r_10[9] ),
    .A1(\cpu.ex.r_14[9] ),
    .S(_10812_),
    .X(_11023_));
 sg13g2_a22oi_1 _17829_ (.Y(_11024_),
    .B1(_11023_),
    .B2(net759),
    .A2(net879),
    .A1(_10310_));
 sg13g2_nor2_1 _17830_ (.A(net878),
    .B(_11024_),
    .Y(_11025_));
 sg13g2_nor4_1 _17831_ (.A(_11014_),
    .B(_11019_),
    .C(_11022_),
    .D(_11025_),
    .Y(_11026_));
 sg13g2_mux2_1 _17832_ (.A0(_11012_),
    .A1(_11026_),
    .S(net620),
    .X(_11027_));
 sg13g2_inv_1 _17833_ (.Y(_11028_),
    .A(_11027_));
 sg13g2_mux2_1 _17834_ (.A0(_11011_),
    .A1(_11028_),
    .S(net279),
    .X(_11029_));
 sg13g2_buf_1 _17835_ (.A(_11029_),
    .X(_11030_));
 sg13g2_inv_1 _17836_ (.Y(_11031_),
    .A(_00273_));
 sg13g2_inv_2 _17837_ (.Y(_11032_),
    .A(_10693_));
 sg13g2_a22oi_1 _17838_ (.Y(_11033_),
    .B1(_10896_),
    .B2(\cpu.ex.r_9[11] ),
    .A2(_10895_),
    .A1(\cpu.ex.r_14[11] ));
 sg13g2_nor2_1 _17839_ (.A(_10823_),
    .B(_11033_),
    .Y(_11034_));
 sg13g2_nor2_1 _17840_ (.A(_00249_),
    .B(_10991_),
    .Y(_11035_));
 sg13g2_and2_1 _17841_ (.A(\cpu.ex.r_lr[11] ),
    .B(_10992_),
    .X(_11036_));
 sg13g2_o21ai_1 _17842_ (.B1(net683),
    .Y(_11037_),
    .A1(_11035_),
    .A2(_11036_));
 sg13g2_a22oi_1 _17843_ (.Y(_11038_),
    .B1(_10953_),
    .B2(\cpu.ex.r_mult[27] ),
    .A2(net621),
    .A1(\cpu.ex.r_epc[11] ));
 sg13g2_nand3_1 _17844_ (.B(net879),
    .C(net764),
    .A(_10697_),
    .Y(_11039_));
 sg13g2_nand3_1 _17845_ (.B(_11038_),
    .C(_11039_),
    .A(_11037_),
    .Y(_11040_));
 sg13g2_a22oi_1 _17846_ (.Y(_11041_),
    .B1(_10900_),
    .B2(\cpu.ex.r_8[11] ),
    .A2(_10859_),
    .A1(\cpu.ex.r_11[11] ));
 sg13g2_a22oi_1 _17847_ (.Y(_11042_),
    .B1(_10862_),
    .B2(\cpu.ex.r_10[11] ),
    .A2(_10855_),
    .A1(\cpu.ex.r_stmp[11] ));
 sg13g2_a22oi_1 _17848_ (.Y(_11043_),
    .B1(_10842_),
    .B2(\cpu.ex.r_12[11] ),
    .A2(_10829_),
    .A1(\cpu.ex.r_13[11] ));
 sg13g2_nand3_1 _17849_ (.B(_11042_),
    .C(_11043_),
    .A(_11041_),
    .Y(_11044_));
 sg13g2_nor4_1 _17850_ (.A(_10967_),
    .B(_11034_),
    .C(_11040_),
    .D(_11044_),
    .Y(_11045_));
 sg13g2_a21oi_1 _17851_ (.A1(_11032_),
    .A2(_10967_),
    .Y(_11046_),
    .B1(_11045_));
 sg13g2_mux2_1 _17852_ (.A0(_11031_),
    .A1(_11046_),
    .S(net279),
    .X(_11047_));
 sg13g2_buf_1 _17853_ (.A(_11047_),
    .X(_11048_));
 sg13g2_mux2_1 _17854_ (.A0(net215),
    .A1(_11048_),
    .S(\cpu.ex.c_mult_off[1] ),
    .X(_11049_));
 sg13g2_a22oi_1 _17855_ (.Y(_11050_),
    .B1(_11010_),
    .B2(_11049_),
    .A2(_11009_),
    .A1(_10965_));
 sg13g2_a22oi_1 _17856_ (.Y(_11051_),
    .B1(_10821_),
    .B2(\cpu.ex.r_9[6] ),
    .A2(net764),
    .A1(\cpu.ex.r_10[6] ));
 sg13g2_nand2b_1 _17857_ (.Y(_11052_),
    .B(net760),
    .A_N(_11051_));
 sg13g2_nand3_1 _17858_ (.B(\cpu.ex.r_8[6] ),
    .C(_10918_),
    .A(net763),
    .Y(_11053_));
 sg13g2_nand3_1 _17859_ (.B(\cpu.ex.r_stmp[6] ),
    .C(net761),
    .A(net880),
    .Y(_11054_));
 sg13g2_a21oi_1 _17860_ (.A1(_11053_),
    .A2(_11054_),
    .Y(_11055_),
    .B1(net683));
 sg13g2_nand3_1 _17861_ (.B(\cpu.ex.r_12[6] ),
    .C(_10840_),
    .A(_10807_),
    .Y(_11056_));
 sg13g2_nand3_1 _17862_ (.B(\cpu.ex.r_lr[6] ),
    .C(net879),
    .A(net683),
    .Y(_11057_));
 sg13g2_a21oi_1 _17863_ (.A1(_11056_),
    .A2(_11057_),
    .Y(_11058_),
    .B1(net880));
 sg13g2_nand3_1 _17864_ (.B(net881),
    .C(net761),
    .A(\cpu.ex.r_mult[22] ),
    .Y(_11059_));
 sg13g2_nand3_1 _17865_ (.B(_10863_),
    .C(_10816_),
    .A(_10354_),
    .Y(_11060_));
 sg13g2_nand2b_1 _17866_ (.Y(_11061_),
    .B(_10334_),
    .A_N(_10831_));
 sg13g2_nand3_1 _17867_ (.B(_11060_),
    .C(_11061_),
    .A(_11059_),
    .Y(_11062_));
 sg13g2_nand3_1 _17868_ (.B(_10840_),
    .C(_10821_),
    .A(\cpu.ex.r_13[6] ),
    .Y(_11063_));
 sg13g2_nand3_1 _17869_ (.B(_10840_),
    .C(_10816_),
    .A(\cpu.ex.r_14[6] ),
    .Y(_11064_));
 sg13g2_nand3_1 _17870_ (.B(_10863_),
    .C(net881),
    .A(\cpu.ex.r_epc[6] ),
    .Y(_11065_));
 sg13g2_nand3_1 _17871_ (.B(net881),
    .C(net760),
    .A(\cpu.ex.r_11[6] ),
    .Y(_11066_));
 sg13g2_nand4_1 _17872_ (.B(_11064_),
    .C(_11065_),
    .A(_11063_),
    .Y(_11067_),
    .D(_11066_));
 sg13g2_nor4_1 _17873_ (.A(_11055_),
    .B(_11058_),
    .C(_11062_),
    .D(_11067_),
    .Y(_11068_));
 sg13g2_nand3_1 _17874_ (.B(_11052_),
    .C(_11068_),
    .A(net620),
    .Y(_11069_));
 sg13g2_o21ai_1 _17875_ (.B1(_11069_),
    .Y(_11070_),
    .A1(_09150_),
    .A2(net619));
 sg13g2_buf_1 _17876_ (.A(_11070_),
    .X(_11071_));
 sg13g2_nor2_1 _17877_ (.A(net886),
    .B(net883),
    .Y(_11072_));
 sg13g2_mux2_1 _17878_ (.A0(\cpu.ex.r_stmp[7] ),
    .A1(\cpu.ex.r_14[7] ),
    .S(_10809_),
    .X(_11073_));
 sg13g2_a22oi_1 _17879_ (.Y(_11074_),
    .B1(_11073_),
    .B2(net880),
    .A2(_11072_),
    .A1(_10458_));
 sg13g2_nand2b_1 _17880_ (.Y(_11075_),
    .B(_10974_),
    .A_N(_11074_));
 sg13g2_and3_1 _17881_ (.X(_11076_),
    .A(net886),
    .B(net883),
    .C(\cpu.ex.r_11[7] ));
 sg13g2_a21o_1 _17882_ (.A2(_11072_),
    .A1(\cpu.ex.r_lr[7] ),
    .B1(_11076_),
    .X(_11077_));
 sg13g2_and3_1 _17883_ (.X(_11078_),
    .A(\cpu.ex.r_12[7] ),
    .B(_10786_),
    .C(_10840_));
 sg13g2_a221oi_1 _17884_ (.B2(_11077_),
    .C1(_11078_),
    .B1(_10975_),
    .A1(\cpu.ex.r_13[7] ),
    .Y(_11079_),
    .A2(_10829_));
 sg13g2_nor2_1 _17885_ (.A(_10813_),
    .B(net878),
    .Y(_11080_));
 sg13g2_mux2_1 _17886_ (.A0(_10460_),
    .A1(\cpu.ex.r_10[7] ),
    .S(net759),
    .X(_11081_));
 sg13g2_nor2_1 _17887_ (.A(_00245_),
    .B(_10831_),
    .Y(_11082_));
 sg13g2_a221oi_1 _17888_ (.B2(_11081_),
    .C1(_11082_),
    .B1(_11080_),
    .A1(\cpu.ex.r_epc[7] ),
    .Y(_11083_),
    .A2(_10838_));
 sg13g2_and3_1 _17889_ (.X(_11084_),
    .A(\cpu.ex.r_9[7] ),
    .B(_10821_),
    .C(net760));
 sg13g2_a221oi_1 _17890_ (.B2(\cpu.ex.r_8[7] ),
    .C1(_11084_),
    .B1(_10900_),
    .A1(\cpu.ex.r_mult[23] ),
    .Y(_11085_),
    .A2(_10953_));
 sg13g2_nand4_1 _17891_ (.B(_11079_),
    .C(_11083_),
    .A(_11075_),
    .Y(_11086_),
    .D(_11085_));
 sg13g2_inv_1 _17892_ (.Y(_11087_),
    .A(_09154_));
 sg13g2_nand2b_1 _17893_ (.Y(_11088_),
    .B(_11087_),
    .A_N(net620));
 sg13g2_o21ai_1 _17894_ (.B1(_11088_),
    .Y(_11089_),
    .A1(_10967_),
    .A2(_11086_));
 sg13g2_buf_1 _17895_ (.A(_11089_),
    .X(_11090_));
 sg13g2_mux4_1 _17896_ (.S0(net239),
    .A0(_10330_),
    .A1(_11071_),
    .A2(_10457_),
    .A3(_11090_),
    .S1(\cpu.ex.c_mult_off[0] ),
    .X(_11091_));
 sg13g2_nor2b_1 _17897_ (.A(_11091_),
    .B_N(_10884_),
    .Y(_11092_));
 sg13g2_nand2_1 _17898_ (.Y(_11093_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_10855_));
 sg13g2_a22oi_1 _17899_ (.Y(_11094_),
    .B1(_10859_),
    .B2(\cpu.ex.r_11[4] ),
    .A2(net621),
    .A1(\cpu.ex.r_epc[4] ));
 sg13g2_nand2_1 _17900_ (.Y(_11095_),
    .A(_11093_),
    .B(_11094_));
 sg13g2_nor2b_1 _17901_ (.A(net765),
    .B_N(net886),
    .Y(_11096_));
 sg13g2_nor2b_2 _17902_ (.A(net1027),
    .B_N(net882),
    .Y(_11097_));
 sg13g2_a221oi_1 _17903_ (.B2(_08285_),
    .C1(net683),
    .B1(_11097_),
    .A1(_10644_),
    .Y(_11098_),
    .A2(_11096_));
 sg13g2_a221oi_1 _17904_ (.B2(\cpu.ex.r_lr[4] ),
    .C1(_10807_),
    .B1(_10803_),
    .A1(\cpu.ex.r_mult[20] ),
    .Y(_11099_),
    .A2(_10800_));
 sg13g2_nor3_1 _17905_ (.A(net759),
    .B(_11098_),
    .C(_11099_),
    .Y(_11100_));
 sg13g2_a22oi_1 _17906_ (.Y(_11101_),
    .B1(_10821_),
    .B2(\cpu.ex.r_9[4] ),
    .A2(net764),
    .A1(\cpu.ex.r_10[4] ));
 sg13g2_nand2b_1 _17907_ (.Y(_11102_),
    .B(net760),
    .A_N(_11101_));
 sg13g2_a22oi_1 _17908_ (.Y(_11103_),
    .B1(_10979_),
    .B2(\cpu.ex.r_8[4] ),
    .A2(_10978_),
    .A1(\cpu.ex.r_13[4] ));
 sg13g2_nand2b_1 _17909_ (.Y(_11104_),
    .B(_10918_),
    .A_N(_11103_));
 sg13g2_nand2b_1 _17910_ (.Y(_11105_),
    .B(net762),
    .A_N(_00242_));
 sg13g2_nand2b_1 _17911_ (.Y(_11106_),
    .B(\cpu.ex.r_14[4] ),
    .A_N(net762));
 sg13g2_a21oi_1 _17912_ (.A1(_11105_),
    .A2(_11106_),
    .Y(_11107_),
    .B1(_10991_));
 sg13g2_a21oi_1 _17913_ (.A1(\cpu.ex.r_12[4] ),
    .A2(net684),
    .Y(_11108_),
    .B1(_11107_));
 sg13g2_nand3_1 _17914_ (.B(_11104_),
    .C(_11108_),
    .A(_11102_),
    .Y(_11109_));
 sg13g2_nor4_1 _17915_ (.A(_10967_),
    .B(_11095_),
    .C(_11100_),
    .D(_11109_),
    .Y(_11110_));
 sg13g2_a21oi_1 _17916_ (.A1(_09318_),
    .A2(_10967_),
    .Y(_11111_),
    .B1(_11110_));
 sg13g2_mux2_1 _17917_ (.A0(_08456_),
    .A1(_11111_),
    .S(net279),
    .X(_11112_));
 sg13g2_buf_1 _17918_ (.A(_11112_),
    .X(_11113_));
 sg13g2_and2_1 _17919_ (.A(_10776_),
    .B(_11113_),
    .X(_11114_));
 sg13g2_a22oi_1 _17920_ (.Y(_11115_),
    .B1(_10840_),
    .B2(\cpu.ex.r_13[5] ),
    .A2(net879),
    .A1(\cpu.ex.r_lr[5] ));
 sg13g2_nor2_1 _17921_ (.A(_10827_),
    .B(_11115_),
    .Y(_11116_));
 sg13g2_mux2_1 _17922_ (.A0(\cpu.ex.r_10[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(_10813_),
    .X(_11117_));
 sg13g2_a22oi_1 _17923_ (.Y(_11118_),
    .B1(_11117_),
    .B2(net759),
    .A2(net761),
    .A1(\cpu.ex.r_stmp[5] ));
 sg13g2_nor2_1 _17924_ (.A(net878),
    .B(_11118_),
    .Y(_11119_));
 sg13g2_nor2_1 _17925_ (.A(_00243_),
    .B(_10831_),
    .Y(_11120_));
 sg13g2_a21oi_1 _17926_ (.A1(\cpu.ex.r_8[5] ),
    .A2(_10900_),
    .Y(_11121_),
    .B1(_11120_));
 sg13g2_mux2_1 _17927_ (.A0(\cpu.ex.r_9[5] ),
    .A1(\cpu.ex.r_11[5] ),
    .S(net886),
    .X(_11122_));
 sg13g2_and2_1 _17928_ (.A(net1025),
    .B(net1024),
    .X(_11123_));
 sg13g2_buf_1 _17929_ (.A(_11123_),
    .X(_11124_));
 sg13g2_and2_1 _17930_ (.A(net763),
    .B(_11124_),
    .X(_11125_));
 sg13g2_a22oi_1 _17931_ (.Y(_11126_),
    .B1(_11122_),
    .B2(_11125_),
    .A2(_10953_),
    .A1(\cpu.ex.r_mult[21] ));
 sg13g2_nand3_1 _17932_ (.B(net879),
    .C(net764),
    .A(_10622_),
    .Y(_11127_));
 sg13g2_a22oi_1 _17933_ (.Y(_11128_),
    .B1(net684),
    .B2(\cpu.ex.r_12[5] ),
    .A2(net621),
    .A1(\cpu.ex.r_epc[5] ));
 sg13g2_nand4_1 _17934_ (.B(_11126_),
    .C(_11127_),
    .A(_11121_),
    .Y(_11129_),
    .D(_11128_));
 sg13g2_or4_1 _17935_ (.A(_10967_),
    .B(_11116_),
    .C(_11119_),
    .D(_11129_),
    .X(_11130_));
 sg13g2_o21ai_1 _17936_ (.B1(_11130_),
    .Y(_11131_),
    .A1(_09907_),
    .A2(net619));
 sg13g2_mux2_1 _17937_ (.A0(_10629_),
    .A1(_11131_),
    .S(net279),
    .X(_11132_));
 sg13g2_buf_1 _17938_ (.A(_11132_),
    .X(_11133_));
 sg13g2_nor2_1 _17939_ (.A(_10940_),
    .B(_11133_),
    .Y(_11134_));
 sg13g2_nor4_1 _17940_ (.A(\cpu.ex.c_mult_off[3] ),
    .B(_11092_),
    .C(_11114_),
    .D(_11134_),
    .Y(_11135_));
 sg13g2_a22oi_1 _17941_ (.Y(_11136_),
    .B1(_10918_),
    .B2(\cpu.ex.r_8[2] ),
    .A2(_10903_),
    .A1(_10524_));
 sg13g2_nand2_1 _17942_ (.Y(_11137_),
    .A(\cpu.ex.r_9[2] ),
    .B(_10954_));
 sg13g2_o21ai_1 _17943_ (.B1(_11137_),
    .Y(_11138_),
    .A1(net683),
    .A2(_11136_));
 sg13g2_mux2_1 _17944_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net882),
    .X(_11139_));
 sg13g2_a22oi_1 _17945_ (.Y(_11140_),
    .B1(_11139_),
    .B2(net759),
    .A2(net761),
    .A1(\cpu.ex.r_stmp[2] ));
 sg13g2_nand2b_1 _17946_ (.Y(_11141_),
    .B(net764),
    .A_N(_11140_));
 sg13g2_mux2_1 _17947_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(net1113),
    .S(net885),
    .X(_11142_));
 sg13g2_a22oi_1 _17948_ (.Y(_11143_),
    .B1(_10969_),
    .B2(_11142_),
    .A2(net684),
    .A1(\cpu.ex.r_12[2] ));
 sg13g2_nor2_1 _17949_ (.A(net884),
    .B(net1024),
    .Y(_11144_));
 sg13g2_a22oi_1 _17950_ (.Y(_11145_),
    .B1(_11144_),
    .B2(net1131),
    .A2(_11124_),
    .A1(\cpu.ex.r_13[2] ));
 sg13g2_nand2b_1 _17951_ (.Y(_11146_),
    .B(_11097_),
    .A_N(_11145_));
 sg13g2_inv_1 _17952_ (.Y(_11147_),
    .A(_00240_));
 sg13g2_a22oi_1 _17953_ (.Y(_11148_),
    .B1(_10840_),
    .B2(_11147_),
    .A2(_10783_),
    .A1(\cpu.ex.r_epc[2] ));
 sg13g2_a22oi_1 _17954_ (.Y(_11149_),
    .B1(net760),
    .B2(\cpu.ex.r_11[2] ),
    .A2(_10849_),
    .A1(\cpu.ex.r_mult[18] ));
 sg13g2_nand2_1 _17955_ (.Y(_11150_),
    .A(net1025),
    .B(net1111));
 sg13g2_a21o_1 _17956_ (.A2(_11149_),
    .A1(_11148_),
    .B1(_11150_),
    .X(_11151_));
 sg13g2_nand4_1 _17957_ (.B(_11143_),
    .C(_11146_),
    .A(_11141_),
    .Y(_11152_),
    .D(_11151_));
 sg13g2_a21oi_1 _17958_ (.A1(_10819_),
    .A2(_11138_),
    .Y(_11153_),
    .B1(_11152_));
 sg13g2_nor2_1 _17959_ (.A(_09140_),
    .B(_10875_),
    .Y(_11154_));
 sg13g2_a21oi_1 _17960_ (.A1(_10941_),
    .A2(_11153_),
    .Y(_11155_),
    .B1(_11154_));
 sg13g2_mux2_1 _17961_ (.A0(_10541_),
    .A1(_11155_),
    .S(net279),
    .X(_11156_));
 sg13g2_buf_2 _17962_ (.A(_11156_),
    .X(_11157_));
 sg13g2_a221oi_1 _17963_ (.B2(_08400_),
    .C1(_08330_),
    .B1(_08398_),
    .A1(_08343_),
    .Y(_11158_),
    .A2(_08362_));
 sg13g2_buf_1 _17964_ (.A(_11158_),
    .X(_11159_));
 sg13g2_nor2_2 _17965_ (.A(_09087_),
    .B(_09135_),
    .Y(_11160_));
 sg13g2_nand2b_1 _17966_ (.Y(_11161_),
    .B(_10791_),
    .A_N(_08286_));
 sg13g2_a21o_1 _17967_ (.A2(_11160_),
    .A1(_11159_),
    .B1(_11161_),
    .X(_11162_));
 sg13g2_nor2_1 _17968_ (.A(net1134),
    .B(_10874_),
    .Y(_11163_));
 sg13g2_inv_1 _17969_ (.Y(_11164_),
    .A(_10561_));
 sg13g2_nand2b_1 _17970_ (.Y(_11165_),
    .B(net1025),
    .A_N(_10782_));
 sg13g2_nand3b_1 _17971_ (.B(_10798_),
    .C(\cpu.ex.r_stmp[0] ),
    .Y(_11166_),
    .A_N(net1025));
 sg13g2_o21ai_1 _17972_ (.B1(_11166_),
    .Y(_11167_),
    .A1(_11164_),
    .A2(_11165_));
 sg13g2_mux2_1 _17973_ (.A0(\cpu.ex.r_8[0] ),
    .A1(\cpu.ex.r_10[0] ),
    .S(net1111),
    .X(_11168_));
 sg13g2_and3_1 _17974_ (.X(_11169_),
    .A(_10818_),
    .B(_10845_),
    .C(_11168_));
 sg13g2_a221oi_1 _17975_ (.B2(_11167_),
    .C1(_11169_),
    .B1(_10903_),
    .A1(\cpu.ex.r_11[0] ),
    .Y(_11170_),
    .A2(_10859_));
 sg13g2_inv_1 _17976_ (.Y(_11171_),
    .A(\cpu.ex.r_14[0] ));
 sg13g2_nand3b_1 _17977_ (.B(\cpu.ex.r_13[0] ),
    .C(net1025),
    .Y(_11172_),
    .A_N(_10797_));
 sg13g2_o21ai_1 _17978_ (.B1(_11172_),
    .Y(_11173_),
    .A1(_11171_),
    .A2(net878));
 sg13g2_nand2_1 _17979_ (.Y(_11174_),
    .A(net1026),
    .B(\cpu.ex.r_12[0] ));
 sg13g2_nand3b_1 _17980_ (.B(\cpu.ex.r_9[0] ),
    .C(_10805_),
    .Y(_11175_),
    .A_N(net1026));
 sg13g2_o21ai_1 _17981_ (.B1(_11175_),
    .Y(_11176_),
    .A1(net884),
    .A2(_11174_));
 sg13g2_a22oi_1 _17982_ (.Y(_11177_),
    .B1(_11176_),
    .B2(_10918_),
    .A2(_11173_),
    .A1(_10840_));
 sg13g2_nand2_1 _17983_ (.Y(_11178_),
    .A(net1024),
    .B(\cpu.ex.r_15[0] ));
 sg13g2_nand2b_1 _17984_ (.Y(_11179_),
    .B(\cpu.ex.r_mult[16] ),
    .A_N(_10808_));
 sg13g2_a21oi_1 _17985_ (.A1(_11178_),
    .A2(_11179_),
    .Y(_11180_),
    .B1(_11150_));
 sg13g2_nor4_1 _17986_ (.A(_09134_),
    .B(_10806_),
    .C(net1027),
    .D(net1024),
    .Y(_11181_));
 sg13g2_o21ai_1 _17987_ (.B1(net885),
    .Y(_11182_),
    .A1(_11180_),
    .A2(_11181_));
 sg13g2_and4_1 _17988_ (.A(_10874_),
    .B(_11170_),
    .C(_11177_),
    .D(_11182_),
    .X(_11183_));
 sg13g2_buf_1 _17989_ (.A(_11183_),
    .X(_11184_));
 sg13g2_nor4_1 _17990_ (.A(_08330_),
    .B(_10789_),
    .C(_11163_),
    .D(_11184_),
    .Y(_11185_));
 sg13g2_nor3_1 _17991_ (.A(_10791_),
    .B(_11163_),
    .C(_11184_),
    .Y(_11186_));
 sg13g2_a21oi_1 _17992_ (.A1(net459),
    .A2(_11185_),
    .Y(_11187_),
    .B1(_11186_));
 sg13g2_nand2_1 _17993_ (.Y(_11188_),
    .A(_11162_),
    .B(_11187_));
 sg13g2_buf_2 _17994_ (.A(_11188_),
    .X(_11189_));
 sg13g2_mux2_1 _17995_ (.A0(_11157_),
    .A1(_11189_),
    .S(_10966_),
    .X(_11190_));
 sg13g2_nor2_1 _17996_ (.A(_09143_),
    .B(net619),
    .Y(_11191_));
 sg13g2_and3_1 _17997_ (.X(_11192_),
    .A(net762),
    .B(net883),
    .C(\cpu.ex.r_13[1] ));
 sg13g2_a21o_1 _17998_ (.A2(_11144_),
    .A1(_10586_),
    .B1(_11192_),
    .X(_11193_));
 sg13g2_or2_1 _17999_ (.X(_11194_),
    .B(net885),
    .A(net886));
 sg13g2_nand3b_1 _18000_ (.B(net765),
    .C(net880),
    .Y(_11195_),
    .A_N(_00239_));
 sg13g2_o21ai_1 _18001_ (.B1(_11195_),
    .Y(_11196_),
    .A1(_10572_),
    .A2(_11194_));
 sg13g2_a22oi_1 _18002_ (.Y(_11197_),
    .B1(_11196_),
    .B2(_11124_),
    .A2(_11193_),
    .A1(_11097_));
 sg13g2_nand2_1 _18003_ (.Y(_11198_),
    .A(net762),
    .B(\cpu.ex.r_11[1] ));
 sg13g2_nand2b_1 _18004_ (.Y(_11199_),
    .B(\cpu.ex.r_10[1] ),
    .A_N(net762));
 sg13g2_nand3b_1 _18005_ (.B(net883),
    .C(net886),
    .Y(_11200_),
    .A_N(net885));
 sg13g2_a21oi_1 _18006_ (.A1(_11198_),
    .A2(_11199_),
    .Y(_11201_),
    .B1(_11200_));
 sg13g2_a221oi_1 _18007_ (.B2(\cpu.ex.r_8[1] ),
    .C1(_11201_),
    .B1(_10900_),
    .A1(\cpu.ex.r_12[1] ),
    .Y(_11202_),
    .A2(net684));
 sg13g2_nand2_1 _18008_ (.Y(_11203_),
    .A(net765),
    .B(\cpu.ex.r_stmp[1] ));
 sg13g2_nand2b_1 _18009_ (.Y(_11204_),
    .B(_10589_),
    .A_N(net885));
 sg13g2_nand3_1 _18010_ (.B(_11203_),
    .C(_11204_),
    .A(_10823_),
    .Y(_11205_));
 sg13g2_nand2_1 _18011_ (.Y(_11206_),
    .A(net765),
    .B(\cpu.ex.r_14[1] ));
 sg13g2_a21oi_1 _18012_ (.A1(net759),
    .A2(_11206_),
    .Y(_11207_),
    .B1(net878));
 sg13g2_mux4_1 _18013_ (.S0(net886),
    .A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.r_epc[1] ),
    .A2(\cpu.ex.mmu_read[1] ),
    .A3(\cpu.ex.r_mult[17] ),
    .S1(net765),
    .X(_11208_));
 sg13g2_a22oi_1 _18014_ (.Y(_11209_),
    .B1(_11208_),
    .B2(_10810_),
    .A2(_11207_),
    .A1(_11205_));
 sg13g2_and4_1 _18015_ (.A(net620),
    .B(_11197_),
    .C(_11202_),
    .D(_11209_),
    .X(_11210_));
 sg13g2_buf_1 _18016_ (.A(_11210_),
    .X(_11211_));
 sg13g2_or2_1 _18017_ (.X(_11212_),
    .B(_11211_),
    .A(_11191_));
 sg13g2_inv_1 _18018_ (.Y(_11213_),
    .A(\cpu.ex.r_11[3] ));
 sg13g2_nor2_1 _18019_ (.A(_11213_),
    .B(_11200_),
    .Y(_11214_));
 sg13g2_inv_1 _18020_ (.Y(_11215_),
    .A(_10505_));
 sg13g2_nor4_1 _18021_ (.A(net880),
    .B(net759),
    .C(net763),
    .D(_11215_),
    .Y(_11216_));
 sg13g2_o21ai_1 _18022_ (.B1(net683),
    .Y(_11217_),
    .A1(_11214_),
    .A2(_11216_));
 sg13g2_a22oi_1 _18023_ (.Y(_11218_),
    .B1(_10930_),
    .B2(\cpu.ex.r_stmp[3] ),
    .A2(_10954_),
    .A1(\cpu.ex.r_13[3] ));
 sg13g2_nand2b_1 _18024_ (.Y(_11219_),
    .B(net765),
    .A_N(_11218_));
 sg13g2_nor2_1 _18025_ (.A(net763),
    .B(_11150_),
    .Y(_11220_));
 sg13g2_mux2_1 _18026_ (.A0(_10496_),
    .A1(\cpu.ex.r_mult[19] ),
    .S(_10823_),
    .X(_11221_));
 sg13g2_a22oi_1 _18027_ (.Y(_11222_),
    .B1(_11220_),
    .B2(_11221_),
    .A2(net684),
    .A1(\cpu.ex.r_12[3] ));
 sg13g2_mux2_1 _18028_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(\cpu.ex.r_9[3] ),
    .S(net883),
    .X(_11223_));
 sg13g2_mux2_1 _18029_ (.A0(_10492_),
    .A1(\cpu.ex.r_10[3] ),
    .S(net883),
    .X(_11224_));
 sg13g2_a22oi_1 _18030_ (.Y(_11225_),
    .B1(_11224_),
    .B2(_11080_),
    .A2(_11223_),
    .A1(_10896_));
 sg13g2_a22oi_1 _18031_ (.Y(_11226_),
    .B1(_10803_),
    .B2(\cpu.ex.r_8[3] ),
    .A2(_10800_),
    .A1(\cpu.ex.r_14[3] ));
 sg13g2_nand2b_1 _18032_ (.Y(_11227_),
    .B(_10845_),
    .A_N(_11226_));
 sg13g2_nor2b_1 _18033_ (.A(net885),
    .B_N(\cpu.ex.r_epc[3] ),
    .Y(_11228_));
 sg13g2_nor2b_1 _18034_ (.A(net762),
    .B_N(net1135),
    .Y(_11229_));
 sg13g2_a22oi_1 _18035_ (.Y(_11230_),
    .B1(_11229_),
    .B2(_11097_),
    .A2(_11228_),
    .A1(net881));
 sg13g2_or2_1 _18036_ (.X(_11231_),
    .B(_11230_),
    .A(net759));
 sg13g2_and4_1 _18037_ (.A(_11222_),
    .B(_11225_),
    .C(_11227_),
    .D(_11231_),
    .X(_11232_));
 sg13g2_nand4_1 _18038_ (.B(_11217_),
    .C(_11219_),
    .A(net619),
    .Y(_11233_),
    .D(_11232_));
 sg13g2_o21ai_1 _18039_ (.B1(_11233_),
    .Y(_11234_),
    .A1(_09163_),
    .A2(net619));
 sg13g2_buf_1 _18040_ (.A(_11234_),
    .X(_11235_));
 sg13g2_mux4_1 _18041_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(_10596_),
    .A1(_10486_),
    .A2(_11212_),
    .A3(_11235_),
    .S1(net239),
    .X(_11236_));
 sg13g2_nor2b_1 _18042_ (.A(_11236_),
    .B_N(_11010_),
    .Y(_11237_));
 sg13g2_a21oi_1 _18043_ (.A1(_10965_),
    .A2(_11190_),
    .Y(_11238_),
    .B1(_11237_));
 sg13g2_a22oi_1 _18044_ (.Y(_11239_),
    .B1(_11135_),
    .B2(_11238_),
    .A2(_11050_),
    .A1(_10964_));
 sg13g2_buf_1 _18045_ (.A(_11239_),
    .X(_11240_));
 sg13g2_a21o_1 _18046_ (.A2(_10595_),
    .A1(_10594_),
    .B1(_10599_),
    .X(_11241_));
 sg13g2_buf_1 _18047_ (.A(_11241_),
    .X(_11242_));
 sg13g2_buf_8 _18048_ (.A(_11242_),
    .X(_11243_));
 sg13g2_buf_1 _18049_ (.A(_00293_),
    .X(_11244_));
 sg13g2_nor2_1 _18050_ (.A(_11244_),
    .B(net505),
    .Y(_11245_));
 sg13g2_nand2_1 _18051_ (.Y(_11246_),
    .A(net236),
    .B(_11245_));
 sg13g2_and4_1 _18052_ (.A(_10519_),
    .B(_10523_),
    .C(_10527_),
    .D(_10536_),
    .X(_11247_));
 sg13g2_nand2_1 _18053_ (.Y(_11248_),
    .A(_09141_),
    .B(_10238_));
 sg13g2_o21ai_1 _18054_ (.B1(_11248_),
    .Y(_11249_),
    .A1(_10172_),
    .A2(_11247_));
 sg13g2_inv_1 _18055_ (.Y(_11250_),
    .A(_10539_));
 sg13g2_a221oi_1 _18056_ (.B2(_11250_),
    .C1(_10543_),
    .B1(_11249_),
    .A1(net1029),
    .Y(_11251_),
    .A2(_10541_));
 sg13g2_buf_2 _18057_ (.A(_11251_),
    .X(_11252_));
 sg13g2_buf_1 _18058_ (.A(_11252_),
    .X(_11253_));
 sg13g2_buf_1 _18059_ (.A(_00292_),
    .X(_11254_));
 sg13g2_nor2_1 _18060_ (.A(_11254_),
    .B(net505),
    .Y(_11255_));
 sg13g2_nand2_1 _18061_ (.Y(_11256_),
    .A(_11253_),
    .B(_11255_));
 sg13g2_nand3_1 _18062_ (.B(_11246_),
    .C(_11256_),
    .A(_10566_),
    .Y(_11257_));
 sg13g2_buf_2 _18063_ (.A(_00288_),
    .X(_11258_));
 sg13g2_buf_1 _18064_ (.A(_00289_),
    .X(_11259_));
 sg13g2_and3_1 _18065_ (.X(_11260_),
    .A(_11258_),
    .B(_11259_),
    .C(net286));
 sg13g2_buf_1 _18066_ (.A(_11259_),
    .X(_11261_));
 sg13g2_xnor2_1 _18067_ (.Y(_11262_),
    .A(net1023),
    .B(_10633_));
 sg13g2_nor2_1 _18068_ (.A(_11258_),
    .B(net573),
    .Y(_11263_));
 sg13g2_inv_1 _18069_ (.Y(_11264_),
    .A(_11263_));
 sg13g2_nor2_1 _18070_ (.A(net286),
    .B(_11264_),
    .Y(_11265_));
 sg13g2_nor2_2 _18071_ (.A(_11259_),
    .B(net573),
    .Y(_11266_));
 sg13g2_nand4_1 _18072_ (.B(_10332_),
    .C(_10362_),
    .A(_11258_),
    .Y(_11267_),
    .D(_11266_));
 sg13g2_and2_1 _18073_ (.A(net573),
    .B(_10631_),
    .X(_11268_));
 sg13g2_nand4_1 _18074_ (.B(_10332_),
    .C(_10362_),
    .A(_10628_),
    .Y(_11269_),
    .D(_11268_));
 sg13g2_o21ai_1 _18075_ (.B1(_11269_),
    .Y(_11270_),
    .A1(_10633_),
    .A2(_11267_));
 sg13g2_a221oi_1 _18076_ (.B2(_11265_),
    .C1(_11270_),
    .B1(_11262_),
    .A1(net241),
    .Y(_11271_),
    .A2(_11260_));
 sg13g2_buf_2 _18077_ (.A(_00290_),
    .X(_11272_));
 sg13g2_nor2_2 _18078_ (.A(_11272_),
    .B(net573),
    .Y(_11273_));
 sg13g2_mux2_1 _18079_ (.A0(_11273_),
    .A1(_11272_),
    .S(net358),
    .X(_11274_));
 sg13g2_buf_1 _18080_ (.A(_00287_),
    .X(_11275_));
 sg13g2_a22oi_1 _18081_ (.Y(_11276_),
    .B1(_11274_),
    .B2(net1110),
    .A2(net358),
    .A1(net505));
 sg13g2_nor2_1 _18082_ (.A(net1110),
    .B(net505),
    .Y(_11277_));
 sg13g2_xnor2_1 _18083_ (.Y(_11278_),
    .A(_11272_),
    .B(net358));
 sg13g2_nand2_1 _18084_ (.Y(_11279_),
    .A(_11277_),
    .B(_11278_));
 sg13g2_nand2b_1 _18085_ (.Y(_11280_),
    .B(net1029),
    .A_N(_10457_));
 sg13g2_o21ai_1 _18086_ (.B1(_11280_),
    .Y(_11281_),
    .A1(net887),
    .A2(_10480_));
 sg13g2_buf_2 _18087_ (.A(_11281_),
    .X(_11282_));
 sg13g2_mux2_1 _18088_ (.A0(_11276_),
    .A1(_11279_),
    .S(_11282_),
    .X(_11283_));
 sg13g2_nand2b_1 _18089_ (.Y(_11284_),
    .B(_10742_),
    .A_N(_11254_));
 sg13g2_buf_1 _18090_ (.A(_11284_),
    .X(_11285_));
 sg13g2_nor2_1 _18091_ (.A(_10546_),
    .B(_11285_),
    .Y(_11286_));
 sg13g2_or2_1 _18092_ (.X(_11287_),
    .B(_11245_),
    .A(_11242_));
 sg13g2_nor2_1 _18093_ (.A(_11286_),
    .B(_11287_),
    .Y(_11288_));
 sg13g2_nor2_1 _18094_ (.A(_10487_),
    .B(_10514_),
    .Y(_11289_));
 sg13g2_buf_2 _18095_ (.A(_11289_),
    .X(_11290_));
 sg13g2_nor2_1 _18096_ (.A(_00291_),
    .B(net505),
    .Y(_11291_));
 sg13g2_buf_1 _18097_ (.A(_11291_),
    .X(_11292_));
 sg13g2_nand2_1 _18098_ (.Y(_11293_),
    .A(net283),
    .B(_11285_));
 sg13g2_o21ai_1 _18099_ (.B1(_11293_),
    .Y(_11294_),
    .A1(_11290_),
    .A2(net403));
 sg13g2_nor4_1 _18100_ (.A(_11271_),
    .B(_11283_),
    .C(_11288_),
    .D(_11294_),
    .Y(_11295_));
 sg13g2_o21ai_1 _18101_ (.B1(_11295_),
    .Y(_11296_),
    .A1(net118),
    .A2(_11257_));
 sg13g2_buf_1 _18102_ (.A(_11296_),
    .X(_11297_));
 sg13g2_nor2_1 _18103_ (.A(net897),
    .B(_10661_),
    .Y(_11298_));
 sg13g2_nor3_2 _18104_ (.A(net887),
    .B(_10663_),
    .C(_10685_),
    .Y(_11299_));
 sg13g2_nor2_2 _18105_ (.A(_11298_),
    .B(_11299_),
    .Y(_11300_));
 sg13g2_inv_1 _18106_ (.Y(_11301_),
    .A(_11272_));
 sg13g2_nand3_1 _18107_ (.B(net241),
    .C(net358),
    .A(_11301_),
    .Y(_11302_));
 sg13g2_a22oi_1 _18108_ (.Y(_11303_),
    .B1(net358),
    .B2(_11301_),
    .A2(_10631_),
    .A1(_10628_));
 sg13g2_or2_1 _18109_ (.X(_11304_),
    .B(_11303_),
    .A(net1023));
 sg13g2_nand2_1 _18110_ (.Y(_11305_),
    .A(_10742_),
    .B(net286));
 sg13g2_and2_1 _18111_ (.A(_11275_),
    .B(_11282_),
    .X(_11306_));
 sg13g2_a221oi_1 _18112_ (.B2(_11264_),
    .C1(_11306_),
    .B1(_11305_),
    .A1(_11302_),
    .Y(_11307_),
    .A2(_11304_));
 sg13g2_nor3_1 _18113_ (.A(_11275_),
    .B(net505),
    .C(_11282_),
    .Y(_11308_));
 sg13g2_nand2_1 _18114_ (.Y(_11309_),
    .A(_10332_),
    .B(_10362_));
 sg13g2_nor3_1 _18115_ (.A(_11309_),
    .B(_11264_),
    .C(_11306_),
    .Y(_11310_));
 sg13g2_or3_1 _18116_ (.A(_11307_),
    .B(_11308_),
    .C(_11310_),
    .X(_11311_));
 sg13g2_buf_1 _18117_ (.A(_11311_),
    .X(_11312_));
 sg13g2_or2_1 _18118_ (.X(_11313_),
    .B(_10514_),
    .A(_10487_));
 sg13g2_buf_2 _18119_ (.A(_11313_),
    .X(_11314_));
 sg13g2_inv_1 _18120_ (.Y(_11315_),
    .A(_00291_));
 sg13g2_buf_1 _18121_ (.A(_10742_),
    .X(_11316_));
 sg13g2_nand2_1 _18122_ (.Y(_11317_),
    .A(_11315_),
    .B(net500));
 sg13g2_nor4_2 _18123_ (.A(_11314_),
    .B(_11271_),
    .C(_11283_),
    .Y(_11318_),
    .D(_11317_));
 sg13g2_nor4_1 _18124_ (.A(_11300_),
    .B(_10773_),
    .C(_11312_),
    .D(_11318_),
    .Y(_11319_));
 sg13g2_a22oi_1 _18125_ (.Y(_11320_),
    .B1(_11297_),
    .B2(_11319_),
    .A2(_10774_),
    .A1(net194));
 sg13g2_buf_1 _18126_ (.A(_00281_),
    .X(_11321_));
 sg13g2_buf_1 _18127_ (.A(_00282_),
    .X(_11322_));
 sg13g2_nand2b_1 _18128_ (.Y(_11323_),
    .B(net500),
    .A_N(_11322_));
 sg13g2_buf_1 _18129_ (.A(_11323_),
    .X(_11324_));
 sg13g2_nor2_1 _18130_ (.A(_11321_),
    .B(_11324_),
    .Y(_11325_));
 sg13g2_nor2_1 _18131_ (.A(_11321_),
    .B(net450),
    .Y(_11326_));
 sg13g2_nand2b_1 _18132_ (.Y(_11327_),
    .B(net887),
    .A_N(_10392_));
 sg13g2_o21ai_1 _18133_ (.B1(_11327_),
    .Y(_11328_),
    .A1(net887),
    .A2(_10423_));
 sg13g2_buf_2 _18134_ (.A(_11328_),
    .X(_11329_));
 sg13g2_nor4_1 _18135_ (.A(_10425_),
    .B(_10773_),
    .C(_11312_),
    .D(_11318_),
    .Y(_11330_));
 sg13g2_nor2_1 _18136_ (.A(net217),
    .B(_11300_),
    .Y(_11331_));
 sg13g2_a221oi_1 _18137_ (.B2(_11330_),
    .C1(_11331_),
    .B1(_11297_),
    .A1(_11329_),
    .Y(_11332_),
    .A2(_10774_));
 sg13g2_a22oi_1 _18138_ (.Y(_11333_),
    .B1(_11326_),
    .B2(_11332_),
    .A2(_11325_),
    .A1(_11320_));
 sg13g2_buf_2 _18139_ (.A(_11333_),
    .X(_11334_));
 sg13g2_nor2_1 _18140_ (.A(_11312_),
    .B(_11318_),
    .Y(_11335_));
 sg13g2_buf_1 _18141_ (.A(_11335_),
    .X(_11336_));
 sg13g2_nor2_1 _18142_ (.A(_11322_),
    .B(net450),
    .Y(_11337_));
 sg13g2_nor2_1 _18143_ (.A(_10773_),
    .B(_11337_),
    .Y(_11338_));
 sg13g2_nand3_1 _18144_ (.B(net97),
    .C(_11338_),
    .A(_11297_),
    .Y(_11339_));
 sg13g2_o21ai_1 _18145_ (.B1(_10774_),
    .Y(_11340_),
    .A1(_10689_),
    .A2(_11324_));
 sg13g2_a22oi_1 _18146_ (.Y(_11341_),
    .B1(_11324_),
    .B2(_10689_),
    .A2(_11319_),
    .A1(_11297_));
 sg13g2_nand4_1 _18147_ (.B(_11339_),
    .C(_11340_),
    .A(net217),
    .Y(_11342_),
    .D(_11341_));
 sg13g2_buf_8 _18148_ (.A(_11342_),
    .X(_11343_));
 sg13g2_buf_1 _18149_ (.A(_00279_),
    .X(_11344_));
 sg13g2_or3_1 _18150_ (.A(net1109),
    .B(net450),
    .C(net168),
    .X(_11345_));
 sg13g2_inv_2 _18151_ (.Y(_11346_),
    .A(_00280_));
 sg13g2_nand2_1 _18152_ (.Y(_11347_),
    .A(_11346_),
    .B(net500));
 sg13g2_or2_1 _18153_ (.X(_11348_),
    .B(_11347_),
    .A(_10247_));
 sg13g2_a22oi_1 _18154_ (.Y(_11349_),
    .B1(_11345_),
    .B2(_11348_),
    .A2(_11343_),
    .A1(_11334_));
 sg13g2_buf_1 _18155_ (.A(_11349_),
    .X(_11350_));
 sg13g2_nand3b_1 _18156_ (.B(_11346_),
    .C(net500),
    .Y(_11351_),
    .A_N(net1109));
 sg13g2_buf_1 _18157_ (.A(_11351_),
    .X(_11352_));
 sg13g2_a21oi_2 _18158_ (.B1(_11352_),
    .Y(_11353_),
    .A2(_11343_),
    .A1(_11334_));
 sg13g2_a21oi_1 _18159_ (.A1(_11348_),
    .A2(_11352_),
    .Y(_11354_),
    .B1(net168));
 sg13g2_nor3_1 _18160_ (.A(_11344_),
    .B(net450),
    .C(_10247_),
    .Y(_11355_));
 sg13g2_or2_1 _18161_ (.X(_11356_),
    .B(_11355_),
    .A(_11354_));
 sg13g2_buf_1 _18162_ (.A(_11356_),
    .X(_11357_));
 sg13g2_a21oi_1 _18163_ (.A1(net897),
    .A2(_10244_),
    .Y(_11358_),
    .B1(_10245_));
 sg13g2_buf_1 _18164_ (.A(_11358_),
    .X(_11359_));
 sg13g2_inv_1 _18165_ (.Y(_11360_),
    .A(_10291_));
 sg13g2_nand2_1 _18166_ (.Y(_11361_),
    .A(net235),
    .B(_11360_));
 sg13g2_a21oi_2 _18167_ (.B1(_11361_),
    .Y(_11362_),
    .A2(_11343_),
    .A1(_11334_));
 sg13g2_nor4_2 _18168_ (.A(_11350_),
    .B(_11353_),
    .C(_11357_),
    .Y(_11363_),
    .D(_11362_));
 sg13g2_buf_8 _18169_ (.A(_11363_),
    .X(_11364_));
 sg13g2_nor2_1 _18170_ (.A(net79),
    .B(net28),
    .Y(_11365_));
 sg13g2_buf_2 _18171_ (.A(_11365_),
    .X(_11366_));
 sg13g2_buf_1 _18172_ (.A(net359),
    .X(_11367_));
 sg13g2_buf_1 _18173_ (.A(net118),
    .X(_11368_));
 sg13g2_buf_1 _18174_ (.A(net96),
    .X(_11369_));
 sg13g2_nand3b_1 _18175_ (.B(net277),
    .C(net87),
    .Y(_11370_),
    .A_N(_10719_));
 sg13g2_buf_1 _18176_ (.A(_11370_),
    .X(_11371_));
 sg13g2_nor2b_1 _18177_ (.A(_11366_),
    .B_N(_11371_),
    .Y(_11372_));
 sg13g2_buf_1 _18178_ (.A(\cpu.ex.r_mult[0] ),
    .X(_11373_));
 sg13g2_inv_1 _18179_ (.Y(_11374_),
    .A(_10140_));
 sg13g2_nor2_1 _18180_ (.A(net1117),
    .B(_11374_),
    .Y(_11375_));
 sg13g2_nand4_1 _18181_ (.B(net1037),
    .C(_10136_),
    .A(net1116),
    .Y(_11376_),
    .D(_11375_));
 sg13g2_buf_1 _18182_ (.A(_11376_),
    .X(_11377_));
 sg13g2_buf_1 _18183_ (.A(_11377_),
    .X(_11378_));
 sg13g2_nor2_1 _18184_ (.A(_09257_),
    .B(net1124),
    .Y(_11379_));
 sg13g2_nand2_1 _18185_ (.Y(_11380_),
    .A(_09271_),
    .B(_11379_));
 sg13g2_buf_2 _18186_ (.A(_11380_),
    .X(_11381_));
 sg13g2_nand2_1 _18187_ (.Y(_11382_),
    .A(net618),
    .B(_11381_));
 sg13g2_buf_2 _18188_ (.A(_11382_),
    .X(_11383_));
 sg13g2_nand2_1 _18189_ (.Y(_11384_),
    .A(_11373_),
    .B(_11383_));
 sg13g2_o21ai_1 _18190_ (.B1(_11384_),
    .Y(\cpu.ex.c_mult[0] ),
    .A1(_10148_),
    .A2(_11372_));
 sg13g2_buf_1 _18191_ (.A(\cpu.dec.load ),
    .X(_11385_));
 sg13g2_nand2_1 _18192_ (.Y(_11386_),
    .A(_08283_),
    .B(_08404_));
 sg13g2_nand2b_1 _18193_ (.Y(_11387_),
    .B(_09081_),
    .A_N(_09273_));
 sg13g2_nand2b_1 _18194_ (.Y(_11388_),
    .B(_11387_),
    .A_N(_11379_));
 sg13g2_buf_1 _18195_ (.A(_11388_),
    .X(_11389_));
 sg13g2_nor2_1 _18196_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11390_));
 sg13g2_nand2_1 _18197_ (.Y(_11391_),
    .A(_10561_),
    .B(\cpu.dec.r_swapsp ));
 sg13g2_nor2_1 _18198_ (.A(\cpu.ex.r_branch_stall ),
    .B(_09261_),
    .Y(_11392_));
 sg13g2_buf_1 _18199_ (.A(_11392_),
    .X(_11393_));
 sg13g2_nand2_1 _18200_ (.Y(_11394_),
    .A(_09081_),
    .B(_11393_));
 sg13g2_buf_1 _18201_ (.A(_11394_),
    .X(_11395_));
 sg13g2_nor2_1 _18202_ (.A(_09146_),
    .B(_11395_),
    .Y(_11396_));
 sg13g2_nand2_1 _18203_ (.Y(_11397_),
    .A(_10791_),
    .B(\cpu.cond[2] ));
 sg13g2_nand2_1 _18204_ (.Y(_11398_),
    .A(_00238_),
    .B(_11397_));
 sg13g2_nand2_1 _18205_ (.Y(_11399_),
    .A(_08336_),
    .B(_11398_));
 sg13g2_o21ai_1 _18206_ (.B1(_11399_),
    .Y(_11400_),
    .A1(_10791_),
    .A2(\cpu.dec.jmp ));
 sg13g2_nand4_1 _18207_ (.B(_11391_),
    .C(_11396_),
    .A(_11390_),
    .Y(_11401_),
    .D(_11400_));
 sg13g2_nand3_1 _18208_ (.B(_11389_),
    .C(_11401_),
    .A(_11386_),
    .Y(_11402_));
 sg13g2_buf_1 _18209_ (.A(_11402_),
    .X(_11403_));
 sg13g2_and2_1 _18210_ (.A(_09081_),
    .B(_11403_),
    .X(_11404_));
 sg13g2_buf_1 _18211_ (.A(_11404_),
    .X(_11405_));
 sg13g2_buf_1 _18212_ (.A(_11405_),
    .X(_11406_));
 sg13g2_nand2_1 _18213_ (.Y(_11407_),
    .A(_00294_),
    .B(net86));
 sg13g2_nand2b_1 _18214_ (.Y(_11408_),
    .B(_09765_),
    .A_N(_09767_));
 sg13g2_a21o_1 _18215_ (.A2(_11408_),
    .A1(_09771_),
    .B1(_09149_),
    .X(_11409_));
 sg13g2_buf_1 _18216_ (.A(_11409_),
    .X(_11410_));
 sg13g2_o21ai_1 _18217_ (.B1(_11407_),
    .Y(_11411_),
    .A1(net86),
    .A2(_11410_));
 sg13g2_nand2_1 _18218_ (.Y(_11412_),
    .A(net1132),
    .B(_11411_));
 sg13g2_o21ai_1 _18219_ (.B1(_11412_),
    .Y(_00054_),
    .A1(_11385_),
    .A2(_11407_));
 sg13g2_inv_1 _18220_ (.Y(_11413_),
    .A(net1124));
 sg13g2_buf_1 _18221_ (.A(_11413_),
    .X(_11414_));
 sg13g2_nand2_1 _18222_ (.Y(_11415_),
    .A(\cpu.dec.mult ),
    .B(net710));
 sg13g2_buf_1 _18223_ (.A(_11415_),
    .X(_11416_));
 sg13g2_buf_1 _18224_ (.A(_11416_),
    .X(_11417_));
 sg13g2_buf_1 _18225_ (.A(net499),
    .X(_11418_));
 sg13g2_buf_1 _18226_ (.A(net445),
    .X(_11419_));
 sg13g2_nand2_1 _18227_ (.Y(_11420_),
    .A(_11373_),
    .B(net402));
 sg13g2_buf_1 _18228_ (.A(net282),
    .X(_11421_));
 sg13g2_and2_1 _18229_ (.A(_11421_),
    .B(net118),
    .X(_11422_));
 sg13g2_mux2_1 _18230_ (.A0(_11420_),
    .A1(_11373_),
    .S(_11422_),
    .X(_11423_));
 sg13g2_buf_1 _18231_ (.A(_09278_),
    .X(_11424_));
 sg13g2_buf_1 _18232_ (.A(net444),
    .X(_11425_));
 sg13g2_a22oi_1 _18233_ (.Y(_11426_),
    .B1(_11422_),
    .B2(net401),
    .A2(_10722_),
    .A1(_11373_));
 sg13g2_o21ai_1 _18234_ (.B1(_11426_),
    .Y(_11427_),
    .A1(net877),
    .A2(_11423_));
 sg13g2_buf_1 _18235_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11428_));
 sg13g2_inv_1 _18236_ (.Y(_11429_),
    .A(_11428_));
 sg13g2_a21oi_1 _18237_ (.A1(_11378_),
    .A2(_11381_),
    .Y(_11430_),
    .B1(_11429_));
 sg13g2_a21o_1 _18238_ (.A2(_11427_),
    .A1(net618),
    .B1(_11430_),
    .X(\cpu.ex.c_mult[1] ));
 sg13g2_nand2_1 _18239_ (.Y(_11431_),
    .A(_11428_),
    .B(net402));
 sg13g2_buf_1 _18240_ (.A(net283),
    .X(_11432_));
 sg13g2_and2_1 _18241_ (.A(_11373_),
    .B(net282),
    .X(_11433_));
 sg13g2_buf_1 _18242_ (.A(_11433_),
    .X(_11434_));
 sg13g2_nand2_1 _18243_ (.Y(_11435_),
    .A(net445),
    .B(_11434_));
 sg13g2_xnor2_1 _18244_ (.Y(_11436_),
    .A(net233),
    .B(_11435_));
 sg13g2_nand2_1 _18245_ (.Y(_11437_),
    .A(net96),
    .B(_11436_));
 sg13g2_mux2_1 _18246_ (.A0(_11428_),
    .A1(_11431_),
    .S(_11437_),
    .X(_11438_));
 sg13g2_buf_1 _18247_ (.A(_10722_),
    .X(_11439_));
 sg13g2_and3_1 _18248_ (.X(_11440_),
    .A(net444),
    .B(net233),
    .C(_11368_));
 sg13g2_a21oi_1 _18249_ (.A1(_11428_),
    .A2(net85),
    .Y(_11441_),
    .B1(_11440_));
 sg13g2_o21ai_1 _18250_ (.B1(_11441_),
    .Y(_11442_),
    .A1(net877),
    .A2(_11438_));
 sg13g2_buf_2 _18251_ (.A(\cpu.ex.r_mult[2] ),
    .X(_11443_));
 sg13g2_and2_1 _18252_ (.A(_11443_),
    .B(_11383_),
    .X(_11444_));
 sg13g2_a21oi_1 _18253_ (.A1(net618),
    .A2(_11442_),
    .Y(_11445_),
    .B1(_11444_));
 sg13g2_inv_1 _18254_ (.Y(\cpu.ex.c_mult[2] ),
    .A(_11445_));
 sg13g2_buf_1 _18255_ (.A(\cpu.ex.r_mult[3] ),
    .X(_11446_));
 sg13g2_buf_1 _18256_ (.A(_11383_),
    .X(_11447_));
 sg13g2_nand2_1 _18257_ (.Y(_11448_),
    .A(_11429_),
    .B(_11252_));
 sg13g2_nor2_1 _18258_ (.A(_11429_),
    .B(_11252_),
    .Y(_11449_));
 sg13g2_a21oi_1 _18259_ (.A1(_11434_),
    .A2(_11448_),
    .Y(_11450_),
    .B1(_11449_));
 sg13g2_buf_1 _18260_ (.A(_11314_),
    .X(_11451_));
 sg13g2_buf_1 _18261_ (.A(net232),
    .X(_11452_));
 sg13g2_nand2_1 _18262_ (.Y(_11453_),
    .A(net213),
    .B(net87));
 sg13g2_buf_1 _18263_ (.A(_11290_),
    .X(_11454_));
 sg13g2_nand3_1 _18264_ (.B(net402),
    .C(net231),
    .A(_11443_),
    .Y(_11455_));
 sg13g2_o21ai_1 _18265_ (.B1(_11455_),
    .Y(_11456_),
    .A1(_11443_),
    .A2(_11453_));
 sg13g2_inv_2 _18266_ (.Y(_11457_),
    .A(net118));
 sg13g2_nand2_1 _18267_ (.Y(_11458_),
    .A(_11443_),
    .B(_11314_));
 sg13g2_nor2_2 _18268_ (.A(_11443_),
    .B(_11314_),
    .Y(_11459_));
 sg13g2_nand2_1 _18269_ (.Y(_11460_),
    .A(net96),
    .B(_11459_));
 sg13g2_a21oi_1 _18270_ (.A1(_11458_),
    .A2(_11460_),
    .Y(_11461_),
    .B1(_11450_));
 sg13g2_a21o_1 _18271_ (.A2(_11457_),
    .A1(_11443_),
    .B1(_11461_),
    .X(_11462_));
 sg13g2_a22oi_1 _18272_ (.Y(_11463_),
    .B1(_11462_),
    .B2(_11419_),
    .A2(_11456_),
    .A1(_11450_));
 sg13g2_and2_1 _18273_ (.A(net444),
    .B(net96),
    .X(_11464_));
 sg13g2_a22oi_1 _18274_ (.Y(_11465_),
    .B1(_11464_),
    .B2(net213),
    .A2(net85),
    .A1(_11443_));
 sg13g2_o21ai_1 _18275_ (.B1(_11465_),
    .Y(_11466_),
    .A1(net877),
    .A2(_11463_));
 sg13g2_buf_1 _18276_ (.A(net618),
    .X(_11467_));
 sg13g2_a22oi_1 _18277_ (.Y(_11468_),
    .B1(_11466_),
    .B2(_11467_),
    .A2(net214),
    .A1(_11446_));
 sg13g2_inv_1 _18278_ (.Y(\cpu.ex.c_mult[3] ),
    .A(_11468_));
 sg13g2_buf_2 _18279_ (.A(\cpu.ex.r_mult[4] ),
    .X(_11469_));
 sg13g2_nand2_1 _18280_ (.Y(_11470_),
    .A(_11446_),
    .B(_11416_));
 sg13g2_a221oi_1 _18281_ (.B2(_11448_),
    .C1(_11449_),
    .B1(_11434_),
    .A1(_11443_),
    .Y(_11471_),
    .A2(net232));
 sg13g2_buf_1 _18282_ (.A(_11471_),
    .X(_11472_));
 sg13g2_nor3_1 _18283_ (.A(net504),
    .B(_11459_),
    .C(_11472_),
    .Y(_11473_));
 sg13g2_xnor2_1 _18284_ (.Y(_11474_),
    .A(net281),
    .B(_11473_));
 sg13g2_nand2_1 _18285_ (.Y(_11475_),
    .A(_11368_),
    .B(_11474_));
 sg13g2_mux2_1 _18286_ (.A0(_11446_),
    .A1(_11470_),
    .S(_11475_),
    .X(_11476_));
 sg13g2_a22oi_1 _18287_ (.Y(_11477_),
    .B1(_11464_),
    .B2(_11474_),
    .A2(_10722_),
    .A1(_11446_));
 sg13g2_o21ai_1 _18288_ (.B1(_11477_),
    .Y(_11478_),
    .A1(net877),
    .A2(_11476_));
 sg13g2_a22oi_1 _18289_ (.Y(_11479_),
    .B1(_11478_),
    .B2(net618),
    .A2(_11383_),
    .A1(_11469_));
 sg13g2_inv_1 _18290_ (.Y(\cpu.ex.c_mult[4] ),
    .A(_11479_));
 sg13g2_nand2_1 _18291_ (.Y(_11480_),
    .A(_11469_),
    .B(_11419_));
 sg13g2_o21ai_1 _18292_ (.B1(net281),
    .Y(_11481_),
    .A1(_11459_),
    .A2(_11472_));
 sg13g2_nor3_1 _18293_ (.A(_10659_),
    .B(_11459_),
    .C(_11472_),
    .Y(_11482_));
 sg13g2_a21oi_1 _18294_ (.A1(_11446_),
    .A2(_11481_),
    .Y(_11483_),
    .B1(_11482_));
 sg13g2_or3_1 _18295_ (.A(net444),
    .B(_10635_),
    .C(_11483_),
    .X(_11484_));
 sg13g2_o21ai_1 _18296_ (.B1(_10635_),
    .Y(_11485_),
    .A1(_11424_),
    .A2(_11483_));
 sg13g2_nand3_1 _18297_ (.B(_11484_),
    .C(_11485_),
    .A(net87),
    .Y(_11486_));
 sg13g2_mux2_1 _18298_ (.A0(_11469_),
    .A1(_11480_),
    .S(_11486_),
    .X(_11487_));
 sg13g2_nor3_1 _18299_ (.A(net402),
    .B(net216),
    .C(_11457_),
    .Y(_11488_));
 sg13g2_a21oi_1 _18300_ (.A1(_11469_),
    .A2(_11439_),
    .Y(_11489_),
    .B1(_11488_));
 sg13g2_o21ai_1 _18301_ (.B1(_11489_),
    .Y(_11490_),
    .A1(net877),
    .A2(_11487_));
 sg13g2_buf_2 _18302_ (.A(\cpu.ex.r_mult[5] ),
    .X(_11491_));
 sg13g2_inv_1 _18303_ (.Y(_11492_),
    .A(_11491_));
 sg13g2_a21oi_1 _18304_ (.A1(_11378_),
    .A2(_11381_),
    .Y(_11493_),
    .B1(_11492_));
 sg13g2_a21oi_1 _18305_ (.A1(net618),
    .A2(_11490_),
    .Y(_11494_),
    .B1(_11493_));
 sg13g2_inv_1 _18306_ (.Y(\cpu.ex.c_mult[5] ),
    .A(_11494_));
 sg13g2_buf_1 _18307_ (.A(\cpu.ex.r_mult[6] ),
    .X(_11495_));
 sg13g2_nand2_1 _18308_ (.Y(_11496_),
    .A(_11491_),
    .B(net445));
 sg13g2_buf_1 _18309_ (.A(_11309_),
    .X(_11497_));
 sg13g2_nand2_1 _18310_ (.Y(_11498_),
    .A(_10628_),
    .B(_10631_));
 sg13g2_buf_2 _18311_ (.A(_11498_),
    .X(_11499_));
 sg13g2_nor2_1 _18312_ (.A(_09269_),
    .B(net358),
    .Y(_11500_));
 sg13g2_o21ai_1 _18313_ (.B1(_11500_),
    .Y(_11501_),
    .A1(_11469_),
    .A2(_11499_));
 sg13g2_inv_1 _18314_ (.Y(_11502_),
    .A(_11469_));
 sg13g2_a21o_1 _18315_ (.A2(net241),
    .A1(_11502_),
    .B1(_11470_),
    .X(_11503_));
 sg13g2_a221oi_1 _18316_ (.B2(_11503_),
    .C1(_11459_),
    .B1(_11501_),
    .A1(_11450_),
    .Y(_11504_),
    .A2(_11458_));
 sg13g2_buf_1 _18317_ (.A(_11504_),
    .X(_11505_));
 sg13g2_nand3_1 _18318_ (.B(_11416_),
    .C(_11499_),
    .A(_11469_),
    .Y(_11506_));
 sg13g2_nor2_1 _18319_ (.A(net358),
    .B(_11470_),
    .Y(_11507_));
 sg13g2_o21ai_1 _18320_ (.B1(_11507_),
    .Y(_11508_),
    .A1(_11469_),
    .A2(_11499_));
 sg13g2_nand2_1 _18321_ (.Y(_11509_),
    .A(_11506_),
    .B(_11508_));
 sg13g2_nor3_1 _18322_ (.A(net276),
    .B(_11505_),
    .C(_11509_),
    .Y(_11510_));
 sg13g2_o21ai_1 _18323_ (.B1(net276),
    .Y(_11511_),
    .A1(_11505_),
    .A2(_11509_));
 sg13g2_nand3b_1 _18324_ (.B(_11511_),
    .C(net96),
    .Y(_11512_),
    .A_N(_11510_));
 sg13g2_mux2_1 _18325_ (.A0(_11491_),
    .A1(_11496_),
    .S(_11512_),
    .X(_11513_));
 sg13g2_buf_1 _18326_ (.A(net276),
    .X(_11514_));
 sg13g2_and3_1 _18327_ (.X(_11515_),
    .A(_11424_),
    .B(net230),
    .C(net96));
 sg13g2_a21oi_1 _18328_ (.A1(_11491_),
    .A2(_10722_),
    .Y(_11516_),
    .B1(_11515_));
 sg13g2_o21ai_1 _18329_ (.B1(_11516_),
    .Y(_11517_),
    .A1(_11414_),
    .A2(_11513_));
 sg13g2_a22oi_1 _18330_ (.Y(_11518_),
    .B1(_11517_),
    .B2(net618),
    .A2(_11383_),
    .A1(_11495_));
 sg13g2_inv_1 _18331_ (.Y(\cpu.ex.c_mult[6] ),
    .A(_11518_));
 sg13g2_o21ai_1 _18332_ (.B1(_11377_),
    .Y(_11519_),
    .A1(net1124),
    .A2(net444));
 sg13g2_buf_1 _18333_ (.A(_11519_),
    .X(_11520_));
 sg13g2_nand2_1 _18334_ (.Y(_11521_),
    .A(net1108),
    .B(net445));
 sg13g2_buf_8 _18335_ (.A(_11282_),
    .X(_11522_));
 sg13g2_o21ai_1 _18336_ (.B1(_11511_),
    .Y(_11523_),
    .A1(_11510_),
    .A2(_11496_));
 sg13g2_buf_1 _18337_ (.A(_11523_),
    .X(_11524_));
 sg13g2_nand2_1 _18338_ (.Y(_11525_),
    .A(net229),
    .B(_11524_));
 sg13g2_nand2b_1 _18339_ (.Y(_11526_),
    .B(net242),
    .A_N(_11524_));
 sg13g2_nand3_1 _18340_ (.B(_11525_),
    .C(_11526_),
    .A(_11369_),
    .Y(_11527_));
 sg13g2_xnor2_1 _18341_ (.Y(_11528_),
    .A(_11521_),
    .B(_11527_));
 sg13g2_buf_1 _18342_ (.A(\cpu.ex.r_mult[7] ),
    .X(_11529_));
 sg13g2_buf_1 _18343_ (.A(_11529_),
    .X(_11530_));
 sg13g2_nor2_1 _18344_ (.A(_10146_),
    .B(_10723_),
    .Y(_11531_));
 sg13g2_buf_2 _18345_ (.A(_11531_),
    .X(_11532_));
 sg13g2_a22oi_1 _18346_ (.Y(_11533_),
    .B1(_11532_),
    .B2(net1108),
    .A2(_11383_),
    .A1(_11530_));
 sg13g2_o21ai_1 _18347_ (.B1(_11533_),
    .Y(\cpu.ex.c_mult[7] ),
    .A1(_11520_),
    .A2(_11528_));
 sg13g2_nand2_1 _18348_ (.Y(_11534_),
    .A(net767),
    .B(_10456_));
 sg13g2_buf_2 _18349_ (.A(_11534_),
    .X(_11535_));
 sg13g2_buf_1 _18350_ (.A(_11535_),
    .X(_11536_));
 sg13g2_nor2_1 _18351_ (.A(_11505_),
    .B(_11509_),
    .Y(_11537_));
 sg13g2_o21ai_1 _18352_ (.B1(_11416_),
    .Y(_11538_),
    .A1(_11491_),
    .A2(net1108));
 sg13g2_nand3_1 _18353_ (.B(net229),
    .C(_11538_),
    .A(net276),
    .Y(_11539_));
 sg13g2_xnor2_1 _18354_ (.Y(_11540_),
    .A(net1108),
    .B(_10482_));
 sg13g2_nand4_1 _18355_ (.B(net499),
    .C(net286),
    .A(_11491_),
    .Y(_11541_),
    .D(_11540_));
 sg13g2_nor2b_1 _18356_ (.A(_11491_),
    .B_N(net1108),
    .Y(_11542_));
 sg13g2_nand4_1 _18357_ (.B(net276),
    .C(_10483_),
    .A(net499),
    .Y(_11543_),
    .D(_11542_));
 sg13g2_and3_1 _18358_ (.X(_11544_),
    .A(_11539_),
    .B(_11541_),
    .C(_11543_));
 sg13g2_nand2_1 _18359_ (.Y(_11545_),
    .A(net1108),
    .B(net229));
 sg13g2_a21oi_1 _18360_ (.A1(_10332_),
    .A2(_10362_),
    .Y(_11546_),
    .B1(_11492_));
 sg13g2_o21ai_1 _18361_ (.B1(_11546_),
    .Y(_11547_),
    .A1(net1108),
    .A2(net229));
 sg13g2_a21o_1 _18362_ (.A2(_11547_),
    .A1(_11545_),
    .B1(_09269_),
    .X(_11548_));
 sg13g2_buf_1 _18363_ (.A(_11548_),
    .X(_11549_));
 sg13g2_o21ai_1 _18364_ (.B1(_11549_),
    .Y(_11550_),
    .A1(_11537_),
    .A2(_11544_));
 sg13g2_xnor2_1 _18365_ (.Y(_11551_),
    .A(_11536_),
    .B(_11550_));
 sg13g2_nor2_1 _18366_ (.A(_11457_),
    .B(_11551_),
    .Y(_11552_));
 sg13g2_a22oi_1 _18367_ (.Y(_11553_),
    .B1(_11552_),
    .B2(net401),
    .A2(net85),
    .A1(_11530_));
 sg13g2_nand2_1 _18368_ (.Y(_11554_),
    .A(net1022),
    .B(net499));
 sg13g2_inv_1 _18369_ (.Y(_11555_),
    .A(_11554_));
 sg13g2_o21ai_1 _18370_ (.B1(_11555_),
    .Y(_11556_),
    .A1(_11457_),
    .A2(_11551_));
 sg13g2_or3_1 _18371_ (.A(net1022),
    .B(_11457_),
    .C(_11551_),
    .X(_11557_));
 sg13g2_a21o_1 _18372_ (.A2(_11557_),
    .A1(_11556_),
    .B1(net877),
    .X(_11558_));
 sg13g2_a21oi_1 _18373_ (.A1(_11553_),
    .A2(_11558_),
    .Y(_11559_),
    .B1(_10147_));
 sg13g2_buf_2 _18374_ (.A(\cpu.ex.r_mult[8] ),
    .X(_11560_));
 sg13g2_nand2_1 _18375_ (.Y(_11561_),
    .A(_11560_),
    .B(net214));
 sg13g2_nand2b_1 _18376_ (.Y(\cpu.ex.c_mult[8] ),
    .B(_11561_),
    .A_N(_11559_));
 sg13g2_buf_1 _18377_ (.A(_10329_),
    .X(_11562_));
 sg13g2_nor2_1 _18378_ (.A(_10719_),
    .B(_10146_),
    .Y(_11563_));
 sg13g2_nand2_1 _18379_ (.Y(_11564_),
    .A(_11560_),
    .B(net499));
 sg13g2_and4_1 _18380_ (.A(net212),
    .B(net87),
    .C(_11563_),
    .D(_11564_),
    .X(_11565_));
 sg13g2_buf_1 _18381_ (.A(_10729_),
    .X(_11566_));
 sg13g2_and4_1 _18382_ (.A(_11566_),
    .B(_11369_),
    .C(_11563_),
    .D(_11564_),
    .X(_11567_));
 sg13g2_a21o_1 _18383_ (.A2(_11524_),
    .A1(net229),
    .B1(_11536_),
    .X(_11568_));
 sg13g2_nor2_1 _18384_ (.A(net1022),
    .B(_11535_),
    .Y(_11569_));
 sg13g2_nor2_1 _18385_ (.A(_11521_),
    .B(_11569_),
    .Y(_11570_));
 sg13g2_and3_1 _18386_ (.X(_11571_),
    .A(net192),
    .B(net229),
    .C(_11524_));
 sg13g2_a221oi_1 _18387_ (.B2(_11526_),
    .C1(_11571_),
    .B1(_11570_),
    .A1(_11555_),
    .Y(_11572_),
    .A2(_11568_));
 sg13g2_mux2_1 _18388_ (.A0(_11565_),
    .A1(_11567_),
    .S(_11572_),
    .X(_11573_));
 sg13g2_or2_1 _18389_ (.X(_11574_),
    .B(_11564_),
    .A(_11520_));
 sg13g2_buf_1 _18390_ (.A(_11574_),
    .X(_11575_));
 sg13g2_nor2_1 _18391_ (.A(_11562_),
    .B(_11575_),
    .Y(_11576_));
 sg13g2_nor2_1 _18392_ (.A(_11566_),
    .B(_11575_),
    .Y(_11577_));
 sg13g2_mux2_1 _18393_ (.A0(_11576_),
    .A1(_11577_),
    .S(_11572_),
    .X(_11578_));
 sg13g2_buf_1 _18394_ (.A(net87),
    .X(_11579_));
 sg13g2_buf_1 _18395_ (.A(\cpu.ex.r_mult[9] ),
    .X(_11580_));
 sg13g2_a22oi_1 _18396_ (.Y(_11581_),
    .B1(_11532_),
    .B2(_11560_),
    .A2(_11383_),
    .A1(_11580_));
 sg13g2_o21ai_1 _18397_ (.B1(_11581_),
    .Y(_11582_),
    .A1(_11579_),
    .A2(_11575_));
 sg13g2_or3_1 _18398_ (.A(_11573_),
    .B(_11578_),
    .C(_11582_),
    .X(\cpu.ex.c_mult[9] ));
 sg13g2_inv_1 _18399_ (.Y(_11583_),
    .A(_11580_));
 sg13g2_nand3_1 _18400_ (.B(_11541_),
    .C(_11543_),
    .A(_11539_),
    .Y(_11584_));
 sg13g2_inv_1 _18401_ (.Y(_11585_),
    .A(_11529_));
 sg13g2_nand3_1 _18402_ (.B(_11560_),
    .C(net243),
    .A(_11585_),
    .Y(_11586_));
 sg13g2_or3_1 _18403_ (.A(_11560_),
    .B(_10294_),
    .C(_10326_),
    .X(_11587_));
 sg13g2_buf_1 _18404_ (.A(_11587_),
    .X(_11588_));
 sg13g2_o21ai_1 _18405_ (.B1(_11560_),
    .Y(_11589_),
    .A1(_10294_),
    .A2(_10326_));
 sg13g2_nand3_1 _18406_ (.B(_11588_),
    .C(_11589_),
    .A(net1022),
    .Y(_11590_));
 sg13g2_mux2_1 _18407_ (.A0(_11586_),
    .A1(_11590_),
    .S(_10747_),
    .X(_11591_));
 sg13g2_o21ai_1 _18408_ (.B1(_11416_),
    .Y(_11592_),
    .A1(net1022),
    .A2(_11560_));
 sg13g2_nand3_1 _18409_ (.B(_11535_),
    .C(_11592_),
    .A(_10729_),
    .Y(_11593_));
 sg13g2_o21ai_1 _18410_ (.B1(_11593_),
    .Y(_11594_),
    .A1(net504),
    .A2(_11591_));
 sg13g2_nand3b_1 _18411_ (.B(_11584_),
    .C(_11594_),
    .Y(_11595_),
    .A_N(_11537_));
 sg13g2_buf_1 _18412_ (.A(_11595_),
    .X(_11596_));
 sg13g2_nand2_1 _18413_ (.Y(_11597_),
    .A(_10729_),
    .B(_11535_));
 sg13g2_nand3_1 _18414_ (.B(_11417_),
    .C(_11588_),
    .A(net1022),
    .Y(_11598_));
 sg13g2_a21oi_1 _18415_ (.A1(_11597_),
    .A2(_11598_),
    .Y(_11599_),
    .B1(_11549_));
 sg13g2_buf_1 _18416_ (.A(_10747_),
    .X(_11600_));
 sg13g2_nor3_1 _18417_ (.A(net191),
    .B(_11549_),
    .C(_11564_),
    .Y(_11601_));
 sg13g2_nand4_1 _18418_ (.B(_11417_),
    .C(_11535_),
    .A(net1022),
    .Y(_11602_),
    .D(_11588_));
 sg13g2_o21ai_1 _18419_ (.B1(_11602_),
    .Y(_11603_),
    .A1(_10329_),
    .A2(_11564_));
 sg13g2_nor3_2 _18420_ (.A(_11599_),
    .B(_11601_),
    .C(_11603_),
    .Y(_11604_));
 sg13g2_nand2_1 _18421_ (.Y(_11605_),
    .A(net285),
    .B(net96));
 sg13g2_a21oi_1 _18422_ (.A1(_11596_),
    .A2(_11604_),
    .Y(_11606_),
    .B1(_11605_));
 sg13g2_or2_1 _18423_ (.X(_11607_),
    .B(_10387_),
    .A(_10366_));
 sg13g2_buf_1 _18424_ (.A(_11607_),
    .X(_11608_));
 sg13g2_buf_1 _18425_ (.A(_11608_),
    .X(_11609_));
 sg13g2_and4_1 _18426_ (.A(net275),
    .B(net96),
    .C(_11596_),
    .D(_11604_),
    .X(_11610_));
 sg13g2_buf_1 _18427_ (.A(_11610_),
    .X(_11611_));
 sg13g2_o21ai_1 _18428_ (.B1(_11425_),
    .Y(_11612_),
    .A1(_11606_),
    .A2(_11611_));
 sg13g2_o21ai_1 _18429_ (.B1(_11612_),
    .Y(_11613_),
    .A1(_11583_),
    .A2(_10723_));
 sg13g2_or4_1 _18430_ (.A(_11583_),
    .B(_11425_),
    .C(_11606_),
    .D(_11611_),
    .X(_11614_));
 sg13g2_o21ai_1 _18431_ (.B1(_11583_),
    .Y(_11615_),
    .A1(_11606_),
    .A2(_11611_));
 sg13g2_a21oi_1 _18432_ (.A1(_11614_),
    .A2(_11615_),
    .Y(_11616_),
    .B1(_11414_));
 sg13g2_o21ai_1 _18433_ (.B1(_11467_),
    .Y(_11617_),
    .A1(_11613_),
    .A2(_11616_));
 sg13g2_buf_1 _18434_ (.A(\cpu.ex.r_mult[10] ),
    .X(_11618_));
 sg13g2_nand2_1 _18435_ (.Y(_11619_),
    .A(_11618_),
    .B(net214));
 sg13g2_nand2_1 _18436_ (.Y(\cpu.ex.c_mult[10] ),
    .A(_11617_),
    .B(_11619_));
 sg13g2_nand2_1 _18437_ (.Y(_11620_),
    .A(net1107),
    .B(_11416_));
 sg13g2_a21oi_1 _18438_ (.A1(_10429_),
    .A2(_10456_),
    .Y(_11621_),
    .B1(_11585_));
 sg13g2_o21ai_1 _18439_ (.B1(net499),
    .Y(_11622_),
    .A1(net1108),
    .A2(_11621_));
 sg13g2_a221oi_1 _18440_ (.B2(net242),
    .C1(net243),
    .B1(_11622_),
    .A1(net191),
    .Y(_11623_),
    .A2(_11554_));
 sg13g2_nand2_1 _18441_ (.Y(_11624_),
    .A(net275),
    .B(_11623_));
 sg13g2_nor2_1 _18442_ (.A(_11583_),
    .B(_09269_),
    .Y(_11625_));
 sg13g2_o21ai_1 _18443_ (.B1(_11625_),
    .Y(_11626_),
    .A1(net275),
    .A2(_11623_));
 sg13g2_a22oi_1 _18444_ (.Y(_11627_),
    .B1(_11622_),
    .B2(net242),
    .A2(_11554_),
    .A1(net191));
 sg13g2_inv_1 _18445_ (.Y(_11628_),
    .A(_11560_));
 sg13g2_nor2_1 _18446_ (.A(_11580_),
    .B(net275),
    .Y(_11629_));
 sg13g2_nor3_1 _18447_ (.A(_11628_),
    .B(net504),
    .C(_11629_),
    .Y(_11630_));
 sg13g2_o21ai_1 _18448_ (.B1(_11630_),
    .Y(_11631_),
    .A1(net228),
    .A2(_11627_));
 sg13g2_nand3_1 _18449_ (.B(_11626_),
    .C(_11631_),
    .A(_11624_),
    .Y(_11632_));
 sg13g2_buf_1 _18450_ (.A(_11632_),
    .X(_11633_));
 sg13g2_o21ai_1 _18451_ (.B1(_11580_),
    .Y(_11634_),
    .A1(_10366_),
    .A2(_10387_));
 sg13g2_o21ai_1 _18452_ (.B1(_11634_),
    .Y(_11635_),
    .A1(_11589_),
    .A2(_11629_));
 sg13g2_nand2_1 _18453_ (.Y(_11636_),
    .A(net1022),
    .B(_11535_));
 sg13g2_a21oi_1 _18454_ (.A1(_11545_),
    .A2(_11636_),
    .Y(_11637_),
    .B1(_11569_));
 sg13g2_o21ai_1 _18455_ (.B1(_11418_),
    .Y(_11638_),
    .A1(_11635_),
    .A2(_11637_));
 sg13g2_nand2b_1 _18456_ (.Y(_11639_),
    .B(_11638_),
    .A_N(_11524_));
 sg13g2_buf_2 _18457_ (.A(_11639_),
    .X(_11640_));
 sg13g2_nand3_1 _18458_ (.B(_11633_),
    .C(_11640_),
    .A(net240),
    .Y(_11641_));
 sg13g2_a21o_1 _18459_ (.A2(_11640_),
    .A1(_11633_),
    .B1(net240),
    .X(_11642_));
 sg13g2_nand3_1 _18460_ (.B(_11641_),
    .C(_11642_),
    .A(net78),
    .Y(_11643_));
 sg13g2_xnor2_1 _18461_ (.Y(_11644_),
    .A(_11620_),
    .B(_11643_));
 sg13g2_buf_1 _18462_ (.A(\cpu.ex.r_mult[11] ),
    .X(_11645_));
 sg13g2_buf_1 _18463_ (.A(_11645_),
    .X(_11646_));
 sg13g2_a22oi_1 _18464_ (.Y(_11647_),
    .B1(_11532_),
    .B2(net1107),
    .A2(net214),
    .A1(_11646_));
 sg13g2_o21ai_1 _18465_ (.B1(_11647_),
    .Y(\cpu.ex.c_mult[11] ),
    .A1(_11520_),
    .A2(_11644_));
 sg13g2_nand2_1 _18466_ (.Y(_11648_),
    .A(net1107),
    .B(_11625_));
 sg13g2_nor2_1 _18467_ (.A(_11609_),
    .B(net240),
    .Y(_11649_));
 sg13g2_a221oi_1 _18468_ (.B2(_11238_),
    .C1(_11649_),
    .B1(_11135_),
    .A1(_10964_),
    .Y(_11650_),
    .A2(_11050_));
 sg13g2_mux2_1 _18469_ (.A0(net1107),
    .A1(_11620_),
    .S(net280),
    .X(_11651_));
 sg13g2_nand2_1 _18470_ (.Y(_11652_),
    .A(net504),
    .B(_10716_));
 sg13g2_o21ai_1 _18471_ (.B1(_11652_),
    .Y(_11653_),
    .A1(_11580_),
    .A2(_11651_));
 sg13g2_and2_1 _18472_ (.A(net285),
    .B(_11625_),
    .X(_11654_));
 sg13g2_nor2_1 _18473_ (.A(net1107),
    .B(net280),
    .Y(_11655_));
 sg13g2_a22oi_1 _18474_ (.Y(_11656_),
    .B1(_11654_),
    .B2(_11655_),
    .A2(_11653_),
    .A1(net275));
 sg13g2_o21ai_1 _18475_ (.B1(_11656_),
    .Y(_11657_),
    .A1(_11648_),
    .A2(_11650_));
 sg13g2_nor3_1 _18476_ (.A(_11585_),
    .B(_11628_),
    .C(_11648_),
    .Y(_11658_));
 sg13g2_mux2_1 _18477_ (.A0(_11658_),
    .A1(_11594_),
    .S(_11240_),
    .X(_11659_));
 sg13g2_nand3_1 _18478_ (.B(_11657_),
    .C(_11659_),
    .A(_11550_),
    .Y(_11660_));
 sg13g2_o21ai_1 _18479_ (.B1(net1107),
    .Y(_11661_),
    .A1(_10691_),
    .A2(_10714_));
 sg13g2_nor3_1 _18480_ (.A(net1107),
    .B(_10691_),
    .C(_10714_),
    .Y(_11662_));
 sg13g2_nor2_1 _18481_ (.A(_11628_),
    .B(net243),
    .Y(_11663_));
 sg13g2_a221oi_1 _18482_ (.B2(net284),
    .C1(_11585_),
    .B1(_10429_),
    .A1(_11628_),
    .Y(_11664_),
    .A2(net243));
 sg13g2_nor3_1 _18483_ (.A(net275),
    .B(_11663_),
    .C(_11664_),
    .Y(_11665_));
 sg13g2_o21ai_1 _18484_ (.B1(net275),
    .Y(_11666_),
    .A1(_11663_),
    .A2(_11664_));
 sg13g2_o21ai_1 _18485_ (.B1(_11666_),
    .Y(_11667_),
    .A1(_11583_),
    .A2(_11665_));
 sg13g2_nand2b_1 _18486_ (.Y(_11668_),
    .B(_11667_),
    .A_N(_11662_));
 sg13g2_a21o_1 _18487_ (.A2(_11668_),
    .A1(_11661_),
    .B1(net444),
    .X(_11669_));
 sg13g2_a21oi_1 _18488_ (.A1(_11660_),
    .A2(_11669_),
    .Y(_11670_),
    .B1(net194));
 sg13g2_and3_1 _18489_ (.X(_11671_),
    .A(net194),
    .B(_11660_),
    .C(_11669_));
 sg13g2_o21ai_1 _18490_ (.B1(_11579_),
    .Y(_11672_),
    .A1(_11670_),
    .A2(_11671_));
 sg13g2_nand2_1 _18491_ (.Y(_11673_),
    .A(net1021),
    .B(net402));
 sg13g2_xnor2_1 _18492_ (.Y(_11674_),
    .A(_11672_),
    .B(_11673_));
 sg13g2_buf_1 _18493_ (.A(\cpu.ex.r_mult[12] ),
    .X(_11675_));
 sg13g2_a22oi_1 _18494_ (.Y(_11676_),
    .B1(_11532_),
    .B2(net1021),
    .A2(_11447_),
    .A1(_11675_));
 sg13g2_o21ai_1 _18495_ (.B1(_11676_),
    .Y(_11677_),
    .A1(_11520_),
    .A2(_11674_));
 sg13g2_buf_1 _18496_ (.A(_11677_),
    .X(\cpu.ex.c_mult[12] ));
 sg13g2_buf_1 _18497_ (.A(\cpu.ex.r_mult[13] ),
    .X(_11678_));
 sg13g2_nor2_1 _18498_ (.A(_11678_),
    .B(net568),
    .Y(_11679_));
 sg13g2_and3_1 _18499_ (.X(_11680_),
    .A(_11645_),
    .B(_10662_),
    .C(_10687_));
 sg13g2_xnor2_1 _18500_ (.Y(_11681_),
    .A(net1021),
    .B(_11300_));
 sg13g2_and2_1 _18501_ (.A(net1107),
    .B(net280),
    .X(_11682_));
 sg13g2_a22oi_1 _18502_ (.Y(_11683_),
    .B1(_11681_),
    .B2(_11682_),
    .A2(_11680_),
    .A1(_11655_));
 sg13g2_o21ai_1 _18503_ (.B1(_11418_),
    .Y(_11684_),
    .A1(_11618_),
    .A2(_11646_));
 sg13g2_nand3_1 _18504_ (.B(net240),
    .C(_11684_),
    .A(net194),
    .Y(_11685_));
 sg13g2_o21ai_1 _18505_ (.B1(_11685_),
    .Y(_11686_),
    .A1(net444),
    .A2(_11683_));
 sg13g2_nand3_1 _18506_ (.B(_11640_),
    .C(_11686_),
    .A(_11633_),
    .Y(_11687_));
 sg13g2_nor3_1 _18507_ (.A(net1021),
    .B(_11298_),
    .C(_11299_),
    .Y(_11688_));
 sg13g2_o21ai_1 _18508_ (.B1(net1021),
    .Y(_11689_),
    .A1(_11298_),
    .A2(_11299_));
 sg13g2_o21ai_1 _18509_ (.B1(_11689_),
    .Y(_11690_),
    .A1(_11661_),
    .A2(_11688_));
 sg13g2_and2_1 _18510_ (.A(net445),
    .B(_11690_),
    .X(_11691_));
 sg13g2_inv_1 _18511_ (.Y(_11692_),
    .A(_11691_));
 sg13g2_nand2_1 _18512_ (.Y(_11693_),
    .A(net217),
    .B(net78));
 sg13g2_a21oi_1 _18513_ (.A1(_11687_),
    .A2(_11692_),
    .Y(_11694_),
    .B1(_11693_));
 sg13g2_buf_1 _18514_ (.A(_11329_),
    .X(_11695_));
 sg13g2_and4_1 _18515_ (.A(net211),
    .B(net87),
    .C(_11687_),
    .D(_11692_),
    .X(_11696_));
 sg13g2_buf_1 _18516_ (.A(_11696_),
    .X(_11697_));
 sg13g2_o21ai_1 _18517_ (.B1(net401),
    .Y(_11698_),
    .A1(_11694_),
    .A2(_11697_));
 sg13g2_and2_1 _18518_ (.A(_09271_),
    .B(_11379_),
    .X(_11699_));
 sg13g2_buf_1 _18519_ (.A(_11699_),
    .X(_11700_));
 sg13g2_a221oi_1 _18520_ (.B2(net1105),
    .C1(net691),
    .B1(_11700_),
    .A1(net1106),
    .Y(_11701_),
    .A2(_11439_));
 sg13g2_nand3_1 _18521_ (.B(net1106),
    .C(net402),
    .A(net1124),
    .Y(_11702_));
 sg13g2_or3_1 _18522_ (.A(_11694_),
    .B(_11697_),
    .C(_11702_),
    .X(_11703_));
 sg13g2_nor2_1 _18523_ (.A(net877),
    .B(net1106),
    .Y(_11704_));
 sg13g2_o21ai_1 _18524_ (.B1(_11704_),
    .Y(_11705_),
    .A1(_11694_),
    .A2(_11697_));
 sg13g2_nand4_1 _18525_ (.B(_11701_),
    .C(_11703_),
    .A(_11698_),
    .Y(_11706_),
    .D(_11705_));
 sg13g2_nor2b_1 _18526_ (.A(_11679_),
    .B_N(_11706_),
    .Y(\cpu.ex.c_mult[13] ));
 sg13g2_buf_1 _18527_ (.A(net168),
    .X(_11707_));
 sg13g2_nand3_1 _18528_ (.B(net142),
    .C(net78),
    .A(net401),
    .Y(_11708_));
 sg13g2_buf_1 _18529_ (.A(_11360_),
    .X(_11709_));
 sg13g2_inv_1 _18530_ (.Y(_11710_),
    .A(\cpu.ex.r_mult[12] ));
 sg13g2_o21ai_1 _18531_ (.B1(_11661_),
    .Y(_11711_),
    .A1(_11634_),
    .A2(_11662_));
 sg13g2_o21ai_1 _18532_ (.B1(_11711_),
    .Y(_11712_),
    .A1(net1021),
    .A2(_10689_));
 sg13g2_a22oi_1 _18533_ (.Y(_11713_),
    .B1(_10689_),
    .B2(net1021),
    .A2(_11329_),
    .A1(net1106));
 sg13g2_a22oi_1 _18534_ (.Y(_11714_),
    .B1(_11712_),
    .B2(_11713_),
    .A2(net217),
    .A1(_11710_));
 sg13g2_buf_1 _18535_ (.A(_11714_),
    .X(_11715_));
 sg13g2_nor4_1 _18536_ (.A(net1105),
    .B(net141),
    .C(_11457_),
    .D(_11715_),
    .Y(_11716_));
 sg13g2_nand2_1 _18537_ (.Y(_11717_),
    .A(net1105),
    .B(net499));
 sg13g2_nor3_1 _18538_ (.A(net142),
    .B(_11715_),
    .C(_11717_),
    .Y(_11718_));
 sg13g2_nor2_1 _18539_ (.A(_10764_),
    .B(_11648_),
    .Y(_11719_));
 sg13g2_a221oi_1 _18540_ (.B2(_11655_),
    .C1(_11719_),
    .B1(_11654_),
    .A1(net275),
    .Y(_11720_),
    .A2(_11653_));
 sg13g2_xnor2_1 _18541_ (.Y(_11721_),
    .A(net1106),
    .B(_10425_));
 sg13g2_nor2_1 _18542_ (.A(_11710_),
    .B(_11329_),
    .Y(_11722_));
 sg13g2_a21oi_1 _18543_ (.A1(_10662_),
    .A2(_10687_),
    .Y(_11723_),
    .B1(net1021));
 sg13g2_a22oi_1 _18544_ (.Y(_11724_),
    .B1(_11722_),
    .B2(_11723_),
    .A2(_11721_),
    .A1(_11680_));
 sg13g2_o21ai_1 _18545_ (.B1(net499),
    .Y(_11725_),
    .A1(_11645_),
    .A2(_11675_));
 sg13g2_nand3_1 _18546_ (.B(_10689_),
    .C(_11725_),
    .A(_11329_),
    .Y(_11726_));
 sg13g2_o21ai_1 _18547_ (.B1(_11726_),
    .Y(_11727_),
    .A1(net504),
    .A2(_11724_));
 sg13g2_nand3b_1 _18548_ (.B(net118),
    .C(_11727_),
    .Y(_11728_),
    .A_N(_11720_));
 sg13g2_a21o_1 _18549_ (.A2(_11604_),
    .A1(_11596_),
    .B1(_11728_),
    .X(_11729_));
 sg13g2_buf_1 _18550_ (.A(_11729_),
    .X(_11730_));
 sg13g2_o21ai_1 _18551_ (.B1(_11730_),
    .Y(_11731_),
    .A1(_11716_),
    .A2(_11718_));
 sg13g2_or2_1 _18552_ (.X(_11732_),
    .B(_11717_),
    .A(net78));
 sg13g2_and3_1 _18553_ (.X(_11733_),
    .A(_11708_),
    .B(_11731_),
    .C(_11732_));
 sg13g2_nand2b_1 _18554_ (.Y(_11734_),
    .B(net142),
    .A_N(_11717_));
 sg13g2_nor2_1 _18555_ (.A(_11730_),
    .B(_11734_),
    .Y(_11735_));
 sg13g2_inv_1 _18556_ (.Y(_11736_),
    .A(net1105));
 sg13g2_nand4_1 _18557_ (.B(net402),
    .C(net141),
    .A(_11736_),
    .Y(_11737_),
    .D(net87));
 sg13g2_inv_1 _18558_ (.Y(_11738_),
    .A(_11715_));
 sg13g2_a21oi_1 _18559_ (.A1(_11734_),
    .A2(_11737_),
    .Y(_11739_),
    .B1(_11738_));
 sg13g2_nor3_1 _18560_ (.A(net1105),
    .B(_11707_),
    .C(_11730_),
    .Y(_11740_));
 sg13g2_nor3_1 _18561_ (.A(_11735_),
    .B(_11739_),
    .C(_11740_),
    .Y(_11741_));
 sg13g2_a21oi_1 _18562_ (.A1(_11733_),
    .A2(_11741_),
    .Y(_11742_),
    .B1(_11520_));
 sg13g2_a22oi_1 _18563_ (.Y(_11743_),
    .B1(_11532_),
    .B2(_11678_),
    .A2(_11447_),
    .A1(\cpu.ex.r_mult[14] ));
 sg13g2_nand2b_1 _18564_ (.Y(\cpu.ex.c_mult[14] ),
    .B(_11743_),
    .A_N(_11742_));
 sg13g2_nor3_1 _18565_ (.A(net1106),
    .B(_11736_),
    .C(net168),
    .Y(_11744_));
 sg13g2_xnor2_1 _18566_ (.Y(_11745_),
    .A(_11736_),
    .B(net168));
 sg13g2_a22oi_1 _18567_ (.Y(_11746_),
    .B1(_11745_),
    .B2(_11722_),
    .A2(_11744_),
    .A1(_11329_));
 sg13g2_o21ai_1 _18568_ (.B1(net445),
    .Y(_11747_),
    .A1(net1106),
    .A2(net1105));
 sg13g2_nand3_1 _18569_ (.B(net168),
    .C(_11747_),
    .A(net211),
    .Y(_11748_));
 sg13g2_o21ai_1 _18570_ (.B1(_11748_),
    .Y(_11749_),
    .A1(net444),
    .A2(_11746_));
 sg13g2_and2_1 _18571_ (.A(_11686_),
    .B(_11749_),
    .X(_11750_));
 sg13g2_nand3_1 _18572_ (.B(_11640_),
    .C(_11750_),
    .A(_11633_),
    .Y(_11751_));
 sg13g2_o21ai_1 _18573_ (.B1(net1106),
    .Y(_11752_),
    .A1(net211),
    .A2(_11690_));
 sg13g2_nand2_1 _18574_ (.Y(_11753_),
    .A(net211),
    .B(_11690_));
 sg13g2_a22oi_1 _18575_ (.Y(_11754_),
    .B1(_11752_),
    .B2(_11753_),
    .A2(net141),
    .A1(_11736_));
 sg13g2_a21oi_1 _18576_ (.A1(net1105),
    .A2(net142),
    .Y(_11755_),
    .B1(_11754_));
 sg13g2_or2_1 _18577_ (.X(_11756_),
    .B(_11755_),
    .A(net401));
 sg13g2_buf_1 _18578_ (.A(_00147_),
    .X(_11757_));
 sg13g2_nor2_1 _18579_ (.A(_11757_),
    .B(_09269_),
    .Y(_11758_));
 sg13g2_buf_1 _18580_ (.A(_11758_),
    .X(_11759_));
 sg13g2_nor2_1 _18581_ (.A(_11520_),
    .B(_11759_),
    .Y(_11760_));
 sg13g2_nand3_1 _18582_ (.B(net78),
    .C(_11760_),
    .A(net235),
    .Y(_11761_));
 sg13g2_nand2_1 _18583_ (.Y(_11762_),
    .A(_11563_),
    .B(_11759_));
 sg13g2_buf_1 _18584_ (.A(_10247_),
    .X(_11763_));
 sg13g2_nand2b_1 _18585_ (.Y(_11764_),
    .B(net210),
    .A_N(_11762_));
 sg13g2_a22oi_1 _18586_ (.Y(_11765_),
    .B1(_11761_),
    .B2(_11764_),
    .A2(_11756_),
    .A1(_11751_));
 sg13g2_and3_1 _18587_ (.X(_11766_),
    .A(_11633_),
    .B(_11640_),
    .C(_11750_));
 sg13g2_nor2_1 _18588_ (.A(net401),
    .B(_11755_),
    .Y(_11767_));
 sg13g2_nand3_1 _18589_ (.B(net78),
    .C(_11760_),
    .A(net210),
    .Y(_11768_));
 sg13g2_nor3_1 _18590_ (.A(_11766_),
    .B(_11767_),
    .C(_11768_),
    .Y(_11769_));
 sg13g2_nor4_1 _18591_ (.A(net210),
    .B(_11766_),
    .C(_11767_),
    .D(_11762_),
    .Y(_11770_));
 sg13g2_inv_1 _18592_ (.Y(_11771_),
    .A(_11757_));
 sg13g2_a22oi_1 _18593_ (.Y(_11772_),
    .B1(_11532_),
    .B2(_11771_),
    .A2(_11383_),
    .A1(\cpu.ex.r_mult[15] ));
 sg13g2_o21ai_1 _18594_ (.B1(_11772_),
    .Y(_11773_),
    .A1(net78),
    .A2(_11762_));
 sg13g2_nor4_2 _18595_ (.A(_11765_),
    .B(_11769_),
    .C(_11770_),
    .Y(_11774_),
    .D(_11773_));
 sg13g2_inv_1 _18596_ (.Y(\cpu.ex.c_mult[15] ),
    .A(_11774_));
 sg13g2_inv_1 _18597_ (.Y(_00000_),
    .A(net2));
 sg13g2_buf_2 _18598_ (.A(\cpu.qspi.r_state[13] ),
    .X(_11775_));
 sg13g2_buf_1 _18599_ (.A(net802),
    .X(_11776_));
 sg13g2_and2_1 _18600_ (.A(_11775_),
    .B(net682),
    .X(_00006_));
 sg13g2_and3_1 _18601_ (.X(_00005_),
    .A(net1122),
    .B(net682),
    .C(_09786_));
 sg13g2_inv_1 _18602_ (.Y(_11777_),
    .A(\cpu.qspi.r_state[11] ));
 sg13g2_nor2_1 _18603_ (.A(_11777_),
    .B(net711),
    .Y(_00004_));
 sg13g2_buf_1 _18604_ (.A(\cpu.qspi.r_state[10] ),
    .X(_11778_));
 sg13g2_inv_1 _18605_ (.Y(_11779_),
    .A(_11778_));
 sg13g2_nor2_1 _18606_ (.A(_11779_),
    .B(net711),
    .Y(_00003_));
 sg13g2_buf_1 _18607_ (.A(\cpu.qspi.r_state[15] ),
    .X(_11780_));
 sg13g2_and2_1 _18608_ (.A(_11780_),
    .B(net682),
    .X(_00002_));
 sg13g2_inv_1 _18609_ (.Y(_11781_),
    .A(_09790_));
 sg13g2_nor3_1 _18610_ (.A(_11781_),
    .B(net796),
    .C(net626),
    .Y(_00001_));
 sg13g2_o21ai_1 _18611_ (.B1(_09815_),
    .Y(_11782_),
    .A1(_09816_),
    .A2(_09818_));
 sg13g2_buf_1 _18612_ (.A(_11782_),
    .X(_11783_));
 sg13g2_and2_1 _18613_ (.A(_11783_),
    .B(_09823_),
    .X(_00007_));
 sg13g2_inv_2 _18614_ (.Y(_11784_),
    .A(_08336_));
 sg13g2_nand3_1 _18615_ (.B(_11212_),
    .C(_11235_),
    .A(_11071_),
    .Y(_11785_));
 sg13g2_nand2_1 _18616_ (.Y(_11786_),
    .A(_11027_),
    .B(_11090_));
 sg13g2_or4_1 _18617_ (.A(_11046_),
    .B(_11155_),
    .C(_11111_),
    .D(_11786_),
    .X(_11787_));
 sg13g2_or2_1 _18618_ (.X(_11788_),
    .B(_11184_),
    .A(_11163_));
 sg13g2_nand4_1 _18619_ (.B(_11006_),
    .C(_11788_),
    .A(_10959_),
    .Y(_11789_),
    .D(_11131_));
 sg13g2_nand2b_1 _18620_ (.Y(_11790_),
    .B(_10911_),
    .A_N(_10885_));
 sg13g2_nand3_1 _18621_ (.B(_11790_),
    .C(_10987_),
    .A(_10876_),
    .Y(_11791_));
 sg13g2_nor4_1 _18622_ (.A(_11785_),
    .B(_11787_),
    .C(_11789_),
    .D(_11791_),
    .Y(_11792_));
 sg13g2_nand2b_1 _18623_ (.Y(_11793_),
    .B(_10934_),
    .A_N(_10916_));
 sg13g2_o21ai_1 _18624_ (.B1(_11793_),
    .Y(_11794_),
    .A1(\cpu.cond[1] ),
    .A2(_11792_));
 sg13g2_xnor2_1 _18625_ (.Y(_11795_),
    .A(_11784_),
    .B(_11794_));
 sg13g2_a21oi_1 _18626_ (.A1(_00254_),
    .A2(_11795_),
    .Y(_11796_),
    .B1(_10792_));
 sg13g2_nor2_1 _18627_ (.A(\cpu.dec.jmp ),
    .B(_11796_),
    .Y(_11797_));
 sg13g2_nor2_1 _18628_ (.A(_11395_),
    .B(_11797_),
    .Y(_00053_));
 sg13g2_buf_1 _18629_ (.A(\cpu.qspi.r_state[3] ),
    .X(_11798_));
 sg13g2_and2_1 _18630_ (.A(_11798_),
    .B(net682),
    .X(_00009_));
 sg13g2_inv_1 _18631_ (.Y(_11799_),
    .A(_09795_));
 sg13g2_nor3_1 _18632_ (.A(_11799_),
    .B(net796),
    .C(_09794_),
    .Y(_00008_));
 sg13g2_buf_2 _18633_ (.A(\cpu.qspi.r_state[6] ),
    .X(_11800_));
 sg13g2_and2_1 _18634_ (.A(_11800_),
    .B(net682),
    .X(_00010_));
 sg13g2_nor2_1 _18635_ (.A(net105),
    .B(net711),
    .Y(_00052_));
 sg13g2_or2_1 _18636_ (.X(_11801_),
    .B(net1126),
    .A(_09173_));
 sg13g2_buf_1 _18637_ (.A(_11801_),
    .X(_11802_));
 sg13g2_nor3_1 _18638_ (.A(net1125),
    .B(_09239_),
    .C(_11802_),
    .Y(_11803_));
 sg13g2_a21oi_1 _18639_ (.A1(_09225_),
    .A2(_11802_),
    .Y(_11804_),
    .B1(_11803_));
 sg13g2_nand2_1 _18640_ (.Y(_11805_),
    .A(_09280_),
    .B(_11804_));
 sg13g2_inv_1 _18641_ (.Y(_11806_),
    .A(_00207_));
 sg13g2_nor3_2 _18642_ (.A(net1126),
    .B(net1125),
    .C(_11806_),
    .Y(_11807_));
 sg13g2_buf_1 _18643_ (.A(\cpu.spi.r_sel[1] ),
    .X(_11808_));
 sg13g2_buf_1 _18644_ (.A(_11808_),
    .X(_11809_));
 sg13g2_buf_1 _18645_ (.A(net1020),
    .X(_11810_));
 sg13g2_buf_1 _18646_ (.A(\cpu.spi.r_src[2] ),
    .X(_11811_));
 sg13g2_inv_1 _18647_ (.Y(_11812_),
    .A(_00263_));
 sg13g2_buf_1 _18648_ (.A(\cpu.spi.r_sel[0] ),
    .X(_11813_));
 sg13g2_buf_1 _18649_ (.A(_11813_),
    .X(_11814_));
 sg13g2_mux2_1 _18650_ (.A0(_11811_),
    .A1(_11812_),
    .S(net1019),
    .X(_11815_));
 sg13g2_buf_1 _18651_ (.A(_11813_),
    .X(_11816_));
 sg13g2_buf_1 _18652_ (.A(_11813_),
    .X(_11817_));
 sg13g2_nand2_1 _18653_ (.Y(_11818_),
    .A(net1017),
    .B(_00264_));
 sg13g2_o21ai_1 _18654_ (.B1(_11818_),
    .Y(_11819_),
    .A1(net1018),
    .A2(_11812_));
 sg13g2_nor2_1 _18655_ (.A(_11809_),
    .B(_11819_),
    .Y(_11820_));
 sg13g2_a21oi_2 _18656_ (.B1(_11820_),
    .Y(_11821_),
    .A2(_11815_),
    .A1(_11810_));
 sg13g2_nor2_1 _18657_ (.A(_11807_),
    .B(_11821_),
    .Y(_11822_));
 sg13g2_nor2_1 _18658_ (.A(net1055),
    .B(_09223_),
    .Y(_11823_));
 sg13g2_inv_2 _18659_ (.Y(_11824_),
    .A(_11808_));
 sg13g2_buf_1 _18660_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_11825_));
 sg13g2_buf_1 _18661_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_11826_));
 sg13g2_buf_1 _18662_ (.A(net1017),
    .X(_11827_));
 sg13g2_mux2_1 _18663_ (.A0(_11825_),
    .A1(_11826_),
    .S(_11827_),
    .X(_11828_));
 sg13g2_nor2_1 _18664_ (.A(_11824_),
    .B(_11813_),
    .Y(_11829_));
 sg13g2_buf_1 _18665_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_11830_));
 sg13g2_a22oi_1 _18666_ (.Y(_11831_),
    .B1(_11829_),
    .B2(_11830_),
    .A2(_11828_),
    .A1(_11824_));
 sg13g2_xnor2_1 _18667_ (.Y(_11832_),
    .A(_11823_),
    .B(_11831_));
 sg13g2_buf_1 _18668_ (.A(net1120),
    .X(_11833_));
 sg13g2_buf_1 _18669_ (.A(net1016),
    .X(_11834_));
 sg13g2_buf_1 _18670_ (.A(net779),
    .X(_11835_));
 sg13g2_nand2_1 _18671_ (.Y(_11836_),
    .A(net779),
    .B(_00264_));
 sg13g2_o21ai_1 _18672_ (.B1(_11836_),
    .Y(_11837_),
    .A1(_11835_),
    .A2(_11812_));
 sg13g2_buf_1 _18673_ (.A(_09319_),
    .X(_11838_));
 sg13g2_buf_1 _18674_ (.A(net758),
    .X(_11839_));
 sg13g2_nand3_1 _18675_ (.B(net680),
    .C(_11811_),
    .A(net874),
    .Y(_11840_));
 sg13g2_o21ai_1 _18676_ (.B1(_11840_),
    .Y(_11841_),
    .A1(net874),
    .A2(_11837_));
 sg13g2_and2_1 _18677_ (.A(_11807_),
    .B(_11841_),
    .X(_11842_));
 sg13g2_buf_1 _18678_ (.A(_11834_),
    .X(_11843_));
 sg13g2_nand2b_1 _18679_ (.Y(_11844_),
    .B(net681),
    .A_N(_11825_));
 sg13g2_o21ai_1 _18680_ (.B1(_11844_),
    .Y(_11845_),
    .A1(net681),
    .A2(_11830_));
 sg13g2_mux2_1 _18681_ (.A0(_11825_),
    .A1(_11826_),
    .S(net681),
    .X(_11846_));
 sg13g2_nor2_1 _18682_ (.A(net874),
    .B(_11846_),
    .Y(_11847_));
 sg13g2_a21oi_1 _18683_ (.A1(net757),
    .A2(_11845_),
    .Y(_11848_),
    .B1(_11847_));
 sg13g2_a22oi_1 _18684_ (.Y(_11849_),
    .B1(_11842_),
    .B2(_11848_),
    .A2(_11832_),
    .A1(_11822_));
 sg13g2_nor2_1 _18685_ (.A(_11822_),
    .B(_11842_),
    .Y(_11850_));
 sg13g2_buf_1 _18686_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_11851_));
 sg13g2_o21ai_1 _18687_ (.B1(_11851_),
    .Y(_11852_),
    .A1(_11805_),
    .A2(_11850_));
 sg13g2_o21ai_1 _18688_ (.B1(_11852_),
    .Y(_00314_),
    .A1(_11805_),
    .A2(_11849_));
 sg13g2_nor2b_1 _18689_ (.A(_11805_),
    .B_N(_11850_),
    .Y(_11853_));
 sg13g2_or3_1 _18690_ (.A(_09216_),
    .B(net1125),
    .C(_11806_),
    .X(_11854_));
 sg13g2_buf_1 _18691_ (.A(_11854_),
    .X(_11855_));
 sg13g2_and2_1 _18692_ (.A(_11807_),
    .B(_11848_),
    .X(_11856_));
 sg13g2_a21oi_1 _18693_ (.A1(net873),
    .A2(_11832_),
    .Y(_11857_),
    .B1(_11856_));
 sg13g2_buf_1 _18694_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_11858_));
 sg13g2_nor2_1 _18695_ (.A(_11858_),
    .B(_11853_),
    .Y(_11859_));
 sg13g2_a21oi_1 _18696_ (.A1(_11853_),
    .A2(_11857_),
    .Y(_00315_),
    .B1(_11859_));
 sg13g2_buf_1 _18697_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_11860_));
 sg13g2_mux2_1 _18698_ (.A0(\cpu.spi.r_out[7] ),
    .A1(net1118),
    .S(_09217_),
    .X(_11861_));
 sg13g2_nor2_1 _18699_ (.A(net1053),
    .B(_09235_),
    .Y(_11862_));
 sg13g2_inv_1 _18700_ (.Y(_11863_),
    .A(_00205_));
 sg13g2_mux2_1 _18701_ (.A0(_11863_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .S(_11813_),
    .X(_11864_));
 sg13g2_a22oi_1 _18702_ (.Y(_11865_),
    .B1(_11864_),
    .B2(_11824_),
    .A2(_11829_),
    .A1(\cpu.spi.r_mode[2][0] ));
 sg13g2_buf_1 _18703_ (.A(_11865_),
    .X(_11866_));
 sg13g2_nand2_1 _18704_ (.Y(_11867_),
    .A(net410),
    .B(_11866_));
 sg13g2_a21o_1 _18705_ (.A2(_09177_),
    .A1(_00201_),
    .B1(net1126),
    .X(_11868_));
 sg13g2_o21ai_1 _18706_ (.B1(net1126),
    .Y(_11869_),
    .A1(_09225_),
    .A2(_11866_));
 sg13g2_nand2b_1 _18707_ (.Y(_11870_),
    .B(_11869_),
    .A_N(_09173_));
 sg13g2_o21ai_1 _18708_ (.B1(_11870_),
    .Y(_11871_),
    .A1(_11867_),
    .A2(_11868_));
 sg13g2_nand2_1 _18709_ (.Y(_11872_),
    .A(_11862_),
    .B(_11871_));
 sg13g2_nor3_1 _18710_ (.A(net1127),
    .B(net1125),
    .C(_11802_),
    .Y(_11873_));
 sg13g2_nor4_1 _18711_ (.A(net507),
    .B(_09234_),
    .C(_09170_),
    .D(_11866_),
    .Y(_11874_));
 sg13g2_nor3_1 _18712_ (.A(_11872_),
    .B(_11873_),
    .C(_11874_),
    .Y(_11875_));
 sg13g2_nor2b_1 _18713_ (.A(_11821_),
    .B_N(_11875_),
    .Y(_11876_));
 sg13g2_mux2_1 _18714_ (.A0(net1102),
    .A1(_11861_),
    .S(_11876_),
    .X(_00316_));
 sg13g2_buf_1 _18715_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_11877_));
 sg13g2_nand2_1 _18716_ (.Y(_11878_),
    .A(_11821_),
    .B(_11875_));
 sg13g2_mux2_1 _18717_ (.A0(_11861_),
    .A1(net1101),
    .S(_11878_),
    .X(_00317_));
 sg13g2_buf_1 _18718_ (.A(net789),
    .X(_11879_));
 sg13g2_nand2_1 _18719_ (.Y(_11880_),
    .A(_11879_),
    .B(_09365_));
 sg13g2_buf_1 _18720_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_11881_));
 sg13g2_buf_1 _18721_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_11882_));
 sg13g2_inv_1 _18722_ (.Y(_11883_),
    .A(_11882_));
 sg13g2_buf_1 _18723_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_11884_));
 sg13g2_inv_1 _18724_ (.Y(_11885_),
    .A(_11884_));
 sg13g2_nor2_1 _18725_ (.A(_11883_),
    .B(_11885_),
    .Y(_11886_));
 sg13g2_buf_2 _18726_ (.A(_11886_),
    .X(_11887_));
 sg13g2_nand3_1 _18727_ (.B(\cpu.d_wstrobe_d ),
    .C(_11887_),
    .A(net1100),
    .Y(_11888_));
 sg13g2_buf_1 _18728_ (.A(_11888_),
    .X(_11889_));
 sg13g2_nor2_1 _18729_ (.A(_09281_),
    .B(_08339_),
    .Y(_11890_));
 sg13g2_nand2_1 _18730_ (.Y(_11891_),
    .A(_09771_),
    .B(_11890_));
 sg13g2_a21o_1 _18731_ (.A2(net617),
    .A1(_09767_),
    .B1(_11891_),
    .X(_11892_));
 sg13g2_buf_1 _18732_ (.A(_11892_),
    .X(_11893_));
 sg13g2_or2_1 _18733_ (.X(_11894_),
    .B(_11893_),
    .A(_11880_));
 sg13g2_buf_1 _18734_ (.A(_11894_),
    .X(_11895_));
 sg13g2_nand2_1 _18735_ (.Y(_11896_),
    .A(_08323_),
    .B(net902));
 sg13g2_buf_1 _18736_ (.A(_11896_),
    .X(_11897_));
 sg13g2_buf_2 _18737_ (.A(_00256_),
    .X(_11898_));
 sg13g2_o21ai_1 _18738_ (.B1(_11898_),
    .Y(_11899_),
    .A1(_08325_),
    .A2(_11897_));
 sg13g2_nor2_1 _18739_ (.A(_11895_),
    .B(_11899_),
    .Y(_11900_));
 sg13g2_buf_2 _18740_ (.A(_11900_),
    .X(_11901_));
 sg13g2_buf_1 _18741_ (.A(_11901_),
    .X(_11902_));
 sg13g2_buf_1 _18742_ (.A(uio_in[0]),
    .X(_11903_));
 sg13g2_buf_1 _18743_ (.A(_11903_),
    .X(_11904_));
 sg13g2_buf_2 _18744_ (.A(net1099),
    .X(_11905_));
 sg13g2_buf_1 _18745_ (.A(_11880_),
    .X(_11906_));
 sg13g2_buf_1 _18746_ (.A(\cpu.d_wstrobe_d ),
    .X(_11907_));
 sg13g2_buf_1 _18747_ (.A(_00257_),
    .X(_11908_));
 sg13g2_buf_1 _18748_ (.A(_11908_),
    .X(_11909_));
 sg13g2_buf_1 _18749_ (.A(_11882_),
    .X(_11910_));
 sg13g2_nor2_1 _18750_ (.A(net1013),
    .B(_11885_),
    .Y(_11911_));
 sg13g2_nand3_1 _18751_ (.B(net1014),
    .C(_11911_),
    .A(net1098),
    .Y(_11912_));
 sg13g2_buf_2 _18752_ (.A(_11912_),
    .X(_11913_));
 sg13g2_nor2_1 _18753_ (.A(net567),
    .B(_11913_),
    .Y(_11914_));
 sg13g2_buf_2 _18754_ (.A(_11914_),
    .X(_11915_));
 sg13g2_nor2b_1 _18755_ (.A(_11915_),
    .B_N(\cpu.dcache.r_data[0][0] ),
    .Y(_11916_));
 sg13g2_a21oi_1 _18756_ (.A1(net1015),
    .A2(_11915_),
    .Y(_11917_),
    .B1(_11916_));
 sg13g2_nand2_1 _18757_ (.Y(_11918_),
    .A(net899),
    .B(net65));
 sg13g2_o21ai_1 _18758_ (.B1(_11918_),
    .Y(_00318_),
    .A1(net65),
    .A2(_11917_));
 sg13g2_inv_1 _18759_ (.Y(_11919_),
    .A(_11898_));
 sg13g2_mux2_1 _18760_ (.A0(_09246_),
    .A1(net1012),
    .S(_08326_),
    .X(_11920_));
 sg13g2_nor3_1 _18761_ (.A(_11895_),
    .B(_11897_),
    .C(_11920_),
    .Y(_11921_));
 sg13g2_buf_2 _18762_ (.A(_11921_),
    .X(_11922_));
 sg13g2_buf_1 _18763_ (.A(_11922_),
    .X(_11923_));
 sg13g2_buf_1 _18764_ (.A(uio_in[2]),
    .X(_11924_));
 sg13g2_buf_1 _18765_ (.A(_11924_),
    .X(_11925_));
 sg13g2_buf_2 _18766_ (.A(net1097),
    .X(_11926_));
 sg13g2_nand3_1 _18767_ (.B(net1014),
    .C(_11887_),
    .A(net1098),
    .Y(_11927_));
 sg13g2_buf_2 _18768_ (.A(_11927_),
    .X(_11928_));
 sg13g2_nor2_1 _18769_ (.A(net567),
    .B(_11928_),
    .Y(_11929_));
 sg13g2_buf_2 _18770_ (.A(_11929_),
    .X(_11930_));
 sg13g2_nor2b_1 _18771_ (.A(_11930_),
    .B_N(\cpu.dcache.r_data[0][10] ),
    .Y(_11931_));
 sg13g2_a21oi_1 _18772_ (.A1(net1011),
    .A2(_11930_),
    .Y(_11932_),
    .B1(_11931_));
 sg13g2_nand3_1 _18773_ (.B(_08325_),
    .C(net902),
    .A(_08323_),
    .Y(_11933_));
 sg13g2_buf_4 _18774_ (.X(_11934_),
    .A(_11933_));
 sg13g2_mux2_1 _18775_ (.A0(_10099_),
    .A1(_10001_),
    .S(_11934_),
    .X(_11935_));
 sg13g2_buf_2 _18776_ (.A(_11935_),
    .X(_11936_));
 sg13g2_buf_1 _18777_ (.A(_11936_),
    .X(_11937_));
 sg13g2_nand2_1 _18778_ (.Y(_11938_),
    .A(net498),
    .B(_11922_));
 sg13g2_o21ai_1 _18779_ (.B1(_11938_),
    .Y(_00319_),
    .A1(net64),
    .A2(_11932_));
 sg13g2_buf_1 _18780_ (.A(uio_in[3]),
    .X(_11939_));
 sg13g2_buf_1 _18781_ (.A(_11939_),
    .X(_11940_));
 sg13g2_buf_2 _18782_ (.A(_11940_),
    .X(_11941_));
 sg13g2_nor2b_1 _18783_ (.A(_11930_),
    .B_N(\cpu.dcache.r_data[0][11] ),
    .Y(_11942_));
 sg13g2_a21oi_1 _18784_ (.A1(net1010),
    .A2(_11930_),
    .Y(_11943_),
    .B1(_11942_));
 sg13g2_mux2_1 _18785_ (.A0(_10105_),
    .A1(_10007_),
    .S(_11934_),
    .X(_11944_));
 sg13g2_buf_2 _18786_ (.A(_11944_),
    .X(_11945_));
 sg13g2_nand2_1 _18787_ (.Y(_11946_),
    .A(net64),
    .B(_11945_));
 sg13g2_o21ai_1 _18788_ (.B1(_11946_),
    .Y(_00320_),
    .A1(net64),
    .A2(_11943_));
 sg13g2_buf_1 _18789_ (.A(_11884_),
    .X(_11947_));
 sg13g2_nor2_1 _18790_ (.A(_11883_),
    .B(net1009),
    .Y(_11948_));
 sg13g2_nand3_1 _18791_ (.B(net1014),
    .C(_11948_),
    .A(net1098),
    .Y(_11949_));
 sg13g2_buf_2 _18792_ (.A(_11949_),
    .X(_11950_));
 sg13g2_nor2_1 _18793_ (.A(_11906_),
    .B(_11950_),
    .Y(_11951_));
 sg13g2_buf_2 _18794_ (.A(_11951_),
    .X(_11952_));
 sg13g2_nor2b_1 _18795_ (.A(_11952_),
    .B_N(\cpu.dcache.r_data[0][12] ),
    .Y(_11953_));
 sg13g2_a21oi_1 _18796_ (.A1(net1015),
    .A2(_11952_),
    .Y(_11954_),
    .B1(_11953_));
 sg13g2_mux2_1 _18797_ (.A0(_10113_),
    .A1(_10013_),
    .S(_11934_),
    .X(_11955_));
 sg13g2_buf_2 _18798_ (.A(_11955_),
    .X(_11956_));
 sg13g2_nand2_1 _18799_ (.Y(_11957_),
    .A(_11923_),
    .B(_11956_));
 sg13g2_o21ai_1 _18800_ (.B1(_11957_),
    .Y(_00321_),
    .A1(net64),
    .A2(_11954_));
 sg13g2_buf_1 _18801_ (.A(uio_in[1]),
    .X(_11958_));
 sg13g2_buf_1 _18802_ (.A(_11958_),
    .X(_11959_));
 sg13g2_buf_2 _18803_ (.A(net1095),
    .X(_11960_));
 sg13g2_nor2b_1 _18804_ (.A(_11952_),
    .B_N(\cpu.dcache.r_data[0][13] ),
    .Y(_11961_));
 sg13g2_a21oi_1 _18805_ (.A1(net1008),
    .A2(_11952_),
    .Y(_11962_),
    .B1(_11961_));
 sg13g2_mux2_1 _18806_ (.A0(_10119_),
    .A1(_10019_),
    .S(_11934_),
    .X(_11963_));
 sg13g2_buf_2 _18807_ (.A(_11963_),
    .X(_11964_));
 sg13g2_nand2_1 _18808_ (.Y(_11965_),
    .A(_11922_),
    .B(_11964_));
 sg13g2_o21ai_1 _18809_ (.B1(_11965_),
    .Y(_00322_),
    .A1(net64),
    .A2(_11962_));
 sg13g2_nor2b_1 _18810_ (.A(_11952_),
    .B_N(\cpu.dcache.r_data[0][14] ),
    .Y(_11966_));
 sg13g2_a21oi_1 _18811_ (.A1(net1011),
    .A2(_11952_),
    .Y(_11967_),
    .B1(_11966_));
 sg13g2_mux2_1 _18812_ (.A0(_10125_),
    .A1(net1119),
    .S(_11934_),
    .X(_11968_));
 sg13g2_buf_2 _18813_ (.A(_11968_),
    .X(_11969_));
 sg13g2_nand2_1 _18814_ (.Y(_11970_),
    .A(_11922_),
    .B(_11969_));
 sg13g2_o21ai_1 _18815_ (.B1(_11970_),
    .Y(_00323_),
    .A1(_11923_),
    .A2(_11967_));
 sg13g2_nor2b_1 _18816_ (.A(_11952_),
    .B_N(\cpu.dcache.r_data[0][15] ),
    .Y(_11971_));
 sg13g2_a21oi_1 _18817_ (.A1(net1010),
    .A2(_11952_),
    .Y(_11972_),
    .B1(_11971_));
 sg13g2_mux2_1 _18818_ (.A0(_10130_),
    .A1(_10033_),
    .S(_11934_),
    .X(_11973_));
 sg13g2_buf_2 _18819_ (.A(_11973_),
    .X(_11974_));
 sg13g2_nand2_1 _18820_ (.Y(_11975_),
    .A(_11922_),
    .B(_11974_));
 sg13g2_o21ai_1 _18821_ (.B1(_11975_),
    .Y(_00324_),
    .A1(net64),
    .A2(_11972_));
 sg13g2_o21ai_1 _18822_ (.B1(net797),
    .Y(_11976_),
    .A1(_08325_),
    .A2(_11897_));
 sg13g2_nor2_1 _18823_ (.A(_11895_),
    .B(_11976_),
    .Y(_11977_));
 sg13g2_buf_2 _18824_ (.A(_11977_),
    .X(_11978_));
 sg13g2_buf_1 _18825_ (.A(_11978_),
    .X(_11979_));
 sg13g2_buf_1 _18826_ (.A(net1100),
    .X(_11980_));
 sg13g2_nand3_1 _18827_ (.B(net1098),
    .C(_11911_),
    .A(net1007),
    .Y(_11981_));
 sg13g2_buf_2 _18828_ (.A(_11981_),
    .X(_11982_));
 sg13g2_nor2_1 _18829_ (.A(net567),
    .B(_11982_),
    .Y(_11983_));
 sg13g2_buf_2 _18830_ (.A(_11983_),
    .X(_11984_));
 sg13g2_nor2b_1 _18831_ (.A(_11984_),
    .B_N(\cpu.dcache.r_data[0][16] ),
    .Y(_11985_));
 sg13g2_a21oi_1 _18832_ (.A1(net1015),
    .A2(_11984_),
    .Y(_11986_),
    .B1(_11985_));
 sg13g2_nand2_1 _18833_ (.Y(_11987_),
    .A(net899),
    .B(net63));
 sg13g2_o21ai_1 _18834_ (.B1(_11987_),
    .Y(_00325_),
    .A1(net63),
    .A2(_11986_));
 sg13g2_nor2b_1 _18835_ (.A(_11984_),
    .B_N(\cpu.dcache.r_data[0][17] ),
    .Y(_11988_));
 sg13g2_a21oi_1 _18836_ (.A1(net1008),
    .A2(_11984_),
    .Y(_11989_),
    .B1(_11988_));
 sg13g2_buf_1 _18837_ (.A(net1046),
    .X(_11990_));
 sg13g2_nand2_1 _18838_ (.Y(_11991_),
    .A(net872),
    .B(_11979_));
 sg13g2_o21ai_1 _18839_ (.B1(_11991_),
    .Y(_00326_),
    .A1(_11979_),
    .A2(_11989_));
 sg13g2_nor2b_1 _18840_ (.A(_11984_),
    .B_N(\cpu.dcache.r_data[0][18] ),
    .Y(_11992_));
 sg13g2_a21oi_1 _18841_ (.A1(net1011),
    .A2(_11984_),
    .Y(_11993_),
    .B1(_11992_));
 sg13g2_buf_1 _18842_ (.A(net1045),
    .X(_11994_));
 sg13g2_nand2_1 _18843_ (.Y(_11995_),
    .A(net871),
    .B(_11978_));
 sg13g2_o21ai_1 _18844_ (.B1(_11995_),
    .Y(_00327_),
    .A1(net63),
    .A2(_11993_));
 sg13g2_inv_2 _18845_ (.Y(_11996_),
    .A(_10007_));
 sg13g2_buf_1 _18846_ (.A(_11996_),
    .X(_11997_));
 sg13g2_buf_1 _18847_ (.A(_11939_),
    .X(_11998_));
 sg13g2_mux2_1 _18848_ (.A0(\cpu.dcache.r_data[0][19] ),
    .A1(net1094),
    .S(_11984_),
    .X(_11999_));
 sg13g2_nor2_1 _18849_ (.A(_11978_),
    .B(_11999_),
    .Y(_12000_));
 sg13g2_a21oi_1 _18850_ (.A1(net870),
    .A2(net63),
    .Y(_00328_),
    .B1(_12000_));
 sg13g2_nor2b_1 _18851_ (.A(_11915_),
    .B_N(\cpu.dcache.r_data[0][1] ),
    .Y(_12001_));
 sg13g2_a21oi_1 _18852_ (.A1(net1008),
    .A2(_11915_),
    .Y(_12002_),
    .B1(_12001_));
 sg13g2_nand2_1 _18853_ (.Y(_12003_),
    .A(net872),
    .B(_11902_));
 sg13g2_o21ai_1 _18854_ (.B1(_12003_),
    .Y(_00329_),
    .A1(net65),
    .A2(_12002_));
 sg13g2_nor2_1 _18855_ (.A(net1013),
    .B(_11884_),
    .Y(_12004_));
 sg13g2_nand3_1 _18856_ (.B(net1098),
    .C(_12004_),
    .A(net1007),
    .Y(_12005_));
 sg13g2_buf_2 _18857_ (.A(_12005_),
    .X(_12006_));
 sg13g2_nor2_1 _18858_ (.A(net567),
    .B(_12006_),
    .Y(_12007_));
 sg13g2_buf_2 _18859_ (.A(_12007_),
    .X(_12008_));
 sg13g2_nor2b_1 _18860_ (.A(_12008_),
    .B_N(\cpu.dcache.r_data[0][20] ),
    .Y(_12009_));
 sg13g2_a21oi_1 _18861_ (.A1(net1015),
    .A2(_12008_),
    .Y(_12010_),
    .B1(_12009_));
 sg13g2_buf_1 _18862_ (.A(_10013_),
    .X(_12011_));
 sg13g2_nand2_1 _18863_ (.Y(_12012_),
    .A(net1006),
    .B(_11978_));
 sg13g2_o21ai_1 _18864_ (.B1(_12012_),
    .Y(_00330_),
    .A1(net63),
    .A2(_12010_));
 sg13g2_nor2b_1 _18865_ (.A(_12008_),
    .B_N(\cpu.dcache.r_data[0][21] ),
    .Y(_12013_));
 sg13g2_a21oi_1 _18866_ (.A1(net1008),
    .A2(_12008_),
    .Y(_12014_),
    .B1(_12013_));
 sg13g2_buf_1 _18867_ (.A(_10019_),
    .X(_12015_));
 sg13g2_nand2_1 _18868_ (.Y(_12016_),
    .A(net1005),
    .B(_11978_));
 sg13g2_o21ai_1 _18869_ (.B1(_12016_),
    .Y(_00331_),
    .A1(net63),
    .A2(_12014_));
 sg13g2_inv_1 _18870_ (.Y(_12017_),
    .A(net1119));
 sg13g2_buf_2 _18871_ (.A(_12017_),
    .X(_12018_));
 sg13g2_buf_1 _18872_ (.A(_12018_),
    .X(_12019_));
 sg13g2_buf_1 _18873_ (.A(_11924_),
    .X(_12020_));
 sg13g2_mux2_1 _18874_ (.A0(\cpu.dcache.r_data[0][22] ),
    .A1(net1093),
    .S(_12008_),
    .X(_12021_));
 sg13g2_nor2_1 _18875_ (.A(_11978_),
    .B(_12021_),
    .Y(_12022_));
 sg13g2_a21oi_1 _18876_ (.A1(net756),
    .A2(net63),
    .Y(_00332_),
    .B1(_12022_));
 sg13g2_inv_1 _18877_ (.Y(_12023_),
    .A(net1118));
 sg13g2_buf_2 _18878_ (.A(_12023_),
    .X(_12024_));
 sg13g2_buf_1 _18879_ (.A(_12024_),
    .X(_12025_));
 sg13g2_mux2_1 _18880_ (.A0(\cpu.dcache.r_data[0][23] ),
    .A1(net1094),
    .S(_12008_),
    .X(_12026_));
 sg13g2_nor2_1 _18881_ (.A(_11978_),
    .B(_12026_),
    .Y(_12027_));
 sg13g2_a21oi_1 _18882_ (.A1(net755),
    .A2(net63),
    .Y(_00333_),
    .B1(_12027_));
 sg13g2_or2_1 _18883_ (.X(_12028_),
    .B(net617),
    .A(net567));
 sg13g2_buf_2 _18884_ (.A(_12028_),
    .X(_12029_));
 sg13g2_buf_1 _18885_ (.A(_12029_),
    .X(_12030_));
 sg13g2_mux2_1 _18886_ (.A0(_11904_),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net400),
    .X(_12031_));
 sg13g2_mux2_1 _18887_ (.A0(_10087_),
    .A1(_09987_),
    .S(_11934_),
    .X(_12032_));
 sg13g2_buf_2 _18888_ (.A(_12032_),
    .X(_12033_));
 sg13g2_buf_1 _18889_ (.A(_12033_),
    .X(_12034_));
 sg13g2_nand2_1 _18890_ (.Y(_12035_),
    .A(_08325_),
    .B(_11898_));
 sg13g2_o21ai_1 _18891_ (.B1(_12035_),
    .Y(_12036_),
    .A1(_08325_),
    .A2(_09246_));
 sg13g2_nor3_2 _18892_ (.A(_11895_),
    .B(_11897_),
    .C(_12036_),
    .Y(_12037_));
 sg13g2_buf_1 _18893_ (.A(_12037_),
    .X(_12038_));
 sg13g2_mux2_1 _18894_ (.A0(_12031_),
    .A1(_12034_),
    .S(_12038_),
    .X(_00334_));
 sg13g2_mux2_1 _18895_ (.A0(_11959_),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(_12029_),
    .X(_12039_));
 sg13g2_mux2_1 _18896_ (.A0(_10094_),
    .A1(_09995_),
    .S(_11934_),
    .X(_12040_));
 sg13g2_buf_2 _18897_ (.A(_12040_),
    .X(_12041_));
 sg13g2_buf_1 _18898_ (.A(_12041_),
    .X(_12042_));
 sg13g2_mux2_1 _18899_ (.A0(_12039_),
    .A1(net496),
    .S(_12038_),
    .X(_00335_));
 sg13g2_buf_2 _18900_ (.A(_11924_),
    .X(_12043_));
 sg13g2_mux2_1 _18901_ (.A0(_12043_),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(_12029_),
    .X(_12044_));
 sg13g2_mux2_1 _18902_ (.A0(_12044_),
    .A1(_11937_),
    .S(net77),
    .X(_00336_));
 sg13g2_mux2_1 _18903_ (.A0(net1094),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(_12029_),
    .X(_12045_));
 sg13g2_buf_1 _18904_ (.A(_11945_),
    .X(_12046_));
 sg13g2_mux2_1 _18905_ (.A0(_12045_),
    .A1(net495),
    .S(net77),
    .X(_00337_));
 sg13g2_nand3_1 _18906_ (.B(net1098),
    .C(_11948_),
    .A(_11980_),
    .Y(_12047_));
 sg13g2_buf_2 _18907_ (.A(_12047_),
    .X(_12048_));
 sg13g2_nor2_1 _18908_ (.A(_11906_),
    .B(_12048_),
    .Y(_12049_));
 sg13g2_buf_2 _18909_ (.A(_12049_),
    .X(_12050_));
 sg13g2_nor2b_1 _18910_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][28] ),
    .Y(_12051_));
 sg13g2_a21oi_1 _18911_ (.A1(net1015),
    .A2(_12050_),
    .Y(_12052_),
    .B1(_12051_));
 sg13g2_buf_1 _18912_ (.A(_11956_),
    .X(_12053_));
 sg13g2_nand2_1 _18913_ (.Y(_12054_),
    .A(net494),
    .B(net77));
 sg13g2_o21ai_1 _18914_ (.B1(_12054_),
    .Y(_00338_),
    .A1(net77),
    .A2(_12052_));
 sg13g2_nor2b_1 _18915_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][29] ),
    .Y(_12055_));
 sg13g2_a21oi_1 _18916_ (.A1(net1008),
    .A2(_12050_),
    .Y(_12056_),
    .B1(_12055_));
 sg13g2_buf_1 _18917_ (.A(_11964_),
    .X(_12057_));
 sg13g2_nand2_1 _18918_ (.Y(_12058_),
    .A(net493),
    .B(net77));
 sg13g2_o21ai_1 _18919_ (.B1(_12058_),
    .Y(_00339_),
    .A1(net77),
    .A2(_12056_));
 sg13g2_nor2b_1 _18920_ (.A(_11915_),
    .B_N(\cpu.dcache.r_data[0][2] ),
    .Y(_12059_));
 sg13g2_a21oi_1 _18921_ (.A1(net1011),
    .A2(_11915_),
    .Y(_12060_),
    .B1(_12059_));
 sg13g2_nand2_1 _18922_ (.Y(_12061_),
    .A(_11994_),
    .B(_11901_));
 sg13g2_o21ai_1 _18923_ (.B1(_12061_),
    .Y(_00340_),
    .A1(_11902_),
    .A2(_12060_));
 sg13g2_nor2b_1 _18924_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][30] ),
    .Y(_12062_));
 sg13g2_a21oi_1 _18925_ (.A1(net1011),
    .A2(_12050_),
    .Y(_12063_),
    .B1(_12062_));
 sg13g2_buf_1 _18926_ (.A(_11969_),
    .X(_12064_));
 sg13g2_nand2_1 _18927_ (.Y(_12065_),
    .A(net492),
    .B(_12037_));
 sg13g2_o21ai_1 _18928_ (.B1(_12065_),
    .Y(_00341_),
    .A1(net77),
    .A2(_12063_));
 sg13g2_nor2b_1 _18929_ (.A(_12050_),
    .B_N(\cpu.dcache.r_data[0][31] ),
    .Y(_12066_));
 sg13g2_a21oi_1 _18930_ (.A1(net1010),
    .A2(_12050_),
    .Y(_12067_),
    .B1(_12066_));
 sg13g2_buf_1 _18931_ (.A(_11974_),
    .X(_12068_));
 sg13g2_nand2_1 _18932_ (.Y(_12069_),
    .A(net491),
    .B(_12037_));
 sg13g2_o21ai_1 _18933_ (.B1(_12069_),
    .Y(_00342_),
    .A1(net77),
    .A2(_12067_));
 sg13g2_mux2_1 _18934_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(net1094),
    .S(_11915_),
    .X(_12070_));
 sg13g2_nor2_1 _18935_ (.A(_11901_),
    .B(_12070_),
    .Y(_12071_));
 sg13g2_a21oi_1 _18936_ (.A1(net870),
    .A2(net65),
    .Y(_00343_),
    .B1(_12071_));
 sg13g2_nand3_1 _18937_ (.B(net1014),
    .C(_12004_),
    .A(net1098),
    .Y(_12072_));
 sg13g2_buf_2 _18938_ (.A(_12072_),
    .X(_12073_));
 sg13g2_nor2_1 _18939_ (.A(net567),
    .B(_12073_),
    .Y(_12074_));
 sg13g2_buf_2 _18940_ (.A(_12074_),
    .X(_12075_));
 sg13g2_nor2b_1 _18941_ (.A(_12075_),
    .B_N(\cpu.dcache.r_data[0][4] ),
    .Y(_12076_));
 sg13g2_a21oi_1 _18942_ (.A1(net1015),
    .A2(_12075_),
    .Y(_12077_),
    .B1(_12076_));
 sg13g2_buf_1 _18943_ (.A(_10013_),
    .X(_12078_));
 sg13g2_nand2_1 _18944_ (.Y(_12079_),
    .A(_12078_),
    .B(_11901_));
 sg13g2_o21ai_1 _18945_ (.B1(_12079_),
    .Y(_00344_),
    .A1(net65),
    .A2(_12077_));
 sg13g2_nor2b_1 _18946_ (.A(_12075_),
    .B_N(\cpu.dcache.r_data[0][5] ),
    .Y(_12080_));
 sg13g2_a21oi_1 _18947_ (.A1(net1008),
    .A2(_12075_),
    .Y(_12081_),
    .B1(_12080_));
 sg13g2_buf_1 _18948_ (.A(_10019_),
    .X(_12082_));
 sg13g2_nand2_1 _18949_ (.Y(_12083_),
    .A(_12082_),
    .B(_11901_));
 sg13g2_o21ai_1 _18950_ (.B1(_12083_),
    .Y(_00345_),
    .A1(net65),
    .A2(_12081_));
 sg13g2_mux2_1 _18951_ (.A0(\cpu.dcache.r_data[0][6] ),
    .A1(net1093),
    .S(_12075_),
    .X(_12084_));
 sg13g2_nor2_1 _18952_ (.A(_11901_),
    .B(_12084_),
    .Y(_12085_));
 sg13g2_a21oi_1 _18953_ (.A1(_12019_),
    .A2(net65),
    .Y(_00346_),
    .B1(_12085_));
 sg13g2_buf_1 _18954_ (.A(net1096),
    .X(_12086_));
 sg13g2_mux2_1 _18955_ (.A0(\cpu.dcache.r_data[0][7] ),
    .A1(net1002),
    .S(_12075_),
    .X(_12087_));
 sg13g2_nor2_1 _18956_ (.A(_11901_),
    .B(_12087_),
    .Y(_12088_));
 sg13g2_a21oi_1 _18957_ (.A1(_12025_),
    .A2(net65),
    .Y(_00347_),
    .B1(_12088_));
 sg13g2_buf_1 _18958_ (.A(net1099),
    .X(_12089_));
 sg13g2_nor2b_1 _18959_ (.A(_11930_),
    .B_N(\cpu.dcache.r_data[0][8] ),
    .Y(_12090_));
 sg13g2_a21oi_1 _18960_ (.A1(net1001),
    .A2(_11930_),
    .Y(_12091_),
    .B1(_12090_));
 sg13g2_nand2_1 _18961_ (.Y(_12092_),
    .A(_11922_),
    .B(_12033_));
 sg13g2_o21ai_1 _18962_ (.B1(_12092_),
    .Y(_00348_),
    .A1(net64),
    .A2(_12091_));
 sg13g2_buf_1 _18963_ (.A(net1095),
    .X(_12093_));
 sg13g2_nor2b_1 _18964_ (.A(_11930_),
    .B_N(\cpu.dcache.r_data[0][9] ),
    .Y(_12094_));
 sg13g2_a21oi_1 _18965_ (.A1(net1000),
    .A2(_11930_),
    .Y(_12095_),
    .B1(_12094_));
 sg13g2_nand2_1 _18966_ (.Y(_12096_),
    .A(_11922_),
    .B(_12041_));
 sg13g2_o21ai_1 _18967_ (.B1(_12096_),
    .Y(_00349_),
    .A1(net64),
    .A2(_12095_));
 sg13g2_buf_1 _18968_ (.A(net572),
    .X(_12097_));
 sg13g2_or2_1 _18969_ (.X(_12098_),
    .B(_11899_),
    .A(_11893_));
 sg13g2_buf_2 _18970_ (.A(_12098_),
    .X(_12099_));
 sg13g2_nor2_1 _18971_ (.A(net490),
    .B(_12099_),
    .Y(_12100_));
 sg13g2_buf_2 _18972_ (.A(_12100_),
    .X(_12101_));
 sg13g2_buf_1 _18973_ (.A(_12101_),
    .X(_12102_));
 sg13g2_nor2_1 _18974_ (.A(net572),
    .B(_11913_),
    .Y(_12103_));
 sg13g2_buf_2 _18975_ (.A(_12103_),
    .X(_12104_));
 sg13g2_nor2b_1 _18976_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[1][0] ),
    .Y(_12105_));
 sg13g2_a21oi_1 _18977_ (.A1(net1001),
    .A2(_12104_),
    .Y(_12106_),
    .B1(_12105_));
 sg13g2_nand2_1 _18978_ (.Y(_12107_),
    .A(net899),
    .B(net62));
 sg13g2_o21ai_1 _18979_ (.B1(_12107_),
    .Y(_00350_),
    .A1(_12102_),
    .A2(_12106_));
 sg13g2_or3_1 _18980_ (.A(_11893_),
    .B(_11897_),
    .C(_11920_),
    .X(_12108_));
 sg13g2_buf_2 _18981_ (.A(_12108_),
    .X(_12109_));
 sg13g2_nor2_1 _18982_ (.A(net490),
    .B(_12109_),
    .Y(_12110_));
 sg13g2_buf_2 _18983_ (.A(_12110_),
    .X(_12111_));
 sg13g2_buf_1 _18984_ (.A(_12111_),
    .X(_12112_));
 sg13g2_nor2_1 _18985_ (.A(net490),
    .B(_11928_),
    .Y(_12113_));
 sg13g2_buf_2 _18986_ (.A(_12113_),
    .X(_12114_));
 sg13g2_nor2b_1 _18987_ (.A(_12114_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12115_));
 sg13g2_a21oi_1 _18988_ (.A1(net1011),
    .A2(_12114_),
    .Y(_12116_),
    .B1(_12115_));
 sg13g2_nand2_1 _18989_ (.Y(_12117_),
    .A(net498),
    .B(net61));
 sg13g2_o21ai_1 _18990_ (.B1(_12117_),
    .Y(_00351_),
    .A1(net61),
    .A2(_12116_));
 sg13g2_nor2b_1 _18991_ (.A(_12114_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12118_));
 sg13g2_a21oi_1 _18992_ (.A1(net1010),
    .A2(_12114_),
    .Y(_12119_),
    .B1(_12118_));
 sg13g2_nand2_1 _18993_ (.Y(_12120_),
    .A(net495),
    .B(net61));
 sg13g2_o21ai_1 _18994_ (.B1(_12120_),
    .Y(_00352_),
    .A1(net61),
    .A2(_12119_));
 sg13g2_nor2_1 _18995_ (.A(net490),
    .B(_11950_),
    .Y(_12121_));
 sg13g2_buf_2 _18996_ (.A(_12121_),
    .X(_12122_));
 sg13g2_nor2b_1 _18997_ (.A(_12122_),
    .B_N(\cpu.dcache.r_data[1][12] ),
    .Y(_12123_));
 sg13g2_a21oi_1 _18998_ (.A1(net1001),
    .A2(_12122_),
    .Y(_12124_),
    .B1(_12123_));
 sg13g2_nand2_1 _18999_ (.Y(_12125_),
    .A(net494),
    .B(_12111_));
 sg13g2_o21ai_1 _19000_ (.B1(_12125_),
    .Y(_00353_),
    .A1(net61),
    .A2(_12124_));
 sg13g2_nor2b_1 _19001_ (.A(_12122_),
    .B_N(\cpu.dcache.r_data[1][13] ),
    .Y(_12126_));
 sg13g2_a21oi_1 _19002_ (.A1(net1000),
    .A2(_12122_),
    .Y(_12127_),
    .B1(_12126_));
 sg13g2_nand2_1 _19003_ (.Y(_12128_),
    .A(net493),
    .B(_12111_));
 sg13g2_o21ai_1 _19004_ (.B1(_12128_),
    .Y(_00354_),
    .A1(_12112_),
    .A2(_12127_));
 sg13g2_buf_1 _19005_ (.A(net1097),
    .X(_12129_));
 sg13g2_nor2b_1 _19006_ (.A(_12122_),
    .B_N(\cpu.dcache.r_data[1][14] ),
    .Y(_12130_));
 sg13g2_a21oi_1 _19007_ (.A1(net999),
    .A2(_12122_),
    .Y(_12131_),
    .B1(_12130_));
 sg13g2_nand2_1 _19008_ (.Y(_12132_),
    .A(net492),
    .B(_12111_));
 sg13g2_o21ai_1 _19009_ (.B1(_12132_),
    .Y(_00355_),
    .A1(_12112_),
    .A2(_12131_));
 sg13g2_nor2b_1 _19010_ (.A(_12122_),
    .B_N(\cpu.dcache.r_data[1][15] ),
    .Y(_12133_));
 sg13g2_a21oi_1 _19011_ (.A1(net1010),
    .A2(_12122_),
    .Y(_12134_),
    .B1(_12133_));
 sg13g2_nand2_1 _19012_ (.Y(_12135_),
    .A(net491),
    .B(_12111_));
 sg13g2_o21ai_1 _19013_ (.B1(_12135_),
    .Y(_00356_),
    .A1(net61),
    .A2(_12134_));
 sg13g2_or2_1 _19014_ (.X(_12136_),
    .B(_11976_),
    .A(_11893_));
 sg13g2_buf_2 _19015_ (.A(_12136_),
    .X(_12137_));
 sg13g2_nor2_1 _19016_ (.A(net490),
    .B(_12137_),
    .Y(_12138_));
 sg13g2_buf_2 _19017_ (.A(_12138_),
    .X(_12139_));
 sg13g2_buf_1 _19018_ (.A(_12139_),
    .X(_12140_));
 sg13g2_nor2_1 _19019_ (.A(net572),
    .B(_11982_),
    .Y(_12141_));
 sg13g2_buf_2 _19020_ (.A(_12141_),
    .X(_12142_));
 sg13g2_nor2b_1 _19021_ (.A(_12142_),
    .B_N(\cpu.dcache.r_data[1][16] ),
    .Y(_12143_));
 sg13g2_a21oi_1 _19022_ (.A1(net1001),
    .A2(_12142_),
    .Y(_12144_),
    .B1(_12143_));
 sg13g2_nand2_1 _19023_ (.Y(_12145_),
    .A(_10049_),
    .B(net60));
 sg13g2_o21ai_1 _19024_ (.B1(_12145_),
    .Y(_00357_),
    .A1(net60),
    .A2(_12144_));
 sg13g2_nor2b_1 _19025_ (.A(_12142_),
    .B_N(\cpu.dcache.r_data[1][17] ),
    .Y(_12146_));
 sg13g2_a21oi_1 _19026_ (.A1(net1000),
    .A2(_12142_),
    .Y(_12147_),
    .B1(_12146_));
 sg13g2_nand2_1 _19027_ (.Y(_12148_),
    .A(net872),
    .B(_12140_));
 sg13g2_o21ai_1 _19028_ (.B1(_12148_),
    .Y(_00358_),
    .A1(_12140_),
    .A2(_12147_));
 sg13g2_nor2b_1 _19029_ (.A(_12142_),
    .B_N(\cpu.dcache.r_data[1][18] ),
    .Y(_12149_));
 sg13g2_a21oi_1 _19030_ (.A1(net999),
    .A2(_12142_),
    .Y(_12150_),
    .B1(_12149_));
 sg13g2_nand2_1 _19031_ (.Y(_12151_),
    .A(net871),
    .B(_12139_));
 sg13g2_o21ai_1 _19032_ (.B1(_12151_),
    .Y(_00359_),
    .A1(net60),
    .A2(_12150_));
 sg13g2_mux2_1 _19033_ (.A0(\cpu.dcache.r_data[1][19] ),
    .A1(net1002),
    .S(_12142_),
    .X(_12152_));
 sg13g2_nor2_1 _19034_ (.A(_12139_),
    .B(_12152_),
    .Y(_12153_));
 sg13g2_a21oi_1 _19035_ (.A1(net870),
    .A2(net60),
    .Y(_00360_),
    .B1(_12153_));
 sg13g2_nor2b_1 _19036_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[1][1] ),
    .Y(_12154_));
 sg13g2_a21oi_1 _19037_ (.A1(net1000),
    .A2(_12104_),
    .Y(_12155_),
    .B1(_12154_));
 sg13g2_nand2_1 _19038_ (.Y(_12156_),
    .A(_11990_),
    .B(_12102_));
 sg13g2_o21ai_1 _19039_ (.B1(_12156_),
    .Y(_00361_),
    .A1(net62),
    .A2(_12155_));
 sg13g2_nor2_1 _19040_ (.A(net490),
    .B(_12006_),
    .Y(_12157_));
 sg13g2_buf_2 _19041_ (.A(_12157_),
    .X(_12158_));
 sg13g2_nor2b_1 _19042_ (.A(_12158_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_12159_));
 sg13g2_a21oi_1 _19043_ (.A1(net1001),
    .A2(_12158_),
    .Y(_12160_),
    .B1(_12159_));
 sg13g2_nand2_1 _19044_ (.Y(_12161_),
    .A(net1004),
    .B(_12139_));
 sg13g2_o21ai_1 _19045_ (.B1(_12161_),
    .Y(_00362_),
    .A1(net60),
    .A2(_12160_));
 sg13g2_nor2b_1 _19046_ (.A(_12158_),
    .B_N(\cpu.dcache.r_data[1][21] ),
    .Y(_12162_));
 sg13g2_a21oi_1 _19047_ (.A1(net1000),
    .A2(_12158_),
    .Y(_12163_),
    .B1(_12162_));
 sg13g2_nand2_1 _19048_ (.Y(_12164_),
    .A(net1003),
    .B(_12139_));
 sg13g2_o21ai_1 _19049_ (.B1(_12164_),
    .Y(_00363_),
    .A1(net60),
    .A2(_12163_));
 sg13g2_mux2_1 _19050_ (.A0(\cpu.dcache.r_data[1][22] ),
    .A1(net1093),
    .S(_12158_),
    .X(_12165_));
 sg13g2_nor2_1 _19051_ (.A(_12139_),
    .B(_12165_),
    .Y(_12166_));
 sg13g2_a21oi_1 _19052_ (.A1(net756),
    .A2(net60),
    .Y(_00364_),
    .B1(_12166_));
 sg13g2_mux2_1 _19053_ (.A0(\cpu.dcache.r_data[1][23] ),
    .A1(net1002),
    .S(_12158_),
    .X(_12167_));
 sg13g2_nor2_1 _19054_ (.A(_12139_),
    .B(_12167_),
    .Y(_12168_));
 sg13g2_a21oi_1 _19055_ (.A1(net755),
    .A2(net60),
    .Y(_00365_),
    .B1(_12168_));
 sg13g2_or3_1 _19056_ (.A(_11893_),
    .B(_11897_),
    .C(_12036_),
    .X(_12169_));
 sg13g2_buf_2 _19057_ (.A(_12169_),
    .X(_12170_));
 sg13g2_nor2_1 _19058_ (.A(_12097_),
    .B(_12170_),
    .Y(_12171_));
 sg13g2_buf_2 _19059_ (.A(_12171_),
    .X(_12172_));
 sg13g2_buf_1 _19060_ (.A(_12172_),
    .X(_12173_));
 sg13g2_nor2_1 _19061_ (.A(_09593_),
    .B(_11889_),
    .Y(_12174_));
 sg13g2_buf_1 _19062_ (.A(_12174_),
    .X(_12175_));
 sg13g2_buf_1 _19063_ (.A(_12175_),
    .X(_12176_));
 sg13g2_nor2b_1 _19064_ (.A(net399),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12177_));
 sg13g2_a21oi_1 _19065_ (.A1(net1001),
    .A2(net399),
    .Y(_12178_),
    .B1(_12177_));
 sg13g2_nand2_1 _19066_ (.Y(_12179_),
    .A(net497),
    .B(_12173_));
 sg13g2_o21ai_1 _19067_ (.B1(_12179_),
    .Y(_00366_),
    .A1(net59),
    .A2(_12178_));
 sg13g2_nor2b_1 _19068_ (.A(net399),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12180_));
 sg13g2_a21oi_1 _19069_ (.A1(net1000),
    .A2(net399),
    .Y(_12181_),
    .B1(_12180_));
 sg13g2_nand2_1 _19070_ (.Y(_12182_),
    .A(net496),
    .B(net59));
 sg13g2_o21ai_1 _19071_ (.B1(_12182_),
    .Y(_00367_),
    .A1(_12173_),
    .A2(_12181_));
 sg13g2_nor2b_1 _19072_ (.A(net399),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12183_));
 sg13g2_a21oi_1 _19073_ (.A1(net999),
    .A2(net399),
    .Y(_12184_),
    .B1(_12183_));
 sg13g2_nand2_1 _19074_ (.Y(_12185_),
    .A(net498),
    .B(_12172_));
 sg13g2_o21ai_1 _19075_ (.B1(_12185_),
    .Y(_00368_),
    .A1(net59),
    .A2(_12184_));
 sg13g2_nor2b_1 _19076_ (.A(_12175_),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12186_));
 sg13g2_a21oi_1 _19077_ (.A1(net1010),
    .A2(net399),
    .Y(_12187_),
    .B1(_12186_));
 sg13g2_nand2_1 _19078_ (.Y(_12188_),
    .A(_12046_),
    .B(_12172_));
 sg13g2_o21ai_1 _19079_ (.B1(_12188_),
    .Y(_00369_),
    .A1(net59),
    .A2(_12187_));
 sg13g2_nor2_1 _19080_ (.A(_12097_),
    .B(_12048_),
    .Y(_12189_));
 sg13g2_buf_2 _19081_ (.A(_12189_),
    .X(_12190_));
 sg13g2_nor2b_1 _19082_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[1][28] ),
    .Y(_12191_));
 sg13g2_a21oi_1 _19083_ (.A1(_12089_),
    .A2(_12190_),
    .Y(_12192_),
    .B1(_12191_));
 sg13g2_nand2_1 _19084_ (.Y(_12193_),
    .A(_12053_),
    .B(_12172_));
 sg13g2_o21ai_1 _19085_ (.B1(_12193_),
    .Y(_00370_),
    .A1(net59),
    .A2(_12192_));
 sg13g2_nor2b_1 _19086_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[1][29] ),
    .Y(_12194_));
 sg13g2_a21oi_1 _19087_ (.A1(_12093_),
    .A2(_12190_),
    .Y(_12195_),
    .B1(_12194_));
 sg13g2_nand2_1 _19088_ (.Y(_12196_),
    .A(_12057_),
    .B(_12172_));
 sg13g2_o21ai_1 _19089_ (.B1(_12196_),
    .Y(_00371_),
    .A1(net59),
    .A2(_12195_));
 sg13g2_nor2b_1 _19090_ (.A(_12104_),
    .B_N(\cpu.dcache.r_data[1][2] ),
    .Y(_12197_));
 sg13g2_a21oi_1 _19091_ (.A1(net999),
    .A2(_12104_),
    .Y(_12198_),
    .B1(_12197_));
 sg13g2_nand2_1 _19092_ (.Y(_12199_),
    .A(_11994_),
    .B(_12101_));
 sg13g2_o21ai_1 _19093_ (.B1(_12199_),
    .Y(_00372_),
    .A1(net62),
    .A2(_12198_));
 sg13g2_nor2b_1 _19094_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[1][30] ),
    .Y(_12200_));
 sg13g2_a21oi_1 _19095_ (.A1(_12129_),
    .A2(_12190_),
    .Y(_12201_),
    .B1(_12200_));
 sg13g2_nand2_1 _19096_ (.Y(_12202_),
    .A(_12064_),
    .B(_12172_));
 sg13g2_o21ai_1 _19097_ (.B1(_12202_),
    .Y(_00373_),
    .A1(net59),
    .A2(_12201_));
 sg13g2_buf_1 _19098_ (.A(net1096),
    .X(_12203_));
 sg13g2_nor2b_1 _19099_ (.A(_12190_),
    .B_N(\cpu.dcache.r_data[1][31] ),
    .Y(_12204_));
 sg13g2_a21oi_1 _19100_ (.A1(net998),
    .A2(_12190_),
    .Y(_12205_),
    .B1(_12204_));
 sg13g2_nand2_1 _19101_ (.Y(_12206_),
    .A(_12068_),
    .B(_12172_));
 sg13g2_o21ai_1 _19102_ (.B1(_12206_),
    .Y(_00374_),
    .A1(net59),
    .A2(_12205_));
 sg13g2_mux2_1 _19103_ (.A0(\cpu.dcache.r_data[1][3] ),
    .A1(_12086_),
    .S(_12104_),
    .X(_12207_));
 sg13g2_nor2_1 _19104_ (.A(_12101_),
    .B(_12207_),
    .Y(_12208_));
 sg13g2_a21oi_1 _19105_ (.A1(net870),
    .A2(net62),
    .Y(_00375_),
    .B1(_12208_));
 sg13g2_nor2_1 _19106_ (.A(net490),
    .B(_12073_),
    .Y(_12209_));
 sg13g2_buf_2 _19107_ (.A(_12209_),
    .X(_12210_));
 sg13g2_nor2b_1 _19108_ (.A(_12210_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12211_));
 sg13g2_a21oi_1 _19109_ (.A1(net1001),
    .A2(_12210_),
    .Y(_12212_),
    .B1(_12211_));
 sg13g2_nand2_1 _19110_ (.Y(_12213_),
    .A(net1004),
    .B(_12101_));
 sg13g2_o21ai_1 _19111_ (.B1(_12213_),
    .Y(_00376_),
    .A1(net62),
    .A2(_12212_));
 sg13g2_nor2b_1 _19112_ (.A(_12210_),
    .B_N(\cpu.dcache.r_data[1][5] ),
    .Y(_12214_));
 sg13g2_a21oi_1 _19113_ (.A1(net1000),
    .A2(_12210_),
    .Y(_12215_),
    .B1(_12214_));
 sg13g2_nand2_1 _19114_ (.Y(_12216_),
    .A(net1003),
    .B(_12101_));
 sg13g2_o21ai_1 _19115_ (.B1(_12216_),
    .Y(_00377_),
    .A1(net62),
    .A2(_12215_));
 sg13g2_mux2_1 _19116_ (.A0(\cpu.dcache.r_data[1][6] ),
    .A1(net1093),
    .S(_12210_),
    .X(_12217_));
 sg13g2_nor2_1 _19117_ (.A(_12101_),
    .B(_12217_),
    .Y(_12218_));
 sg13g2_a21oi_1 _19118_ (.A1(net756),
    .A2(net62),
    .Y(_00378_),
    .B1(_12218_));
 sg13g2_mux2_1 _19119_ (.A0(\cpu.dcache.r_data[1][7] ),
    .A1(_12086_),
    .S(_12210_),
    .X(_12219_));
 sg13g2_nor2_1 _19120_ (.A(_12101_),
    .B(_12219_),
    .Y(_12220_));
 sg13g2_a21oi_1 _19121_ (.A1(net755),
    .A2(net62),
    .Y(_00379_),
    .B1(_12220_));
 sg13g2_nor2b_1 _19122_ (.A(_12114_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12221_));
 sg13g2_a21oi_1 _19123_ (.A1(_12089_),
    .A2(_12114_),
    .Y(_12222_),
    .B1(_12221_));
 sg13g2_nand2_1 _19124_ (.Y(_12223_),
    .A(net497),
    .B(_12111_));
 sg13g2_o21ai_1 _19125_ (.B1(_12223_),
    .Y(_00380_),
    .A1(net61),
    .A2(_12222_));
 sg13g2_nor2b_1 _19126_ (.A(_12114_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12224_));
 sg13g2_a21oi_1 _19127_ (.A1(_12093_),
    .A2(_12114_),
    .Y(_12225_),
    .B1(_12224_));
 sg13g2_nand2_1 _19128_ (.Y(_12226_),
    .A(net496),
    .B(_12111_));
 sg13g2_o21ai_1 _19129_ (.B1(_12226_),
    .Y(_00381_),
    .A1(net61),
    .A2(_12225_));
 sg13g2_buf_1 _19130_ (.A(_09390_),
    .X(_12227_));
 sg13g2_nor2_1 _19131_ (.A(net678),
    .B(_12099_),
    .Y(_12228_));
 sg13g2_buf_1 _19132_ (.A(_12228_),
    .X(_12229_));
 sg13g2_buf_1 _19133_ (.A(_12229_),
    .X(_12230_));
 sg13g2_nor2_1 _19134_ (.A(_09390_),
    .B(_11913_),
    .Y(_12231_));
 sg13g2_buf_2 _19135_ (.A(_12231_),
    .X(_12232_));
 sg13g2_nor2b_1 _19136_ (.A(_12232_),
    .B_N(\cpu.dcache.r_data[2][0] ),
    .Y(_12233_));
 sg13g2_a21oi_1 _19137_ (.A1(net1001),
    .A2(_12232_),
    .Y(_12234_),
    .B1(_12233_));
 sg13g2_nand2_1 _19138_ (.Y(_12235_),
    .A(_10049_),
    .B(net58));
 sg13g2_o21ai_1 _19139_ (.B1(_12235_),
    .Y(_00382_),
    .A1(net58),
    .A2(_12234_));
 sg13g2_nor2_1 _19140_ (.A(net678),
    .B(_12109_),
    .Y(_12236_));
 sg13g2_buf_2 _19141_ (.A(_12236_),
    .X(_12237_));
 sg13g2_buf_1 _19142_ (.A(_12237_),
    .X(_12238_));
 sg13g2_nor2_1 _19143_ (.A(net678),
    .B(_11928_),
    .Y(_12239_));
 sg13g2_buf_2 _19144_ (.A(_12239_),
    .X(_12240_));
 sg13g2_nor2b_1 _19145_ (.A(_12240_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12241_));
 sg13g2_a21oi_1 _19146_ (.A1(net999),
    .A2(_12240_),
    .Y(_12242_),
    .B1(_12241_));
 sg13g2_nand2_1 _19147_ (.Y(_12243_),
    .A(net498),
    .B(net57));
 sg13g2_o21ai_1 _19148_ (.B1(_12243_),
    .Y(_00383_),
    .A1(net57),
    .A2(_12242_));
 sg13g2_nor2b_1 _19149_ (.A(_12240_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12244_));
 sg13g2_a21oi_1 _19150_ (.A1(net998),
    .A2(_12240_),
    .Y(_12245_),
    .B1(_12244_));
 sg13g2_nand2_1 _19151_ (.Y(_12246_),
    .A(net495),
    .B(net57));
 sg13g2_o21ai_1 _19152_ (.B1(_12246_),
    .Y(_00384_),
    .A1(net57),
    .A2(_12245_));
 sg13g2_buf_1 _19153_ (.A(net1099),
    .X(_12247_));
 sg13g2_nor2_1 _19154_ (.A(net678),
    .B(_11950_),
    .Y(_12248_));
 sg13g2_buf_2 _19155_ (.A(_12248_),
    .X(_12249_));
 sg13g2_nor2b_1 _19156_ (.A(_12249_),
    .B_N(\cpu.dcache.r_data[2][12] ),
    .Y(_12250_));
 sg13g2_a21oi_1 _19157_ (.A1(net997),
    .A2(_12249_),
    .Y(_12251_),
    .B1(_12250_));
 sg13g2_nand2_1 _19158_ (.Y(_12252_),
    .A(net494),
    .B(_12237_));
 sg13g2_o21ai_1 _19159_ (.B1(_12252_),
    .Y(_00385_),
    .A1(net57),
    .A2(_12251_));
 sg13g2_nor2b_1 _19160_ (.A(_12249_),
    .B_N(\cpu.dcache.r_data[2][13] ),
    .Y(_12253_));
 sg13g2_a21oi_1 _19161_ (.A1(net1000),
    .A2(_12249_),
    .Y(_12254_),
    .B1(_12253_));
 sg13g2_nand2_1 _19162_ (.Y(_12255_),
    .A(net493),
    .B(_12237_));
 sg13g2_o21ai_1 _19163_ (.B1(_12255_),
    .Y(_00386_),
    .A1(net57),
    .A2(_12254_));
 sg13g2_nor2b_1 _19164_ (.A(_12249_),
    .B_N(\cpu.dcache.r_data[2][14] ),
    .Y(_12256_));
 sg13g2_a21oi_1 _19165_ (.A1(net999),
    .A2(_12249_),
    .Y(_12257_),
    .B1(_12256_));
 sg13g2_nand2_1 _19166_ (.Y(_12258_),
    .A(net492),
    .B(_12237_));
 sg13g2_o21ai_1 _19167_ (.B1(_12258_),
    .Y(_00387_),
    .A1(net57),
    .A2(_12257_));
 sg13g2_nor2b_1 _19168_ (.A(_12249_),
    .B_N(\cpu.dcache.r_data[2][15] ),
    .Y(_12259_));
 sg13g2_a21oi_1 _19169_ (.A1(net998),
    .A2(_12249_),
    .Y(_12260_),
    .B1(_12259_));
 sg13g2_nand2_1 _19170_ (.Y(_12261_),
    .A(net491),
    .B(_12237_));
 sg13g2_o21ai_1 _19171_ (.B1(_12261_),
    .Y(_00388_),
    .A1(net57),
    .A2(_12260_));
 sg13g2_nor2_1 _19172_ (.A(net678),
    .B(_12137_),
    .Y(_12262_));
 sg13g2_buf_1 _19173_ (.A(_12262_),
    .X(_12263_));
 sg13g2_buf_1 _19174_ (.A(_12263_),
    .X(_12264_));
 sg13g2_nor2_1 _19175_ (.A(_09390_),
    .B(_11982_),
    .Y(_12265_));
 sg13g2_buf_2 _19176_ (.A(_12265_),
    .X(_12266_));
 sg13g2_nor2b_1 _19177_ (.A(_12266_),
    .B_N(\cpu.dcache.r_data[2][16] ),
    .Y(_12267_));
 sg13g2_a21oi_1 _19178_ (.A1(net997),
    .A2(_12266_),
    .Y(_12268_),
    .B1(_12267_));
 sg13g2_buf_1 _19179_ (.A(net1047),
    .X(_12269_));
 sg13g2_nand2_1 _19180_ (.Y(_12270_),
    .A(net869),
    .B(net56));
 sg13g2_o21ai_1 _19181_ (.B1(_12270_),
    .Y(_00389_),
    .A1(net56),
    .A2(_12268_));
 sg13g2_buf_1 _19182_ (.A(net1095),
    .X(_12271_));
 sg13g2_nor2b_1 _19183_ (.A(_12266_),
    .B_N(\cpu.dcache.r_data[2][17] ),
    .Y(_12272_));
 sg13g2_a21oi_1 _19184_ (.A1(net996),
    .A2(_12266_),
    .Y(_12273_),
    .B1(_12272_));
 sg13g2_nand2_1 _19185_ (.Y(_12274_),
    .A(_11990_),
    .B(net56));
 sg13g2_o21ai_1 _19186_ (.B1(_12274_),
    .Y(_00390_),
    .A1(_12264_),
    .A2(_12273_));
 sg13g2_nor2b_1 _19187_ (.A(_12266_),
    .B_N(\cpu.dcache.r_data[2][18] ),
    .Y(_12275_));
 sg13g2_a21oi_1 _19188_ (.A1(net999),
    .A2(_12266_),
    .Y(_12276_),
    .B1(_12275_));
 sg13g2_nand2_1 _19189_ (.Y(_12277_),
    .A(net871),
    .B(_12263_));
 sg13g2_o21ai_1 _19190_ (.B1(_12277_),
    .Y(_00391_),
    .A1(_12264_),
    .A2(_12276_));
 sg13g2_mux2_1 _19191_ (.A0(\cpu.dcache.r_data[2][19] ),
    .A1(net1002),
    .S(_12266_),
    .X(_12278_));
 sg13g2_nor2_1 _19192_ (.A(_12263_),
    .B(_12278_),
    .Y(_12279_));
 sg13g2_a21oi_1 _19193_ (.A1(net870),
    .A2(net56),
    .Y(_00392_),
    .B1(_12279_));
 sg13g2_nor2b_1 _19194_ (.A(_12232_),
    .B_N(\cpu.dcache.r_data[2][1] ),
    .Y(_12280_));
 sg13g2_a21oi_1 _19195_ (.A1(net996),
    .A2(_12232_),
    .Y(_12281_),
    .B1(_12280_));
 sg13g2_buf_1 _19196_ (.A(_09996_),
    .X(_12282_));
 sg13g2_nand2_1 _19197_ (.Y(_12283_),
    .A(net868),
    .B(net58));
 sg13g2_o21ai_1 _19198_ (.B1(_12283_),
    .Y(_00393_),
    .A1(_12230_),
    .A2(_12281_));
 sg13g2_nor2_1 _19199_ (.A(net678),
    .B(_12006_),
    .Y(_12284_));
 sg13g2_buf_2 _19200_ (.A(_12284_),
    .X(_12285_));
 sg13g2_nor2b_1 _19201_ (.A(_12285_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12286_));
 sg13g2_a21oi_1 _19202_ (.A1(net997),
    .A2(_12285_),
    .Y(_12287_),
    .B1(_12286_));
 sg13g2_nand2_1 _19203_ (.Y(_12288_),
    .A(net1004),
    .B(_12263_));
 sg13g2_o21ai_1 _19204_ (.B1(_12288_),
    .Y(_00394_),
    .A1(net56),
    .A2(_12287_));
 sg13g2_nor2b_1 _19205_ (.A(_12285_),
    .B_N(\cpu.dcache.r_data[2][21] ),
    .Y(_12289_));
 sg13g2_a21oi_1 _19206_ (.A1(net996),
    .A2(_12285_),
    .Y(_12290_),
    .B1(_12289_));
 sg13g2_nand2_1 _19207_ (.Y(_12291_),
    .A(net1003),
    .B(_12263_));
 sg13g2_o21ai_1 _19208_ (.B1(_12291_),
    .Y(_00395_),
    .A1(net56),
    .A2(_12290_));
 sg13g2_mux2_1 _19209_ (.A0(\cpu.dcache.r_data[2][22] ),
    .A1(net1093),
    .S(_12285_),
    .X(_12292_));
 sg13g2_nor2_1 _19210_ (.A(_12263_),
    .B(_12292_),
    .Y(_12293_));
 sg13g2_a21oi_1 _19211_ (.A1(net756),
    .A2(net56),
    .Y(_00396_),
    .B1(_12293_));
 sg13g2_mux2_1 _19212_ (.A0(\cpu.dcache.r_data[2][23] ),
    .A1(net1002),
    .S(_12285_),
    .X(_12294_));
 sg13g2_nor2_1 _19213_ (.A(_12263_),
    .B(_12294_),
    .Y(_12295_));
 sg13g2_a21oi_1 _19214_ (.A1(net755),
    .A2(net56),
    .Y(_00397_),
    .B1(_12295_));
 sg13g2_nor2_1 _19215_ (.A(_12227_),
    .B(_12170_),
    .Y(_12296_));
 sg13g2_buf_2 _19216_ (.A(_12296_),
    .X(_12297_));
 sg13g2_buf_1 _19217_ (.A(_12297_),
    .X(_12298_));
 sg13g2_nor2_1 _19218_ (.A(net678),
    .B(net617),
    .Y(_12299_));
 sg13g2_buf_1 _19219_ (.A(_12299_),
    .X(_12300_));
 sg13g2_nor2b_1 _19220_ (.A(net489),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12301_));
 sg13g2_a21oi_1 _19221_ (.A1(net997),
    .A2(net489),
    .Y(_12302_),
    .B1(_12301_));
 sg13g2_nand2_1 _19222_ (.Y(_12303_),
    .A(net497),
    .B(_12298_));
 sg13g2_o21ai_1 _19223_ (.B1(_12303_),
    .Y(_00398_),
    .A1(net55),
    .A2(_12302_));
 sg13g2_nor2b_1 _19224_ (.A(net489),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12304_));
 sg13g2_a21oi_1 _19225_ (.A1(net996),
    .A2(net489),
    .Y(_12305_),
    .B1(_12304_));
 sg13g2_nand2_1 _19226_ (.Y(_12306_),
    .A(_12042_),
    .B(net55));
 sg13g2_o21ai_1 _19227_ (.B1(_12306_),
    .Y(_00399_),
    .A1(_12298_),
    .A2(_12305_));
 sg13g2_nor2b_1 _19228_ (.A(net489),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12307_));
 sg13g2_a21oi_1 _19229_ (.A1(_12129_),
    .A2(net489),
    .Y(_12308_),
    .B1(_12307_));
 sg13g2_nand2_1 _19230_ (.Y(_12309_),
    .A(net498),
    .B(_12297_));
 sg13g2_o21ai_1 _19231_ (.B1(_12309_),
    .Y(_00400_),
    .A1(net55),
    .A2(_12308_));
 sg13g2_nor2b_1 _19232_ (.A(net489),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12310_));
 sg13g2_a21oi_1 _19233_ (.A1(_12203_),
    .A2(net489),
    .Y(_12311_),
    .B1(_12310_));
 sg13g2_nand2_1 _19234_ (.Y(_12312_),
    .A(net495),
    .B(_12297_));
 sg13g2_o21ai_1 _19235_ (.B1(_12312_),
    .Y(_00401_),
    .A1(net55),
    .A2(_12311_));
 sg13g2_nor2_1 _19236_ (.A(_12227_),
    .B(_12048_),
    .Y(_12313_));
 sg13g2_buf_2 _19237_ (.A(_12313_),
    .X(_12314_));
 sg13g2_nor2b_1 _19238_ (.A(_12314_),
    .B_N(\cpu.dcache.r_data[2][28] ),
    .Y(_12315_));
 sg13g2_a21oi_1 _19239_ (.A1(net997),
    .A2(_12314_),
    .Y(_12316_),
    .B1(_12315_));
 sg13g2_nand2_1 _19240_ (.Y(_12317_),
    .A(net494),
    .B(_12297_));
 sg13g2_o21ai_1 _19241_ (.B1(_12317_),
    .Y(_00402_),
    .A1(net55),
    .A2(_12316_));
 sg13g2_nor2b_1 _19242_ (.A(_12314_),
    .B_N(\cpu.dcache.r_data[2][29] ),
    .Y(_12318_));
 sg13g2_a21oi_1 _19243_ (.A1(net996),
    .A2(_12314_),
    .Y(_12319_),
    .B1(_12318_));
 sg13g2_nand2_1 _19244_ (.Y(_12320_),
    .A(net493),
    .B(_12297_));
 sg13g2_o21ai_1 _19245_ (.B1(_12320_),
    .Y(_00403_),
    .A1(net55),
    .A2(_12319_));
 sg13g2_nor2b_1 _19246_ (.A(_12232_),
    .B_N(\cpu.dcache.r_data[2][2] ),
    .Y(_12321_));
 sg13g2_a21oi_1 _19247_ (.A1(net999),
    .A2(_12232_),
    .Y(_12322_),
    .B1(_12321_));
 sg13g2_nand2_1 _19248_ (.Y(_12323_),
    .A(net871),
    .B(_12229_));
 sg13g2_o21ai_1 _19249_ (.B1(_12323_),
    .Y(_00404_),
    .A1(_12230_),
    .A2(_12322_));
 sg13g2_buf_1 _19250_ (.A(net1097),
    .X(_12324_));
 sg13g2_nor2b_1 _19251_ (.A(_12314_),
    .B_N(\cpu.dcache.r_data[2][30] ),
    .Y(_12325_));
 sg13g2_a21oi_1 _19252_ (.A1(net995),
    .A2(_12314_),
    .Y(_12326_),
    .B1(_12325_));
 sg13g2_nand2_1 _19253_ (.Y(_12327_),
    .A(net492),
    .B(_12297_));
 sg13g2_o21ai_1 _19254_ (.B1(_12327_),
    .Y(_00405_),
    .A1(net55),
    .A2(_12326_));
 sg13g2_nor2b_1 _19255_ (.A(_12314_),
    .B_N(\cpu.dcache.r_data[2][31] ),
    .Y(_12328_));
 sg13g2_a21oi_1 _19256_ (.A1(_12203_),
    .A2(_12314_),
    .Y(_12329_),
    .B1(_12328_));
 sg13g2_nand2_1 _19257_ (.Y(_12330_),
    .A(net491),
    .B(_12297_));
 sg13g2_o21ai_1 _19258_ (.B1(_12330_),
    .Y(_00406_),
    .A1(net55),
    .A2(_12329_));
 sg13g2_mux2_1 _19259_ (.A0(\cpu.dcache.r_data[2][3] ),
    .A1(net1002),
    .S(_12232_),
    .X(_12331_));
 sg13g2_nor2_1 _19260_ (.A(_12229_),
    .B(_12331_),
    .Y(_12332_));
 sg13g2_a21oi_1 _19261_ (.A1(net870),
    .A2(net58),
    .Y(_00407_),
    .B1(_12332_));
 sg13g2_nor2_1 _19262_ (.A(_09390_),
    .B(_12073_),
    .Y(_12333_));
 sg13g2_buf_2 _19263_ (.A(_12333_),
    .X(_12334_));
 sg13g2_nor2b_1 _19264_ (.A(_12334_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12335_));
 sg13g2_a21oi_1 _19265_ (.A1(net997),
    .A2(_12334_),
    .Y(_12336_),
    .B1(_12335_));
 sg13g2_nand2_1 _19266_ (.Y(_12337_),
    .A(net1004),
    .B(_12229_));
 sg13g2_o21ai_1 _19267_ (.B1(_12337_),
    .Y(_00408_),
    .A1(net58),
    .A2(_12336_));
 sg13g2_nor2b_1 _19268_ (.A(_12334_),
    .B_N(\cpu.dcache.r_data[2][5] ),
    .Y(_12338_));
 sg13g2_a21oi_1 _19269_ (.A1(net996),
    .A2(_12334_),
    .Y(_12339_),
    .B1(_12338_));
 sg13g2_nand2_1 _19270_ (.Y(_12340_),
    .A(net1003),
    .B(_12229_));
 sg13g2_o21ai_1 _19271_ (.B1(_12340_),
    .Y(_00409_),
    .A1(net58),
    .A2(_12339_));
 sg13g2_mux2_1 _19272_ (.A0(\cpu.dcache.r_data[2][6] ),
    .A1(net1093),
    .S(_12334_),
    .X(_12341_));
 sg13g2_nor2_1 _19273_ (.A(_12229_),
    .B(_12341_),
    .Y(_12342_));
 sg13g2_a21oi_1 _19274_ (.A1(net756),
    .A2(net58),
    .Y(_00410_),
    .B1(_12342_));
 sg13g2_mux2_1 _19275_ (.A0(\cpu.dcache.r_data[2][7] ),
    .A1(net1002),
    .S(_12334_),
    .X(_12343_));
 sg13g2_nor2_1 _19276_ (.A(_12229_),
    .B(_12343_),
    .Y(_12344_));
 sg13g2_a21oi_1 _19277_ (.A1(net755),
    .A2(net58),
    .Y(_00411_),
    .B1(_12344_));
 sg13g2_nor2b_1 _19278_ (.A(_12240_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12345_));
 sg13g2_a21oi_1 _19279_ (.A1(_12247_),
    .A2(_12240_),
    .Y(_12346_),
    .B1(_12345_));
 sg13g2_nand2_1 _19280_ (.Y(_12347_),
    .A(net497),
    .B(_12237_));
 sg13g2_o21ai_1 _19281_ (.B1(_12347_),
    .Y(_00412_),
    .A1(_12238_),
    .A2(_12346_));
 sg13g2_nor2b_1 _19282_ (.A(_12240_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12348_));
 sg13g2_a21oi_1 _19283_ (.A1(_12271_),
    .A2(_12240_),
    .Y(_12349_),
    .B1(_12348_));
 sg13g2_nand2_1 _19284_ (.Y(_12350_),
    .A(net496),
    .B(_12237_));
 sg13g2_o21ai_1 _19285_ (.B1(_12350_),
    .Y(_00413_),
    .A1(_12238_),
    .A2(_12349_));
 sg13g2_nand2_2 _19286_ (.Y(_12351_),
    .A(net1050),
    .B(net693));
 sg13g2_buf_1 _19287_ (.A(_12351_),
    .X(_12352_));
 sg13g2_nor2_1 _19288_ (.A(net566),
    .B(_12099_),
    .Y(_12353_));
 sg13g2_buf_1 _19289_ (.A(_12353_),
    .X(_12354_));
 sg13g2_buf_1 _19290_ (.A(_12354_),
    .X(_12355_));
 sg13g2_nor2_1 _19291_ (.A(net566),
    .B(_11913_),
    .Y(_12356_));
 sg13g2_buf_2 _19292_ (.A(_12356_),
    .X(_12357_));
 sg13g2_nor2b_1 _19293_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[3][0] ),
    .Y(_12358_));
 sg13g2_a21oi_1 _19294_ (.A1(net997),
    .A2(_12357_),
    .Y(_12359_),
    .B1(_12358_));
 sg13g2_nand2_1 _19295_ (.Y(_12360_),
    .A(_12269_),
    .B(net54));
 sg13g2_o21ai_1 _19296_ (.B1(_12360_),
    .Y(_00414_),
    .A1(net54),
    .A2(_12359_));
 sg13g2_nor2_1 _19297_ (.A(net566),
    .B(_12109_),
    .Y(_12361_));
 sg13g2_buf_2 _19298_ (.A(_12361_),
    .X(_12362_));
 sg13g2_buf_1 _19299_ (.A(_12362_),
    .X(_12363_));
 sg13g2_nor2_1 _19300_ (.A(net566),
    .B(_11928_),
    .Y(_12364_));
 sg13g2_buf_2 _19301_ (.A(_12364_),
    .X(_12365_));
 sg13g2_nor2b_1 _19302_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12366_));
 sg13g2_a21oi_1 _19303_ (.A1(net995),
    .A2(_12365_),
    .Y(_12367_),
    .B1(_12366_));
 sg13g2_nand2_1 _19304_ (.Y(_12368_),
    .A(net498),
    .B(net53));
 sg13g2_o21ai_1 _19305_ (.B1(_12368_),
    .Y(_00415_),
    .A1(net53),
    .A2(_12367_));
 sg13g2_nor2b_1 _19306_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12369_));
 sg13g2_a21oi_1 _19307_ (.A1(net998),
    .A2(_12365_),
    .Y(_12370_),
    .B1(_12369_));
 sg13g2_nand2_1 _19308_ (.Y(_12371_),
    .A(net495),
    .B(net53));
 sg13g2_o21ai_1 _19309_ (.B1(_12371_),
    .Y(_00416_),
    .A1(net53),
    .A2(_12370_));
 sg13g2_nor2_1 _19310_ (.A(net566),
    .B(_11950_),
    .Y(_12372_));
 sg13g2_buf_2 _19311_ (.A(_12372_),
    .X(_12373_));
 sg13g2_nor2b_1 _19312_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[3][12] ),
    .Y(_12374_));
 sg13g2_a21oi_1 _19313_ (.A1(_12247_),
    .A2(_12373_),
    .Y(_12375_),
    .B1(_12374_));
 sg13g2_nand2_1 _19314_ (.Y(_12376_),
    .A(net494),
    .B(_12362_));
 sg13g2_o21ai_1 _19315_ (.B1(_12376_),
    .Y(_00417_),
    .A1(net53),
    .A2(_12375_));
 sg13g2_nor2b_1 _19316_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[3][13] ),
    .Y(_12377_));
 sg13g2_a21oi_1 _19317_ (.A1(_12271_),
    .A2(_12373_),
    .Y(_12378_),
    .B1(_12377_));
 sg13g2_nand2_1 _19318_ (.Y(_12379_),
    .A(net493),
    .B(_12362_));
 sg13g2_o21ai_1 _19319_ (.B1(_12379_),
    .Y(_00418_),
    .A1(net53),
    .A2(_12378_));
 sg13g2_nor2b_1 _19320_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[3][14] ),
    .Y(_12380_));
 sg13g2_a21oi_1 _19321_ (.A1(net995),
    .A2(_12373_),
    .Y(_12381_),
    .B1(_12380_));
 sg13g2_nand2_1 _19322_ (.Y(_12382_),
    .A(net492),
    .B(_12362_));
 sg13g2_o21ai_1 _19323_ (.B1(_12382_),
    .Y(_00419_),
    .A1(_12363_),
    .A2(_12381_));
 sg13g2_nor2b_1 _19324_ (.A(_12373_),
    .B_N(\cpu.dcache.r_data[3][15] ),
    .Y(_12383_));
 sg13g2_a21oi_1 _19325_ (.A1(net998),
    .A2(_12373_),
    .Y(_12384_),
    .B1(_12383_));
 sg13g2_nand2_1 _19326_ (.Y(_12385_),
    .A(net491),
    .B(_12362_));
 sg13g2_o21ai_1 _19327_ (.B1(_12385_),
    .Y(_00420_),
    .A1(_12363_),
    .A2(_12384_));
 sg13g2_nor2_1 _19328_ (.A(net566),
    .B(_12137_),
    .Y(_12386_));
 sg13g2_buf_1 _19329_ (.A(_12386_),
    .X(_12387_));
 sg13g2_buf_1 _19330_ (.A(_12387_),
    .X(_12388_));
 sg13g2_nor2_1 _19331_ (.A(net566),
    .B(_11982_),
    .Y(_12389_));
 sg13g2_buf_2 _19332_ (.A(_12389_),
    .X(_12390_));
 sg13g2_nor2b_1 _19333_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[3][16] ),
    .Y(_12391_));
 sg13g2_a21oi_1 _19334_ (.A1(net997),
    .A2(_12390_),
    .Y(_12392_),
    .B1(_12391_));
 sg13g2_nand2_1 _19335_ (.Y(_12393_),
    .A(net869),
    .B(net52));
 sg13g2_o21ai_1 _19336_ (.B1(_12393_),
    .Y(_00421_),
    .A1(net52),
    .A2(_12392_));
 sg13g2_nor2b_1 _19337_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[3][17] ),
    .Y(_12394_));
 sg13g2_a21oi_1 _19338_ (.A1(net996),
    .A2(_12390_),
    .Y(_12395_),
    .B1(_12394_));
 sg13g2_nand2_1 _19339_ (.Y(_12396_),
    .A(net868),
    .B(net52));
 sg13g2_o21ai_1 _19340_ (.B1(_12396_),
    .Y(_00422_),
    .A1(_12388_),
    .A2(_12395_));
 sg13g2_nor2b_1 _19341_ (.A(_12390_),
    .B_N(\cpu.dcache.r_data[3][18] ),
    .Y(_12397_));
 sg13g2_a21oi_1 _19342_ (.A1(net995),
    .A2(_12390_),
    .Y(_12398_),
    .B1(_12397_));
 sg13g2_buf_1 _19343_ (.A(_10002_),
    .X(_12399_));
 sg13g2_nand2_1 _19344_ (.Y(_12400_),
    .A(net867),
    .B(_12387_));
 sg13g2_o21ai_1 _19345_ (.B1(_12400_),
    .Y(_00423_),
    .A1(_12388_),
    .A2(_12398_));
 sg13g2_mux2_1 _19346_ (.A0(\cpu.dcache.r_data[3][19] ),
    .A1(net1002),
    .S(_12390_),
    .X(_12401_));
 sg13g2_nor2_1 _19347_ (.A(_12387_),
    .B(_12401_),
    .Y(_12402_));
 sg13g2_a21oi_1 _19348_ (.A1(net870),
    .A2(net52),
    .Y(_00424_),
    .B1(_12402_));
 sg13g2_nor2b_1 _19349_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[3][1] ),
    .Y(_12403_));
 sg13g2_a21oi_1 _19350_ (.A1(net996),
    .A2(_12357_),
    .Y(_12404_),
    .B1(_12403_));
 sg13g2_nand2_1 _19351_ (.Y(_12405_),
    .A(_12282_),
    .B(net54));
 sg13g2_o21ai_1 _19352_ (.B1(_12405_),
    .Y(_00425_),
    .A1(net54),
    .A2(_12404_));
 sg13g2_or2_1 _19353_ (.X(_12406_),
    .B(_12006_),
    .A(_12351_));
 sg13g2_buf_1 _19354_ (.A(_12406_),
    .X(_12407_));
 sg13g2_mux2_1 _19355_ (.A0(net1099),
    .A1(\cpu.dcache.r_data[3][20] ),
    .S(_12407_),
    .X(_12408_));
 sg13g2_buf_1 _19356_ (.A(_10013_),
    .X(_12409_));
 sg13g2_mux2_1 _19357_ (.A0(_12408_),
    .A1(net994),
    .S(net52),
    .X(_00426_));
 sg13g2_mux2_1 _19358_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[3][21] ),
    .S(_12407_),
    .X(_12410_));
 sg13g2_buf_1 _19359_ (.A(_10019_),
    .X(_12411_));
 sg13g2_mux2_1 _19360_ (.A0(_12410_),
    .A1(net993),
    .S(net52),
    .X(_00427_));
 sg13g2_mux2_1 _19361_ (.A0(net1093),
    .A1(\cpu.dcache.r_data[3][22] ),
    .S(_12407_),
    .X(_12412_));
 sg13g2_nor2_1 _19362_ (.A(_12387_),
    .B(_12412_),
    .Y(_12413_));
 sg13g2_a21oi_1 _19363_ (.A1(net756),
    .A2(net52),
    .Y(_00428_),
    .B1(_12413_));
 sg13g2_mux2_1 _19364_ (.A0(net1094),
    .A1(\cpu.dcache.r_data[3][23] ),
    .S(_12407_),
    .X(_12414_));
 sg13g2_nor2_1 _19365_ (.A(_12387_),
    .B(_12414_),
    .Y(_12415_));
 sg13g2_a21oi_1 _19366_ (.A1(net755),
    .A2(net52),
    .Y(_00429_),
    .B1(_12415_));
 sg13g2_nor2_1 _19367_ (.A(_12352_),
    .B(_12170_),
    .Y(_12416_));
 sg13g2_buf_2 _19368_ (.A(_12416_),
    .X(_12417_));
 sg13g2_buf_1 _19369_ (.A(_12417_),
    .X(_12418_));
 sg13g2_buf_1 _19370_ (.A(net1099),
    .X(_12419_));
 sg13g2_nor2_1 _19371_ (.A(_12351_),
    .B(net617),
    .Y(_12420_));
 sg13g2_buf_1 _19372_ (.A(_12420_),
    .X(_12421_));
 sg13g2_nor2b_1 _19373_ (.A(net488),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12422_));
 sg13g2_a21oi_1 _19374_ (.A1(net992),
    .A2(net488),
    .Y(_12423_),
    .B1(_12422_));
 sg13g2_nand2_1 _19375_ (.Y(_12424_),
    .A(net497),
    .B(net51));
 sg13g2_o21ai_1 _19376_ (.B1(_12424_),
    .Y(_00430_),
    .A1(net51),
    .A2(_12423_));
 sg13g2_buf_1 _19377_ (.A(net1095),
    .X(_12425_));
 sg13g2_nor2b_1 _19378_ (.A(net488),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12426_));
 sg13g2_a21oi_1 _19379_ (.A1(net991),
    .A2(net488),
    .Y(_12427_),
    .B1(_12426_));
 sg13g2_nand2_1 _19380_ (.Y(_12428_),
    .A(net496),
    .B(net51));
 sg13g2_o21ai_1 _19381_ (.B1(_12428_),
    .Y(_00431_),
    .A1(net51),
    .A2(_12427_));
 sg13g2_nor2b_1 _19382_ (.A(net488),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12429_));
 sg13g2_a21oi_1 _19383_ (.A1(net995),
    .A2(net488),
    .Y(_12430_),
    .B1(_12429_));
 sg13g2_nand2_1 _19384_ (.Y(_12431_),
    .A(net498),
    .B(_12417_));
 sg13g2_o21ai_1 _19385_ (.B1(_12431_),
    .Y(_00432_),
    .A1(_12418_),
    .A2(_12430_));
 sg13g2_nor2b_1 _19386_ (.A(net488),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12432_));
 sg13g2_a21oi_1 _19387_ (.A1(net998),
    .A2(net488),
    .Y(_12433_),
    .B1(_12432_));
 sg13g2_nand2_1 _19388_ (.Y(_12434_),
    .A(_12046_),
    .B(_12417_));
 sg13g2_o21ai_1 _19389_ (.B1(_12434_),
    .Y(_00433_),
    .A1(net51),
    .A2(_12433_));
 sg13g2_nor2_1 _19390_ (.A(_12352_),
    .B(_12048_),
    .Y(_12435_));
 sg13g2_buf_2 _19391_ (.A(_12435_),
    .X(_12436_));
 sg13g2_nor2b_1 _19392_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[3][28] ),
    .Y(_12437_));
 sg13g2_a21oi_1 _19393_ (.A1(net992),
    .A2(_12436_),
    .Y(_12438_),
    .B1(_12437_));
 sg13g2_nand2_1 _19394_ (.Y(_12439_),
    .A(_12053_),
    .B(_12417_));
 sg13g2_o21ai_1 _19395_ (.B1(_12439_),
    .Y(_00434_),
    .A1(net51),
    .A2(_12438_));
 sg13g2_nor2b_1 _19396_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[3][29] ),
    .Y(_12440_));
 sg13g2_a21oi_1 _19397_ (.A1(net991),
    .A2(_12436_),
    .Y(_12441_),
    .B1(_12440_));
 sg13g2_nand2_1 _19398_ (.Y(_12442_),
    .A(_12057_),
    .B(_12417_));
 sg13g2_o21ai_1 _19399_ (.B1(_12442_),
    .Y(_00435_),
    .A1(_12418_),
    .A2(_12441_));
 sg13g2_nor2b_1 _19400_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[3][2] ),
    .Y(_12443_));
 sg13g2_a21oi_1 _19401_ (.A1(net995),
    .A2(_12357_),
    .Y(_12444_),
    .B1(_12443_));
 sg13g2_nand2_1 _19402_ (.Y(_12445_),
    .A(_12399_),
    .B(_12354_));
 sg13g2_o21ai_1 _19403_ (.B1(_12445_),
    .Y(_00436_),
    .A1(_12355_),
    .A2(_12444_));
 sg13g2_nor2b_1 _19404_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[3][30] ),
    .Y(_12446_));
 sg13g2_a21oi_1 _19405_ (.A1(_12324_),
    .A2(_12436_),
    .Y(_12447_),
    .B1(_12446_));
 sg13g2_nand2_1 _19406_ (.Y(_12448_),
    .A(_12064_),
    .B(_12417_));
 sg13g2_o21ai_1 _19407_ (.B1(_12448_),
    .Y(_00437_),
    .A1(net51),
    .A2(_12447_));
 sg13g2_nor2b_1 _19408_ (.A(_12436_),
    .B_N(\cpu.dcache.r_data[3][31] ),
    .Y(_12449_));
 sg13g2_a21oi_1 _19409_ (.A1(net998),
    .A2(_12436_),
    .Y(_12450_),
    .B1(_12449_));
 sg13g2_nand2_1 _19410_ (.Y(_12451_),
    .A(_12068_),
    .B(_12417_));
 sg13g2_o21ai_1 _19411_ (.B1(_12451_),
    .Y(_00438_),
    .A1(net51),
    .A2(_12450_));
 sg13g2_buf_1 _19412_ (.A(_11939_),
    .X(_12452_));
 sg13g2_mux2_1 _19413_ (.A0(\cpu.dcache.r_data[3][3] ),
    .A1(net1092),
    .S(_12357_),
    .X(_12453_));
 sg13g2_nor2_1 _19414_ (.A(_12354_),
    .B(_12453_),
    .Y(_12454_));
 sg13g2_a21oi_1 _19415_ (.A1(_11997_),
    .A2(_12355_),
    .Y(_00439_),
    .B1(_12454_));
 sg13g2_or2_1 _19416_ (.X(_12455_),
    .B(_12073_),
    .A(_12351_));
 sg13g2_buf_1 _19417_ (.A(_12455_),
    .X(_12456_));
 sg13g2_mux2_1 _19418_ (.A0(net1099),
    .A1(\cpu.dcache.r_data[3][4] ),
    .S(_12456_),
    .X(_12457_));
 sg13g2_mux2_1 _19419_ (.A0(_12457_),
    .A1(net994),
    .S(net54),
    .X(_00440_));
 sg13g2_mux2_1 _19420_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[3][5] ),
    .S(_12456_),
    .X(_12458_));
 sg13g2_mux2_1 _19421_ (.A0(_12458_),
    .A1(net993),
    .S(net54),
    .X(_00441_));
 sg13g2_mux2_1 _19422_ (.A0(_12020_),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(_12456_),
    .X(_12459_));
 sg13g2_nor2_1 _19423_ (.A(_12354_),
    .B(_12459_),
    .Y(_12460_));
 sg13g2_a21oi_1 _19424_ (.A1(_12019_),
    .A2(net54),
    .Y(_00442_),
    .B1(_12460_));
 sg13g2_mux2_1 _19425_ (.A0(net1094),
    .A1(\cpu.dcache.r_data[3][7] ),
    .S(_12456_),
    .X(_12461_));
 sg13g2_nor2_1 _19426_ (.A(_12354_),
    .B(_12461_),
    .Y(_12462_));
 sg13g2_a21oi_1 _19427_ (.A1(_12025_),
    .A2(net54),
    .Y(_00443_),
    .B1(_12462_));
 sg13g2_nor2b_1 _19428_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12463_));
 sg13g2_a21oi_1 _19429_ (.A1(net992),
    .A2(_12365_),
    .Y(_12464_),
    .B1(_12463_));
 sg13g2_nand2_1 _19430_ (.Y(_12465_),
    .A(net497),
    .B(_12362_));
 sg13g2_o21ai_1 _19431_ (.B1(_12465_),
    .Y(_00444_),
    .A1(net53),
    .A2(_12464_));
 sg13g2_nor2b_1 _19432_ (.A(_12365_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12466_));
 sg13g2_a21oi_1 _19433_ (.A1(net991),
    .A2(_12365_),
    .Y(_12467_),
    .B1(_12466_));
 sg13g2_nand2_1 _19434_ (.Y(_12468_),
    .A(net496),
    .B(_12362_));
 sg13g2_o21ai_1 _19435_ (.B1(_12468_),
    .Y(_00445_),
    .A1(net53),
    .A2(_12467_));
 sg13g2_buf_1 _19436_ (.A(_10042_),
    .X(_12469_));
 sg13g2_nor2_1 _19437_ (.A(net565),
    .B(_12099_),
    .Y(_12470_));
 sg13g2_buf_2 _19438_ (.A(_12470_),
    .X(_12471_));
 sg13g2_buf_1 _19439_ (.A(_12471_),
    .X(_12472_));
 sg13g2_nor2_1 _19440_ (.A(net565),
    .B(_11913_),
    .Y(_12473_));
 sg13g2_buf_2 _19441_ (.A(_12473_),
    .X(_12474_));
 sg13g2_nor2b_1 _19442_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[4][0] ),
    .Y(_12475_));
 sg13g2_a21oi_1 _19443_ (.A1(net992),
    .A2(_12474_),
    .Y(_12476_),
    .B1(_12475_));
 sg13g2_nand2_1 _19444_ (.Y(_12477_),
    .A(net869),
    .B(net50));
 sg13g2_o21ai_1 _19445_ (.B1(_12477_),
    .Y(_00446_),
    .A1(net50),
    .A2(_12476_));
 sg13g2_nor2_1 _19446_ (.A(net565),
    .B(_12109_),
    .Y(_12478_));
 sg13g2_buf_2 _19447_ (.A(_12478_),
    .X(_12479_));
 sg13g2_buf_1 _19448_ (.A(_12479_),
    .X(_12480_));
 sg13g2_nor2_1 _19449_ (.A(_12469_),
    .B(_11928_),
    .Y(_12481_));
 sg13g2_buf_2 _19450_ (.A(_12481_),
    .X(_12482_));
 sg13g2_nor2b_1 _19451_ (.A(_12482_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12483_));
 sg13g2_a21oi_1 _19452_ (.A1(net995),
    .A2(_12482_),
    .Y(_12484_),
    .B1(_12483_));
 sg13g2_nand2_1 _19453_ (.Y(_12485_),
    .A(net498),
    .B(net49));
 sg13g2_o21ai_1 _19454_ (.B1(_12485_),
    .Y(_00447_),
    .A1(net49),
    .A2(_12484_));
 sg13g2_nor2b_1 _19455_ (.A(_12482_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12486_));
 sg13g2_a21oi_1 _19456_ (.A1(net998),
    .A2(_12482_),
    .Y(_12487_),
    .B1(_12486_));
 sg13g2_nand2_1 _19457_ (.Y(_12488_),
    .A(net495),
    .B(net49));
 sg13g2_o21ai_1 _19458_ (.B1(_12488_),
    .Y(_00448_),
    .A1(net49),
    .A2(_12487_));
 sg13g2_nor2_1 _19459_ (.A(net565),
    .B(_11950_),
    .Y(_12489_));
 sg13g2_buf_2 _19460_ (.A(_12489_),
    .X(_12490_));
 sg13g2_nor2b_1 _19461_ (.A(_12490_),
    .B_N(\cpu.dcache.r_data[4][12] ),
    .Y(_12491_));
 sg13g2_a21oi_1 _19462_ (.A1(net992),
    .A2(_12490_),
    .Y(_12492_),
    .B1(_12491_));
 sg13g2_nand2_1 _19463_ (.Y(_12493_),
    .A(net494),
    .B(_12479_));
 sg13g2_o21ai_1 _19464_ (.B1(_12493_),
    .Y(_00449_),
    .A1(net49),
    .A2(_12492_));
 sg13g2_nor2b_1 _19465_ (.A(_12490_),
    .B_N(\cpu.dcache.r_data[4][13] ),
    .Y(_12494_));
 sg13g2_a21oi_1 _19466_ (.A1(net991),
    .A2(_12490_),
    .Y(_12495_),
    .B1(_12494_));
 sg13g2_nand2_1 _19467_ (.Y(_12496_),
    .A(net493),
    .B(_12479_));
 sg13g2_o21ai_1 _19468_ (.B1(_12496_),
    .Y(_00450_),
    .A1(_12480_),
    .A2(_12495_));
 sg13g2_nor2b_1 _19469_ (.A(_12490_),
    .B_N(\cpu.dcache.r_data[4][14] ),
    .Y(_12497_));
 sg13g2_a21oi_1 _19470_ (.A1(_12324_),
    .A2(_12490_),
    .Y(_12498_),
    .B1(_12497_));
 sg13g2_nand2_1 _19471_ (.Y(_12499_),
    .A(net492),
    .B(_12479_));
 sg13g2_o21ai_1 _19472_ (.B1(_12499_),
    .Y(_00451_),
    .A1(net49),
    .A2(_12498_));
 sg13g2_buf_1 _19473_ (.A(net1096),
    .X(_12500_));
 sg13g2_nor2b_1 _19474_ (.A(_12490_),
    .B_N(\cpu.dcache.r_data[4][15] ),
    .Y(_12501_));
 sg13g2_a21oi_1 _19475_ (.A1(net990),
    .A2(_12490_),
    .Y(_12502_),
    .B1(_12501_));
 sg13g2_nand2_1 _19476_ (.Y(_12503_),
    .A(net491),
    .B(_12479_));
 sg13g2_o21ai_1 _19477_ (.B1(_12503_),
    .Y(_00452_),
    .A1(_12480_),
    .A2(_12502_));
 sg13g2_nor2_1 _19478_ (.A(net565),
    .B(_12137_),
    .Y(_12504_));
 sg13g2_buf_1 _19479_ (.A(_12504_),
    .X(_12505_));
 sg13g2_buf_1 _19480_ (.A(_12505_),
    .X(_12506_));
 sg13g2_nor2_1 _19481_ (.A(_10042_),
    .B(_11982_),
    .Y(_12507_));
 sg13g2_buf_2 _19482_ (.A(_12507_),
    .X(_12508_));
 sg13g2_nor2b_1 _19483_ (.A(_12508_),
    .B_N(\cpu.dcache.r_data[4][16] ),
    .Y(_12509_));
 sg13g2_a21oi_1 _19484_ (.A1(net992),
    .A2(_12508_),
    .Y(_12510_),
    .B1(_12509_));
 sg13g2_nand2_1 _19485_ (.Y(_12511_),
    .A(net869),
    .B(net48));
 sg13g2_o21ai_1 _19486_ (.B1(_12511_),
    .Y(_00453_),
    .A1(net48),
    .A2(_12510_));
 sg13g2_nor2b_1 _19487_ (.A(_12508_),
    .B_N(\cpu.dcache.r_data[4][17] ),
    .Y(_12512_));
 sg13g2_a21oi_1 _19488_ (.A1(net991),
    .A2(_12508_),
    .Y(_12513_),
    .B1(_12512_));
 sg13g2_nand2_1 _19489_ (.Y(_12514_),
    .A(net868),
    .B(net48));
 sg13g2_o21ai_1 _19490_ (.B1(_12514_),
    .Y(_00454_),
    .A1(_12506_),
    .A2(_12513_));
 sg13g2_nor2b_1 _19491_ (.A(_12508_),
    .B_N(\cpu.dcache.r_data[4][18] ),
    .Y(_12515_));
 sg13g2_a21oi_1 _19492_ (.A1(net995),
    .A2(_12508_),
    .Y(_12516_),
    .B1(_12515_));
 sg13g2_nand2_1 _19493_ (.Y(_12517_),
    .A(net867),
    .B(_12505_));
 sg13g2_o21ai_1 _19494_ (.B1(_12517_),
    .Y(_00455_),
    .A1(_12506_),
    .A2(_12516_));
 sg13g2_mux2_1 _19495_ (.A0(\cpu.dcache.r_data[4][19] ),
    .A1(net1092),
    .S(_12508_),
    .X(_12518_));
 sg13g2_nor2_1 _19496_ (.A(_12505_),
    .B(_12518_),
    .Y(_12519_));
 sg13g2_a21oi_1 _19497_ (.A1(net870),
    .A2(net48),
    .Y(_00456_),
    .B1(_12519_));
 sg13g2_nor2b_1 _19498_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[4][1] ),
    .Y(_12520_));
 sg13g2_a21oi_1 _19499_ (.A1(net991),
    .A2(_12474_),
    .Y(_12521_),
    .B1(_12520_));
 sg13g2_nand2_1 _19500_ (.Y(_12522_),
    .A(net868),
    .B(net50));
 sg13g2_o21ai_1 _19501_ (.B1(_12522_),
    .Y(_00457_),
    .A1(_12472_),
    .A2(_12521_));
 sg13g2_nor2_1 _19502_ (.A(net565),
    .B(_12006_),
    .Y(_12523_));
 sg13g2_buf_2 _19503_ (.A(_12523_),
    .X(_12524_));
 sg13g2_nor2b_1 _19504_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12525_));
 sg13g2_a21oi_1 _19505_ (.A1(net992),
    .A2(_12524_),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nand2_1 _19506_ (.Y(_12527_),
    .A(net1004),
    .B(_12505_));
 sg13g2_o21ai_1 _19507_ (.B1(_12527_),
    .Y(_00458_),
    .A1(net48),
    .A2(_12526_));
 sg13g2_nor2b_1 _19508_ (.A(_12524_),
    .B_N(\cpu.dcache.r_data[4][21] ),
    .Y(_12528_));
 sg13g2_a21oi_1 _19509_ (.A1(net991),
    .A2(_12524_),
    .Y(_12529_),
    .B1(_12528_));
 sg13g2_nand2_1 _19510_ (.Y(_12530_),
    .A(net1003),
    .B(_12505_));
 sg13g2_o21ai_1 _19511_ (.B1(_12530_),
    .Y(_00459_),
    .A1(net48),
    .A2(_12529_));
 sg13g2_mux2_1 _19512_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(net1097),
    .S(_12524_),
    .X(_12531_));
 sg13g2_nor2_1 _19513_ (.A(_12505_),
    .B(_12531_),
    .Y(_12532_));
 sg13g2_a21oi_1 _19514_ (.A1(net756),
    .A2(net48),
    .Y(_00460_),
    .B1(_12532_));
 sg13g2_mux2_1 _19515_ (.A0(\cpu.dcache.r_data[4][23] ),
    .A1(net1092),
    .S(_12524_),
    .X(_12533_));
 sg13g2_nor2_1 _19516_ (.A(_12505_),
    .B(_12533_),
    .Y(_12534_));
 sg13g2_a21oi_1 _19517_ (.A1(net755),
    .A2(net48),
    .Y(_00461_),
    .B1(_12534_));
 sg13g2_or2_1 _19518_ (.X(_12535_),
    .B(net617),
    .A(_10042_));
 sg13g2_buf_2 _19519_ (.A(_12535_),
    .X(_12536_));
 sg13g2_mux2_1 _19520_ (.A0(_11904_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(_12536_),
    .X(_12537_));
 sg13g2_nor2_1 _19521_ (.A(_12469_),
    .B(_12170_),
    .Y(_12538_));
 sg13g2_buf_2 _19522_ (.A(_12538_),
    .X(_12539_));
 sg13g2_mux2_1 _19523_ (.A0(_12537_),
    .A1(_12034_),
    .S(net76),
    .X(_00462_));
 sg13g2_mux2_1 _19524_ (.A0(_11959_),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(_12536_),
    .X(_12540_));
 sg13g2_mux2_1 _19525_ (.A0(_12540_),
    .A1(_12042_),
    .S(_12539_),
    .X(_00463_));
 sg13g2_mux2_1 _19526_ (.A0(_12043_),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(_12536_),
    .X(_12541_));
 sg13g2_mux2_1 _19527_ (.A0(_12541_),
    .A1(_11937_),
    .S(_12539_),
    .X(_00464_));
 sg13g2_mux2_1 _19528_ (.A0(_11998_),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(_12536_),
    .X(_12542_));
 sg13g2_mux2_1 _19529_ (.A0(_12542_),
    .A1(net495),
    .S(net76),
    .X(_00465_));
 sg13g2_nor2_1 _19530_ (.A(net565),
    .B(_12048_),
    .Y(_12543_));
 sg13g2_buf_2 _19531_ (.A(_12543_),
    .X(_12544_));
 sg13g2_nor2b_1 _19532_ (.A(_12544_),
    .B_N(\cpu.dcache.r_data[4][28] ),
    .Y(_12545_));
 sg13g2_a21oi_1 _19533_ (.A1(_12419_),
    .A2(_12544_),
    .Y(_12546_),
    .B1(_12545_));
 sg13g2_nand2_1 _19534_ (.Y(_12547_),
    .A(net494),
    .B(net76));
 sg13g2_o21ai_1 _19535_ (.B1(_12547_),
    .Y(_00466_),
    .A1(net76),
    .A2(_12546_));
 sg13g2_nor2b_1 _19536_ (.A(_12544_),
    .B_N(\cpu.dcache.r_data[4][29] ),
    .Y(_12548_));
 sg13g2_a21oi_1 _19537_ (.A1(_12425_),
    .A2(_12544_),
    .Y(_12549_),
    .B1(_12548_));
 sg13g2_nand2_1 _19538_ (.Y(_12550_),
    .A(net493),
    .B(net76));
 sg13g2_o21ai_1 _19539_ (.B1(_12550_),
    .Y(_00467_),
    .A1(net76),
    .A2(_12549_));
 sg13g2_buf_1 _19540_ (.A(net1097),
    .X(_12551_));
 sg13g2_nor2b_1 _19541_ (.A(_12474_),
    .B_N(\cpu.dcache.r_data[4][2] ),
    .Y(_12552_));
 sg13g2_a21oi_1 _19542_ (.A1(net989),
    .A2(_12474_),
    .Y(_12553_),
    .B1(_12552_));
 sg13g2_nand2_1 _19543_ (.Y(_12554_),
    .A(_12399_),
    .B(_12471_));
 sg13g2_o21ai_1 _19544_ (.B1(_12554_),
    .Y(_00468_),
    .A1(_12472_),
    .A2(_12553_));
 sg13g2_nor2b_1 _19545_ (.A(_12544_),
    .B_N(\cpu.dcache.r_data[4][30] ),
    .Y(_12555_));
 sg13g2_a21oi_1 _19546_ (.A1(net989),
    .A2(_12544_),
    .Y(_12556_),
    .B1(_12555_));
 sg13g2_nand2_1 _19547_ (.Y(_12557_),
    .A(net492),
    .B(_12538_));
 sg13g2_o21ai_1 _19548_ (.B1(_12557_),
    .Y(_00469_),
    .A1(net76),
    .A2(_12556_));
 sg13g2_nor2b_1 _19549_ (.A(_12544_),
    .B_N(\cpu.dcache.r_data[4][31] ),
    .Y(_12558_));
 sg13g2_a21oi_1 _19550_ (.A1(net990),
    .A2(_12544_),
    .Y(_12559_),
    .B1(_12558_));
 sg13g2_nand2_1 _19551_ (.Y(_12560_),
    .A(net491),
    .B(_12538_));
 sg13g2_o21ai_1 _19552_ (.B1(_12560_),
    .Y(_00470_),
    .A1(net76),
    .A2(_12559_));
 sg13g2_mux2_1 _19553_ (.A0(\cpu.dcache.r_data[4][3] ),
    .A1(net1092),
    .S(_12474_),
    .X(_12561_));
 sg13g2_nor2_1 _19554_ (.A(_12471_),
    .B(_12561_),
    .Y(_12562_));
 sg13g2_a21oi_1 _19555_ (.A1(_11997_),
    .A2(net50),
    .Y(_00471_),
    .B1(_12562_));
 sg13g2_nor2_1 _19556_ (.A(net565),
    .B(_12073_),
    .Y(_12563_));
 sg13g2_buf_2 _19557_ (.A(_12563_),
    .X(_12564_));
 sg13g2_nor2b_1 _19558_ (.A(_12564_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_12565_));
 sg13g2_a21oi_1 _19559_ (.A1(net992),
    .A2(_12564_),
    .Y(_12566_),
    .B1(_12565_));
 sg13g2_nand2_1 _19560_ (.Y(_12567_),
    .A(net1004),
    .B(_12471_));
 sg13g2_o21ai_1 _19561_ (.B1(_12567_),
    .Y(_00472_),
    .A1(net50),
    .A2(_12566_));
 sg13g2_nor2b_1 _19562_ (.A(_12564_),
    .B_N(\cpu.dcache.r_data[4][5] ),
    .Y(_12568_));
 sg13g2_a21oi_1 _19563_ (.A1(net991),
    .A2(_12564_),
    .Y(_12569_),
    .B1(_12568_));
 sg13g2_nand2_1 _19564_ (.Y(_12570_),
    .A(net1003),
    .B(_12471_));
 sg13g2_o21ai_1 _19565_ (.B1(_12570_),
    .Y(_00473_),
    .A1(net50),
    .A2(_12569_));
 sg13g2_mux2_1 _19566_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(_11925_),
    .S(_12564_),
    .X(_12571_));
 sg13g2_nor2_1 _19567_ (.A(_12471_),
    .B(_12571_),
    .Y(_12572_));
 sg13g2_a21oi_1 _19568_ (.A1(net756),
    .A2(net50),
    .Y(_00474_),
    .B1(_12572_));
 sg13g2_mux2_1 _19569_ (.A0(\cpu.dcache.r_data[4][7] ),
    .A1(_12452_),
    .S(_12564_),
    .X(_12573_));
 sg13g2_nor2_1 _19570_ (.A(_12471_),
    .B(_12573_),
    .Y(_12574_));
 sg13g2_a21oi_1 _19571_ (.A1(net755),
    .A2(net50),
    .Y(_00475_),
    .B1(_12574_));
 sg13g2_nor2b_1 _19572_ (.A(_12482_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_12575_));
 sg13g2_a21oi_1 _19573_ (.A1(_12419_),
    .A2(_12482_),
    .Y(_12576_),
    .B1(_12575_));
 sg13g2_nand2_1 _19574_ (.Y(_12577_),
    .A(net497),
    .B(_12479_));
 sg13g2_o21ai_1 _19575_ (.B1(_12577_),
    .Y(_00476_),
    .A1(net49),
    .A2(_12576_));
 sg13g2_nor2b_1 _19576_ (.A(_12482_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_12578_));
 sg13g2_a21oi_1 _19577_ (.A1(_12425_),
    .A2(_12482_),
    .Y(_12579_),
    .B1(_12578_));
 sg13g2_nand2_1 _19578_ (.Y(_12580_),
    .A(net496),
    .B(_12479_));
 sg13g2_o21ai_1 _19579_ (.B1(_12580_),
    .Y(_00477_),
    .A1(net49),
    .A2(_12579_));
 sg13g2_buf_1 _19580_ (.A(_09395_),
    .X(_12581_));
 sg13g2_nor2_1 _19581_ (.A(net754),
    .B(_12099_),
    .Y(_12582_));
 sg13g2_buf_2 _19582_ (.A(_12582_),
    .X(_12583_));
 sg13g2_buf_1 _19583_ (.A(_12583_),
    .X(_12584_));
 sg13g2_buf_1 _19584_ (.A(_11903_),
    .X(_12585_));
 sg13g2_nor2_1 _19585_ (.A(_09395_),
    .B(_11913_),
    .Y(_12586_));
 sg13g2_buf_2 _19586_ (.A(_12586_),
    .X(_12587_));
 sg13g2_nor2b_1 _19587_ (.A(_12587_),
    .B_N(\cpu.dcache.r_data[5][0] ),
    .Y(_12588_));
 sg13g2_a21oi_1 _19588_ (.A1(net1091),
    .A2(_12587_),
    .Y(_12589_),
    .B1(_12588_));
 sg13g2_nand2_1 _19589_ (.Y(_12590_),
    .A(_12269_),
    .B(_12584_));
 sg13g2_o21ai_1 _19590_ (.B1(_12590_),
    .Y(_00478_),
    .A1(_12584_),
    .A2(_12589_));
 sg13g2_nor2_1 _19591_ (.A(net754),
    .B(_12109_),
    .Y(_12591_));
 sg13g2_buf_2 _19592_ (.A(_12591_),
    .X(_12592_));
 sg13g2_buf_1 _19593_ (.A(_12592_),
    .X(_12593_));
 sg13g2_nor2_1 _19594_ (.A(_12581_),
    .B(_11928_),
    .Y(_12594_));
 sg13g2_buf_2 _19595_ (.A(_12594_),
    .X(_12595_));
 sg13g2_nor2b_1 _19596_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_12596_));
 sg13g2_a21oi_1 _19597_ (.A1(net989),
    .A2(_12595_),
    .Y(_12597_),
    .B1(_12596_));
 sg13g2_nand2_1 _19598_ (.Y(_12598_),
    .A(_11936_),
    .B(net46));
 sg13g2_o21ai_1 _19599_ (.B1(_12598_),
    .Y(_00479_),
    .A1(net46),
    .A2(_12597_));
 sg13g2_nor2b_1 _19600_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_12599_));
 sg13g2_a21oi_1 _19601_ (.A1(net990),
    .A2(_12595_),
    .Y(_12600_),
    .B1(_12599_));
 sg13g2_nand2_1 _19602_ (.Y(_12601_),
    .A(net495),
    .B(net46));
 sg13g2_o21ai_1 _19603_ (.B1(_12601_),
    .Y(_00480_),
    .A1(net46),
    .A2(_12600_));
 sg13g2_nor2_1 _19604_ (.A(_12581_),
    .B(_11950_),
    .Y(_12602_));
 sg13g2_buf_2 _19605_ (.A(_12602_),
    .X(_12603_));
 sg13g2_nor2b_1 _19606_ (.A(_12603_),
    .B_N(\cpu.dcache.r_data[5][12] ),
    .Y(_12604_));
 sg13g2_a21oi_1 _19607_ (.A1(net1091),
    .A2(_12603_),
    .Y(_12605_),
    .B1(_12604_));
 sg13g2_nand2_1 _19608_ (.Y(_12606_),
    .A(net494),
    .B(_12592_));
 sg13g2_o21ai_1 _19609_ (.B1(_12606_),
    .Y(_00481_),
    .A1(net46),
    .A2(_12605_));
 sg13g2_buf_1 _19610_ (.A(_11958_),
    .X(_12607_));
 sg13g2_nor2b_1 _19611_ (.A(_12603_),
    .B_N(\cpu.dcache.r_data[5][13] ),
    .Y(_12608_));
 sg13g2_a21oi_1 _19612_ (.A1(net1090),
    .A2(_12603_),
    .Y(_12609_),
    .B1(_12608_));
 sg13g2_nand2_1 _19613_ (.Y(_12610_),
    .A(net493),
    .B(_12592_));
 sg13g2_o21ai_1 _19614_ (.B1(_12610_),
    .Y(_00482_),
    .A1(_12593_),
    .A2(_12609_));
 sg13g2_nor2b_1 _19615_ (.A(_12603_),
    .B_N(\cpu.dcache.r_data[5][14] ),
    .Y(_12611_));
 sg13g2_a21oi_1 _19616_ (.A1(net989),
    .A2(_12603_),
    .Y(_12612_),
    .B1(_12611_));
 sg13g2_nand2_1 _19617_ (.Y(_12613_),
    .A(net492),
    .B(_12592_));
 sg13g2_o21ai_1 _19618_ (.B1(_12613_),
    .Y(_00483_),
    .A1(net46),
    .A2(_12612_));
 sg13g2_nor2b_1 _19619_ (.A(_12603_),
    .B_N(\cpu.dcache.r_data[5][15] ),
    .Y(_12614_));
 sg13g2_a21oi_1 _19620_ (.A1(net990),
    .A2(_12603_),
    .Y(_12615_),
    .B1(_12614_));
 sg13g2_nand2_1 _19621_ (.Y(_12616_),
    .A(net491),
    .B(_12592_));
 sg13g2_o21ai_1 _19622_ (.B1(_12616_),
    .Y(_00484_),
    .A1(_12593_),
    .A2(_12615_));
 sg13g2_nor2_1 _19623_ (.A(net754),
    .B(_12137_),
    .Y(_12617_));
 sg13g2_buf_2 _19624_ (.A(_12617_),
    .X(_12618_));
 sg13g2_buf_1 _19625_ (.A(_12618_),
    .X(_12619_));
 sg13g2_nor2_1 _19626_ (.A(_09395_),
    .B(_11982_),
    .Y(_12620_));
 sg13g2_buf_2 _19627_ (.A(_12620_),
    .X(_12621_));
 sg13g2_nor2b_1 _19628_ (.A(_12621_),
    .B_N(\cpu.dcache.r_data[5][16] ),
    .Y(_12622_));
 sg13g2_a21oi_1 _19629_ (.A1(net1091),
    .A2(_12621_),
    .Y(_12623_),
    .B1(_12622_));
 sg13g2_nand2_1 _19630_ (.Y(_12624_),
    .A(net869),
    .B(_12619_));
 sg13g2_o21ai_1 _19631_ (.B1(_12624_),
    .Y(_00485_),
    .A1(net45),
    .A2(_12623_));
 sg13g2_nor2b_1 _19632_ (.A(_12621_),
    .B_N(\cpu.dcache.r_data[5][17] ),
    .Y(_12625_));
 sg13g2_a21oi_1 _19633_ (.A1(net1090),
    .A2(_12621_),
    .Y(_12626_),
    .B1(_12625_));
 sg13g2_nand2_1 _19634_ (.Y(_12627_),
    .A(net868),
    .B(net45));
 sg13g2_o21ai_1 _19635_ (.B1(_12627_),
    .Y(_00486_),
    .A1(net45),
    .A2(_12626_));
 sg13g2_nor2b_1 _19636_ (.A(_12621_),
    .B_N(\cpu.dcache.r_data[5][18] ),
    .Y(_12628_));
 sg13g2_a21oi_1 _19637_ (.A1(net989),
    .A2(_12621_),
    .Y(_12629_),
    .B1(_12628_));
 sg13g2_nand2_1 _19638_ (.Y(_12630_),
    .A(net867),
    .B(_12618_));
 sg13g2_o21ai_1 _19639_ (.B1(_12630_),
    .Y(_00487_),
    .A1(net45),
    .A2(_12629_));
 sg13g2_buf_1 _19640_ (.A(_11996_),
    .X(_12631_));
 sg13g2_mux2_1 _19641_ (.A0(\cpu.dcache.r_data[5][19] ),
    .A1(net1092),
    .S(_12621_),
    .X(_12632_));
 sg13g2_nor2_1 _19642_ (.A(_12618_),
    .B(_12632_),
    .Y(_12633_));
 sg13g2_a21oi_1 _19643_ (.A1(net866),
    .A2(_12619_),
    .Y(_00488_),
    .B1(_12633_));
 sg13g2_nor2b_1 _19644_ (.A(_12587_),
    .B_N(\cpu.dcache.r_data[5][1] ),
    .Y(_12634_));
 sg13g2_a21oi_1 _19645_ (.A1(net1090),
    .A2(_12587_),
    .Y(_12635_),
    .B1(_12634_));
 sg13g2_nand2_1 _19646_ (.Y(_12636_),
    .A(net868),
    .B(net47));
 sg13g2_o21ai_1 _19647_ (.B1(_12636_),
    .Y(_00489_),
    .A1(net47),
    .A2(_12635_));
 sg13g2_nor2_1 _19648_ (.A(net754),
    .B(_12006_),
    .Y(_12637_));
 sg13g2_buf_2 _19649_ (.A(_12637_),
    .X(_12638_));
 sg13g2_nor2b_1 _19650_ (.A(_12638_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_12639_));
 sg13g2_a21oi_1 _19651_ (.A1(net1091),
    .A2(_12638_),
    .Y(_12640_),
    .B1(_12639_));
 sg13g2_nand2_1 _19652_ (.Y(_12641_),
    .A(net1004),
    .B(_12618_));
 sg13g2_o21ai_1 _19653_ (.B1(_12641_),
    .Y(_00490_),
    .A1(net45),
    .A2(_12640_));
 sg13g2_nor2b_1 _19654_ (.A(_12638_),
    .B_N(\cpu.dcache.r_data[5][21] ),
    .Y(_12642_));
 sg13g2_a21oi_1 _19655_ (.A1(net1090),
    .A2(_12638_),
    .Y(_12643_),
    .B1(_12642_));
 sg13g2_nand2_1 _19656_ (.Y(_12644_),
    .A(net1003),
    .B(_12618_));
 sg13g2_o21ai_1 _19657_ (.B1(_12644_),
    .Y(_00491_),
    .A1(net45),
    .A2(_12643_));
 sg13g2_buf_1 _19658_ (.A(_12018_),
    .X(_12645_));
 sg13g2_mux2_1 _19659_ (.A0(\cpu.dcache.r_data[5][22] ),
    .A1(net1097),
    .S(_12638_),
    .X(_12646_));
 sg13g2_nor2_1 _19660_ (.A(_12618_),
    .B(_12646_),
    .Y(_12647_));
 sg13g2_a21oi_1 _19661_ (.A1(net753),
    .A2(net45),
    .Y(_00492_),
    .B1(_12647_));
 sg13g2_buf_1 _19662_ (.A(_12024_),
    .X(_12648_));
 sg13g2_mux2_1 _19663_ (.A0(\cpu.dcache.r_data[5][23] ),
    .A1(net1092),
    .S(_12638_),
    .X(_12649_));
 sg13g2_nor2_1 _19664_ (.A(_12618_),
    .B(_12649_),
    .Y(_12650_));
 sg13g2_a21oi_1 _19665_ (.A1(net752),
    .A2(net45),
    .Y(_00493_),
    .B1(_12650_));
 sg13g2_nor2_1 _19666_ (.A(net754),
    .B(_12170_),
    .Y(_12651_));
 sg13g2_buf_2 _19667_ (.A(_12651_),
    .X(_12652_));
 sg13g2_buf_1 _19668_ (.A(_12652_),
    .X(_12653_));
 sg13g2_nor2_1 _19669_ (.A(net754),
    .B(net617),
    .Y(_12654_));
 sg13g2_buf_1 _19670_ (.A(_12654_),
    .X(_12655_));
 sg13g2_nor2b_1 _19671_ (.A(net487),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_12656_));
 sg13g2_a21oi_1 _19672_ (.A1(net1091),
    .A2(net487),
    .Y(_12657_),
    .B1(_12656_));
 sg13g2_nand2_1 _19673_ (.Y(_12658_),
    .A(net497),
    .B(net44));
 sg13g2_o21ai_1 _19674_ (.B1(_12658_),
    .Y(_00494_),
    .A1(net44),
    .A2(_12657_));
 sg13g2_nor2b_1 _19675_ (.A(net487),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_12659_));
 sg13g2_a21oi_1 _19676_ (.A1(net1090),
    .A2(net487),
    .Y(_12660_),
    .B1(_12659_));
 sg13g2_nand2_1 _19677_ (.Y(_12661_),
    .A(net496),
    .B(net44));
 sg13g2_o21ai_1 _19678_ (.B1(_12661_),
    .Y(_00495_),
    .A1(net44),
    .A2(_12660_));
 sg13g2_nor2b_1 _19679_ (.A(net487),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_12662_));
 sg13g2_a21oi_1 _19680_ (.A1(net989),
    .A2(net487),
    .Y(_12663_),
    .B1(_12662_));
 sg13g2_nand2_1 _19681_ (.Y(_12664_),
    .A(_11936_),
    .B(_12652_));
 sg13g2_o21ai_1 _19682_ (.B1(_12664_),
    .Y(_00496_),
    .A1(net44),
    .A2(_12663_));
 sg13g2_nor2b_1 _19683_ (.A(net487),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_12665_));
 sg13g2_a21oi_1 _19684_ (.A1(net990),
    .A2(net487),
    .Y(_12666_),
    .B1(_12665_));
 sg13g2_nand2_1 _19685_ (.Y(_12667_),
    .A(_11945_),
    .B(_12652_));
 sg13g2_o21ai_1 _19686_ (.B1(_12667_),
    .Y(_00497_),
    .A1(net44),
    .A2(_12666_));
 sg13g2_nor2_1 _19687_ (.A(net754),
    .B(_12048_),
    .Y(_12668_));
 sg13g2_buf_2 _19688_ (.A(_12668_),
    .X(_12669_));
 sg13g2_nor2b_1 _19689_ (.A(_12669_),
    .B_N(\cpu.dcache.r_data[5][28] ),
    .Y(_12670_));
 sg13g2_a21oi_1 _19690_ (.A1(net1091),
    .A2(_12669_),
    .Y(_12671_),
    .B1(_12670_));
 sg13g2_nand2_1 _19691_ (.Y(_12672_),
    .A(_11956_),
    .B(_12652_));
 sg13g2_o21ai_1 _19692_ (.B1(_12672_),
    .Y(_00498_),
    .A1(_12653_),
    .A2(_12671_));
 sg13g2_nor2b_1 _19693_ (.A(_12669_),
    .B_N(\cpu.dcache.r_data[5][29] ),
    .Y(_12673_));
 sg13g2_a21oi_1 _19694_ (.A1(net1090),
    .A2(_12669_),
    .Y(_12674_),
    .B1(_12673_));
 sg13g2_nand2_1 _19695_ (.Y(_12675_),
    .A(_11964_),
    .B(_12652_));
 sg13g2_o21ai_1 _19696_ (.B1(_12675_),
    .Y(_00499_),
    .A1(net44),
    .A2(_12674_));
 sg13g2_nor2b_1 _19697_ (.A(_12587_),
    .B_N(\cpu.dcache.r_data[5][2] ),
    .Y(_12676_));
 sg13g2_a21oi_1 _19698_ (.A1(net989),
    .A2(_12587_),
    .Y(_12677_),
    .B1(_12676_));
 sg13g2_nand2_1 _19699_ (.Y(_12678_),
    .A(net867),
    .B(_12583_));
 sg13g2_o21ai_1 _19700_ (.B1(_12678_),
    .Y(_00500_),
    .A1(net47),
    .A2(_12677_));
 sg13g2_nor2b_1 _19701_ (.A(_12669_),
    .B_N(\cpu.dcache.r_data[5][30] ),
    .Y(_12679_));
 sg13g2_a21oi_1 _19702_ (.A1(_12551_),
    .A2(_12669_),
    .Y(_12680_),
    .B1(_12679_));
 sg13g2_nand2_1 _19703_ (.Y(_12681_),
    .A(_11969_),
    .B(_12652_));
 sg13g2_o21ai_1 _19704_ (.B1(_12681_),
    .Y(_00501_),
    .A1(_12653_),
    .A2(_12680_));
 sg13g2_nor2b_1 _19705_ (.A(_12669_),
    .B_N(\cpu.dcache.r_data[5][31] ),
    .Y(_12682_));
 sg13g2_a21oi_1 _19706_ (.A1(net990),
    .A2(_12669_),
    .Y(_12683_),
    .B1(_12682_));
 sg13g2_nand2_1 _19707_ (.Y(_12684_),
    .A(_11974_),
    .B(_12652_));
 sg13g2_o21ai_1 _19708_ (.B1(_12684_),
    .Y(_00502_),
    .A1(net44),
    .A2(_12683_));
 sg13g2_mux2_1 _19709_ (.A0(\cpu.dcache.r_data[5][3] ),
    .A1(net1092),
    .S(_12587_),
    .X(_12685_));
 sg13g2_nor2_1 _19710_ (.A(_12583_),
    .B(_12685_),
    .Y(_12686_));
 sg13g2_a21oi_1 _19711_ (.A1(net866),
    .A2(net47),
    .Y(_00503_),
    .B1(_12686_));
 sg13g2_nor2_1 _19712_ (.A(_09395_),
    .B(_12073_),
    .Y(_12687_));
 sg13g2_buf_2 _19713_ (.A(_12687_),
    .X(_12688_));
 sg13g2_nor2b_1 _19714_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_12689_));
 sg13g2_a21oi_1 _19715_ (.A1(net1091),
    .A2(_12688_),
    .Y(_12690_),
    .B1(_12689_));
 sg13g2_nand2_1 _19716_ (.Y(_12691_),
    .A(_12078_),
    .B(_12583_));
 sg13g2_o21ai_1 _19717_ (.B1(_12691_),
    .Y(_00504_),
    .A1(net47),
    .A2(_12690_));
 sg13g2_nor2b_1 _19718_ (.A(_12688_),
    .B_N(\cpu.dcache.r_data[5][5] ),
    .Y(_12692_));
 sg13g2_a21oi_1 _19719_ (.A1(net1090),
    .A2(_12688_),
    .Y(_12693_),
    .B1(_12692_));
 sg13g2_nand2_1 _19720_ (.Y(_12694_),
    .A(_12082_),
    .B(_12583_));
 sg13g2_o21ai_1 _19721_ (.B1(_12694_),
    .Y(_00505_),
    .A1(net47),
    .A2(_12693_));
 sg13g2_mux2_1 _19722_ (.A0(\cpu.dcache.r_data[5][6] ),
    .A1(net1097),
    .S(_12688_),
    .X(_12695_));
 sg13g2_nor2_1 _19723_ (.A(_12583_),
    .B(_12695_),
    .Y(_12696_));
 sg13g2_a21oi_1 _19724_ (.A1(net753),
    .A2(net47),
    .Y(_00506_),
    .B1(_12696_));
 sg13g2_mux2_1 _19725_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(_12452_),
    .S(_12688_),
    .X(_12697_));
 sg13g2_nor2_1 _19726_ (.A(_12583_),
    .B(_12697_),
    .Y(_12698_));
 sg13g2_a21oi_1 _19727_ (.A1(net752),
    .A2(net47),
    .Y(_00507_),
    .B1(_12698_));
 sg13g2_nor2b_1 _19728_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_12699_));
 sg13g2_a21oi_1 _19729_ (.A1(_12585_),
    .A2(_12595_),
    .Y(_12700_),
    .B1(_12699_));
 sg13g2_nand2_1 _19730_ (.Y(_12701_),
    .A(_12033_),
    .B(_12592_));
 sg13g2_o21ai_1 _19731_ (.B1(_12701_),
    .Y(_00508_),
    .A1(net46),
    .A2(_12700_));
 sg13g2_nor2b_1 _19732_ (.A(_12595_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_12702_));
 sg13g2_a21oi_1 _19733_ (.A1(_12607_),
    .A2(_12595_),
    .Y(_12703_),
    .B1(_12702_));
 sg13g2_nand2_1 _19734_ (.Y(_12704_),
    .A(_12041_),
    .B(_12592_));
 sg13g2_o21ai_1 _19735_ (.B1(_12704_),
    .Y(_00509_),
    .A1(net46),
    .A2(_12703_));
 sg13g2_buf_1 _19736_ (.A(_09400_),
    .X(_12705_));
 sg13g2_nor2_1 _19737_ (.A(net677),
    .B(_12099_),
    .Y(_12706_));
 sg13g2_buf_1 _19738_ (.A(_12706_),
    .X(_12707_));
 sg13g2_buf_1 _19739_ (.A(_12707_),
    .X(_12708_));
 sg13g2_nor2_1 _19740_ (.A(_09400_),
    .B(_11913_),
    .Y(_12709_));
 sg13g2_buf_2 _19741_ (.A(_12709_),
    .X(_12710_));
 sg13g2_nor2b_1 _19742_ (.A(_12710_),
    .B_N(\cpu.dcache.r_data[6][0] ),
    .Y(_12711_));
 sg13g2_a21oi_1 _19743_ (.A1(net1091),
    .A2(_12710_),
    .Y(_12712_),
    .B1(_12711_));
 sg13g2_nand2_1 _19744_ (.Y(_12713_),
    .A(net869),
    .B(_12708_));
 sg13g2_o21ai_1 _19745_ (.B1(_12713_),
    .Y(_00510_),
    .A1(net43),
    .A2(_12712_));
 sg13g2_nor2_1 _19746_ (.A(net677),
    .B(_12109_),
    .Y(_12714_));
 sg13g2_buf_2 _19747_ (.A(_12714_),
    .X(_12715_));
 sg13g2_buf_1 _19748_ (.A(_12715_),
    .X(_12716_));
 sg13g2_nor2_1 _19749_ (.A(_12705_),
    .B(_11928_),
    .Y(_12717_));
 sg13g2_buf_2 _19750_ (.A(_12717_),
    .X(_12718_));
 sg13g2_nor2b_1 _19751_ (.A(_12718_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_12719_));
 sg13g2_a21oi_1 _19752_ (.A1(net989),
    .A2(_12718_),
    .Y(_12720_),
    .B1(_12719_));
 sg13g2_nand2_1 _19753_ (.Y(_12721_),
    .A(_11936_),
    .B(net42));
 sg13g2_o21ai_1 _19754_ (.B1(_12721_),
    .Y(_00511_),
    .A1(net42),
    .A2(_12720_));
 sg13g2_nor2b_1 _19755_ (.A(_12718_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_12722_));
 sg13g2_a21oi_1 _19756_ (.A1(net990),
    .A2(_12718_),
    .Y(_12723_),
    .B1(_12722_));
 sg13g2_nand2_1 _19757_ (.Y(_12724_),
    .A(_11945_),
    .B(net42));
 sg13g2_o21ai_1 _19758_ (.B1(_12724_),
    .Y(_00512_),
    .A1(net42),
    .A2(_12723_));
 sg13g2_nor2_1 _19759_ (.A(net677),
    .B(_11950_),
    .Y(_12725_));
 sg13g2_buf_2 _19760_ (.A(_12725_),
    .X(_12726_));
 sg13g2_nor2b_1 _19761_ (.A(_12726_),
    .B_N(\cpu.dcache.r_data[6][12] ),
    .Y(_12727_));
 sg13g2_a21oi_1 _19762_ (.A1(_12585_),
    .A2(_12726_),
    .Y(_12728_),
    .B1(_12727_));
 sg13g2_nand2_1 _19763_ (.Y(_12729_),
    .A(_11956_),
    .B(_12715_));
 sg13g2_o21ai_1 _19764_ (.B1(_12729_),
    .Y(_00513_),
    .A1(net42),
    .A2(_12728_));
 sg13g2_nor2b_1 _19765_ (.A(_12726_),
    .B_N(\cpu.dcache.r_data[6][13] ),
    .Y(_12730_));
 sg13g2_a21oi_1 _19766_ (.A1(_12607_),
    .A2(_12726_),
    .Y(_12731_),
    .B1(_12730_));
 sg13g2_nand2_1 _19767_ (.Y(_12732_),
    .A(_11964_),
    .B(_12715_));
 sg13g2_o21ai_1 _19768_ (.B1(_12732_),
    .Y(_00514_),
    .A1(net42),
    .A2(_12731_));
 sg13g2_nor2b_1 _19769_ (.A(_12726_),
    .B_N(\cpu.dcache.r_data[6][14] ),
    .Y(_12733_));
 sg13g2_a21oi_1 _19770_ (.A1(_12551_),
    .A2(_12726_),
    .Y(_12734_),
    .B1(_12733_));
 sg13g2_nand2_1 _19771_ (.Y(_12735_),
    .A(_11969_),
    .B(_12715_));
 sg13g2_o21ai_1 _19772_ (.B1(_12735_),
    .Y(_00515_),
    .A1(_12716_),
    .A2(_12734_));
 sg13g2_nor2b_1 _19773_ (.A(_12726_),
    .B_N(\cpu.dcache.r_data[6][15] ),
    .Y(_12736_));
 sg13g2_a21oi_1 _19774_ (.A1(net990),
    .A2(_12726_),
    .Y(_12737_),
    .B1(_12736_));
 sg13g2_nand2_1 _19775_ (.Y(_12738_),
    .A(_11974_),
    .B(_12715_));
 sg13g2_o21ai_1 _19776_ (.B1(_12738_),
    .Y(_00516_),
    .A1(_12716_),
    .A2(_12737_));
 sg13g2_nor2_1 _19777_ (.A(net677),
    .B(_12137_),
    .Y(_12739_));
 sg13g2_buf_1 _19778_ (.A(_12739_),
    .X(_12740_));
 sg13g2_buf_1 _19779_ (.A(_12740_),
    .X(_02676_));
 sg13g2_buf_1 _19780_ (.A(_11903_),
    .X(_02677_));
 sg13g2_nor2_1 _19781_ (.A(_09400_),
    .B(_11982_),
    .Y(_02678_));
 sg13g2_buf_2 _19782_ (.A(_02678_),
    .X(_02679_));
 sg13g2_nor2b_1 _19783_ (.A(_02679_),
    .B_N(\cpu.dcache.r_data[6][16] ),
    .Y(_02680_));
 sg13g2_a21oi_1 _19784_ (.A1(net1089),
    .A2(_02679_),
    .Y(_02681_),
    .B1(_02680_));
 sg13g2_nand2_1 _19785_ (.Y(_02682_),
    .A(net869),
    .B(net41));
 sg13g2_o21ai_1 _19786_ (.B1(_02682_),
    .Y(_00517_),
    .A1(net41),
    .A2(_02681_));
 sg13g2_nor2b_1 _19787_ (.A(_02679_),
    .B_N(\cpu.dcache.r_data[6][17] ),
    .Y(_02683_));
 sg13g2_a21oi_1 _19788_ (.A1(net1090),
    .A2(_02679_),
    .Y(_02684_),
    .B1(_02683_));
 sg13g2_nand2_1 _19789_ (.Y(_02685_),
    .A(net868),
    .B(_02676_));
 sg13g2_o21ai_1 _19790_ (.B1(_02685_),
    .Y(_00518_),
    .A1(_02676_),
    .A2(_02684_));
 sg13g2_buf_1 _19791_ (.A(_11924_),
    .X(_02686_));
 sg13g2_nor2b_1 _19792_ (.A(_02679_),
    .B_N(\cpu.dcache.r_data[6][18] ),
    .Y(_02687_));
 sg13g2_a21oi_1 _19793_ (.A1(net1088),
    .A2(_02679_),
    .Y(_02688_),
    .B1(_02687_));
 sg13g2_nand2_1 _19794_ (.Y(_02689_),
    .A(net867),
    .B(_12740_));
 sg13g2_o21ai_1 _19795_ (.B1(_02689_),
    .Y(_00519_),
    .A1(net41),
    .A2(_02688_));
 sg13g2_mux2_1 _19796_ (.A0(\cpu.dcache.r_data[6][19] ),
    .A1(net1092),
    .S(_02679_),
    .X(_02690_));
 sg13g2_nor2_1 _19797_ (.A(_12740_),
    .B(_02690_),
    .Y(_02691_));
 sg13g2_a21oi_1 _19798_ (.A1(net866),
    .A2(net41),
    .Y(_00520_),
    .B1(_02691_));
 sg13g2_buf_1 _19799_ (.A(_11958_),
    .X(_02692_));
 sg13g2_nor2b_1 _19800_ (.A(_12710_),
    .B_N(\cpu.dcache.r_data[6][1] ),
    .Y(_02693_));
 sg13g2_a21oi_1 _19801_ (.A1(net1087),
    .A2(_12710_),
    .Y(_02694_),
    .B1(_02693_));
 sg13g2_nand2_1 _19802_ (.Y(_02695_),
    .A(_12282_),
    .B(net43));
 sg13g2_o21ai_1 _19803_ (.B1(_02695_),
    .Y(_00521_),
    .A1(net43),
    .A2(_02694_));
 sg13g2_nor2_1 _19804_ (.A(net677),
    .B(_12006_),
    .Y(_02696_));
 sg13g2_buf_2 _19805_ (.A(_02696_),
    .X(_02697_));
 sg13g2_nor2b_1 _19806_ (.A(_02697_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02698_));
 sg13g2_a21oi_1 _19807_ (.A1(net1089),
    .A2(_02697_),
    .Y(_02699_),
    .B1(_02698_));
 sg13g2_nand2_1 _19808_ (.Y(_02700_),
    .A(net1004),
    .B(_12740_));
 sg13g2_o21ai_1 _19809_ (.B1(_02700_),
    .Y(_00522_),
    .A1(net41),
    .A2(_02699_));
 sg13g2_nor2b_1 _19810_ (.A(_02697_),
    .B_N(\cpu.dcache.r_data[6][21] ),
    .Y(_02701_));
 sg13g2_a21oi_1 _19811_ (.A1(net1087),
    .A2(_02697_),
    .Y(_02702_),
    .B1(_02701_));
 sg13g2_nand2_1 _19812_ (.Y(_02703_),
    .A(net1003),
    .B(_12740_));
 sg13g2_o21ai_1 _19813_ (.B1(_02703_),
    .Y(_00523_),
    .A1(net41),
    .A2(_02702_));
 sg13g2_mux2_1 _19814_ (.A0(\cpu.dcache.r_data[6][22] ),
    .A1(net1097),
    .S(_02697_),
    .X(_02704_));
 sg13g2_nor2_1 _19815_ (.A(_12740_),
    .B(_02704_),
    .Y(_02705_));
 sg13g2_a21oi_1 _19816_ (.A1(net753),
    .A2(net41),
    .Y(_00524_),
    .B1(_02705_));
 sg13g2_mux2_1 _19817_ (.A0(\cpu.dcache.r_data[6][23] ),
    .A1(net1096),
    .S(_02697_),
    .X(_02706_));
 sg13g2_nor2_1 _19818_ (.A(_12740_),
    .B(_02706_),
    .Y(_02707_));
 sg13g2_a21oi_1 _19819_ (.A1(_12648_),
    .A2(net41),
    .Y(_00525_),
    .B1(_02707_));
 sg13g2_nor2_1 _19820_ (.A(net677),
    .B(_12170_),
    .Y(_02708_));
 sg13g2_buf_2 _19821_ (.A(_02708_),
    .X(_02709_));
 sg13g2_buf_1 _19822_ (.A(_02709_),
    .X(_02710_));
 sg13g2_nor2_1 _19823_ (.A(net677),
    .B(net617),
    .Y(_02711_));
 sg13g2_buf_1 _19824_ (.A(_02711_),
    .X(_02712_));
 sg13g2_nor2b_1 _19825_ (.A(net486),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02713_));
 sg13g2_a21oi_1 _19826_ (.A1(net1089),
    .A2(net486),
    .Y(_02714_),
    .B1(_02713_));
 sg13g2_nand2_1 _19827_ (.Y(_02715_),
    .A(_12033_),
    .B(net40));
 sg13g2_o21ai_1 _19828_ (.B1(_02715_),
    .Y(_00526_),
    .A1(net40),
    .A2(_02714_));
 sg13g2_nor2b_1 _19829_ (.A(net486),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02716_));
 sg13g2_a21oi_1 _19830_ (.A1(net1087),
    .A2(net486),
    .Y(_02717_),
    .B1(_02716_));
 sg13g2_nand2_1 _19831_ (.Y(_02718_),
    .A(_12041_),
    .B(_02710_));
 sg13g2_o21ai_1 _19832_ (.B1(_02718_),
    .Y(_00527_),
    .A1(net40),
    .A2(_02717_));
 sg13g2_nor2b_1 _19833_ (.A(net486),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02719_));
 sg13g2_a21oi_1 _19834_ (.A1(net1088),
    .A2(net486),
    .Y(_02720_),
    .B1(_02719_));
 sg13g2_nand2_1 _19835_ (.Y(_02721_),
    .A(_11936_),
    .B(_02709_));
 sg13g2_o21ai_1 _19836_ (.B1(_02721_),
    .Y(_00528_),
    .A1(net40),
    .A2(_02720_));
 sg13g2_nor2b_1 _19837_ (.A(net486),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02722_));
 sg13g2_a21oi_1 _19838_ (.A1(_12500_),
    .A2(net486),
    .Y(_02723_),
    .B1(_02722_));
 sg13g2_nand2_1 _19839_ (.Y(_02724_),
    .A(_11945_),
    .B(_02709_));
 sg13g2_o21ai_1 _19840_ (.B1(_02724_),
    .Y(_00529_),
    .A1(net40),
    .A2(_02723_));
 sg13g2_nor2_1 _19841_ (.A(_12705_),
    .B(_12048_),
    .Y(_02725_));
 sg13g2_buf_2 _19842_ (.A(_02725_),
    .X(_02726_));
 sg13g2_nor2b_1 _19843_ (.A(_02726_),
    .B_N(\cpu.dcache.r_data[6][28] ),
    .Y(_02727_));
 sg13g2_a21oi_1 _19844_ (.A1(net1089),
    .A2(_02726_),
    .Y(_02728_),
    .B1(_02727_));
 sg13g2_nand2_1 _19845_ (.Y(_02729_),
    .A(_11956_),
    .B(_02709_));
 sg13g2_o21ai_1 _19846_ (.B1(_02729_),
    .Y(_00530_),
    .A1(_02710_),
    .A2(_02728_));
 sg13g2_nor2b_1 _19847_ (.A(_02726_),
    .B_N(\cpu.dcache.r_data[6][29] ),
    .Y(_02730_));
 sg13g2_a21oi_1 _19848_ (.A1(net1087),
    .A2(_02726_),
    .Y(_02731_),
    .B1(_02730_));
 sg13g2_nand2_1 _19849_ (.Y(_02732_),
    .A(_11964_),
    .B(_02709_));
 sg13g2_o21ai_1 _19850_ (.B1(_02732_),
    .Y(_00531_),
    .A1(net40),
    .A2(_02731_));
 sg13g2_nor2b_1 _19851_ (.A(_12710_),
    .B_N(\cpu.dcache.r_data[6][2] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _19852_ (.A1(net1088),
    .A2(_12710_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2_1 _19853_ (.Y(_02735_),
    .A(net867),
    .B(_12707_));
 sg13g2_o21ai_1 _19854_ (.B1(_02735_),
    .Y(_00532_),
    .A1(_12708_),
    .A2(_02734_));
 sg13g2_nor2b_1 _19855_ (.A(_02726_),
    .B_N(\cpu.dcache.r_data[6][30] ),
    .Y(_02736_));
 sg13g2_a21oi_1 _19856_ (.A1(net1088),
    .A2(_02726_),
    .Y(_02737_),
    .B1(_02736_));
 sg13g2_nand2_1 _19857_ (.Y(_02738_),
    .A(_11969_),
    .B(_02709_));
 sg13g2_o21ai_1 _19858_ (.B1(_02738_),
    .Y(_00533_),
    .A1(net40),
    .A2(_02737_));
 sg13g2_nor2b_1 _19859_ (.A(_02726_),
    .B_N(\cpu.dcache.r_data[6][31] ),
    .Y(_02739_));
 sg13g2_a21oi_1 _19860_ (.A1(_12500_),
    .A2(_02726_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_nand2_1 _19861_ (.Y(_02741_),
    .A(_11974_),
    .B(_02709_));
 sg13g2_o21ai_1 _19862_ (.B1(_02741_),
    .Y(_00534_),
    .A1(net40),
    .A2(_02740_));
 sg13g2_mux2_1 _19863_ (.A0(\cpu.dcache.r_data[6][3] ),
    .A1(net1096),
    .S(_12710_),
    .X(_02742_));
 sg13g2_nor2_1 _19864_ (.A(_12707_),
    .B(_02742_),
    .Y(_02743_));
 sg13g2_a21oi_1 _19865_ (.A1(net866),
    .A2(net43),
    .Y(_00535_),
    .B1(_02743_));
 sg13g2_nor2_1 _19866_ (.A(_09400_),
    .B(_12073_),
    .Y(_02744_));
 sg13g2_buf_2 _19867_ (.A(_02744_),
    .X(_02745_));
 sg13g2_nor2b_1 _19868_ (.A(_02745_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02746_));
 sg13g2_a21oi_1 _19869_ (.A1(net1089),
    .A2(_02745_),
    .Y(_02747_),
    .B1(_02746_));
 sg13g2_nand2_1 _19870_ (.Y(_02748_),
    .A(net1043),
    .B(_12707_));
 sg13g2_o21ai_1 _19871_ (.B1(_02748_),
    .Y(_00536_),
    .A1(net43),
    .A2(_02747_));
 sg13g2_nor2b_1 _19872_ (.A(_02745_),
    .B_N(\cpu.dcache.r_data[6][5] ),
    .Y(_02749_));
 sg13g2_a21oi_1 _19873_ (.A1(net1087),
    .A2(_02745_),
    .Y(_02750_),
    .B1(_02749_));
 sg13g2_nand2_1 _19874_ (.Y(_02751_),
    .A(net1042),
    .B(_12707_));
 sg13g2_o21ai_1 _19875_ (.B1(_02751_),
    .Y(_00537_),
    .A1(net43),
    .A2(_02750_));
 sg13g2_mux2_1 _19876_ (.A0(\cpu.dcache.r_data[6][6] ),
    .A1(_11925_),
    .S(_02745_),
    .X(_02752_));
 sg13g2_nor2_1 _19877_ (.A(_12707_),
    .B(_02752_),
    .Y(_02753_));
 sg13g2_a21oi_1 _19878_ (.A1(net753),
    .A2(net43),
    .Y(_00538_),
    .B1(_02753_));
 sg13g2_mux2_1 _19879_ (.A0(\cpu.dcache.r_data[6][7] ),
    .A1(net1096),
    .S(_02745_),
    .X(_02754_));
 sg13g2_nor2_1 _19880_ (.A(_12707_),
    .B(_02754_),
    .Y(_02755_));
 sg13g2_a21oi_1 _19881_ (.A1(net752),
    .A2(net43),
    .Y(_00539_),
    .B1(_02755_));
 sg13g2_nor2b_1 _19882_ (.A(_12718_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02756_));
 sg13g2_a21oi_1 _19883_ (.A1(net1089),
    .A2(_12718_),
    .Y(_02757_),
    .B1(_02756_));
 sg13g2_nand2_1 _19884_ (.Y(_02758_),
    .A(_12033_),
    .B(_12715_));
 sg13g2_o21ai_1 _19885_ (.B1(_02758_),
    .Y(_00540_),
    .A1(net42),
    .A2(_02757_));
 sg13g2_nor2b_1 _19886_ (.A(_12718_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02759_));
 sg13g2_a21oi_1 _19887_ (.A1(net1087),
    .A2(_12718_),
    .Y(_02760_),
    .B1(_02759_));
 sg13g2_nand2_1 _19888_ (.Y(_02761_),
    .A(_12041_),
    .B(_12715_));
 sg13g2_o21ai_1 _19889_ (.B1(_02761_),
    .Y(_00541_),
    .A1(net42),
    .A2(_02760_));
 sg13g2_buf_1 _19890_ (.A(_09906_),
    .X(_02762_));
 sg13g2_nor2_1 _19891_ (.A(net485),
    .B(_12099_),
    .Y(_02763_));
 sg13g2_buf_1 _19892_ (.A(_02763_),
    .X(_02764_));
 sg13g2_buf_1 _19893_ (.A(_02764_),
    .X(_02765_));
 sg13g2_nor2_1 _19894_ (.A(net485),
    .B(_11913_),
    .Y(_02766_));
 sg13g2_buf_2 _19895_ (.A(_02766_),
    .X(_02767_));
 sg13g2_nor2b_1 _19896_ (.A(_02767_),
    .B_N(\cpu.dcache.r_data[7][0] ),
    .Y(_02768_));
 sg13g2_a21oi_1 _19897_ (.A1(net1089),
    .A2(_02767_),
    .Y(_02769_),
    .B1(_02768_));
 sg13g2_nand2_1 _19898_ (.Y(_02770_),
    .A(net869),
    .B(_02765_));
 sg13g2_o21ai_1 _19899_ (.B1(_02770_),
    .Y(_00542_),
    .A1(net39),
    .A2(_02769_));
 sg13g2_nor2_1 _19900_ (.A(net485),
    .B(_12109_),
    .Y(_02771_));
 sg13g2_buf_2 _19901_ (.A(_02771_),
    .X(_02772_));
 sg13g2_buf_1 _19902_ (.A(_02772_),
    .X(_02773_));
 sg13g2_nor2_1 _19903_ (.A(_02762_),
    .B(_11928_),
    .Y(_02774_));
 sg13g2_buf_2 _19904_ (.A(_02774_),
    .X(_02775_));
 sg13g2_nor2b_1 _19905_ (.A(_02775_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02776_));
 sg13g2_a21oi_1 _19906_ (.A1(net1088),
    .A2(_02775_),
    .Y(_02777_),
    .B1(_02776_));
 sg13g2_nand2_1 _19907_ (.Y(_02778_),
    .A(_11936_),
    .B(net38));
 sg13g2_o21ai_1 _19908_ (.B1(_02778_),
    .Y(_00543_),
    .A1(net38),
    .A2(_02777_));
 sg13g2_buf_1 _19909_ (.A(_11940_),
    .X(_02779_));
 sg13g2_nor2b_1 _19910_ (.A(_02775_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02780_));
 sg13g2_a21oi_1 _19911_ (.A1(net988),
    .A2(_02775_),
    .Y(_02781_),
    .B1(_02780_));
 sg13g2_nand2_1 _19912_ (.Y(_02782_),
    .A(_11945_),
    .B(net38));
 sg13g2_o21ai_1 _19913_ (.B1(_02782_),
    .Y(_00544_),
    .A1(net38),
    .A2(_02781_));
 sg13g2_nor2_1 _19914_ (.A(net485),
    .B(_11950_),
    .Y(_02783_));
 sg13g2_buf_2 _19915_ (.A(_02783_),
    .X(_02784_));
 sg13g2_nor2b_1 _19916_ (.A(_02784_),
    .B_N(\cpu.dcache.r_data[7][12] ),
    .Y(_02785_));
 sg13g2_a21oi_1 _19917_ (.A1(_02677_),
    .A2(_02784_),
    .Y(_02786_),
    .B1(_02785_));
 sg13g2_nand2_1 _19918_ (.Y(_02787_),
    .A(_11956_),
    .B(_02772_));
 sg13g2_o21ai_1 _19919_ (.B1(_02787_),
    .Y(_00545_),
    .A1(net38),
    .A2(_02786_));
 sg13g2_nor2b_1 _19920_ (.A(_02784_),
    .B_N(\cpu.dcache.r_data[7][13] ),
    .Y(_02788_));
 sg13g2_a21oi_1 _19921_ (.A1(_02692_),
    .A2(_02784_),
    .Y(_02789_),
    .B1(_02788_));
 sg13g2_nand2_1 _19922_ (.Y(_02790_),
    .A(_11964_),
    .B(_02772_));
 sg13g2_o21ai_1 _19923_ (.B1(_02790_),
    .Y(_00546_),
    .A1(_02773_),
    .A2(_02789_));
 sg13g2_nor2b_1 _19924_ (.A(_02784_),
    .B_N(\cpu.dcache.r_data[7][14] ),
    .Y(_02791_));
 sg13g2_a21oi_1 _19925_ (.A1(net1088),
    .A2(_02784_),
    .Y(_02792_),
    .B1(_02791_));
 sg13g2_nand2_1 _19926_ (.Y(_02793_),
    .A(_11969_),
    .B(_02772_));
 sg13g2_o21ai_1 _19927_ (.B1(_02793_),
    .Y(_00547_),
    .A1(_02773_),
    .A2(_02792_));
 sg13g2_nor2b_1 _19928_ (.A(_02784_),
    .B_N(\cpu.dcache.r_data[7][15] ),
    .Y(_02794_));
 sg13g2_a21oi_1 _19929_ (.A1(net988),
    .A2(_02784_),
    .Y(_02795_),
    .B1(_02794_));
 sg13g2_nand2_1 _19930_ (.Y(_02796_),
    .A(_11974_),
    .B(_02772_));
 sg13g2_o21ai_1 _19931_ (.B1(_02796_),
    .Y(_00548_),
    .A1(net38),
    .A2(_02795_));
 sg13g2_nor2_1 _19932_ (.A(net485),
    .B(_12137_),
    .Y(_02797_));
 sg13g2_buf_1 _19933_ (.A(_02797_),
    .X(_02798_));
 sg13g2_buf_1 _19934_ (.A(_02798_),
    .X(_02799_));
 sg13g2_nor2_1 _19935_ (.A(net485),
    .B(_11982_),
    .Y(_02800_));
 sg13g2_buf_2 _19936_ (.A(_02800_),
    .X(_02801_));
 sg13g2_nor2b_1 _19937_ (.A(_02801_),
    .B_N(\cpu.dcache.r_data[7][16] ),
    .Y(_02802_));
 sg13g2_a21oi_1 _19938_ (.A1(net1089),
    .A2(_02801_),
    .Y(_02803_),
    .B1(_02802_));
 sg13g2_buf_1 _19939_ (.A(_09988_),
    .X(_02804_));
 sg13g2_nand2_1 _19940_ (.Y(_02805_),
    .A(_02804_),
    .B(net37));
 sg13g2_o21ai_1 _19941_ (.B1(_02805_),
    .Y(_00549_),
    .A1(net37),
    .A2(_02803_));
 sg13g2_nor2b_1 _19942_ (.A(_02801_),
    .B_N(\cpu.dcache.r_data[7][17] ),
    .Y(_02806_));
 sg13g2_a21oi_1 _19943_ (.A1(net1087),
    .A2(_02801_),
    .Y(_02807_),
    .B1(_02806_));
 sg13g2_nand2_1 _19944_ (.Y(_02808_),
    .A(net868),
    .B(_02799_));
 sg13g2_o21ai_1 _19945_ (.B1(_02808_),
    .Y(_00550_),
    .A1(net37),
    .A2(_02807_));
 sg13g2_nor2b_1 _19946_ (.A(_02801_),
    .B_N(\cpu.dcache.r_data[7][18] ),
    .Y(_02809_));
 sg13g2_a21oi_1 _19947_ (.A1(net1088),
    .A2(_02801_),
    .Y(_02810_),
    .B1(_02809_));
 sg13g2_nand2_1 _19948_ (.Y(_02811_),
    .A(net867),
    .B(_02798_));
 sg13g2_o21ai_1 _19949_ (.B1(_02811_),
    .Y(_00551_),
    .A1(_02799_),
    .A2(_02810_));
 sg13g2_mux2_1 _19950_ (.A0(\cpu.dcache.r_data[7][19] ),
    .A1(net1096),
    .S(_02801_),
    .X(_02812_));
 sg13g2_nor2_1 _19951_ (.A(_02798_),
    .B(_02812_),
    .Y(_02813_));
 sg13g2_a21oi_1 _19952_ (.A1(net866),
    .A2(net37),
    .Y(_00552_),
    .B1(_02813_));
 sg13g2_nor2b_1 _19953_ (.A(_02767_),
    .B_N(\cpu.dcache.r_data[7][1] ),
    .Y(_02814_));
 sg13g2_a21oi_1 _19954_ (.A1(net1087),
    .A2(_02767_),
    .Y(_02815_),
    .B1(_02814_));
 sg13g2_nand2_1 _19955_ (.Y(_02816_),
    .A(net1040),
    .B(net39));
 sg13g2_o21ai_1 _19956_ (.B1(_02816_),
    .Y(_00553_),
    .A1(net39),
    .A2(_02815_));
 sg13g2_or2_1 _19957_ (.X(_02817_),
    .B(_12006_),
    .A(_09906_));
 sg13g2_buf_1 _19958_ (.A(_02817_),
    .X(_02818_));
 sg13g2_mux2_1 _19959_ (.A0(net1099),
    .A1(\cpu.dcache.r_data[7][20] ),
    .S(_02818_),
    .X(_02819_));
 sg13g2_mux2_1 _19960_ (.A0(_02819_),
    .A1(net1006),
    .S(net37),
    .X(_00554_));
 sg13g2_mux2_1 _19961_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[7][21] ),
    .S(_02818_),
    .X(_02820_));
 sg13g2_mux2_1 _19962_ (.A0(_02820_),
    .A1(net1005),
    .S(net37),
    .X(_00555_));
 sg13g2_mux2_1 _19963_ (.A0(net1093),
    .A1(\cpu.dcache.r_data[7][22] ),
    .S(_02818_),
    .X(_02821_));
 sg13g2_nor2_1 _19964_ (.A(_02798_),
    .B(_02821_),
    .Y(_02822_));
 sg13g2_a21oi_1 _19965_ (.A1(net753),
    .A2(net37),
    .Y(_00556_),
    .B1(_02822_));
 sg13g2_mux2_1 _19966_ (.A0(net1094),
    .A1(\cpu.dcache.r_data[7][23] ),
    .S(_02818_),
    .X(_02823_));
 sg13g2_nor2_1 _19967_ (.A(_02798_),
    .B(_02823_),
    .Y(_02824_));
 sg13g2_a21oi_1 _19968_ (.A1(net752),
    .A2(net37),
    .Y(_00557_),
    .B1(_02824_));
 sg13g2_nor2_1 _19969_ (.A(net485),
    .B(_12170_),
    .Y(_02825_));
 sg13g2_buf_2 _19970_ (.A(_02825_),
    .X(_02826_));
 sg13g2_buf_1 _19971_ (.A(_02826_),
    .X(_02827_));
 sg13g2_nor2_1 _19972_ (.A(_09906_),
    .B(net617),
    .Y(_02828_));
 sg13g2_buf_1 _19973_ (.A(_02828_),
    .X(_02829_));
 sg13g2_nor2b_1 _19974_ (.A(net443),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02830_));
 sg13g2_a21oi_1 _19975_ (.A1(_02677_),
    .A2(net443),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_nand2_1 _19976_ (.Y(_02832_),
    .A(_12033_),
    .B(net36));
 sg13g2_o21ai_1 _19977_ (.B1(_02832_),
    .Y(_00558_),
    .A1(net36),
    .A2(_02831_));
 sg13g2_nor2b_1 _19978_ (.A(net443),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02833_));
 sg13g2_a21oi_1 _19979_ (.A1(_02692_),
    .A2(net443),
    .Y(_02834_),
    .B1(_02833_));
 sg13g2_nand2_1 _19980_ (.Y(_02835_),
    .A(_12041_),
    .B(_02827_));
 sg13g2_o21ai_1 _19981_ (.B1(_02835_),
    .Y(_00559_),
    .A1(_02827_),
    .A2(_02834_));
 sg13g2_nor2b_1 _19982_ (.A(net443),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02836_));
 sg13g2_a21oi_1 _19983_ (.A1(_02686_),
    .A2(net443),
    .Y(_02837_),
    .B1(_02836_));
 sg13g2_nand2_1 _19984_ (.Y(_02838_),
    .A(_11936_),
    .B(_02826_));
 sg13g2_o21ai_1 _19985_ (.B1(_02838_),
    .Y(_00560_),
    .A1(net36),
    .A2(_02837_));
 sg13g2_nor2b_1 _19986_ (.A(_02829_),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02839_));
 sg13g2_a21oi_1 _19987_ (.A1(net988),
    .A2(_02829_),
    .Y(_02840_),
    .B1(_02839_));
 sg13g2_nand2_1 _19988_ (.Y(_02841_),
    .A(_11945_),
    .B(_02826_));
 sg13g2_o21ai_1 _19989_ (.B1(_02841_),
    .Y(_00561_),
    .A1(net36),
    .A2(_02840_));
 sg13g2_buf_2 _19990_ (.A(_11903_),
    .X(_02842_));
 sg13g2_nor2_1 _19991_ (.A(_02762_),
    .B(_12048_),
    .Y(_02843_));
 sg13g2_buf_2 _19992_ (.A(_02843_),
    .X(_02844_));
 sg13g2_nor2b_1 _19993_ (.A(_02844_),
    .B_N(\cpu.dcache.r_data[7][28] ),
    .Y(_02845_));
 sg13g2_a21oi_1 _19994_ (.A1(_02842_),
    .A2(_02844_),
    .Y(_02846_),
    .B1(_02845_));
 sg13g2_nand2_1 _19995_ (.Y(_02847_),
    .A(_11956_),
    .B(_02826_));
 sg13g2_o21ai_1 _19996_ (.B1(_02847_),
    .Y(_00562_),
    .A1(net36),
    .A2(_02846_));
 sg13g2_buf_2 _19997_ (.A(_11958_),
    .X(_02848_));
 sg13g2_nor2b_1 _19998_ (.A(_02844_),
    .B_N(\cpu.dcache.r_data[7][29] ),
    .Y(_02849_));
 sg13g2_a21oi_1 _19999_ (.A1(_02848_),
    .A2(_02844_),
    .Y(_02850_),
    .B1(_02849_));
 sg13g2_nand2_1 _20000_ (.Y(_02851_),
    .A(_11964_),
    .B(_02826_));
 sg13g2_o21ai_1 _20001_ (.B1(_02851_),
    .Y(_00563_),
    .A1(net36),
    .A2(_02850_));
 sg13g2_nor2b_1 _20002_ (.A(_02767_),
    .B_N(\cpu.dcache.r_data[7][2] ),
    .Y(_02852_));
 sg13g2_a21oi_1 _20003_ (.A1(net1088),
    .A2(_02767_),
    .Y(_02853_),
    .B1(_02852_));
 sg13g2_nand2_1 _20004_ (.Y(_02854_),
    .A(net867),
    .B(_02764_));
 sg13g2_o21ai_1 _20005_ (.B1(_02854_),
    .Y(_00564_),
    .A1(_02765_),
    .A2(_02853_));
 sg13g2_nor2b_1 _20006_ (.A(_02844_),
    .B_N(\cpu.dcache.r_data[7][30] ),
    .Y(_02855_));
 sg13g2_a21oi_1 _20007_ (.A1(_02686_),
    .A2(_02844_),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_nand2_1 _20008_ (.Y(_02857_),
    .A(_11969_),
    .B(_02826_));
 sg13g2_o21ai_1 _20009_ (.B1(_02857_),
    .Y(_00565_),
    .A1(net36),
    .A2(_02856_));
 sg13g2_nor2b_1 _20010_ (.A(_02844_),
    .B_N(\cpu.dcache.r_data[7][31] ),
    .Y(_02858_));
 sg13g2_a21oi_1 _20011_ (.A1(net988),
    .A2(_02844_),
    .Y(_02859_),
    .B1(_02858_));
 sg13g2_nand2_1 _20012_ (.Y(_02860_),
    .A(_11974_),
    .B(_02826_));
 sg13g2_o21ai_1 _20013_ (.B1(_02860_),
    .Y(_00566_),
    .A1(net36),
    .A2(_02859_));
 sg13g2_mux2_1 _20014_ (.A0(\cpu.dcache.r_data[7][3] ),
    .A1(net1096),
    .S(_02767_),
    .X(_02861_));
 sg13g2_nor2_1 _20015_ (.A(_02764_),
    .B(_02861_),
    .Y(_02862_));
 sg13g2_a21oi_1 _20016_ (.A1(_12631_),
    .A2(net39),
    .Y(_00567_),
    .B1(_02862_));
 sg13g2_or2_1 _20017_ (.X(_02863_),
    .B(_12073_),
    .A(_09906_));
 sg13g2_buf_1 _20018_ (.A(_02863_),
    .X(_02864_));
 sg13g2_mux2_1 _20019_ (.A0(net1099),
    .A1(\cpu.dcache.r_data[7][4] ),
    .S(_02864_),
    .X(_02865_));
 sg13g2_mux2_1 _20020_ (.A0(_02865_),
    .A1(net1006),
    .S(net39),
    .X(_00568_));
 sg13g2_mux2_1 _20021_ (.A0(net1095),
    .A1(\cpu.dcache.r_data[7][5] ),
    .S(_02864_),
    .X(_02866_));
 sg13g2_mux2_1 _20022_ (.A0(_02866_),
    .A1(net1005),
    .S(net39),
    .X(_00569_));
 sg13g2_mux2_1 _20023_ (.A0(_12020_),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(_02864_),
    .X(_02867_));
 sg13g2_nor2_1 _20024_ (.A(_02764_),
    .B(_02867_),
    .Y(_02868_));
 sg13g2_a21oi_1 _20025_ (.A1(net753),
    .A2(net39),
    .Y(_00570_),
    .B1(_02868_));
 sg13g2_mux2_1 _20026_ (.A0(net1094),
    .A1(\cpu.dcache.r_data[7][7] ),
    .S(_02864_),
    .X(_02869_));
 sg13g2_nor2_1 _20027_ (.A(_02764_),
    .B(_02869_),
    .Y(_02870_));
 sg13g2_a21oi_1 _20028_ (.A1(net752),
    .A2(net39),
    .Y(_00571_),
    .B1(_02870_));
 sg13g2_nor2b_1 _20029_ (.A(_02775_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_02871_));
 sg13g2_a21oi_1 _20030_ (.A1(_02842_),
    .A2(_02775_),
    .Y(_02872_),
    .B1(_02871_));
 sg13g2_nand2_1 _20031_ (.Y(_02873_),
    .A(_12033_),
    .B(_02772_));
 sg13g2_o21ai_1 _20032_ (.B1(_02873_),
    .Y(_00572_),
    .A1(net38),
    .A2(_02872_));
 sg13g2_nor2b_1 _20033_ (.A(_02775_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_02874_));
 sg13g2_a21oi_1 _20034_ (.A1(_02848_),
    .A2(_02775_),
    .Y(_02875_),
    .B1(_02874_));
 sg13g2_nand2_1 _20035_ (.Y(_02876_),
    .A(_12041_),
    .B(_02772_));
 sg13g2_o21ai_1 _20036_ (.B1(_02876_),
    .Y(_00573_),
    .A1(net38),
    .A2(_02875_));
 sg13g2_buf_1 _20037_ (.A(_08321_),
    .X(_02877_));
 sg13g2_buf_1 _20038_ (.A(\cpu.d_rstrobe_d ),
    .X(_02878_));
 sg13g2_nor2_1 _20039_ (.A(_02877_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_nand3_1 _20040_ (.B(_11890_),
    .C(_02879_),
    .A(_11907_),
    .Y(_02880_));
 sg13g2_o21ai_1 _20041_ (.B1(_02880_),
    .Y(_02881_),
    .A1(_09767_),
    .A2(_11891_));
 sg13g2_buf_2 _20042_ (.A(_02881_),
    .X(_02882_));
 sg13g2_xor2_1 _20043_ (.B(net1098),
    .A(_02878_),
    .X(_02883_));
 sg13g2_nand3_1 _20044_ (.B(_11887_),
    .C(_02883_),
    .A(net1007),
    .Y(_02884_));
 sg13g2_o21ai_1 _20045_ (.B1(_02884_),
    .Y(_02885_),
    .A1(_09767_),
    .A2(_11891_));
 sg13g2_buf_2 _20046_ (.A(_02885_),
    .X(_02886_));
 sg13g2_nor2b_1 _20047_ (.A(net567),
    .B_N(_02886_),
    .Y(_02887_));
 sg13g2_mux2_1 _20048_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_02882_),
    .S(_02887_),
    .X(_00574_));
 sg13g2_buf_1 _20049_ (.A(net627),
    .X(_02888_));
 sg13g2_buf_1 _20050_ (.A(net564),
    .X(_02889_));
 sg13g2_nand2_1 _20051_ (.Y(_02890_),
    .A(net484),
    .B(_02886_));
 sg13g2_mux2_1 _20052_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[1] ),
    .S(_02890_),
    .X(_00575_));
 sg13g2_buf_1 _20053_ (.A(net629),
    .X(_02891_));
 sg13g2_buf_1 _20054_ (.A(net563),
    .X(_02892_));
 sg13g2_nand2_1 _20055_ (.Y(_02893_),
    .A(net483),
    .B(_02886_));
 sg13g2_mux2_1 _20056_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[2] ),
    .S(_02893_),
    .X(_00576_));
 sg13g2_buf_1 _20057_ (.A(net698),
    .X(_02894_));
 sg13g2_buf_1 _20058_ (.A(net616),
    .X(_02895_));
 sg13g2_buf_1 _20059_ (.A(_02895_),
    .X(_02896_));
 sg13g2_nand2_1 _20060_ (.Y(_02897_),
    .A(net482),
    .B(_02886_));
 sg13g2_mux2_1 _20061_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[3] ),
    .S(_02897_),
    .X(_00577_));
 sg13g2_nand2_1 _20062_ (.Y(_02898_),
    .A(net503),
    .B(_02886_));
 sg13g2_mux2_1 _20063_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[4] ),
    .S(_02898_),
    .X(_00578_));
 sg13g2_buf_1 _20064_ (.A(net700),
    .X(_02899_));
 sg13g2_buf_1 _20065_ (.A(_02899_),
    .X(_02900_));
 sg13g2_nand2_1 _20066_ (.Y(_02901_),
    .A(_02900_),
    .B(_02886_));
 sg13g2_mux2_1 _20067_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[5] ),
    .S(_02901_),
    .X(_00579_));
 sg13g2_buf_1 _20068_ (.A(_09336_),
    .X(_02902_));
 sg13g2_buf_1 _20069_ (.A(net560),
    .X(_02903_));
 sg13g2_buf_1 _20070_ (.A(_02903_),
    .X(_02904_));
 sg13g2_nand2_1 _20071_ (.Y(_02905_),
    .A(net442),
    .B(_02886_));
 sg13g2_mux2_1 _20072_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[6] ),
    .S(_02905_),
    .X(_00580_));
 sg13g2_buf_1 _20073_ (.A(net697),
    .X(_02906_));
 sg13g2_buf_1 _20074_ (.A(_02906_),
    .X(_02907_));
 sg13g2_nand2_1 _20075_ (.Y(_02908_),
    .A(_02907_),
    .B(_02886_));
 sg13g2_mux2_1 _20076_ (.A0(_02882_),
    .A1(\cpu.dcache.r_dirty[7] ),
    .S(_02908_),
    .X(_00581_));
 sg13g2_buf_1 _20077_ (.A(net757),
    .X(_02909_));
 sg13g2_buf_2 _20078_ (.A(net676),
    .X(_02910_));
 sg13g2_buf_1 _20079_ (.A(_02910_),
    .X(_02911_));
 sg13g2_buf_1 _20080_ (.A(net400),
    .X(_02912_));
 sg13g2_mux2_1 _20081_ (.A0(net558),
    .A1(\cpu.dcache.r_tag[0][5] ),
    .S(net357),
    .X(_00585_));
 sg13g2_nand2_1 _20082_ (.Y(_02913_),
    .A(_09438_),
    .B(_09447_));
 sg13g2_buf_1 _20083_ (.A(_02913_),
    .X(_02914_));
 sg13g2_mux2_1 _20084_ (.A0(net356),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(_02912_),
    .X(_00586_));
 sg13g2_buf_1 _20085_ (.A(_12029_),
    .X(_02915_));
 sg13g2_mux2_1 _20086_ (.A0(net405),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net398),
    .X(_00587_));
 sg13g2_mux2_1 _20087_ (.A0(_09385_),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(net398),
    .X(_00588_));
 sg13g2_mux2_1 _20088_ (.A0(net448),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net398),
    .X(_00589_));
 sg13g2_mux2_1 _20089_ (.A0(net409),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net398),
    .X(_00590_));
 sg13g2_mux2_1 _20090_ (.A0(net406),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(net398),
    .X(_00591_));
 sg13g2_nand2_1 _20091_ (.Y(_02916_),
    .A(\cpu.dcache.r_tag[0][21] ),
    .B(net398));
 sg13g2_o21ai_1 _20092_ (.B1(_02916_),
    .Y(_00592_),
    .A1(_09618_),
    .A2(net357));
 sg13g2_nand2_1 _20093_ (.Y(_02917_),
    .A(\cpu.dcache.r_tag[0][22] ),
    .B(_12030_));
 sg13g2_o21ai_1 _20094_ (.B1(_02917_),
    .Y(_00593_),
    .A1(_09422_),
    .A2(net357));
 sg13g2_mux2_1 _20095_ (.A0(net404),
    .A1(\cpu.dcache.r_tag[0][23] ),
    .S(net398),
    .X(_00594_));
 sg13g2_inv_1 _20096_ (.Y(_02918_),
    .A(net1058));
 sg13g2_buf_1 _20097_ (.A(_02918_),
    .X(_02919_));
 sg13g2_buf_1 _20098_ (.A(_02919_),
    .X(_02920_));
 sg13g2_nand2_1 _20099_ (.Y(_02921_),
    .A(\cpu.dcache.r_tag[0][6] ),
    .B(net400));
 sg13g2_o21ai_1 _20100_ (.B1(_02921_),
    .Y(_00595_),
    .A1(net675),
    .A2(net357));
 sg13g2_buf_1 _20101_ (.A(_11087_),
    .X(_02922_));
 sg13g2_buf_1 _20102_ (.A(net864),
    .X(_02923_));
 sg13g2_nand2_1 _20103_ (.Y(_02924_),
    .A(\cpu.dcache.r_tag[0][7] ),
    .B(net400));
 sg13g2_o21ai_1 _20104_ (.B1(_02924_),
    .Y(_00596_),
    .A1(_02923_),
    .A2(net357));
 sg13g2_buf_1 _20105_ (.A(_09153_),
    .X(_02925_));
 sg13g2_buf_1 _20106_ (.A(_02925_),
    .X(_02926_));
 sg13g2_nand2_1 _20107_ (.Y(_02927_),
    .A(\cpu.dcache.r_tag[0][8] ),
    .B(net400));
 sg13g2_o21ai_1 _20108_ (.B1(_02927_),
    .Y(_00597_),
    .A1(net749),
    .A2(net357));
 sg13g2_buf_1 _20109_ (.A(_11012_),
    .X(_02928_));
 sg13g2_buf_1 _20110_ (.A(_02928_),
    .X(_02929_));
 sg13g2_nand2_1 _20111_ (.Y(_02930_),
    .A(\cpu.dcache.r_tag[0][9] ),
    .B(net400));
 sg13g2_o21ai_1 _20112_ (.B1(_02930_),
    .Y(_00598_),
    .A1(net748),
    .A2(net357));
 sg13g2_inv_1 _20113_ (.Y(_02931_),
    .A(_10368_));
 sg13g2_buf_1 _20114_ (.A(_02931_),
    .X(_02932_));
 sg13g2_buf_1 _20115_ (.A(_02932_),
    .X(_02933_));
 sg13g2_nand2_1 _20116_ (.Y(_02934_),
    .A(\cpu.dcache.r_tag[0][10] ),
    .B(net400));
 sg13g2_o21ai_1 _20117_ (.B1(_02934_),
    .Y(_00599_),
    .A1(net747),
    .A2(_02912_));
 sg13g2_nand2_1 _20118_ (.Y(_02935_),
    .A(\cpu.dcache.r_tag[0][11] ),
    .B(_12030_));
 sg13g2_o21ai_1 _20119_ (.B1(_02935_),
    .Y(_00600_),
    .A1(_11032_),
    .A2(net357));
 sg13g2_mux2_1 _20120_ (.A0(net407),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net398),
    .X(_00601_));
 sg13g2_mux2_1 _20121_ (.A0(net408),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(_02915_),
    .X(_00602_));
 sg13g2_nand2_1 _20122_ (.Y(_02936_),
    .A(_09500_),
    .B(_09506_));
 sg13g2_buf_1 _20123_ (.A(_02936_),
    .X(_02937_));
 sg13g2_mux2_1 _20124_ (.A0(net355),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(_02915_),
    .X(_00603_));
 sg13g2_buf_1 _20125_ (.A(net613),
    .X(_02938_));
 sg13g2_buf_1 _20126_ (.A(_12176_),
    .X(_02939_));
 sg13g2_mux2_1 _20127_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net557),
    .S(_02939_),
    .X(_00604_));
 sg13g2_mux2_1 _20128_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net356),
    .S(net354),
    .X(_00605_));
 sg13g2_mux2_1 _20129_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net405),
    .S(net354),
    .X(_00606_));
 sg13g2_mux2_1 _20130_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(_09385_),
    .S(_02939_),
    .X(_00607_));
 sg13g2_mux2_1 _20131_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net448),
    .S(net354),
    .X(_00608_));
 sg13g2_mux2_1 _20132_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(_09307_),
    .S(net354),
    .X(_00609_));
 sg13g2_mux2_1 _20133_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net406),
    .S(net354),
    .X(_00610_));
 sg13g2_buf_1 _20134_ (.A(_12175_),
    .X(_02940_));
 sg13g2_nand2_1 _20135_ (.Y(_02941_),
    .A(_09616_),
    .B(net397));
 sg13g2_o21ai_1 _20136_ (.B1(_02941_),
    .Y(_00611_),
    .A1(_09620_),
    .A2(net354));
 sg13g2_nor2b_1 _20137_ (.A(net1065),
    .B_N(_09420_),
    .Y(_02942_));
 sg13g2_buf_1 _20138_ (.A(_02942_),
    .X(_02943_));
 sg13g2_nand2_1 _20139_ (.Y(_02944_),
    .A(_02943_),
    .B(_12176_));
 sg13g2_o21ai_1 _20140_ (.B1(_02944_),
    .Y(_00612_),
    .A1(_09406_),
    .A2(net354));
 sg13g2_mux2_1 _20141_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(net404),
    .S(net354),
    .X(_00613_));
 sg13g2_buf_1 _20142_ (.A(net1058),
    .X(_02945_));
 sg13g2_buf_1 _20143_ (.A(net860),
    .X(_02946_));
 sg13g2_mux2_1 _20144_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net746),
    .S(net397),
    .X(_00614_));
 sg13g2_buf_1 _20145_ (.A(net1057),
    .X(_02947_));
 sg13g2_buf_1 _20146_ (.A(net859),
    .X(_02948_));
 sg13g2_mux2_1 _20147_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net745),
    .S(net397),
    .X(_00615_));
 sg13g2_buf_1 _20148_ (.A(_09152_),
    .X(_02949_));
 sg13g2_buf_1 _20149_ (.A(net986),
    .X(_02950_));
 sg13g2_mux2_1 _20150_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net858),
    .S(net397),
    .X(_00616_));
 sg13g2_buf_1 _20151_ (.A(_10297_),
    .X(_02951_));
 sg13g2_buf_1 _20152_ (.A(net985),
    .X(_02952_));
 sg13g2_mux2_1 _20153_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net857),
    .S(_02940_),
    .X(_00617_));
 sg13g2_buf_1 _20154_ (.A(_10368_),
    .X(_02953_));
 sg13g2_buf_1 _20155_ (.A(_02953_),
    .X(_02954_));
 sg13g2_mux2_1 _20156_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net856),
    .S(net397),
    .X(_00618_));
 sg13g2_buf_2 _20157_ (.A(_10693_),
    .X(_02955_));
 sg13g2_buf_1 _20158_ (.A(_02955_),
    .X(_02956_));
 sg13g2_mux2_1 _20159_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net855),
    .S(net397),
    .X(_00619_));
 sg13g2_mux2_1 _20160_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net407),
    .S(net397),
    .X(_00620_));
 sg13g2_mux2_1 _20161_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net408),
    .S(net397),
    .X(_00621_));
 sg13g2_mux2_1 _20162_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net355),
    .S(_02940_),
    .X(_00622_));
 sg13g2_buf_1 _20163_ (.A(_12300_),
    .X(_02957_));
 sg13g2_mux2_1 _20164_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net557),
    .S(net441),
    .X(_00623_));
 sg13g2_mux2_1 _20165_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net356),
    .S(net441),
    .X(_00624_));
 sg13g2_mux2_1 _20166_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net405),
    .S(net441),
    .X(_00625_));
 sg13g2_mux2_1 _20167_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net449),
    .S(_02957_),
    .X(_00626_));
 sg13g2_mux2_1 _20168_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net448),
    .S(net441),
    .X(_00627_));
 sg13g2_mux2_1 _20169_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net409),
    .S(net441),
    .X(_00628_));
 sg13g2_mux2_1 _20170_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net406),
    .S(net441),
    .X(_00629_));
 sg13g2_mux2_1 _20171_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(_09616_),
    .S(_02957_),
    .X(_00630_));
 sg13g2_buf_1 _20172_ (.A(_12299_),
    .X(_02958_));
 sg13g2_nand2_1 _20173_ (.Y(_02959_),
    .A(_02943_),
    .B(net480));
 sg13g2_o21ai_1 _20174_ (.B1(_02959_),
    .Y(_00631_),
    .A1(_09388_),
    .A2(net441));
 sg13g2_mux2_1 _20175_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(net404),
    .S(net441),
    .X(_00632_));
 sg13g2_mux2_1 _20176_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net746),
    .S(net480),
    .X(_00633_));
 sg13g2_mux2_1 _20177_ (.A0(\cpu.dcache.r_tag[2][7] ),
    .A1(net745),
    .S(net480),
    .X(_00634_));
 sg13g2_mux2_1 _20178_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net858),
    .S(net480),
    .X(_00635_));
 sg13g2_mux2_1 _20179_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net857),
    .S(net480),
    .X(_00636_));
 sg13g2_mux2_1 _20180_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net856),
    .S(net480),
    .X(_00637_));
 sg13g2_mux2_1 _20181_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net855),
    .S(net480),
    .X(_00638_));
 sg13g2_mux2_1 _20182_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net407),
    .S(net480),
    .X(_00639_));
 sg13g2_mux2_1 _20183_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net408),
    .S(_02958_),
    .X(_00640_));
 sg13g2_mux2_1 _20184_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net355),
    .S(_02958_),
    .X(_00641_));
 sg13g2_buf_1 _20185_ (.A(_12421_),
    .X(_02960_));
 sg13g2_mux2_1 _20186_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net557),
    .S(net440),
    .X(_00642_));
 sg13g2_mux2_1 _20187_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(net356),
    .S(net440),
    .X(_00643_));
 sg13g2_mux2_1 _20188_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net405),
    .S(net440),
    .X(_00644_));
 sg13g2_mux2_1 _20189_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net449),
    .S(_02960_),
    .X(_00645_));
 sg13g2_mux2_1 _20190_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net448),
    .S(net440),
    .X(_00646_));
 sg13g2_mux2_1 _20191_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(_09307_),
    .S(net440),
    .X(_00647_));
 sg13g2_mux2_1 _20192_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(net406),
    .S(net440),
    .X(_00648_));
 sg13g2_mux2_1 _20193_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(_09616_),
    .S(_02960_),
    .X(_00649_));
 sg13g2_mux2_1 _20194_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(_02943_),
    .S(net440),
    .X(_00650_));
 sg13g2_mux2_1 _20195_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(net404),
    .S(net440),
    .X(_00651_));
 sg13g2_buf_1 _20196_ (.A(_12421_),
    .X(_02961_));
 sg13g2_mux2_1 _20197_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net746),
    .S(net439),
    .X(_00652_));
 sg13g2_mux2_1 _20198_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net745),
    .S(net439),
    .X(_00653_));
 sg13g2_mux2_1 _20199_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net858),
    .S(net439),
    .X(_00654_));
 sg13g2_mux2_1 _20200_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net857),
    .S(net439),
    .X(_00655_));
 sg13g2_mux2_1 _20201_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net856),
    .S(net439),
    .X(_00656_));
 sg13g2_mux2_1 _20202_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net855),
    .S(_02961_),
    .X(_00657_));
 sg13g2_mux2_1 _20203_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net407),
    .S(net439),
    .X(_00658_));
 sg13g2_mux2_1 _20204_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net408),
    .S(net439),
    .X(_00659_));
 sg13g2_mux2_1 _20205_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net355),
    .S(net439),
    .X(_00660_));
 sg13g2_buf_1 _20206_ (.A(_12536_),
    .X(_02962_));
 sg13g2_buf_1 _20207_ (.A(net438),
    .X(_02963_));
 sg13g2_mux2_1 _20208_ (.A0(net558),
    .A1(\cpu.dcache.r_tag[4][5] ),
    .S(net396),
    .X(_00661_));
 sg13g2_buf_1 _20209_ (.A(net438),
    .X(_02964_));
 sg13g2_mux2_1 _20210_ (.A0(net356),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(_02964_),
    .X(_00662_));
 sg13g2_mux2_1 _20211_ (.A0(net405),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net395),
    .X(_00663_));
 sg13g2_mux2_1 _20212_ (.A0(net449),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(net395),
    .X(_00664_));
 sg13g2_mux2_1 _20213_ (.A0(net448),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net395),
    .X(_00665_));
 sg13g2_mux2_1 _20214_ (.A0(net409),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net395),
    .X(_00666_));
 sg13g2_mux2_1 _20215_ (.A0(net406),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(net395),
    .X(_00667_));
 sg13g2_nand2_1 _20216_ (.Y(_02965_),
    .A(\cpu.dcache.r_tag[4][21] ),
    .B(net438));
 sg13g2_o21ai_1 _20217_ (.B1(_02965_),
    .Y(_00668_),
    .A1(_09618_),
    .A2(net396));
 sg13g2_nand2_1 _20218_ (.Y(_02966_),
    .A(\cpu.dcache.r_tag[4][22] ),
    .B(net438));
 sg13g2_o21ai_1 _20219_ (.B1(_02966_),
    .Y(_00669_),
    .A1(_09422_),
    .A2(net396));
 sg13g2_mux2_1 _20220_ (.A0(net404),
    .A1(\cpu.dcache.r_tag[4][23] ),
    .S(net395),
    .X(_00670_));
 sg13g2_nand2_1 _20221_ (.Y(_02967_),
    .A(\cpu.dcache.r_tag[4][6] ),
    .B(net438));
 sg13g2_o21ai_1 _20222_ (.B1(_02967_),
    .Y(_00671_),
    .A1(net675),
    .A2(_02963_));
 sg13g2_nand2_1 _20223_ (.Y(_02968_),
    .A(\cpu.dcache.r_tag[4][7] ),
    .B(net438));
 sg13g2_o21ai_1 _20224_ (.B1(_02968_),
    .Y(_00672_),
    .A1(_02923_),
    .A2(net396));
 sg13g2_nand2_1 _20225_ (.Y(_02969_),
    .A(\cpu.dcache.r_tag[4][8] ),
    .B(net438));
 sg13g2_o21ai_1 _20226_ (.B1(_02969_),
    .Y(_00673_),
    .A1(net749),
    .A2(net396));
 sg13g2_nand2_1 _20227_ (.Y(_02970_),
    .A(\cpu.dcache.r_tag[4][9] ),
    .B(_02962_));
 sg13g2_o21ai_1 _20228_ (.B1(_02970_),
    .Y(_00674_),
    .A1(net748),
    .A2(net396));
 sg13g2_nand2_1 _20229_ (.Y(_02971_),
    .A(\cpu.dcache.r_tag[4][10] ),
    .B(net438));
 sg13g2_o21ai_1 _20230_ (.B1(_02971_),
    .Y(_00675_),
    .A1(net747),
    .A2(net396));
 sg13g2_nand2_1 _20231_ (.Y(_02972_),
    .A(\cpu.dcache.r_tag[4][11] ),
    .B(_02962_));
 sg13g2_o21ai_1 _20232_ (.B1(_02972_),
    .Y(_00676_),
    .A1(_11032_),
    .A2(_02963_));
 sg13g2_mux2_1 _20233_ (.A0(net407),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net395),
    .X(_00677_));
 sg13g2_mux2_1 _20234_ (.A0(net408),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net395),
    .X(_00678_));
 sg13g2_mux2_1 _20235_ (.A0(net355),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(_02964_),
    .X(_00679_));
 sg13g2_buf_1 _20236_ (.A(_12655_),
    .X(_02973_));
 sg13g2_mux2_1 _20237_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net557),
    .S(net437),
    .X(_00680_));
 sg13g2_mux2_1 _20238_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net356),
    .S(_02973_),
    .X(_00681_));
 sg13g2_mux2_1 _20239_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(net405),
    .S(net437),
    .X(_00682_));
 sg13g2_mux2_1 _20240_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(net449),
    .S(_02973_),
    .X(_00683_));
 sg13g2_mux2_1 _20241_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net448),
    .S(net437),
    .X(_00684_));
 sg13g2_mux2_1 _20242_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net409),
    .S(net437),
    .X(_00685_));
 sg13g2_mux2_1 _20243_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net406),
    .S(net437),
    .X(_00686_));
 sg13g2_mux2_1 _20244_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(_09616_),
    .S(net437),
    .X(_00687_));
 sg13g2_buf_1 _20245_ (.A(_12654_),
    .X(_02974_));
 sg13g2_nand2_1 _20246_ (.Y(_02975_),
    .A(_02943_),
    .B(net479));
 sg13g2_o21ai_1 _20247_ (.B1(_02975_),
    .Y(_00688_),
    .A1(_09393_),
    .A2(net437));
 sg13g2_mux2_1 _20248_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(net404),
    .S(net437),
    .X(_00689_));
 sg13g2_mux2_1 _20249_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(net746),
    .S(net479),
    .X(_00690_));
 sg13g2_mux2_1 _20250_ (.A0(\cpu.dcache.r_tag[5][7] ),
    .A1(net745),
    .S(net479),
    .X(_00691_));
 sg13g2_mux2_1 _20251_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net858),
    .S(net479),
    .X(_00692_));
 sg13g2_mux2_1 _20252_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(net857),
    .S(net479),
    .X(_00693_));
 sg13g2_mux2_1 _20253_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(net856),
    .S(_02974_),
    .X(_00694_));
 sg13g2_mux2_1 _20254_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net855),
    .S(_02974_),
    .X(_00695_));
 sg13g2_mux2_1 _20255_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net407),
    .S(net479),
    .X(_00696_));
 sg13g2_mux2_1 _20256_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net408),
    .S(net479),
    .X(_00697_));
 sg13g2_mux2_1 _20257_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net355),
    .S(net479),
    .X(_00698_));
 sg13g2_buf_1 _20258_ (.A(_02712_),
    .X(_02976_));
 sg13g2_mux2_1 _20259_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net557),
    .S(_02976_),
    .X(_00699_));
 sg13g2_mux2_1 _20260_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net356),
    .S(_02976_),
    .X(_00700_));
 sg13g2_mux2_1 _20261_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(net405),
    .S(net436),
    .X(_00701_));
 sg13g2_mux2_1 _20262_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(net449),
    .S(net436),
    .X(_00702_));
 sg13g2_mux2_1 _20263_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net448),
    .S(net436),
    .X(_00703_));
 sg13g2_mux2_1 _20264_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(net409),
    .S(net436),
    .X(_00704_));
 sg13g2_mux2_1 _20265_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net406),
    .S(net436),
    .X(_00705_));
 sg13g2_mux2_1 _20266_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(_09616_),
    .S(net436),
    .X(_00706_));
 sg13g2_buf_1 _20267_ (.A(_02711_),
    .X(_02977_));
 sg13g2_nand2_1 _20268_ (.Y(_02978_),
    .A(_02943_),
    .B(net478));
 sg13g2_o21ai_1 _20269_ (.B1(_02978_),
    .Y(_00707_),
    .A1(_09398_),
    .A2(net436));
 sg13g2_mux2_1 _20270_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(net404),
    .S(net436),
    .X(_00708_));
 sg13g2_mux2_1 _20271_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net746),
    .S(net478),
    .X(_00709_));
 sg13g2_mux2_1 _20272_ (.A0(\cpu.dcache.r_tag[6][7] ),
    .A1(net745),
    .S(net478),
    .X(_00710_));
 sg13g2_mux2_1 _20273_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net858),
    .S(net478),
    .X(_00711_));
 sg13g2_mux2_1 _20274_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net857),
    .S(_02977_),
    .X(_00712_));
 sg13g2_mux2_1 _20275_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(net856),
    .S(_02977_),
    .X(_00713_));
 sg13g2_mux2_1 _20276_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net855),
    .S(net478),
    .X(_00714_));
 sg13g2_mux2_1 _20277_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net407),
    .S(net478),
    .X(_00715_));
 sg13g2_mux2_1 _20278_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(net408),
    .S(net478),
    .X(_00716_));
 sg13g2_mux2_1 _20279_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net355),
    .S(net478),
    .X(_00717_));
 sg13g2_buf_1 _20280_ (.A(net613),
    .X(_02979_));
 sg13g2_buf_1 _20281_ (.A(net443),
    .X(_02980_));
 sg13g2_mux2_1 _20282_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(_02979_),
    .S(net394),
    .X(_00718_));
 sg13g2_mux2_1 _20283_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(_02914_),
    .S(_02980_),
    .X(_00719_));
 sg13g2_mux2_1 _20284_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net405),
    .S(net394),
    .X(_00720_));
 sg13g2_mux2_1 _20285_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net449),
    .S(_02980_),
    .X(_00721_));
 sg13g2_mux2_1 _20286_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(net448),
    .S(net394),
    .X(_00722_));
 sg13g2_mux2_1 _20287_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net409),
    .S(net394),
    .X(_00723_));
 sg13g2_mux2_1 _20288_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(_09636_),
    .S(net394),
    .X(_00724_));
 sg13g2_mux2_1 _20289_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(_09616_),
    .S(net394),
    .X(_00725_));
 sg13g2_mux2_1 _20290_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(_02943_),
    .S(net394),
    .X(_00726_));
 sg13g2_mux2_1 _20291_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(net404),
    .S(net394),
    .X(_00727_));
 sg13g2_buf_1 _20292_ (.A(net443),
    .X(_02981_));
 sg13g2_mux2_1 _20293_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net746),
    .S(net393),
    .X(_00728_));
 sg13g2_mux2_1 _20294_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net745),
    .S(net393),
    .X(_00729_));
 sg13g2_mux2_1 _20295_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net858),
    .S(net393),
    .X(_00730_));
 sg13g2_mux2_1 _20296_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net857),
    .S(_02981_),
    .X(_00731_));
 sg13g2_mux2_1 _20297_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net856),
    .S(_02981_),
    .X(_00732_));
 sg13g2_mux2_1 _20298_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net855),
    .S(net393),
    .X(_00733_));
 sg13g2_mux2_1 _20299_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net407),
    .S(net393),
    .X(_00734_));
 sg13g2_mux2_1 _20300_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net408),
    .S(net393),
    .X(_00735_));
 sg13g2_mux2_1 _20301_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(_02937_),
    .S(net393),
    .X(_00736_));
 sg13g2_buf_1 _20302_ (.A(net221),
    .X(_02982_));
 sg13g2_nand2_1 _20303_ (.Y(_02983_),
    .A(net220),
    .B(net190));
 sg13g2_buf_1 _20304_ (.A(_02983_),
    .X(_02984_));
 sg13g2_inv_2 _20305_ (.Y(_02985_),
    .A(_08969_));
 sg13g2_nand2_1 _20306_ (.Y(_02986_),
    .A(_08953_),
    .B(_02985_));
 sg13g2_nor2_1 _20307_ (.A(_02985_),
    .B(_08985_),
    .Y(_02987_));
 sg13g2_nand2_1 _20308_ (.Y(_02988_),
    .A(net221),
    .B(_02987_));
 sg13g2_a21o_1 _20309_ (.A2(_02988_),
    .A1(_02986_),
    .B1(_09056_),
    .X(_02989_));
 sg13g2_buf_1 _20310_ (.A(_02989_),
    .X(_02990_));
 sg13g2_o21ai_1 _20311_ (.B1(_02990_),
    .Y(_02991_),
    .A1(net199),
    .A2(_02984_));
 sg13g2_nor2_1 _20312_ (.A(net120),
    .B(_02991_),
    .Y(_02992_));
 sg13g2_a21oi_1 _20313_ (.A1(_10792_),
    .A2(_09836_),
    .Y(_00745_),
    .B1(_02992_));
 sg13g2_buf_1 _20314_ (.A(_08969_),
    .X(_02993_));
 sg13g2_buf_1 _20315_ (.A(net274),
    .X(_02994_));
 sg13g2_buf_1 _20316_ (.A(_08914_),
    .X(_02995_));
 sg13g2_buf_1 _20317_ (.A(net189),
    .X(_02996_));
 sg13g2_a21oi_1 _20318_ (.A1(_08991_),
    .A2(_09033_),
    .Y(_02997_),
    .B1(_09041_));
 sg13g2_buf_1 _20319_ (.A(_02997_),
    .X(_02998_));
 sg13g2_buf_1 _20320_ (.A(_02998_),
    .X(_02999_));
 sg13g2_nor2_1 _20321_ (.A(_02982_),
    .B(net188),
    .Y(_03000_));
 sg13g2_buf_1 _20322_ (.A(_08985_),
    .X(_03001_));
 sg13g2_nand2_1 _20323_ (.Y(_03002_),
    .A(_08932_),
    .B(net273));
 sg13g2_o21ai_1 _20324_ (.B1(_03002_),
    .Y(_03003_),
    .A1(net167),
    .A2(_03000_));
 sg13g2_nand2_1 _20325_ (.Y(_03004_),
    .A(net189),
    .B(_09051_));
 sg13g2_nor2_1 _20326_ (.A(_08969_),
    .B(_08985_),
    .Y(_03005_));
 sg13g2_buf_1 _20327_ (.A(_03005_),
    .X(_03006_));
 sg13g2_buf_1 _20328_ (.A(_09854_),
    .X(_03007_));
 sg13g2_nor2_1 _20329_ (.A(net209),
    .B(_03004_),
    .Y(_03008_));
 sg13g2_a221oi_1 _20330_ (.B2(_03006_),
    .C1(_03008_),
    .B1(_03004_),
    .A1(net227),
    .Y(_03009_),
    .A2(_03003_));
 sg13g2_buf_1 _20331_ (.A(net1133),
    .X(_03010_));
 sg13g2_buf_1 _20332_ (.A(_03010_),
    .X(_03011_));
 sg13g2_nand2_1 _20333_ (.Y(_03012_),
    .A(_03011_),
    .B(net121));
 sg13g2_o21ai_1 _20334_ (.B1(_03012_),
    .Y(_00746_),
    .A1(net107),
    .A2(_03009_));
 sg13g2_nand2_1 _20335_ (.Y(_03013_),
    .A(_08914_),
    .B(_09854_));
 sg13g2_buf_2 _20336_ (.A(_03013_),
    .X(_03014_));
 sg13g2_buf_1 _20337_ (.A(_02986_),
    .X(_03015_));
 sg13g2_nor3_1 _20338_ (.A(net122),
    .B(_03014_),
    .C(net187),
    .Y(_03016_));
 sg13g2_a21o_1 _20339_ (.A2(net108),
    .A1(\cpu.cond[1] ),
    .B1(_03016_),
    .X(_00747_));
 sg13g2_buf_1 _20340_ (.A(_09051_),
    .X(_03017_));
 sg13g2_nor2_1 _20341_ (.A(net208),
    .B(net274),
    .Y(_03018_));
 sg13g2_nor2_1 _20342_ (.A(net167),
    .B(net227),
    .Y(_03019_));
 sg13g2_nor4_1 _20343_ (.A(net123),
    .B(net209),
    .C(_03018_),
    .D(_03019_),
    .Y(_03020_));
 sg13g2_a21o_1 _20344_ (.A2(net108),
    .A1(\cpu.cond[2] ),
    .B1(_03020_),
    .X(_00748_));
 sg13g2_nor4_1 _20345_ (.A(net123),
    .B(net188),
    .C(_09060_),
    .D(_09076_),
    .Y(_03021_));
 sg13g2_a21o_1 _20346_ (.A2(net108),
    .A1(\cpu.dec.div ),
    .B1(_03021_),
    .X(_00749_));
 sg13g2_or2_1 _20347_ (.X(_03022_),
    .B(net195),
    .A(_03014_));
 sg13g2_buf_1 _20348_ (.A(_03022_),
    .X(_03023_));
 sg13g2_inv_1 _20349_ (.Y(_03024_),
    .A(_00158_));
 sg13g2_a22oi_1 _20350_ (.Y(_03025_),
    .B1(net639),
    .B2(\cpu.icache.r_data[2][9] ),
    .A2(net641),
    .A1(\cpu.icache.r_data[1][9] ));
 sg13g2_mux4_1 _20351_ (.S0(net1067),
    .A0(\cpu.icache.r_data[4][9] ),
    .A1(\cpu.icache.r_data[5][9] ),
    .A2(\cpu.icache.r_data[6][9] ),
    .A3(\cpu.icache.r_data[7][9] ),
    .S1(_08462_),
    .X(_03026_));
 sg13g2_a22oi_1 _20352_ (.Y(_03027_),
    .B1(_03026_),
    .B2(net929),
    .A2(net640),
    .A1(\cpu.icache.r_data[3][9] ));
 sg13g2_nand3_1 _20353_ (.B(_03025_),
    .C(_03027_),
    .A(net576),
    .Y(_03028_));
 sg13g2_o21ai_1 _20354_ (.B1(_03028_),
    .Y(_03029_),
    .A1(_03024_),
    .A2(net576));
 sg13g2_nand2_1 _20355_ (.Y(_03030_),
    .A(\cpu.icache.r_data[1][25] ),
    .B(net641));
 sg13g2_a22oi_1 _20356_ (.Y(_03031_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][25] ),
    .A2(_08485_),
    .A1(\cpu.icache.r_data[2][25] ));
 sg13g2_a22oi_1 _20357_ (.Y(_03032_),
    .B1(_08558_),
    .B2(\cpu.icache.r_data[6][25] ),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[3][25] ));
 sg13g2_a22oi_1 _20358_ (.Y(_03033_),
    .B1(_08562_),
    .B2(\cpu.icache.r_data[5][25] ),
    .A2(_08553_),
    .A1(\cpu.icache.r_data[7][25] ));
 sg13g2_nand4_1 _20359_ (.B(_03031_),
    .C(_03032_),
    .A(_03030_),
    .Y(_03034_),
    .D(_03033_));
 sg13g2_nor2_1 _20360_ (.A(_00159_),
    .B(net576),
    .Y(_03035_));
 sg13g2_o21ai_1 _20361_ (.B1(_08857_),
    .Y(_03036_),
    .A1(_03034_),
    .A2(_03035_));
 sg13g2_o21ai_1 _20362_ (.B1(_03036_),
    .Y(_03037_),
    .A1(_08857_),
    .A2(_03029_));
 sg13g2_buf_2 _20363_ (.A(_03037_),
    .X(_03038_));
 sg13g2_inv_1 _20364_ (.Y(_03039_),
    .A(_00148_));
 sg13g2_mux4_1 _20365_ (.S0(net1067),
    .A0(\cpu.icache.r_data[4][7] ),
    .A1(\cpu.icache.r_data[5][7] ),
    .A2(\cpu.icache.r_data[6][7] ),
    .A3(\cpu.icache.r_data[7][7] ),
    .S1(net927),
    .X(_03040_));
 sg13g2_nand2_1 _20366_ (.Y(_03041_),
    .A(net929),
    .B(_03040_));
 sg13g2_nand2_1 _20367_ (.Y(_03042_),
    .A(\cpu.icache.r_data[1][7] ),
    .B(_08470_));
 sg13g2_a22oi_1 _20368_ (.Y(_03043_),
    .B1(_08485_),
    .B2(\cpu.icache.r_data[2][7] ),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[3][7] ));
 sg13g2_nand4_1 _20369_ (.B(_03041_),
    .C(_03042_),
    .A(net643),
    .Y(_03044_),
    .D(_03043_));
 sg13g2_o21ai_1 _20370_ (.B1(_03044_),
    .Y(_03045_),
    .A1(_03039_),
    .A2(net576));
 sg13g2_mux4_1 _20371_ (.S0(net1067),
    .A0(\cpu.icache.r_data[4][23] ),
    .A1(\cpu.icache.r_data[5][23] ),
    .A2(\cpu.icache.r_data[6][23] ),
    .A3(\cpu.icache.r_data[7][23] ),
    .S1(net923),
    .X(_03046_));
 sg13g2_and2_1 _20372_ (.A(net929),
    .B(_03046_),
    .X(_03047_));
 sg13g2_and2_1 _20373_ (.A(\cpu.icache.r_data[3][23] ),
    .B(_08479_),
    .X(_03048_));
 sg13g2_a221oi_1 _20374_ (.B2(\cpu.icache.r_data[2][23] ),
    .C1(_03048_),
    .B1(_08485_),
    .A1(\cpu.icache.r_data[1][23] ),
    .Y(_03049_),
    .A2(_08470_));
 sg13g2_o21ai_1 _20375_ (.B1(_03049_),
    .Y(_03050_),
    .A1(_00149_),
    .A2(_08452_));
 sg13g2_o21ai_1 _20376_ (.B1(_08857_),
    .Y(_03051_),
    .A1(_03047_),
    .A2(_03050_));
 sg13g2_o21ai_1 _20377_ (.B1(_03051_),
    .Y(_03052_),
    .A1(_08857_),
    .A2(_03045_));
 sg13g2_buf_1 _20378_ (.A(_03052_),
    .X(_03053_));
 sg13g2_or2_1 _20379_ (.X(_03054_),
    .B(net353),
    .A(_03038_));
 sg13g2_buf_1 _20380_ (.A(_03054_),
    .X(_03055_));
 sg13g2_a22oi_1 _20381_ (.Y(_03056_),
    .B1(net636),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(net578),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_a22oi_1 _20382_ (.Y(_03057_),
    .B1(net508),
    .B2(\cpu.icache.r_data[3][8] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(net923),
    .X(_03058_));
 sg13g2_a22oi_1 _20384_ (.Y(_03059_),
    .B1(_03058_),
    .B2(_08607_),
    .A2(net805),
    .A1(\cpu.icache.r_data[7][8] ));
 sg13g2_or2_1 _20385_ (.X(_03060_),
    .B(_03059_),
    .A(net925));
 sg13g2_and4_1 _20386_ (.A(net509),
    .B(_03056_),
    .C(_03057_),
    .D(_03060_),
    .X(_03061_));
 sg13g2_a21oi_1 _20387_ (.A1(_00156_),
    .A2(net635),
    .Y(_03062_),
    .B1(_03061_));
 sg13g2_mux4_1 _20388_ (.S0(net816),
    .A0(\cpu.icache.r_data[4][24] ),
    .A1(\cpu.icache.r_data[5][24] ),
    .A2(\cpu.icache.r_data[6][24] ),
    .A3(\cpu.icache.r_data[7][24] ),
    .S1(net723),
    .X(_03063_));
 sg13g2_and2_1 _20389_ (.A(\cpu.icache.r_data[3][24] ),
    .B(_08480_),
    .X(_03064_));
 sg13g2_a221oi_1 _20390_ (.B2(\cpu.icache.r_data[2][24] ),
    .C1(_03064_),
    .B1(_08550_),
    .A1(\cpu.icache.r_data[1][24] ),
    .Y(_03065_),
    .A2(net581));
 sg13g2_o21ai_1 _20391_ (.B1(_03065_),
    .Y(_03066_),
    .A1(_00157_),
    .A2(net509));
 sg13g2_a21oi_1 _20392_ (.A1(net817),
    .A2(_03063_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_nand2_1 _20393_ (.Y(_03068_),
    .A(_08858_),
    .B(_03067_));
 sg13g2_o21ai_1 _20394_ (.B1(_03068_),
    .Y(_03069_),
    .A1(_08897_),
    .A2(_03062_));
 sg13g2_buf_1 _20395_ (.A(_03069_),
    .X(_03070_));
 sg13g2_buf_1 _20396_ (.A(_03070_),
    .X(_03071_));
 sg13g2_nor2b_1 _20397_ (.A(_03055_),
    .B_N(net207),
    .Y(_03072_));
 sg13g2_nand4_1 _20398_ (.B(_09027_),
    .C(_09043_),
    .A(_09011_),
    .Y(_03073_),
    .D(_03072_));
 sg13g2_buf_1 _20399_ (.A(_03073_),
    .X(_03074_));
 sg13g2_and2_1 _20400_ (.A(net927),
    .B(\cpu.icache.r_data[6][4] ),
    .X(_03075_));
 sg13g2_a21oi_1 _20401_ (.A1(_08441_),
    .A2(\cpu.icache.r_data[4][4] ),
    .Y(_03076_),
    .B1(_03075_));
 sg13g2_a22oi_1 _20402_ (.Y(_03077_),
    .B1(net926),
    .B2(\cpu.icache.r_data[7][4] ),
    .A2(_08658_),
    .A1(\cpu.icache.r_data[5][4] ));
 sg13g2_o21ai_1 _20403_ (.B1(_03077_),
    .Y(_03078_),
    .A1(net928),
    .A2(_03076_));
 sg13g2_nand2_1 _20404_ (.Y(_03079_),
    .A(net929),
    .B(_03078_));
 sg13g2_nand2_1 _20405_ (.Y(_03080_),
    .A(\cpu.icache.r_data[1][4] ),
    .B(net581));
 sg13g2_a22oi_1 _20406_ (.Y(_03081_),
    .B1(net578),
    .B2(\cpu.icache.r_data[2][4] ),
    .A2(net580),
    .A1(\cpu.icache.r_data[3][4] ));
 sg13g2_and4_1 _20407_ (.A(net582),
    .B(_03079_),
    .C(_03080_),
    .D(_03081_),
    .X(_03082_));
 sg13g2_a21oi_1 _20408_ (.A1(_00154_),
    .A2(net635),
    .Y(_03083_),
    .B1(_03082_));
 sg13g2_nor2_1 _20409_ (.A(_00155_),
    .B(net582),
    .Y(_03084_));
 sg13g2_mux2_1 _20410_ (.A0(\cpu.icache.r_data[5][20] ),
    .A1(\cpu.icache.r_data[7][20] ),
    .S(net815),
    .X(_03085_));
 sg13g2_a22oi_1 _20411_ (.Y(_03086_),
    .B1(_03085_),
    .B2(net816),
    .A2(net812),
    .A1(\cpu.icache.r_data[6][20] ));
 sg13g2_nor2_1 _20412_ (.A(net813),
    .B(_03086_),
    .Y(_03087_));
 sg13g2_a22oi_1 _20413_ (.Y(_03088_),
    .B1(net578),
    .B2(\cpu.icache.r_data[2][20] ),
    .A2(net581),
    .A1(\cpu.icache.r_data[1][20] ));
 sg13g2_a22oi_1 _20414_ (.Y(_03089_),
    .B1(net814),
    .B2(\cpu.icache.r_data[4][20] ),
    .A2(net580),
    .A1(\cpu.icache.r_data[3][20] ));
 sg13g2_nand2_1 _20415_ (.Y(_03090_),
    .A(_03088_),
    .B(_03089_));
 sg13g2_or4_1 _20416_ (.A(_08868_),
    .B(_03084_),
    .C(_03087_),
    .D(_03090_),
    .X(_03091_));
 sg13g2_o21ai_1 _20417_ (.B1(_03091_),
    .Y(_03092_),
    .A1(net1062),
    .A2(_03083_));
 sg13g2_buf_1 _20418_ (.A(_03092_),
    .X(_03093_));
 sg13g2_inv_2 _20419_ (.Y(_03094_),
    .A(_03093_));
 sg13g2_nor4_1 _20420_ (.A(_09076_),
    .B(_03023_),
    .C(_03074_),
    .D(_03094_),
    .Y(_03095_));
 sg13g2_buf_1 _20421_ (.A(net123),
    .X(_03096_));
 sg13g2_mux2_1 _20422_ (.A0(_03095_),
    .A1(\cpu.dec.do_flush_all ),
    .S(net95),
    .X(_00750_));
 sg13g2_buf_1 _20423_ (.A(_08953_),
    .X(_03097_));
 sg13g2_buf_1 _20424_ (.A(_02987_),
    .X(_03098_));
 sg13g2_nand2_1 _20425_ (.Y(_03099_),
    .A(net206),
    .B(net205));
 sg13g2_nor3_1 _20426_ (.A(net122),
    .B(_03014_),
    .C(_03099_),
    .Y(_03100_));
 sg13g2_a21o_1 _20427_ (.A2(_03096_),
    .A1(\cpu.dec.do_flush_write ),
    .B1(_03100_),
    .X(_00751_));
 sg13g2_nor2_1 _20428_ (.A(_08914_),
    .B(_09854_),
    .Y(_03101_));
 sg13g2_buf_2 _20429_ (.A(_03101_),
    .X(_03102_));
 sg13g2_nor2_1 _20430_ (.A(_03014_),
    .B(net195),
    .Y(_03103_));
 sg13g2_inv_1 _20431_ (.Y(_03104_),
    .A(_00150_));
 sg13g2_a22oi_1 _20432_ (.Y(_03105_),
    .B1(net636),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(net579),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_a22oi_1 _20433_ (.Y(_03106_),
    .B1(net508),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(net516),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_mux2_1 _20434_ (.A0(\cpu.icache.r_data[4][2] ),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(net815),
    .X(_03107_));
 sg13g2_a22oi_1 _20435_ (.Y(_03108_),
    .B1(_03107_),
    .B2(net717),
    .A2(net805),
    .A1(\cpu.icache.r_data[7][2] ));
 sg13g2_or2_1 _20436_ (.X(_03109_),
    .B(_03108_),
    .A(net813));
 sg13g2_nand4_1 _20437_ (.B(_03105_),
    .C(_03106_),
    .A(net513),
    .Y(_03110_),
    .D(_03109_));
 sg13g2_o21ai_1 _20438_ (.B1(_03110_),
    .Y(_03111_),
    .A1(_03104_),
    .A2(net517));
 sg13g2_nor2_1 _20439_ (.A(_00151_),
    .B(net513),
    .Y(_03112_));
 sg13g2_mux2_1 _20440_ (.A0(\cpu.icache.r_data[4][18] ),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(net815),
    .X(_03113_));
 sg13g2_a22oi_1 _20441_ (.Y(_03114_),
    .B1(_03113_),
    .B2(_08608_),
    .A2(net805),
    .A1(\cpu.icache.r_data[7][18] ));
 sg13g2_nor2_1 _20442_ (.A(net721),
    .B(_03114_),
    .Y(_03115_));
 sg13g2_a22oi_1 _20443_ (.Y(_03116_),
    .B1(net512),
    .B2(\cpu.icache.r_data[2][18] ),
    .A2(net511),
    .A1(\cpu.icache.r_data[1][18] ));
 sg13g2_a22oi_1 _20444_ (.Y(_03117_),
    .B1(net577),
    .B2(\cpu.icache.r_data[5][18] ),
    .A2(net508),
    .A1(\cpu.icache.r_data[3][18] ));
 sg13g2_nand2_1 _20445_ (.Y(_03118_),
    .A(_03116_),
    .B(_03117_));
 sg13g2_nor4_1 _20446_ (.A(net921),
    .B(_03112_),
    .C(_03115_),
    .D(_03118_),
    .Y(_03119_));
 sg13g2_a21oi_1 _20447_ (.A1(net921),
    .A2(_03111_),
    .Y(_03120_),
    .B1(_03119_));
 sg13g2_buf_2 _20448_ (.A(_03120_),
    .X(_03121_));
 sg13g2_nand2_1 _20449_ (.Y(_03122_),
    .A(net220),
    .B(net274));
 sg13g2_nor2_1 _20450_ (.A(net208),
    .B(_02985_),
    .Y(_03123_));
 sg13g2_buf_1 _20451_ (.A(net273),
    .X(_03124_));
 sg13g2_o21ai_1 _20452_ (.B1(net225),
    .Y(_03125_),
    .A1(_03008_),
    .A2(_03123_));
 sg13g2_a21oi_1 _20453_ (.A1(_03122_),
    .A2(_03125_),
    .Y(_03126_),
    .B1(net287));
 sg13g2_a21oi_1 _20454_ (.A1(_03103_),
    .A2(_03121_),
    .Y(_03127_),
    .B1(_03126_));
 sg13g2_buf_1 _20455_ (.A(net220),
    .X(_03128_));
 sg13g2_buf_1 _20456_ (.A(_03093_),
    .X(_03129_));
 sg13g2_nand2b_1 _20457_ (.Y(_03130_),
    .B(net190),
    .A_N(_08878_));
 sg13g2_o21ai_1 _20458_ (.B1(_03130_),
    .Y(_03131_),
    .A1(net190),
    .A2(net204));
 sg13g2_nand3_1 _20459_ (.B(net226),
    .C(_03131_),
    .A(net186),
    .Y(_03132_));
 sg13g2_o21ai_1 _20460_ (.B1(_03132_),
    .Y(_03133_),
    .A1(_03102_),
    .A2(_03127_));
 sg13g2_mux2_1 _20461_ (.A0(_03133_),
    .A1(_10550_),
    .S(net95),
    .X(_00752_));
 sg13g2_inv_1 _20462_ (.Y(_03134_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_and2_1 _20463_ (.A(_09051_),
    .B(_03001_),
    .X(_03135_));
 sg13g2_a21oi_1 _20464_ (.A1(_03129_),
    .A2(_03135_),
    .Y(_03136_),
    .B1(_08935_));
 sg13g2_buf_2 _20465_ (.A(_03136_),
    .X(_03137_));
 sg13g2_nand2b_1 _20466_ (.Y(_03138_),
    .B(net274),
    .A_N(net273));
 sg13g2_nor2_1 _20467_ (.A(_09043_),
    .B(_03015_),
    .Y(_03139_));
 sg13g2_buf_2 _20468_ (.A(_03139_),
    .X(_03140_));
 sg13g2_nor2_1 _20469_ (.A(_03135_),
    .B(_03140_),
    .Y(_03141_));
 sg13g2_o21ai_1 _20470_ (.B1(_03141_),
    .Y(_03142_),
    .A1(_03138_),
    .A2(net207));
 sg13g2_nand2_1 _20471_ (.Y(_03143_),
    .A(_09051_),
    .B(net226));
 sg13g2_buf_1 _20472_ (.A(_03143_),
    .X(_03144_));
 sg13g2_and2_1 _20473_ (.A(_09058_),
    .B(net195),
    .X(_03145_));
 sg13g2_buf_1 _20474_ (.A(_03145_),
    .X(_03146_));
 sg13g2_nand2_1 _20475_ (.Y(_03147_),
    .A(_03140_),
    .B(net117));
 sg13g2_o21ai_1 _20476_ (.B1(_03147_),
    .Y(_03148_),
    .A1(net204),
    .A2(net185));
 sg13g2_nand2_1 _20477_ (.Y(_03149_),
    .A(_09058_),
    .B(net195));
 sg13g2_nand2_1 _20478_ (.Y(_03150_),
    .A(_08935_),
    .B(_03149_));
 sg13g2_a22oi_1 _20479_ (.Y(_03151_),
    .B1(_03148_),
    .B2(_03150_),
    .A2(_03142_),
    .A1(_03137_));
 sg13g2_nor2_1 _20480_ (.A(_02995_),
    .B(net204),
    .Y(_03152_));
 sg13g2_nand2_1 _20481_ (.Y(_03153_),
    .A(_09051_),
    .B(_02987_));
 sg13g2_buf_1 _20482_ (.A(_03153_),
    .X(_03154_));
 sg13g2_nand2_1 _20483_ (.Y(_03155_),
    .A(_08933_),
    .B(_09054_));
 sg13g2_o21ai_1 _20484_ (.B1(_03155_),
    .Y(_03156_),
    .A1(net190),
    .A2(_03154_));
 sg13g2_a21oi_1 _20485_ (.A1(_03152_),
    .A2(_03156_),
    .Y(_03157_),
    .B1(_08853_));
 sg13g2_buf_2 _20486_ (.A(_03157_),
    .X(_03158_));
 sg13g2_a22oi_1 _20487_ (.Y(_00753_),
    .B1(_03151_),
    .B2(_03158_),
    .A2(net105),
    .A1(_03134_));
 sg13g2_inv_1 _20488_ (.Y(_03159_),
    .A(\cpu.dec.imm[11] ));
 sg13g2_nor2_1 _20489_ (.A(net287),
    .B(net185),
    .Y(_03160_));
 sg13g2_o21ai_1 _20490_ (.B1(net117),
    .Y(_03161_),
    .A1(_03140_),
    .A2(_03160_));
 sg13g2_nor2_2 _20491_ (.A(_08953_),
    .B(_08969_),
    .Y(_03162_));
 sg13g2_inv_1 _20492_ (.Y(_03163_),
    .A(_03162_));
 sg13g2_a21oi_1 _20493_ (.A1(_02999_),
    .A2(_03163_),
    .Y(_03164_),
    .B1(net225));
 sg13g2_a21oi_1 _20494_ (.A1(_09052_),
    .A2(net188),
    .Y(_03165_),
    .B1(_03017_));
 sg13g2_nor2_1 _20495_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sg13g2_or3_1 _20496_ (.A(_09026_),
    .B(_03070_),
    .C(_03055_),
    .X(_03167_));
 sg13g2_buf_2 _20497_ (.A(_03167_),
    .X(_03168_));
 sg13g2_nor3_1 _20498_ (.A(_09026_),
    .B(_03071_),
    .C(_03055_),
    .Y(_03169_));
 sg13g2_buf_1 _20499_ (.A(_03169_),
    .X(_03170_));
 sg13g2_a21o_1 _20500_ (.A2(_03170_),
    .A1(net204),
    .B1(_03143_),
    .X(_03171_));
 sg13g2_buf_1 _20501_ (.A(_03171_),
    .X(_03172_));
 sg13g2_a21oi_1 _20502_ (.A1(net287),
    .A2(_03168_),
    .Y(_03173_),
    .B1(_03172_));
 sg13g2_o21ai_1 _20503_ (.B1(_03137_),
    .Y(_03174_),
    .A1(_03166_),
    .A2(_03173_));
 sg13g2_and2_1 _20504_ (.A(_03161_),
    .B(_03174_),
    .X(_03175_));
 sg13g2_a22oi_1 _20505_ (.Y(_00754_),
    .B1(_03158_),
    .B2(_03175_),
    .A2(net105),
    .A1(_03159_));
 sg13g2_inv_1 _20506_ (.Y(_03176_),
    .A(\cpu.dec.imm[12] ));
 sg13g2_nor2_1 _20507_ (.A(_08894_),
    .B(net185),
    .Y(_03177_));
 sg13g2_o21ai_1 _20508_ (.B1(net117),
    .Y(_03178_),
    .A1(_03140_),
    .A2(_03177_));
 sg13g2_a21oi_1 _20509_ (.A1(_08894_),
    .A2(_03168_),
    .Y(_03179_),
    .B1(_03172_));
 sg13g2_o21ai_1 _20510_ (.B1(_03137_),
    .Y(_03180_),
    .A1(_03166_),
    .A2(_03179_));
 sg13g2_and2_1 _20511_ (.A(_03178_),
    .B(_03180_),
    .X(_03181_));
 sg13g2_a22oi_1 _20512_ (.Y(_00755_),
    .B1(_03158_),
    .B2(_03181_),
    .A2(_09836_),
    .A1(_03176_));
 sg13g2_a21oi_1 _20513_ (.A1(net187),
    .A2(net185),
    .Y(_03182_),
    .B1(_09044_));
 sg13g2_a21oi_1 _20514_ (.A1(net198),
    .A2(_03168_),
    .Y(_03183_),
    .B1(_03172_));
 sg13g2_or2_1 _20515_ (.X(_03184_),
    .B(_03183_),
    .A(_03166_));
 sg13g2_a22oi_1 _20516_ (.Y(_03185_),
    .B1(_03184_),
    .B2(_03137_),
    .A2(_03182_),
    .A1(net117));
 sg13g2_a22oi_1 _20517_ (.Y(_00756_),
    .B1(_03158_),
    .B2(_03185_),
    .A2(net105),
    .A1(_10421_));
 sg13g2_inv_1 _20518_ (.Y(_03186_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_nor2_1 _20519_ (.A(_09063_),
    .B(_03144_),
    .Y(_03187_));
 sg13g2_o21ai_1 _20520_ (.B1(net117),
    .Y(_03188_),
    .A1(_03140_),
    .A2(_03187_));
 sg13g2_a21oi_1 _20521_ (.A1(_09063_),
    .A2(_03168_),
    .Y(_03189_),
    .B1(_03172_));
 sg13g2_o21ai_1 _20522_ (.B1(_03137_),
    .Y(_03190_),
    .A1(_03166_),
    .A2(_03189_));
 sg13g2_and2_1 _20523_ (.A(_03158_),
    .B(_03190_),
    .X(_03191_));
 sg13g2_a22oi_1 _20524_ (.Y(_00757_),
    .B1(_03188_),
    .B2(_03191_),
    .A2(net105),
    .A1(_03186_));
 sg13g2_inv_1 _20525_ (.Y(_03192_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_inv_1 _20526_ (.Y(_03193_),
    .A(net196));
 sg13g2_nor2_1 _20527_ (.A(_03193_),
    .B(net185),
    .Y(_03194_));
 sg13g2_o21ai_1 _20528_ (.B1(_03146_),
    .Y(_03195_),
    .A1(_03140_),
    .A2(_03194_));
 sg13g2_a22oi_1 _20529_ (.Y(_00758_),
    .B1(_03191_),
    .B2(_03195_),
    .A2(net107),
    .A1(_03192_));
 sg13g2_nor2_1 _20530_ (.A(_08969_),
    .B(_03168_),
    .Y(_03196_));
 sg13g2_o21ai_1 _20531_ (.B1(net221),
    .Y(_03197_),
    .A1(net273),
    .A2(_03196_));
 sg13g2_inv_1 _20532_ (.Y(_03198_),
    .A(_03197_));
 sg13g2_nand2_1 _20533_ (.Y(_03199_),
    .A(_02985_),
    .B(net273));
 sg13g2_nand2_1 _20534_ (.Y(_03200_),
    .A(_09854_),
    .B(_02987_));
 sg13g2_nand2_1 _20535_ (.Y(_03201_),
    .A(_03199_),
    .B(_03200_));
 sg13g2_buf_1 _20536_ (.A(net208),
    .X(_03202_));
 sg13g2_o21ai_1 _20537_ (.B1(net184),
    .Y(_03203_),
    .A1(_03198_),
    .A2(_03201_));
 sg13g2_nand3_1 _20538_ (.B(net199),
    .C(_03203_),
    .A(net167),
    .Y(_03204_));
 sg13g2_nand2_1 _20539_ (.Y(_03205_),
    .A(_02990_),
    .B(_03023_));
 sg13g2_inv_1 _20540_ (.Y(_03206_),
    .A(_00152_));
 sg13g2_a22oi_1 _20541_ (.Y(_03207_),
    .B1(net722),
    .B2(\cpu.icache.r_data[4][3] ),
    .A2(net511),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_a22oi_1 _20542_ (.Y(_03208_),
    .B1(net577),
    .B2(\cpu.icache.r_data[5][3] ),
    .A2(net637),
    .A1(\cpu.icache.r_data[6][3] ));
 sg13g2_mux2_1 _20543_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(net813),
    .X(_03209_));
 sg13g2_a22oi_1 _20544_ (.Y(_03210_),
    .B1(_03209_),
    .B2(net716),
    .A2(net512),
    .A1(\cpu.icache.r_data[2][3] ));
 sg13g2_nand4_1 _20545_ (.B(_03207_),
    .C(_03208_),
    .A(net456),
    .Y(_03211_),
    .D(_03210_));
 sg13g2_o21ai_1 _20546_ (.B1(_03211_),
    .Y(_03212_),
    .A1(_03206_),
    .A2(net456));
 sg13g2_nor2_1 _20547_ (.A(_00153_),
    .B(net517),
    .Y(_03213_));
 sg13g2_mux2_1 _20548_ (.A0(\cpu.icache.r_data[4][19] ),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(net723),
    .X(_03214_));
 sg13g2_a22oi_1 _20549_ (.Y(_03215_),
    .B1(_03214_),
    .B2(_08608_),
    .A2(net716),
    .A1(\cpu.icache.r_data[7][19] ));
 sg13g2_nor2_1 _20550_ (.A(net721),
    .B(_03215_),
    .Y(_03216_));
 sg13g2_a22oi_1 _20551_ (.Y(_03217_),
    .B1(net577),
    .B2(\cpu.icache.r_data[5][19] ),
    .A2(net457),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_a22oi_1 _20552_ (.Y(_03218_),
    .B1(net514),
    .B2(\cpu.icache.r_data[2][19] ),
    .A2(net515),
    .A1(\cpu.icache.r_data[3][19] ));
 sg13g2_nand2_1 _20553_ (.Y(_03219_),
    .A(_03217_),
    .B(_03218_));
 sg13g2_nor4_1 _20554_ (.A(net921),
    .B(_03213_),
    .C(_03216_),
    .D(_03219_),
    .Y(_03220_));
 sg13g2_a21oi_2 _20555_ (.B1(_03220_),
    .Y(_03221_),
    .A2(_03212_),
    .A1(net921));
 sg13g2_buf_1 _20556_ (.A(_03221_),
    .X(_03222_));
 sg13g2_and2_1 _20557_ (.A(_02984_),
    .B(net203),
    .X(_03223_));
 sg13g2_a22oi_1 _20558_ (.Y(_03224_),
    .B1(_03205_),
    .B2(_03223_),
    .A2(_03204_),
    .A1(_08893_));
 sg13g2_nand2_1 _20559_ (.Y(_03225_),
    .A(_10597_),
    .B(net120));
 sg13g2_o21ai_1 _20560_ (.B1(_03225_),
    .Y(_00759_),
    .A1(net107),
    .A2(_03224_));
 sg13g2_inv_1 _20561_ (.Y(_03226_),
    .A(_03002_));
 sg13g2_a21oi_1 _20562_ (.A1(net189),
    .A2(_03201_),
    .Y(_03227_),
    .B1(_03226_));
 sg13g2_o21ai_1 _20563_ (.B1(_02984_),
    .Y(_03228_),
    .A1(net206),
    .A2(_03227_));
 sg13g2_nand2_1 _20564_ (.Y(_03229_),
    .A(net219),
    .B(_03228_));
 sg13g2_and2_1 _20565_ (.A(net197),
    .B(net203),
    .X(_03230_));
 sg13g2_inv_1 _20566_ (.Y(_03231_),
    .A(_08935_));
 sg13g2_nand2_1 _20567_ (.Y(_03232_),
    .A(_09051_),
    .B(net273));
 sg13g2_nand2_1 _20568_ (.Y(_03233_),
    .A(_03231_),
    .B(_03232_));
 sg13g2_nor4_1 _20569_ (.A(net287),
    .B(net185),
    .C(_03168_),
    .D(_03233_),
    .Y(_03234_));
 sg13g2_nand2_1 _20570_ (.Y(_03235_),
    .A(_03149_),
    .B(_03233_));
 sg13g2_o21ai_1 _20571_ (.B1(_03235_),
    .Y(_03236_),
    .A1(_03230_),
    .A2(_03234_));
 sg13g2_nand2_1 _20572_ (.Y(_03237_),
    .A(net274),
    .B(net203));
 sg13g2_o21ai_1 _20573_ (.B1(_03237_),
    .Y(_03238_),
    .A1(_08878_),
    .A2(net274));
 sg13g2_nand2_1 _20574_ (.Y(_03239_),
    .A(_03154_),
    .B(_03238_));
 sg13g2_o21ai_1 _20575_ (.B1(_03239_),
    .Y(_03240_),
    .A1(_09027_),
    .A2(_03154_));
 sg13g2_nor2_1 _20576_ (.A(net189),
    .B(net221),
    .Y(_03241_));
 sg13g2_buf_1 _20577_ (.A(_03241_),
    .X(_03242_));
 sg13g2_a22oi_1 _20578_ (.Y(_03243_),
    .B1(_03240_),
    .B2(net140),
    .A2(_03205_),
    .A1(_03094_));
 sg13g2_nand3_1 _20579_ (.B(_03236_),
    .C(_03243_),
    .A(_03229_),
    .Y(_03244_));
 sg13g2_mux2_1 _20580_ (.A0(_03244_),
    .A1(_10542_),
    .S(net95),
    .X(_00760_));
 sg13g2_nand2_1 _20581_ (.Y(_03245_),
    .A(_02985_),
    .B(_03170_));
 sg13g2_o21ai_1 _20582_ (.B1(_03200_),
    .Y(_03246_),
    .A1(_03007_),
    .A2(_03245_));
 sg13g2_a22oi_1 _20583_ (.Y(_03247_),
    .B1(_03232_),
    .B2(_02996_),
    .A2(net227),
    .A1(_03007_));
 sg13g2_a21oi_1 _20584_ (.A1(_03202_),
    .A2(_03246_),
    .Y(_03248_),
    .B1(_03247_));
 sg13g2_nand2b_1 _20585_ (.Y(_03249_),
    .B(net208),
    .A_N(net273));
 sg13g2_nor3_1 _20586_ (.A(net189),
    .B(net190),
    .C(net204),
    .Y(_03250_));
 sg13g2_mux2_1 _20587_ (.A0(net273),
    .A1(_03232_),
    .S(_09854_),
    .X(_03251_));
 sg13g2_nor3_1 _20588_ (.A(_08878_),
    .B(net220),
    .C(_03251_),
    .Y(_03252_));
 sg13g2_a21o_1 _20589_ (.A2(_03250_),
    .A1(_03249_),
    .B1(_03252_),
    .X(_03253_));
 sg13g2_nand2_1 _20590_ (.Y(_03254_),
    .A(net197),
    .B(_03094_));
 sg13g2_o21ai_1 _20591_ (.B1(_03254_),
    .Y(_03255_),
    .A1(_09027_),
    .A2(net187));
 sg13g2_a22oi_1 _20592_ (.Y(_03256_),
    .B1(_03255_),
    .B2(_03235_),
    .A2(_03253_),
    .A1(net227));
 sg13g2_o21ai_1 _20593_ (.B1(_03256_),
    .Y(_03257_),
    .A1(net196),
    .A2(_03248_));
 sg13g2_buf_1 _20594_ (.A(_08853_),
    .X(_03258_));
 sg13g2_mux2_1 _20595_ (.A0(_03257_),
    .A1(_10488_),
    .S(_03258_),
    .X(_00761_));
 sg13g2_or3_1 _20596_ (.A(net198),
    .B(_03168_),
    .C(_03249_),
    .X(_03259_));
 sg13g2_o21ai_1 _20597_ (.B1(_03259_),
    .Y(_03260_),
    .A1(net184),
    .A2(net196));
 sg13g2_a22oi_1 _20598_ (.Y(_03261_),
    .B1(_03260_),
    .B2(_02985_),
    .A2(net205),
    .A1(_03193_));
 sg13g2_nor2_1 _20599_ (.A(net209),
    .B(_03097_),
    .Y(_03262_));
 sg13g2_o21ai_1 _20600_ (.B1(net225),
    .Y(_03263_),
    .A1(_03123_),
    .A2(_03262_));
 sg13g2_nand2_1 _20601_ (.Y(_03264_),
    .A(net167),
    .B(_03263_));
 sg13g2_nor2_1 _20602_ (.A(net196),
    .B(net187),
    .Y(_03265_));
 sg13g2_a22oi_1 _20603_ (.Y(_03266_),
    .B1(_03265_),
    .B2(net117),
    .A2(_03264_),
    .A1(net188));
 sg13g2_o21ai_1 _20604_ (.B1(_03266_),
    .Y(_03267_),
    .A1(_03233_),
    .A2(_03261_));
 sg13g2_mux2_1 _20605_ (.A0(_03267_),
    .A1(\cpu.dec.imm[4] ),
    .S(net116),
    .X(_00762_));
 sg13g2_o21ai_1 _20606_ (.B1(net199),
    .Y(_03268_),
    .A1(net287),
    .A2(net226));
 sg13g2_o21ai_1 _20607_ (.B1(_03268_),
    .Y(_03269_),
    .A1(net199),
    .A2(_03121_));
 sg13g2_o21ai_1 _20608_ (.B1(net209),
    .Y(_03270_),
    .A1(_03017_),
    .A2(net205));
 sg13g2_o21ai_1 _20609_ (.B1(_03270_),
    .Y(_03271_),
    .A1(net185),
    .A2(_03170_));
 sg13g2_inv_2 _20610_ (.Y(_03272_),
    .A(_03121_));
 sg13g2_a21oi_1 _20611_ (.A1(net167),
    .A2(_03271_),
    .Y(_03273_),
    .B1(_03272_));
 sg13g2_nor2_1 _20612_ (.A(_03102_),
    .B(_03273_),
    .Y(_03274_));
 sg13g2_a21oi_1 _20613_ (.A1(_03102_),
    .A2(_03269_),
    .Y(_03275_),
    .B1(_03274_));
 sg13g2_mux2_1 _20614_ (.A0(_03275_),
    .A1(\cpu.dec.imm[5] ),
    .S(net116),
    .X(_00763_));
 sg13g2_and4_1 _20615_ (.A(_03231_),
    .B(net205),
    .C(net353),
    .D(_03232_),
    .X(_03276_));
 sg13g2_nor3_1 _20616_ (.A(net287),
    .B(net186),
    .C(_03015_),
    .Y(_03277_));
 sg13g2_o21ai_1 _20617_ (.B1(_03197_),
    .Y(_03278_),
    .A1(net225),
    .A2(_09856_));
 sg13g2_a22oi_1 _20618_ (.Y(_03279_),
    .B1(_03278_),
    .B2(net184),
    .A2(net140),
    .A1(_02985_));
 sg13g2_nor2b_1 _20619_ (.A(_03279_),
    .B_N(net203),
    .Y(_03280_));
 sg13g2_nor4_1 _20620_ (.A(_03102_),
    .B(_03276_),
    .C(_03277_),
    .D(_03280_),
    .Y(_03281_));
 sg13g2_nand2_1 _20621_ (.Y(_03282_),
    .A(_02993_),
    .B(_08988_));
 sg13g2_inv_1 _20622_ (.Y(_03283_),
    .A(_03282_));
 sg13g2_a221oi_1 _20623_ (.B2(net353),
    .C1(_02984_),
    .B1(_03283_),
    .A1(net197),
    .Y(_03284_),
    .A2(net203));
 sg13g2_nor3_1 _20624_ (.A(net122),
    .B(_03281_),
    .C(_03284_),
    .Y(_03285_));
 sg13g2_a21o_1 _20625_ (.A2(net95),
    .A1(\cpu.dec.imm[6] ),
    .B1(_03285_),
    .X(_00764_));
 sg13g2_inv_1 _20626_ (.Y(_03286_),
    .A(_03199_));
 sg13g2_nand2_1 _20627_ (.Y(_03287_),
    .A(net140),
    .B(net205));
 sg13g2_o21ai_1 _20628_ (.B1(_03287_),
    .Y(_03288_),
    .A1(net186),
    .A2(_03197_));
 sg13g2_a22oi_1 _20629_ (.Y(_03289_),
    .B1(_03288_),
    .B2(net184),
    .A2(_03286_),
    .A1(_03242_));
 sg13g2_inv_1 _20630_ (.Y(_03290_),
    .A(_02990_));
 sg13g2_o21ai_1 _20631_ (.B1(_03254_),
    .Y(_03291_),
    .A1(net207),
    .A2(_03282_));
 sg13g2_a22oi_1 _20632_ (.Y(_03292_),
    .B1(_03102_),
    .B2(_03291_),
    .A2(_03290_),
    .A1(_08893_));
 sg13g2_o21ai_1 _20633_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net204),
    .A2(_03289_));
 sg13g2_mux2_1 _20634_ (.A0(_03293_),
    .A1(\cpu.dec.imm[7] ),
    .S(net116),
    .X(_00765_));
 sg13g2_inv_1 _20635_ (.Y(_03294_),
    .A(\cpu.dec.imm[8] ));
 sg13g2_a21oi_1 _20636_ (.A1(_03129_),
    .A2(_03170_),
    .Y(_03295_),
    .B1(_03144_));
 sg13g2_o21ai_1 _20637_ (.B1(_03295_),
    .Y(_03296_),
    .A1(_03121_),
    .A2(_03170_));
 sg13g2_nand2_1 _20638_ (.Y(_03297_),
    .A(net205),
    .B(_03038_));
 sg13g2_nand3_1 _20639_ (.B(_03296_),
    .C(_03297_),
    .A(_03141_),
    .Y(_03298_));
 sg13g2_nand2_1 _20640_ (.Y(_03299_),
    .A(_03102_),
    .B(_03038_));
 sg13g2_nor2_1 _20641_ (.A(_03272_),
    .B(net185),
    .Y(_03300_));
 sg13g2_o21ai_1 _20642_ (.B1(net117),
    .Y(_03301_),
    .A1(_03140_),
    .A2(_03300_));
 sg13g2_o21ai_1 _20643_ (.B1(_03301_),
    .Y(_03302_),
    .A1(_03282_),
    .A2(_03299_));
 sg13g2_a21oi_1 _20644_ (.A1(_03137_),
    .A2(_03298_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_a22oi_1 _20645_ (.Y(_00766_),
    .B1(_03158_),
    .B2(_03303_),
    .A2(net107),
    .A1(_03294_));
 sg13g2_inv_1 _20646_ (.Y(_03304_),
    .A(\cpu.dec.imm[9] ));
 sg13g2_o21ai_1 _20647_ (.B1(_03295_),
    .Y(_03305_),
    .A1(_03170_),
    .A2(_03222_));
 sg13g2_nand2_1 _20648_ (.Y(_03306_),
    .A(net219),
    .B(_03098_));
 sg13g2_nand3_1 _20649_ (.B(_03305_),
    .C(_03306_),
    .A(_03141_),
    .Y(_03307_));
 sg13g2_nand3_1 _20650_ (.B(net226),
    .C(_03222_),
    .A(net184),
    .Y(_03308_));
 sg13g2_o21ai_1 _20651_ (.B1(_03308_),
    .Y(_03309_),
    .A1(_09044_),
    .A2(net187));
 sg13g2_a22oi_1 _20652_ (.Y(_03310_),
    .B1(_03309_),
    .B2(net117),
    .A2(_03307_),
    .A1(_03137_));
 sg13g2_a22oi_1 _20653_ (.Y(_00767_),
    .B1(_03158_),
    .B2(_03310_),
    .A2(net107),
    .A1(_03304_));
 sg13g2_nor4_1 _20654_ (.A(net819),
    .B(_08894_),
    .C(_03023_),
    .D(_03074_),
    .Y(_03311_));
 sg13g2_buf_1 _20655_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03312_));
 sg13g2_mux2_1 _20656_ (.A0(_03311_),
    .A1(_03312_),
    .S(net116),
    .X(_00768_));
 sg13g2_nor4_1 _20657_ (.A(net206),
    .B(_08987_),
    .C(_03014_),
    .D(net226),
    .Y(_03313_));
 sg13g2_mux2_1 _20658_ (.A0(_03313_),
    .A1(\cpu.dec.io ),
    .S(net116),
    .X(_00769_));
 sg13g2_or4_1 _20659_ (.A(_08896_),
    .B(_03094_),
    .C(_03121_),
    .D(_03221_),
    .X(_03314_));
 sg13g2_buf_2 _20660_ (.A(_03314_),
    .X(_03315_));
 sg13g2_nor3_1 _20661_ (.A(net199),
    .B(_09856_),
    .C(_03315_),
    .Y(_03316_));
 sg13g2_mux2_1 _20662_ (.A0(_03316_),
    .A1(\cpu.dec.jmp ),
    .S(net116),
    .X(_00770_));
 sg13g2_nand2_1 _20663_ (.Y(_03317_),
    .A(net209),
    .B(_03124_));
 sg13g2_a21oi_1 _20664_ (.A1(net167),
    .A2(_03317_),
    .Y(_03318_),
    .B1(_03163_));
 sg13g2_mux2_1 _20665_ (.A0(_03318_),
    .A1(_11385_),
    .S(net116),
    .X(_00771_));
 sg13g2_nor4_1 _20666_ (.A(net123),
    .B(_08896_),
    .C(net188),
    .D(_09060_),
    .Y(_03319_));
 sg13g2_a21o_1 _20667_ (.A2(net95),
    .A1(\cpu.dec.mult ),
    .B1(_03319_),
    .X(_00772_));
 sg13g2_a21oi_1 _20668_ (.A1(net196),
    .A2(net198),
    .Y(_03320_),
    .B1(_09838_));
 sg13g2_nor3_1 _20669_ (.A(net167),
    .B(net206),
    .C(net188),
    .Y(_03321_));
 sg13g2_nor3_1 _20670_ (.A(net186),
    .B(_03202_),
    .C(_09028_),
    .Y(_03322_));
 sg13g2_nor4_1 _20671_ (.A(_02982_),
    .B(_09052_),
    .C(_03321_),
    .D(_03322_),
    .Y(_03323_));
 sg13g2_a21oi_1 _20672_ (.A1(_08990_),
    .A2(_03320_),
    .Y(_03324_),
    .B1(_03323_));
 sg13g2_nand2_1 _20673_ (.Y(_03325_),
    .A(net890),
    .B(net120));
 sg13g2_o21ai_1 _20674_ (.B1(_03325_),
    .Y(_00773_),
    .A1(net107),
    .A2(_03324_));
 sg13g2_a21o_1 _20675_ (.A2(_03315_),
    .A1(_08987_),
    .B1(net208),
    .X(_03326_));
 sg13g2_and2_1 _20676_ (.A(net186),
    .B(net353),
    .X(_03327_));
 sg13g2_nor2_1 _20677_ (.A(_03001_),
    .B(net353),
    .Y(_03328_));
 sg13g2_a21oi_1 _20678_ (.A1(net225),
    .A2(_03272_),
    .Y(_03329_),
    .B1(_03328_));
 sg13g2_and2_1 _20679_ (.A(_03124_),
    .B(_03053_),
    .X(_03330_));
 sg13g2_a22oi_1 _20680_ (.Y(_03331_),
    .B1(_03330_),
    .B2(_03123_),
    .A2(_03329_),
    .A1(_03162_));
 sg13g2_o21ai_1 _20681_ (.B1(net353),
    .Y(_03332_),
    .A1(net208),
    .A2(_08987_));
 sg13g2_a21o_1 _20682_ (.A2(_03332_),
    .A1(_03154_),
    .B1(_08935_),
    .X(_03333_));
 sg13g2_o21ai_1 _20683_ (.B1(_03333_),
    .Y(_03334_),
    .A1(_03014_),
    .A2(_03331_));
 sg13g2_a221oi_1 _20684_ (.B2(_03327_),
    .C1(_03334_),
    .B1(_03326_),
    .A1(net188),
    .Y(_03335_),
    .A2(_03316_));
 sg13g2_a21oi_1 _20685_ (.A1(net184),
    .A2(_03272_),
    .Y(_03336_),
    .B1(net205));
 sg13g2_a21oi_1 _20686_ (.A1(net187),
    .A2(_03336_),
    .Y(_03337_),
    .B1(_02984_));
 sg13g2_a21oi_1 _20687_ (.A1(_02984_),
    .A2(_03335_),
    .Y(_03338_),
    .B1(_03337_));
 sg13g2_mux2_1 _20688_ (.A0(_03338_),
    .A1(\cpu.dec.r_rd[0] ),
    .S(_03258_),
    .X(_00774_));
 sg13g2_o21ai_1 _20689_ (.B1(net208),
    .Y(_03339_),
    .A1(_03226_),
    .A2(net226));
 sg13g2_nand2_1 _20690_ (.Y(_03340_),
    .A(net199),
    .B(_03339_));
 sg13g2_a22oi_1 _20691_ (.Y(_03341_),
    .B1(_03340_),
    .B2(_02995_),
    .A2(_03326_),
    .A1(net140));
 sg13g2_nand2_1 _20692_ (.Y(_03342_),
    .A(_03138_),
    .B(_03102_));
 sg13g2_nand2_1 _20693_ (.Y(_03343_),
    .A(_09058_),
    .B(_03286_));
 sg13g2_a21oi_1 _20694_ (.A1(_03342_),
    .A2(_03343_),
    .Y(_03344_),
    .B1(net206));
 sg13g2_or4_1 _20695_ (.A(_08896_),
    .B(_03023_),
    .C(_03074_),
    .D(net204),
    .X(_03345_));
 sg13g2_nand2_1 _20696_ (.Y(_03346_),
    .A(_03272_),
    .B(_03221_));
 sg13g2_nor2_1 _20697_ (.A(_03345_),
    .B(_03346_),
    .Y(_03347_));
 sg13g2_a21oi_1 _20698_ (.A1(net203),
    .A2(_03344_),
    .Y(_03348_),
    .B1(_03347_));
 sg13g2_o21ai_1 _20699_ (.B1(_03348_),
    .Y(_03349_),
    .A1(net207),
    .A2(_03341_));
 sg13g2_mux2_1 _20700_ (.A0(_03349_),
    .A1(\cpu.dec.r_rd[1] ),
    .S(net116),
    .X(_00775_));
 sg13g2_nand2_1 _20701_ (.Y(_03350_),
    .A(_03094_),
    .B(_03344_));
 sg13g2_nand2b_1 _20702_ (.Y(_03351_),
    .B(_03038_),
    .A_N(_03341_));
 sg13g2_a21oi_1 _20703_ (.A1(_03350_),
    .A2(_03351_),
    .Y(_03352_),
    .B1(net120));
 sg13g2_a21o_1 _20704_ (.A2(net95),
    .A1(\cpu.dec.r_rd[2] ),
    .B1(_03352_),
    .X(_00776_));
 sg13g2_o21ai_1 _20705_ (.B1(net225),
    .Y(_03353_),
    .A1(_03097_),
    .A2(_03014_));
 sg13g2_o21ai_1 _20706_ (.B1(_09854_),
    .Y(_03354_),
    .A1(_02993_),
    .A2(_09026_));
 sg13g2_o21ai_1 _20707_ (.B1(net274),
    .Y(_03355_),
    .A1(net189),
    .A2(net219));
 sg13g2_a22oi_1 _20708_ (.Y(_03356_),
    .B1(_03355_),
    .B2(net206),
    .A2(_03354_),
    .A1(_09056_));
 sg13g2_o21ai_1 _20709_ (.B1(_03356_),
    .Y(_03357_),
    .A1(net225),
    .A2(net219));
 sg13g2_a21o_1 _20710_ (.A2(_03353_),
    .A1(net227),
    .B1(_03357_),
    .X(_03358_));
 sg13g2_nor2_1 _20711_ (.A(net167),
    .B(_03315_),
    .Y(_03359_));
 sg13g2_a21o_1 _20712_ (.A2(_03358_),
    .A1(_03342_),
    .B1(net206),
    .X(_03360_));
 sg13g2_o21ai_1 _20713_ (.B1(_03360_),
    .Y(_03361_),
    .A1(_03358_),
    .A2(_03359_));
 sg13g2_mux2_1 _20714_ (.A0(_03361_),
    .A1(\cpu.dec.r_rd[3] ),
    .S(net121),
    .X(_00777_));
 sg13g2_o21ai_1 _20715_ (.B1(net190),
    .Y(_03362_),
    .A1(_03098_),
    .A2(_03162_));
 sg13g2_a21oi_1 _20716_ (.A1(_03143_),
    .A2(_03362_),
    .Y(_03363_),
    .B1(net220));
 sg13g2_a21oi_1 _20717_ (.A1(net189),
    .A2(net195),
    .Y(_03364_),
    .B1(net190));
 sg13g2_a21oi_1 _20718_ (.A1(_09043_),
    .A2(_03315_),
    .Y(_03365_),
    .B1(_08988_));
 sg13g2_o21ai_1 _20719_ (.B1(net140),
    .Y(_03366_),
    .A1(_03283_),
    .A2(_03365_));
 sg13g2_o21ai_1 _20720_ (.B1(_03366_),
    .Y(_03367_),
    .A1(_03363_),
    .A2(_03364_));
 sg13g2_nand2_1 _20721_ (.Y(_03368_),
    .A(net227),
    .B(_03102_));
 sg13g2_nand3_1 _20722_ (.B(_03367_),
    .C(_03368_),
    .A(net353),
    .Y(_03369_));
 sg13g2_o21ai_1 _20723_ (.B1(_03369_),
    .Y(_03370_),
    .A1(net199),
    .A2(_02984_));
 sg13g2_mux2_1 _20724_ (.A0(_03370_),
    .A1(_10886_),
    .S(net121),
    .X(_00778_));
 sg13g2_nand2_1 _20725_ (.Y(_03371_),
    .A(net189),
    .B(net226));
 sg13g2_o21ai_1 _20726_ (.B1(_03122_),
    .Y(_03372_),
    .A1(_03168_),
    .A2(_03371_));
 sg13g2_o21ai_1 _20727_ (.B1(_03138_),
    .Y(_03373_),
    .A1(_02994_),
    .A2(_03071_));
 sg13g2_a22oi_1 _20728_ (.Y(_03374_),
    .B1(_03373_),
    .B2(net186),
    .A2(_03372_),
    .A1(net184));
 sg13g2_a21oi_1 _20729_ (.A1(net227),
    .A2(net207),
    .Y(_03375_),
    .B1(_09856_));
 sg13g2_nand3_1 _20730_ (.B(net198),
    .C(_03315_),
    .A(net197),
    .Y(_03376_));
 sg13g2_nand2_1 _20731_ (.Y(_03377_),
    .A(net221),
    .B(net274));
 sg13g2_nor2b_1 _20732_ (.A(_03162_),
    .B_N(_03377_),
    .Y(_03378_));
 sg13g2_a21oi_1 _20733_ (.A1(net221),
    .A2(_03162_),
    .Y(_03379_),
    .B1(net220));
 sg13g2_o21ai_1 _20734_ (.B1(_03379_),
    .Y(_03380_),
    .A1(net225),
    .A2(_03378_));
 sg13g2_a21oi_1 _20735_ (.A1(_03023_),
    .A2(net207),
    .Y(_03381_),
    .B1(_03380_));
 sg13g2_a21oi_1 _20736_ (.A1(_03375_),
    .A2(_03376_),
    .Y(_03382_),
    .B1(_03381_));
 sg13g2_o21ai_1 _20737_ (.B1(_03382_),
    .Y(_03383_),
    .A1(net209),
    .A2(_03374_));
 sg13g2_mux2_1 _20738_ (.A0(_03383_),
    .A1(net880),
    .S(net121),
    .X(_00779_));
 sg13g2_nand2_1 _20739_ (.Y(_03384_),
    .A(_03366_),
    .B(_03380_));
 sg13g2_o21ai_1 _20740_ (.B1(_03384_),
    .Y(_03385_),
    .A1(_03103_),
    .A2(_03038_));
 sg13g2_o21ai_1 _20741_ (.B1(_03385_),
    .Y(_03386_),
    .A1(net227),
    .A2(_03299_));
 sg13g2_nor2_1 _20742_ (.A(net120),
    .B(_03386_),
    .Y(_03387_));
 sg13g2_a21oi_1 _20743_ (.A1(net763),
    .A2(net105),
    .Y(_00780_),
    .B1(_03387_));
 sg13g2_nand2_1 _20744_ (.Y(_03388_),
    .A(_09064_),
    .B(_03365_));
 sg13g2_nand3_1 _20745_ (.B(_03282_),
    .C(_03388_),
    .A(net186),
    .Y(_03389_));
 sg13g2_o21ai_1 _20746_ (.B1(_03389_),
    .Y(_03390_),
    .A1(_09052_),
    .A2(_03004_));
 sg13g2_o21ai_1 _20747_ (.B1(_03377_),
    .Y(_03391_),
    .A1(net190),
    .A2(_03249_));
 sg13g2_nand3_1 _20748_ (.B(net184),
    .C(_03317_),
    .A(_02996_),
    .Y(_03392_));
 sg13g2_o21ai_1 _20749_ (.B1(_02988_),
    .Y(_03393_),
    .A1(_02994_),
    .A2(_03392_));
 sg13g2_a221oi_1 _20750_ (.B2(net186),
    .C1(_03393_),
    .B1(_03391_),
    .A1(net209),
    .Y(_03394_),
    .A2(_03390_));
 sg13g2_mux2_1 _20751_ (.A0(_03394_),
    .A1(_10892_),
    .S(net121),
    .X(_00781_));
 sg13g2_a22oi_1 _20752_ (.Y(_03395_),
    .B1(_03121_),
    .B2(net197),
    .A2(net353),
    .A1(_03018_));
 sg13g2_nand3_1 _20753_ (.B(_09028_),
    .C(_02998_),
    .A(_08893_),
    .Y(_03396_));
 sg13g2_nand2_1 _20754_ (.Y(_03397_),
    .A(_09053_),
    .B(_03396_));
 sg13g2_nand3_1 _20755_ (.B(_03154_),
    .C(_03397_),
    .A(_09058_),
    .Y(_03398_));
 sg13g2_inv_1 _20756_ (.Y(_03399_),
    .A(_03398_));
 sg13g2_a21oi_1 _20757_ (.A1(net140),
    .A2(_03018_),
    .Y(_03400_),
    .B1(_03399_));
 sg13g2_nand2_1 _20758_ (.Y(_03401_),
    .A(_03121_),
    .B(_03400_));
 sg13g2_o21ai_1 _20759_ (.B1(_03401_),
    .Y(_03402_),
    .A1(_09856_),
    .A2(_03395_));
 sg13g2_mux2_1 _20760_ (.A0(_03402_),
    .A1(_10224_),
    .S(net121),
    .X(_00782_));
 sg13g2_nor2_1 _20761_ (.A(net187),
    .B(net207),
    .Y(_03403_));
 sg13g2_or2_1 _20762_ (.X(_03404_),
    .B(_03403_),
    .A(_03230_));
 sg13g2_a221oi_1 _20763_ (.B2(net140),
    .C1(_09837_),
    .B1(_03404_),
    .A1(net203),
    .Y(_03405_),
    .A2(_03400_));
 sg13g2_a21oi_1 _20764_ (.A1(net1035),
    .A2(net105),
    .Y(_00783_),
    .B1(_03405_));
 sg13g2_a22oi_1 _20765_ (.Y(_03406_),
    .B1(_03094_),
    .B2(net197),
    .A2(_03038_),
    .A1(_03018_));
 sg13g2_nand2_1 _20766_ (.Y(_03407_),
    .A(_03094_),
    .B(_03400_));
 sg13g2_o21ai_1 _20767_ (.B1(_03407_),
    .Y(_03408_),
    .A1(_09856_),
    .A2(_03406_));
 sg13g2_mux2_1 _20768_ (.A0(_03408_),
    .A1(_10213_),
    .S(net121),
    .X(_00784_));
 sg13g2_and2_1 _20769_ (.A(_08878_),
    .B(_09053_),
    .X(_03409_));
 sg13g2_nor2_1 _20770_ (.A(net219),
    .B(net187),
    .Y(_03410_));
 sg13g2_o21ai_1 _20771_ (.B1(net140),
    .Y(_03411_),
    .A1(_03409_),
    .A2(_03410_));
 sg13g2_nand2_1 _20772_ (.Y(_03412_),
    .A(_03398_),
    .B(_03411_));
 sg13g2_nand2_1 _20773_ (.Y(_03413_),
    .A(_10179_),
    .B(net120));
 sg13g2_o21ai_1 _20774_ (.B1(_03413_),
    .Y(_00785_),
    .A1(net107),
    .A2(_03412_));
 sg13g2_nor4_1 _20775_ (.A(net123),
    .B(net198),
    .C(_09060_),
    .D(_09076_),
    .Y(_03414_));
 sg13g2_a21o_1 _20776_ (.A2(net95),
    .A1(net887),
    .B1(_03414_),
    .X(_00786_));
 sg13g2_a22oi_1 _20777_ (.Y(_03415_),
    .B1(_03019_),
    .B2(net206),
    .A2(net205),
    .A1(_09058_));
 sg13g2_buf_1 _20778_ (.A(\cpu.dec.r_store ),
    .X(_03416_));
 sg13g2_nand2_1 _20779_ (.Y(_03417_),
    .A(_03416_),
    .B(net120));
 sg13g2_o21ai_1 _20780_ (.B1(_03417_),
    .Y(_00787_),
    .A1(net107),
    .A2(_03415_));
 sg13g2_mux2_1 _20781_ (.A0(_03347_),
    .A1(\cpu.dec.r_swapsp ),
    .S(_09067_),
    .X(_00788_));
 sg13g2_nor4_1 _20782_ (.A(net123),
    .B(_03272_),
    .C(net203),
    .D(_03345_),
    .Y(_03418_));
 sg13g2_a21o_1 _20783_ (.A2(net95),
    .A1(\cpu.dec.r_sys_call ),
    .B1(_03418_),
    .X(_00789_));
 sg13g2_nor2_1 _20784_ (.A(_08896_),
    .B(_09043_),
    .Y(_03419_));
 sg13g2_a21oi_1 _20785_ (.A1(_09043_),
    .A2(_03272_),
    .Y(_03420_),
    .B1(_03419_));
 sg13g2_a22oi_1 _20786_ (.Y(_03421_),
    .B1(_03420_),
    .B2(_09011_),
    .A2(_02999_),
    .A1(_09028_));
 sg13g2_o21ai_1 _20787_ (.B1(_03231_),
    .Y(_03422_),
    .A1(_08989_),
    .A2(_03421_));
 sg13g2_nor4_1 _20788_ (.A(_08286_),
    .B(_02998_),
    .C(_09832_),
    .D(_03315_),
    .Y(_03423_));
 sg13g2_buf_1 _20789_ (.A(_08364_),
    .X(_03424_));
 sg13g2_or2_1 _20790_ (.X(_03425_),
    .B(_10458_),
    .A(net982));
 sg13g2_o21ai_1 _20791_ (.B1(_09052_),
    .Y(_03426_),
    .A1(net226),
    .A2(_03425_));
 sg13g2_a221oi_1 _20792_ (.B2(net208),
    .C1(_08933_),
    .B1(_03426_),
    .A1(_08987_),
    .Y(_03427_),
    .A2(_09011_));
 sg13g2_o21ai_1 _20793_ (.B1(_03427_),
    .Y(_03428_),
    .A1(_03099_),
    .A2(_03423_));
 sg13g2_nor2b_1 _20794_ (.A(net207),
    .B_N(_03053_),
    .Y(_03429_));
 sg13g2_xnor2_1 _20795_ (.Y(_03430_),
    .A(_03038_),
    .B(_03429_));
 sg13g2_nor4_1 _20796_ (.A(net982),
    .B(_09064_),
    .C(_03143_),
    .D(_03430_),
    .Y(_03431_));
 sg13g2_a21o_1 _20797_ (.A2(_03428_),
    .A1(_03422_),
    .B1(_03431_),
    .X(_03432_));
 sg13g2_nor2_1 _20798_ (.A(_03093_),
    .B(_03346_),
    .Y(_03433_));
 sg13g2_mux2_1 _20799_ (.A0(net204),
    .A1(_03433_),
    .S(_08878_),
    .X(_03434_));
 sg13g2_nor2_1 _20800_ (.A(_08893_),
    .B(_03434_),
    .Y(_03435_));
 sg13g2_nor4_1 _20801_ (.A(_08428_),
    .B(net195),
    .C(_03074_),
    .D(_03435_),
    .Y(_03436_));
 sg13g2_o21ai_1 _20802_ (.B1(net209),
    .Y(_03437_),
    .A1(_03128_),
    .A2(_03436_));
 sg13g2_nor2_1 _20803_ (.A(net982),
    .B(_03430_),
    .Y(_03438_));
 sg13g2_o21ai_1 _20804_ (.B1(_09027_),
    .Y(_03439_),
    .A1(_02985_),
    .A2(_03365_));
 sg13g2_nand2_1 _20805_ (.Y(_03440_),
    .A(_03154_),
    .B(_03439_));
 sg13g2_nand2_1 _20806_ (.Y(_03441_),
    .A(_03438_),
    .B(_03440_));
 sg13g2_nand2_1 _20807_ (.Y(_03442_),
    .A(_03121_),
    .B(_03221_));
 sg13g2_xnor2_1 _20808_ (.Y(_03443_),
    .A(_03094_),
    .B(_03442_));
 sg13g2_nor2_1 _20809_ (.A(_08286_),
    .B(_02998_),
    .Y(_03444_));
 sg13g2_a21oi_1 _20810_ (.A1(net982),
    .A2(net188),
    .Y(_03445_),
    .B1(_03444_));
 sg13g2_nand3_1 _20811_ (.B(_03443_),
    .C(_03445_),
    .A(_03409_),
    .Y(_03446_));
 sg13g2_nand2b_1 _20812_ (.Y(_03447_),
    .B(_03420_),
    .A_N(net195));
 sg13g2_nand4_1 _20813_ (.B(_03441_),
    .C(_03446_),
    .A(_03099_),
    .Y(_03448_),
    .D(_03447_));
 sg13g2_a22oi_1 _20814_ (.Y(_03449_),
    .B1(_03448_),
    .B2(_03128_),
    .A2(_03437_),
    .A1(_03432_));
 sg13g2_nand2_1 _20815_ (.Y(_03450_),
    .A(net287),
    .B(_03072_));
 sg13g2_nor3_1 _20816_ (.A(_09832_),
    .B(_09852_),
    .C(_03315_),
    .Y(_03451_));
 sg13g2_a221oi_1 _20817_ (.B2(_03072_),
    .C1(_03342_),
    .B1(_03451_),
    .A1(_09054_),
    .Y(_03452_),
    .A2(_03450_));
 sg13g2_nor3_1 _20818_ (.A(net122),
    .B(_03449_),
    .C(_03452_),
    .Y(_03453_));
 sg13g2_a21o_1 _20819_ (.A2(_03096_),
    .A1(_09087_),
    .B1(_03453_),
    .X(_00790_));
 sg13g2_buf_1 _20820_ (.A(net1134),
    .X(_03454_));
 sg13g2_buf_1 _20821_ (.A(net981),
    .X(_03455_));
 sg13g2_nand2b_1 _20822_ (.Y(_03456_),
    .B(net1116),
    .A_N(net1037));
 sg13g2_buf_1 _20823_ (.A(_03456_),
    .X(_03457_));
 sg13g2_nand3_1 _20824_ (.B(_11374_),
    .C(_10136_),
    .A(net1117),
    .Y(_03458_));
 sg13g2_buf_1 _20825_ (.A(_03458_),
    .X(_03459_));
 sg13g2_nor2_1 _20826_ (.A(_03457_),
    .B(_03459_),
    .Y(_03460_));
 sg13g2_buf_1 _20827_ (.A(_03460_),
    .X(_03461_));
 sg13g2_buf_1 _20828_ (.A(net612),
    .X(_03462_));
 sg13g2_mux2_1 _20829_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net853),
    .S(net555),
    .X(_00795_));
 sg13g2_mux2_1 _20830_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net856),
    .S(net555),
    .X(_00796_));
 sg13g2_buf_1 _20831_ (.A(_10693_),
    .X(_03463_));
 sg13g2_nand2_1 _20832_ (.Y(_03464_),
    .A(_03463_),
    .B(net612));
 sg13g2_o21ai_1 _20833_ (.B1(_03464_),
    .Y(_00797_),
    .A1(_10706_),
    .A2(net555));
 sg13g2_buf_1 _20834_ (.A(net695),
    .X(_03465_));
 sg13g2_buf_1 _20835_ (.A(net611),
    .X(_03466_));
 sg13g2_mux2_1 _20836_ (.A0(\cpu.ex.r_10[12] ),
    .A1(net554),
    .S(net555),
    .X(_00798_));
 sg13g2_buf_1 _20837_ (.A(net696),
    .X(_03467_));
 sg13g2_buf_1 _20838_ (.A(net610),
    .X(_03468_));
 sg13g2_mux2_1 _20839_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net553),
    .S(net555),
    .X(_00799_));
 sg13g2_buf_1 _20840_ (.A(_09492_),
    .X(_03469_));
 sg13g2_mux2_1 _20841_ (.A0(\cpu.ex.r_10[14] ),
    .A1(_03469_),
    .S(_03462_),
    .X(_00800_));
 sg13g2_buf_1 _20842_ (.A(net904),
    .X(_03470_));
 sg13g2_mux2_1 _20843_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net744),
    .S(_03462_),
    .X(_00801_));
 sg13g2_buf_1 _20844_ (.A(net797),
    .X(_03471_));
 sg13g2_buf_1 _20845_ (.A(net673),
    .X(_03472_));
 sg13g2_buf_1 _20846_ (.A(net609),
    .X(_03473_));
 sg13g2_mux2_1 _20847_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net552),
    .S(net555),
    .X(_00802_));
 sg13g2_nand2_1 _20848_ (.Y(_03474_),
    .A(net506),
    .B(net612));
 sg13g2_o21ai_1 _20849_ (.B1(_03474_),
    .Y(_00803_),
    .A1(_10521_),
    .A2(net555));
 sg13g2_buf_1 _20850_ (.A(net507),
    .X(_03475_));
 sg13g2_nand2_1 _20851_ (.Y(_03476_),
    .A(net435),
    .B(net612));
 sg13g2_o21ai_1 _20852_ (.B1(_03476_),
    .Y(_00804_),
    .A1(_10508_),
    .A2(net555));
 sg13g2_buf_1 _20853_ (.A(net681),
    .X(_03477_));
 sg13g2_buf_2 _20854_ (.A(net608),
    .X(_03478_));
 sg13g2_buf_1 _20855_ (.A(net551),
    .X(_03479_));
 sg13g2_mux2_1 _20856_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net477),
    .S(net612),
    .X(_00805_));
 sg13g2_mux2_1 _20857_ (.A0(\cpu.ex.r_10[5] ),
    .A1(net556),
    .S(net612),
    .X(_00806_));
 sg13g2_mux2_1 _20858_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net746),
    .S(_03461_),
    .X(_00807_));
 sg13g2_mux2_1 _20859_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net745),
    .S(net612),
    .X(_00808_));
 sg13g2_mux2_1 _20860_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net858),
    .S(net612),
    .X(_00809_));
 sg13g2_mux2_1 _20861_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net857),
    .S(_03461_),
    .X(_00810_));
 sg13g2_nor2_1 _20862_ (.A(_10145_),
    .B(_03459_),
    .Y(_03480_));
 sg13g2_buf_2 _20863_ (.A(_03480_),
    .X(_03481_));
 sg13g2_buf_1 _20864_ (.A(_03481_),
    .X(_03482_));
 sg13g2_mux2_1 _20865_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net853),
    .S(net550),
    .X(_00811_));
 sg13g2_mux2_1 _20866_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net856),
    .S(net550),
    .X(_00812_));
 sg13g2_mux2_1 _20867_ (.A0(\cpu.ex.r_11[11] ),
    .A1(_02956_),
    .S(net550),
    .X(_00813_));
 sg13g2_mux2_1 _20868_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net554),
    .S(net550),
    .X(_00814_));
 sg13g2_mux2_1 _20869_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net553),
    .S(net550),
    .X(_00815_));
 sg13g2_mux2_1 _20870_ (.A0(\cpu.ex.r_11[14] ),
    .A1(net674),
    .S(_03482_),
    .X(_00816_));
 sg13g2_mux2_1 _20871_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net744),
    .S(_03482_),
    .X(_00817_));
 sg13g2_mux2_1 _20872_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net552),
    .S(net550),
    .X(_00818_));
 sg13g2_buf_1 _20873_ (.A(net506),
    .X(_03483_));
 sg13g2_mux2_1 _20874_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net434),
    .S(net550),
    .X(_00819_));
 sg13g2_nand2_1 _20875_ (.Y(_03484_),
    .A(net435),
    .B(_03481_));
 sg13g2_o21ai_1 _20876_ (.B1(_03484_),
    .Y(_00820_),
    .A1(_11213_),
    .A2(net550));
 sg13g2_mux2_1 _20877_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net477),
    .S(_03481_),
    .X(_00821_));
 sg13g2_mux2_1 _20878_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net556),
    .S(_03481_),
    .X(_00822_));
 sg13g2_mux2_1 _20879_ (.A0(\cpu.ex.r_11[6] ),
    .A1(net746),
    .S(_03481_),
    .X(_00823_));
 sg13g2_mux2_1 _20880_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net745),
    .S(_03481_),
    .X(_00824_));
 sg13g2_mux2_1 _20881_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net858),
    .S(_03481_),
    .X(_00825_));
 sg13g2_mux2_1 _20882_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net857),
    .S(_03481_),
    .X(_00826_));
 sg13g2_nand3_1 _20883_ (.B(_10140_),
    .C(_10136_),
    .A(net1117),
    .Y(_03485_));
 sg13g2_buf_1 _20884_ (.A(_03485_),
    .X(_03486_));
 sg13g2_nor3_1 _20885_ (.A(net1116),
    .B(net1037),
    .C(_03486_),
    .Y(_03487_));
 sg13g2_buf_2 _20886_ (.A(_03487_),
    .X(_03488_));
 sg13g2_buf_1 _20887_ (.A(_03488_),
    .X(_03489_));
 sg13g2_mux2_1 _20888_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net853),
    .S(net607),
    .X(_00827_));
 sg13g2_mux2_1 _20889_ (.A0(\cpu.ex.r_12[10] ),
    .A1(_02954_),
    .S(net607),
    .X(_00828_));
 sg13g2_mux2_1 _20890_ (.A0(\cpu.ex.r_12[11] ),
    .A1(_02956_),
    .S(net607),
    .X(_00829_));
 sg13g2_mux2_1 _20891_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net554),
    .S(net607),
    .X(_00830_));
 sg13g2_mux2_1 _20892_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net553),
    .S(net607),
    .X(_00831_));
 sg13g2_mux2_1 _20893_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net674),
    .S(_03489_),
    .X(_00832_));
 sg13g2_mux2_1 _20894_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net744),
    .S(_03489_),
    .X(_00833_));
 sg13g2_mux2_1 _20895_ (.A0(\cpu.ex.r_12[1] ),
    .A1(_03473_),
    .S(net607),
    .X(_00834_));
 sg13g2_mux2_1 _20896_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net434),
    .S(net607),
    .X(_00835_));
 sg13g2_mux2_1 _20897_ (.A0(\cpu.ex.r_12[3] ),
    .A1(net435),
    .S(net607),
    .X(_00836_));
 sg13g2_mux2_1 _20898_ (.A0(\cpu.ex.r_12[4] ),
    .A1(_03479_),
    .S(_03488_),
    .X(_00837_));
 sg13g2_mux2_1 _20899_ (.A0(\cpu.ex.r_12[5] ),
    .A1(net556),
    .S(_03488_),
    .X(_00838_));
 sg13g2_mux2_1 _20900_ (.A0(\cpu.ex.r_12[6] ),
    .A1(_02946_),
    .S(_03488_),
    .X(_00839_));
 sg13g2_mux2_1 _20901_ (.A0(\cpu.ex.r_12[7] ),
    .A1(_02948_),
    .S(_03488_),
    .X(_00840_));
 sg13g2_mux2_1 _20902_ (.A0(\cpu.ex.r_12[8] ),
    .A1(_02950_),
    .S(_03488_),
    .X(_00841_));
 sg13g2_mux2_1 _20903_ (.A0(\cpu.ex.r_12[9] ),
    .A1(_02952_),
    .S(_03488_),
    .X(_00842_));
 sg13g2_inv_1 _20904_ (.Y(_03490_),
    .A(net1116));
 sg13g2_nand2_1 _20905_ (.Y(_03491_),
    .A(_03490_),
    .B(net1037));
 sg13g2_nor2_1 _20906_ (.A(_03486_),
    .B(_03491_),
    .Y(_03492_));
 sg13g2_buf_2 _20907_ (.A(_03492_),
    .X(_03493_));
 sg13g2_buf_1 _20908_ (.A(_03493_),
    .X(_03494_));
 sg13g2_mux2_1 _20909_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net853),
    .S(net606),
    .X(_00843_));
 sg13g2_mux2_1 _20910_ (.A0(\cpu.ex.r_13[10] ),
    .A1(_02954_),
    .S(net606),
    .X(_00844_));
 sg13g2_buf_1 _20911_ (.A(_02955_),
    .X(_03495_));
 sg13g2_mux2_1 _20912_ (.A0(\cpu.ex.r_13[11] ),
    .A1(net852),
    .S(net606),
    .X(_00845_));
 sg13g2_inv_1 _20913_ (.Y(_03496_),
    .A(\cpu.ex.r_13[12] ));
 sg13g2_nand2_1 _20914_ (.Y(_03497_),
    .A(net611),
    .B(_03493_));
 sg13g2_o21ai_1 _20915_ (.B1(_03497_),
    .Y(_00846_),
    .A1(_03496_),
    .A2(net606));
 sg13g2_mux2_1 _20916_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net553),
    .S(net606),
    .X(_00847_));
 sg13g2_mux2_1 _20917_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net674),
    .S(_03494_),
    .X(_00848_));
 sg13g2_mux2_1 _20918_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net744),
    .S(_03494_),
    .X(_00849_));
 sg13g2_mux2_1 _20919_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net552),
    .S(net606),
    .X(_00850_));
 sg13g2_mux2_1 _20920_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net434),
    .S(net606),
    .X(_00851_));
 sg13g2_mux2_1 _20921_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net435),
    .S(net606),
    .X(_00852_));
 sg13g2_mux2_1 _20922_ (.A0(\cpu.ex.r_13[4] ),
    .A1(_03479_),
    .S(_03493_),
    .X(_00853_));
 sg13g2_mux2_1 _20923_ (.A0(\cpu.ex.r_13[5] ),
    .A1(_02979_),
    .S(_03493_),
    .X(_00854_));
 sg13g2_mux2_1 _20924_ (.A0(\cpu.ex.r_13[6] ),
    .A1(_02946_),
    .S(_03493_),
    .X(_00855_));
 sg13g2_mux2_1 _20925_ (.A0(\cpu.ex.r_13[7] ),
    .A1(_02948_),
    .S(_03493_),
    .X(_00856_));
 sg13g2_mux2_1 _20926_ (.A0(\cpu.ex.r_13[8] ),
    .A1(_02950_),
    .S(_03493_),
    .X(_00857_));
 sg13g2_mux2_1 _20927_ (.A0(\cpu.ex.r_13[9] ),
    .A1(_02952_),
    .S(_03493_),
    .X(_00858_));
 sg13g2_nor2_1 _20928_ (.A(_03457_),
    .B(_03486_),
    .Y(_03498_));
 sg13g2_buf_1 _20929_ (.A(_03498_),
    .X(_03499_));
 sg13g2_buf_1 _20930_ (.A(_03498_),
    .X(_03500_));
 sg13g2_nand2_1 _20931_ (.Y(_03501_),
    .A(net853),
    .B(net604));
 sg13g2_o21ai_1 _20932_ (.B1(_03501_),
    .Y(_00859_),
    .A1(_11171_),
    .A2(net605));
 sg13g2_buf_1 _20933_ (.A(net984),
    .X(_03502_));
 sg13g2_mux2_1 _20934_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net851),
    .S(_03499_),
    .X(_00860_));
 sg13g2_mux2_1 _20935_ (.A0(\cpu.ex.r_14[11] ),
    .A1(net852),
    .S(net605),
    .X(_00861_));
 sg13g2_mux2_1 _20936_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net554),
    .S(net605),
    .X(_00862_));
 sg13g2_mux2_1 _20937_ (.A0(\cpu.ex.r_14[13] ),
    .A1(net553),
    .S(net605),
    .X(_00863_));
 sg13g2_nand2_1 _20938_ (.Y(_03503_),
    .A(net783),
    .B(net604));
 sg13g2_o21ai_1 _20939_ (.B1(_03503_),
    .Y(_00864_),
    .A1(_10272_),
    .A2(net605));
 sg13g2_mux2_1 _20940_ (.A0(\cpu.ex.r_14[15] ),
    .A1(_03470_),
    .S(net605),
    .X(_00865_));
 sg13g2_nand2_1 _20941_ (.Y(_03504_),
    .A(net552),
    .B(net604));
 sg13g2_o21ai_1 _20942_ (.B1(_03504_),
    .Y(_00866_),
    .A1(_10576_),
    .A2(net605));
 sg13g2_mux2_1 _20943_ (.A0(\cpu.ex.r_14[2] ),
    .A1(_03483_),
    .S(net605),
    .X(_00867_));
 sg13g2_mux2_1 _20944_ (.A0(\cpu.ex.r_14[3] ),
    .A1(_03475_),
    .S(net604),
    .X(_00868_));
 sg13g2_mux2_1 _20945_ (.A0(\cpu.ex.r_14[4] ),
    .A1(net477),
    .S(net604),
    .X(_00869_));
 sg13g2_nand2_1 _20946_ (.Y(_03505_),
    .A(net613),
    .B(net604));
 sg13g2_o21ai_1 _20947_ (.B1(_03505_),
    .Y(_00870_),
    .A1(_10619_),
    .A2(_03499_));
 sg13g2_buf_1 _20948_ (.A(net860),
    .X(_03506_));
 sg13g2_mux2_1 _20949_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net743),
    .S(_03500_),
    .X(_00871_));
 sg13g2_buf_1 _20950_ (.A(net859),
    .X(_03507_));
 sg13g2_mux2_1 _20951_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net742),
    .S(net604),
    .X(_00872_));
 sg13g2_buf_1 _20952_ (.A(net986),
    .X(_03508_));
 sg13g2_mux2_1 _20953_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net850),
    .S(net604),
    .X(_00873_));
 sg13g2_buf_1 _20954_ (.A(net985),
    .X(_03509_));
 sg13g2_mux2_1 _20955_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net849),
    .S(_03500_),
    .X(_00874_));
 sg13g2_nor2_1 _20956_ (.A(_10145_),
    .B(_03486_),
    .Y(_03510_));
 sg13g2_buf_2 _20957_ (.A(_03510_),
    .X(_03511_));
 sg13g2_buf_1 _20958_ (.A(_03511_),
    .X(_03512_));
 sg13g2_mux2_1 _20959_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net853),
    .S(net603),
    .X(_00875_));
 sg13g2_mux2_1 _20960_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net851),
    .S(net603),
    .X(_00876_));
 sg13g2_mux2_1 _20961_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net852),
    .S(net603),
    .X(_00877_));
 sg13g2_mux2_1 _20962_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net554),
    .S(net603),
    .X(_00878_));
 sg13g2_mux2_1 _20963_ (.A0(\cpu.ex.r_15[13] ),
    .A1(net553),
    .S(net603),
    .X(_00879_));
 sg13g2_mux2_1 _20964_ (.A0(\cpu.ex.r_15[14] ),
    .A1(net674),
    .S(_03512_),
    .X(_00880_));
 sg13g2_mux2_1 _20965_ (.A0(\cpu.ex.r_15[15] ),
    .A1(net744),
    .S(net603),
    .X(_00881_));
 sg13g2_mux2_1 _20966_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net552),
    .S(net603),
    .X(_00882_));
 sg13g2_mux2_1 _20967_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net434),
    .S(_03512_),
    .X(_00883_));
 sg13g2_mux2_1 _20968_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net435),
    .S(net603),
    .X(_00884_));
 sg13g2_mux2_1 _20969_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net477),
    .S(_03511_),
    .X(_00885_));
 sg13g2_mux2_1 _20970_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net556),
    .S(_03511_),
    .X(_00886_));
 sg13g2_mux2_1 _20971_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net743),
    .S(_03511_),
    .X(_00887_));
 sg13g2_mux2_1 _20972_ (.A0(\cpu.ex.r_15[7] ),
    .A1(net742),
    .S(_03511_),
    .X(_00888_));
 sg13g2_mux2_1 _20973_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net850),
    .S(_03511_),
    .X(_00889_));
 sg13g2_mux2_1 _20974_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net849),
    .S(_03511_),
    .X(_00890_));
 sg13g2_nor3_1 _20975_ (.A(net1116),
    .B(net1037),
    .C(_03459_),
    .Y(_03513_));
 sg13g2_buf_2 _20976_ (.A(_03513_),
    .X(_03514_));
 sg13g2_buf_1 _20977_ (.A(_03514_),
    .X(_03515_));
 sg13g2_mux2_1 _20978_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net853),
    .S(net549),
    .X(_00891_));
 sg13g2_mux2_1 _20979_ (.A0(\cpu.ex.r_8[10] ),
    .A1(net851),
    .S(net549),
    .X(_00892_));
 sg13g2_mux2_1 _20980_ (.A0(\cpu.ex.r_8[11] ),
    .A1(net852),
    .S(net549),
    .X(_00893_));
 sg13g2_mux2_1 _20981_ (.A0(\cpu.ex.r_8[12] ),
    .A1(net554),
    .S(net549),
    .X(_00894_));
 sg13g2_mux2_1 _20982_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net553),
    .S(net549),
    .X(_00895_));
 sg13g2_mux2_1 _20983_ (.A0(\cpu.ex.r_8[14] ),
    .A1(net674),
    .S(_03515_),
    .X(_00896_));
 sg13g2_mux2_1 _20984_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net744),
    .S(_03515_),
    .X(_00897_));
 sg13g2_mux2_1 _20985_ (.A0(\cpu.ex.r_8[1] ),
    .A1(_03473_),
    .S(net549),
    .X(_00898_));
 sg13g2_mux2_1 _20986_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net434),
    .S(net549),
    .X(_00899_));
 sg13g2_nand2_1 _20987_ (.Y(_03516_),
    .A(_03475_),
    .B(_03514_));
 sg13g2_o21ai_1 _20988_ (.B1(_03516_),
    .Y(_00900_),
    .A1(_10491_),
    .A2(net549));
 sg13g2_mux2_1 _20989_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net477),
    .S(_03514_),
    .X(_00901_));
 sg13g2_mux2_1 _20990_ (.A0(\cpu.ex.r_8[5] ),
    .A1(net556),
    .S(_03514_),
    .X(_00902_));
 sg13g2_mux2_1 _20991_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net743),
    .S(_03514_),
    .X(_00903_));
 sg13g2_mux2_1 _20992_ (.A0(\cpu.ex.r_8[7] ),
    .A1(net742),
    .S(_03514_),
    .X(_00904_));
 sg13g2_mux2_1 _20993_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net850),
    .S(_03514_),
    .X(_00905_));
 sg13g2_mux2_1 _20994_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net849),
    .S(_03514_),
    .X(_00906_));
 sg13g2_nor2_1 _20995_ (.A(_03459_),
    .B(_03491_),
    .Y(_03517_));
 sg13g2_buf_2 _20996_ (.A(_03517_),
    .X(_03518_));
 sg13g2_buf_1 _20997_ (.A(_03518_),
    .X(_03519_));
 sg13g2_mux2_1 _20998_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net853),
    .S(net548),
    .X(_00907_));
 sg13g2_mux2_1 _20999_ (.A0(\cpu.ex.r_9[10] ),
    .A1(net851),
    .S(net548),
    .X(_00908_));
 sg13g2_mux2_1 _21000_ (.A0(\cpu.ex.r_9[11] ),
    .A1(net852),
    .S(net548),
    .X(_00909_));
 sg13g2_mux2_1 _21001_ (.A0(\cpu.ex.r_9[12] ),
    .A1(net554),
    .S(net548),
    .X(_00910_));
 sg13g2_buf_1 _21002_ (.A(net610),
    .X(_03520_));
 sg13g2_mux2_1 _21003_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net547),
    .S(net548),
    .X(_00911_));
 sg13g2_mux2_1 _21004_ (.A0(\cpu.ex.r_9[14] ),
    .A1(net674),
    .S(_03519_),
    .X(_00912_));
 sg13g2_mux2_1 _21005_ (.A0(\cpu.ex.r_9[15] ),
    .A1(_03470_),
    .S(_03519_),
    .X(_00913_));
 sg13g2_nand2_1 _21006_ (.Y(_03521_),
    .A(net552),
    .B(_03518_));
 sg13g2_o21ai_1 _21007_ (.B1(_03521_),
    .Y(_00914_),
    .A1(_10572_),
    .A2(net548));
 sg13g2_mux2_1 _21008_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net434),
    .S(net548),
    .X(_00915_));
 sg13g2_mux2_1 _21009_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net435),
    .S(net548),
    .X(_00916_));
 sg13g2_mux2_1 _21010_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net477),
    .S(_03518_),
    .X(_00917_));
 sg13g2_mux2_1 _21011_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net556),
    .S(_03518_),
    .X(_00918_));
 sg13g2_mux2_1 _21012_ (.A0(\cpu.ex.r_9[6] ),
    .A1(net743),
    .S(_03518_),
    .X(_00919_));
 sg13g2_mux2_1 _21013_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net742),
    .S(_03518_),
    .X(_00920_));
 sg13g2_mux2_1 _21014_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net850),
    .S(_03518_),
    .X(_00921_));
 sg13g2_mux2_1 _21015_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net849),
    .S(_03518_),
    .X(_00922_));
 sg13g2_nand4_1 _21016_ (.B(_10144_),
    .C(_10136_),
    .A(_10142_),
    .Y(_03522_),
    .D(_10163_));
 sg13g2_nor2_1 _21017_ (.A(_08286_),
    .B(_03522_),
    .Y(_03523_));
 sg13g2_buf_2 _21018_ (.A(_03523_),
    .X(_03524_));
 sg13g2_buf_1 _21019_ (.A(_03524_),
    .X(_03525_));
 sg13g2_mux2_1 _21020_ (.A0(\cpu.ex.r_epc[1] ),
    .A1(net552),
    .S(net602),
    .X(_00924_));
 sg13g2_mux2_1 _21021_ (.A0(\cpu.ex.r_epc[11] ),
    .A1(net852),
    .S(net602),
    .X(_00925_));
 sg13g2_mux2_1 _21022_ (.A0(\cpu.ex.r_epc[12] ),
    .A1(net554),
    .S(net602),
    .X(_00926_));
 sg13g2_mux2_1 _21023_ (.A0(\cpu.ex.r_epc[13] ),
    .A1(net547),
    .S(net602),
    .X(_00927_));
 sg13g2_mux2_1 _21024_ (.A0(\cpu.ex.r_epc[14] ),
    .A1(net674),
    .S(_03525_),
    .X(_00928_));
 sg13g2_mux2_1 _21025_ (.A0(\cpu.ex.r_epc[15] ),
    .A1(net744),
    .S(_03525_),
    .X(_00929_));
 sg13g2_mux2_1 _21026_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(net434),
    .S(net602),
    .X(_00930_));
 sg13g2_mux2_1 _21027_ (.A0(\cpu.ex.r_epc[3] ),
    .A1(net435),
    .S(net602),
    .X(_00931_));
 sg13g2_mux2_1 _21028_ (.A0(\cpu.ex.r_epc[4] ),
    .A1(net477),
    .S(net602),
    .X(_00932_));
 sg13g2_mux2_1 _21029_ (.A0(\cpu.ex.r_epc[5] ),
    .A1(net556),
    .S(net602),
    .X(_00933_));
 sg13g2_mux2_1 _21030_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net743),
    .S(_03524_),
    .X(_00934_));
 sg13g2_mux2_1 _21031_ (.A0(\cpu.ex.r_epc[7] ),
    .A1(net742),
    .S(_03524_),
    .X(_00935_));
 sg13g2_mux2_1 _21032_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net850),
    .S(_03524_),
    .X(_00936_));
 sg13g2_mux2_1 _21033_ (.A0(\cpu.ex.r_epc[9] ),
    .A1(net849),
    .S(_03524_),
    .X(_00937_));
 sg13g2_mux2_1 _21034_ (.A0(\cpu.ex.r_epc[10] ),
    .A1(net851),
    .S(_03524_),
    .X(_00938_));
 sg13g2_buf_1 _21035_ (.A(net780),
    .X(_03526_));
 sg13g2_buf_1 _21036_ (.A(net672),
    .X(_03527_));
 sg13g2_nand4_1 _21037_ (.B(net1037),
    .C(_10136_),
    .A(_03490_),
    .Y(_03528_),
    .D(_10163_));
 sg13g2_buf_1 _21038_ (.A(_03528_),
    .X(_03529_));
 sg13g2_buf_1 _21039_ (.A(net741),
    .X(_03530_));
 sg13g2_buf_1 _21040_ (.A(net741),
    .X(_03531_));
 sg13g2_nand2_1 _21041_ (.Y(_03532_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net670));
 sg13g2_o21ai_1 _21042_ (.B1(_03532_),
    .Y(_00944_),
    .A1(net601),
    .A2(net671));
 sg13g2_nand2_1 _21043_ (.Y(_03533_),
    .A(\cpu.ex.r_lr[11] ),
    .B(net670));
 sg13g2_o21ai_1 _21044_ (.B1(_03533_),
    .Y(_00945_),
    .A1(_11032_),
    .A2(_03530_));
 sg13g2_nand2_1 _21045_ (.Y(_03534_),
    .A(\cpu.ex.r_lr[12] ),
    .B(_03531_));
 sg13g2_o21ai_1 _21046_ (.B1(_03534_),
    .Y(_00946_),
    .A1(_09576_),
    .A2(_03530_));
 sg13g2_buf_1 _21047_ (.A(net610),
    .X(_03535_));
 sg13g2_mux2_1 _21048_ (.A0(net546),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net670),
    .X(_00947_));
 sg13g2_buf_1 _21049_ (.A(_09493_),
    .X(_03536_));
 sg13g2_buf_1 _21050_ (.A(net600),
    .X(_03537_));
 sg13g2_nand2_1 _21051_ (.Y(_03538_),
    .A(\cpu.ex.r_lr[14] ),
    .B(net670));
 sg13g2_o21ai_1 _21052_ (.B1(_03538_),
    .Y(_00948_),
    .A1(net545),
    .A2(net671));
 sg13g2_buf_1 _21053_ (.A(net630),
    .X(_03539_));
 sg13g2_nand2_1 _21054_ (.Y(_03540_),
    .A(\cpu.ex.r_lr[15] ),
    .B(net670));
 sg13g2_o21ai_1 _21055_ (.B1(_03540_),
    .Y(_00949_),
    .A1(net544),
    .A2(net671));
 sg13g2_buf_2 _21056_ (.A(net782),
    .X(_03541_));
 sg13g2_nand2_1 _21057_ (.Y(_03542_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net741));
 sg13g2_o21ai_1 _21058_ (.B1(_03542_),
    .Y(_00950_),
    .A1(net669),
    .A2(net671));
 sg13g2_nand2_1 _21059_ (.Y(_03543_),
    .A(\cpu.ex.r_lr[3] ),
    .B(net741));
 sg13g2_o21ai_1 _21060_ (.B1(_03543_),
    .Y(_00951_),
    .A1(net679),
    .A2(net671));
 sg13g2_buf_1 _21061_ (.A(net680),
    .X(_03544_));
 sg13g2_buf_1 _21062_ (.A(_03544_),
    .X(_03545_));
 sg13g2_nand2_1 _21063_ (.Y(_03546_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net741));
 sg13g2_o21ai_1 _21064_ (.B1(_03546_),
    .Y(_00952_),
    .A1(net543),
    .A2(net671));
 sg13g2_mux2_1 _21065_ (.A0(net558),
    .A1(\cpu.ex.r_lr[5] ),
    .S(net670),
    .X(_00953_));
 sg13g2_nand2_1 _21066_ (.Y(_03547_),
    .A(\cpu.ex.r_lr[6] ),
    .B(net741));
 sg13g2_o21ai_1 _21067_ (.B1(_03547_),
    .Y(_00954_),
    .A1(net675),
    .A2(net671));
 sg13g2_nand2_1 _21068_ (.Y(_03548_),
    .A(\cpu.ex.r_lr[7] ),
    .B(net741));
 sg13g2_o21ai_1 _21069_ (.B1(_03548_),
    .Y(_00955_),
    .A1(net750),
    .A2(net671));
 sg13g2_nand2_1 _21070_ (.Y(_03549_),
    .A(\cpu.ex.r_lr[8] ),
    .B(net741));
 sg13g2_o21ai_1 _21071_ (.B1(_03549_),
    .Y(_00956_),
    .A1(_02926_),
    .A2(net670));
 sg13g2_nand2_1 _21072_ (.Y(_03550_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_03529_));
 sg13g2_o21ai_1 _21073_ (.B1(_03550_),
    .Y(_00957_),
    .A1(net748),
    .A2(_03531_));
 sg13g2_nand2_1 _21074_ (.Y(_03551_),
    .A(\cpu.ex.r_lr[10] ),
    .B(_03529_));
 sg13g2_o21ai_1 _21075_ (.B1(_03551_),
    .Y(_00958_),
    .A1(net747),
    .A2(net670));
 sg13g2_inv_1 _21076_ (.Y(_03552_),
    .A(net1134));
 sg13g2_buf_1 _21077_ (.A(net625),
    .X(_03553_));
 sg13g2_or4_1 _21078_ (.A(_11350_),
    .B(_11353_),
    .C(_11357_),
    .D(_11362_),
    .X(_03554_));
 sg13g2_buf_2 _21079_ (.A(_03554_),
    .X(_03555_));
 sg13g2_a21oi_1 _21080_ (.A1(net277),
    .A2(_03555_),
    .Y(_03556_),
    .B1(_11457_));
 sg13g2_or3_1 _21081_ (.A(_10540_),
    .B(_10551_),
    .C(_10565_),
    .X(_03557_));
 sg13g2_buf_1 _21082_ (.A(_03557_),
    .X(_03558_));
 sg13g2_buf_1 _21083_ (.A(_03558_),
    .X(_03559_));
 sg13g2_nor3_1 _21084_ (.A(net272),
    .B(net78),
    .C(net28),
    .Y(_03560_));
 sg13g2_buf_1 _21085_ (.A(net85),
    .X(_03561_));
 sg13g2_o21ai_1 _21086_ (.B1(_03561_),
    .Y(_03562_),
    .A1(_03556_),
    .A2(_03560_));
 sg13g2_buf_1 _21087_ (.A(_11700_),
    .X(_03563_));
 sg13g2_nand2_1 _21088_ (.Y(_03564_),
    .A(\cpu.ex.r_mult[15] ),
    .B(net445));
 sg13g2_nand2_1 _21089_ (.Y(_03565_),
    .A(net1105),
    .B(_11759_));
 sg13g2_a21o_1 _21090_ (.A2(net118),
    .A1(_11361_),
    .B1(_03565_),
    .X(_03566_));
 sg13g2_mux2_1 _21091_ (.A0(_11757_),
    .A1(_11759_),
    .S(net235),
    .X(_03567_));
 sg13g2_a22oi_1 _21092_ (.Y(_03568_),
    .B1(_03567_),
    .B2(_11736_),
    .A2(_10247_),
    .A1(_09278_));
 sg13g2_nor2_1 _21093_ (.A(net141),
    .B(_03568_),
    .Y(_03569_));
 sg13g2_nor4_1 _21094_ (.A(_11771_),
    .B(net235),
    .C(_10291_),
    .D(_11717_),
    .Y(_03570_));
 sg13g2_o21ai_1 _21095_ (.B1(net118),
    .Y(_03571_),
    .A1(_03569_),
    .A2(_03570_));
 sg13g2_a221oi_1 _21096_ (.B2(_03571_),
    .C1(_11728_),
    .B1(_03566_),
    .A1(_11596_),
    .Y(_03572_),
    .A2(_11604_));
 sg13g2_buf_1 _21097_ (.A(_03572_),
    .X(_03573_));
 sg13g2_a21oi_1 _21098_ (.A1(_11757_),
    .A2(net235),
    .Y(_03574_),
    .B1(_11717_));
 sg13g2_and2_1 _21099_ (.A(_10291_),
    .B(_11759_),
    .X(_03575_));
 sg13g2_o21ai_1 _21100_ (.B1(_11715_),
    .Y(_03576_),
    .A1(_03574_),
    .A2(_03575_));
 sg13g2_nor3_1 _21101_ (.A(net504),
    .B(net235),
    .C(net141),
    .Y(_03577_));
 sg13g2_and2_1 _21102_ (.A(_10291_),
    .B(_03574_),
    .X(_03578_));
 sg13g2_a221oi_1 _21103_ (.B2(_11715_),
    .C1(_03578_),
    .B1(_03577_),
    .A1(_10247_),
    .Y(_03579_),
    .A2(_11759_));
 sg13g2_a21oi_1 _21104_ (.A1(_03576_),
    .A2(_03579_),
    .Y(_03580_),
    .B1(_11457_));
 sg13g2_nor2_1 _21105_ (.A(_03573_),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_xor2_1 _21106_ (.B(_03581_),
    .A(_03564_),
    .X(_03582_));
 sg13g2_a221oi_1 _21107_ (.B2(_09277_),
    .C1(net625),
    .B1(_03582_),
    .A1(\cpu.ex.r_mult[16] ),
    .Y(_03583_),
    .A2(net271));
 sg13g2_a22oi_1 _21108_ (.Y(_00959_),
    .B1(_03562_),
    .B2(_03583_),
    .A2(_03553_),
    .A1(_03552_));
 sg13g2_nor2_1 _21109_ (.A(net79),
    .B(_03555_),
    .Y(_03584_));
 sg13g2_buf_1 _21110_ (.A(net236),
    .X(_03585_));
 sg13g2_nor2_1 _21111_ (.A(net272),
    .B(net118),
    .Y(_03586_));
 sg13g2_xnor2_1 _21112_ (.Y(_03587_),
    .A(_03585_),
    .B(_03586_));
 sg13g2_nand2b_1 _21113_ (.Y(_03588_),
    .B(_03587_),
    .A_N(_11245_));
 sg13g2_or3_1 _21114_ (.A(_11244_),
    .B(net450),
    .C(_03587_),
    .X(_03589_));
 sg13g2_o21ai_1 _21115_ (.B1(_03589_),
    .Y(_03590_),
    .A1(_11364_),
    .A2(_03588_));
 sg13g2_nand2_1 _21116_ (.Y(_03591_),
    .A(_09277_),
    .B(net402));
 sg13g2_o21ai_1 _21117_ (.B1(\cpu.ex.r_mult[15] ),
    .Y(_03592_),
    .A1(_03573_),
    .A2(_03580_));
 sg13g2_buf_2 _21118_ (.A(_03592_),
    .X(_03593_));
 sg13g2_xnor2_1 _21119_ (.Y(_03594_),
    .A(_11244_),
    .B(_03593_));
 sg13g2_a21oi_1 _21120_ (.A1(\cpu.ex.r_mult[17] ),
    .A2(net271),
    .Y(_03595_),
    .B1(_10147_));
 sg13g2_o21ai_1 _21121_ (.B1(_03595_),
    .Y(_03596_),
    .A1(_03591_),
    .A2(_03594_));
 sg13g2_a221oi_1 _21122_ (.B2(net75),
    .C1(_03596_),
    .B1(_03590_),
    .A1(_11245_),
    .Y(_03597_),
    .A2(_03584_));
 sg13g2_a21oi_1 _21123_ (.A1(net601),
    .A2(_03553_),
    .Y(_00960_),
    .B1(_03597_));
 sg13g2_o21ai_1 _21124_ (.B1(_11287_),
    .Y(_03598_),
    .A1(net272),
    .A2(net87));
 sg13g2_and2_1 _21125_ (.A(_11246_),
    .B(_03598_),
    .X(_03599_));
 sg13g2_xnor2_1 _21126_ (.Y(_03600_),
    .A(net233),
    .B(_03599_));
 sg13g2_nor2_1 _21127_ (.A(_11255_),
    .B(_03600_),
    .Y(_03601_));
 sg13g2_nor2_1 _21128_ (.A(net877),
    .B(net401),
    .Y(_03602_));
 sg13g2_buf_1 _21129_ (.A(_03602_),
    .X(_03603_));
 sg13g2_nor2_1 _21130_ (.A(_11254_),
    .B(_11244_),
    .Y(_03604_));
 sg13g2_nand2b_1 _21131_ (.Y(_03605_),
    .B(_03604_),
    .A_N(_03593_));
 sg13g2_o21ai_1 _21132_ (.B1(_11254_),
    .Y(_03606_),
    .A1(_11244_),
    .A2(_03593_));
 sg13g2_nand3_1 _21133_ (.B(_03605_),
    .C(_03606_),
    .A(_03603_),
    .Y(_03607_));
 sg13g2_a21oi_1 _21134_ (.A1(\cpu.ex.r_mult[18] ),
    .A2(_03563_),
    .Y(_03608_),
    .B1(net691));
 sg13g2_nand2_1 _21135_ (.Y(_03609_),
    .A(_03607_),
    .B(_03608_));
 sg13g2_a21oi_1 _21136_ (.A1(_11366_),
    .A2(_03601_),
    .Y(_03610_),
    .B1(_03609_));
 sg13g2_nor2_1 _21137_ (.A(_10724_),
    .B(_11285_),
    .Y(_03611_));
 sg13g2_a22oi_1 _21138_ (.Y(_03612_),
    .B1(_03600_),
    .B2(_03611_),
    .A2(_03584_),
    .A1(_11255_));
 sg13g2_a22oi_1 _21139_ (.Y(_00961_),
    .B1(_03610_),
    .B2(_03612_),
    .A2(net542),
    .A1(net669));
 sg13g2_buf_1 _21140_ (.A(_03603_),
    .X(_03613_));
 sg13g2_xnor2_1 _21141_ (.Y(_03614_),
    .A(_11315_),
    .B(_03605_));
 sg13g2_and2_1 _21142_ (.A(_11246_),
    .B(_11256_),
    .X(_03615_));
 sg13g2_a221oi_1 _21143_ (.B2(_03586_),
    .C1(_11288_),
    .B1(_03615_),
    .A1(net233),
    .Y(_03616_),
    .A2(_11285_));
 sg13g2_buf_1 _21144_ (.A(_03616_),
    .X(_03617_));
 sg13g2_xnor2_1 _21145_ (.Y(_03618_),
    .A(net231),
    .B(_03617_));
 sg13g2_nor2_1 _21146_ (.A(net403),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_mux2_1 _21147_ (.A0(net403),
    .A1(_03619_),
    .S(_03555_),
    .X(_03620_));
 sg13g2_nand3_1 _21148_ (.B(net403),
    .C(_03618_),
    .A(net75),
    .Y(_03621_));
 sg13g2_a21oi_1 _21149_ (.A1(\cpu.ex.r_mult[19] ),
    .A2(_03563_),
    .Y(_03622_),
    .B1(net691));
 sg13g2_nand2_1 _21150_ (.Y(_03623_),
    .A(_03621_),
    .B(_03622_));
 sg13g2_a221oi_1 _21151_ (.B2(net75),
    .C1(_03623_),
    .B1(_03620_),
    .A1(net224),
    .Y(_03624_),
    .A2(_03614_));
 sg13g2_a21oi_1 _21152_ (.A1(net679),
    .A2(net542),
    .Y(_00962_),
    .B1(_03624_));
 sg13g2_inv_1 _21153_ (.Y(_03625_),
    .A(net281));
 sg13g2_a21o_1 _21154_ (.A2(_03617_),
    .A1(net403),
    .B1(net231),
    .X(_03626_));
 sg13g2_o21ai_1 _21155_ (.B1(_03626_),
    .Y(_03627_),
    .A1(net403),
    .A2(_03617_));
 sg13g2_xnor2_1 _21156_ (.Y(_03628_),
    .A(_03625_),
    .B(_03627_));
 sg13g2_and2_1 _21157_ (.A(_03561_),
    .B(_11273_),
    .X(_03629_));
 sg13g2_o21ai_1 _21158_ (.B1(_03629_),
    .Y(_03630_),
    .A1(net28),
    .A2(_03628_));
 sg13g2_nor3_1 _21159_ (.A(net79),
    .B(_11273_),
    .C(_03628_),
    .Y(_03631_));
 sg13g2_nor2_1 _21160_ (.A(_00291_),
    .B(_03605_),
    .Y(_03632_));
 sg13g2_xnor2_1 _21161_ (.Y(_03633_),
    .A(_11272_),
    .B(_03632_));
 sg13g2_a221oi_1 _21162_ (.B2(_03613_),
    .C1(net214),
    .B1(_03633_),
    .A1(_03555_),
    .Y(_03634_),
    .A2(_03631_));
 sg13g2_nor3_1 _21163_ (.A(\cpu.ex.r_mult[20] ),
    .B(_10148_),
    .C(_11381_),
    .Y(_03635_));
 sg13g2_a221oi_1 _21164_ (.B2(_03634_),
    .C1(_03635_),
    .B1(_03630_),
    .A1(net599),
    .Y(_00963_),
    .A2(net625));
 sg13g2_nand2_1 _21165_ (.Y(_03636_),
    .A(net281),
    .B(_11273_));
 sg13g2_or2_1 _21166_ (.X(_03637_),
    .B(_11273_),
    .A(net281));
 sg13g2_nand3_1 _21167_ (.B(net403),
    .C(_03637_),
    .A(net231),
    .Y(_03638_));
 sg13g2_nand2_1 _21168_ (.Y(_03639_),
    .A(_03636_),
    .B(_03638_));
 sg13g2_xnor2_1 _21169_ (.Y(_03640_),
    .A(net213),
    .B(net403));
 sg13g2_and3_1 _21170_ (.X(_03641_),
    .A(_03637_),
    .B(_03636_),
    .C(_03640_));
 sg13g2_and2_1 _21171_ (.A(_03617_),
    .B(_03641_),
    .X(_03642_));
 sg13g2_nor2_1 _21172_ (.A(_03639_),
    .B(_03642_),
    .Y(_03643_));
 sg13g2_xnor2_1 _21173_ (.Y(_03644_),
    .A(net216),
    .B(_03643_));
 sg13g2_nand3b_1 _21174_ (.B(_11366_),
    .C(_03644_),
    .Y(_03645_),
    .A_N(_11266_));
 sg13g2_nor3_2 _21175_ (.A(_11350_),
    .B(_11353_),
    .C(_11357_),
    .Y(_03646_));
 sg13g2_and4_1 _21176_ (.A(net75),
    .B(_11334_),
    .C(_11343_),
    .D(_03646_),
    .X(_03647_));
 sg13g2_buf_1 _21177_ (.A(_03647_),
    .X(_03648_));
 sg13g2_a21oi_1 _21178_ (.A1(net210),
    .A2(_11352_),
    .Y(_03649_),
    .B1(net142));
 sg13g2_or4_1 _21179_ (.A(_11350_),
    .B(_11353_),
    .C(_11355_),
    .D(_03649_),
    .X(_03650_));
 sg13g2_buf_1 _21180_ (.A(_03650_),
    .X(_03651_));
 sg13g2_nand2_1 _21181_ (.Y(_03652_),
    .A(_03644_),
    .B(_03651_));
 sg13g2_and2_1 _21182_ (.A(net75),
    .B(_11266_),
    .X(_03653_));
 sg13g2_nor2_1 _21183_ (.A(net1023),
    .B(net401),
    .Y(_03654_));
 sg13g2_nand3_1 _21184_ (.B(_11315_),
    .C(_03604_),
    .A(_11301_),
    .Y(_03655_));
 sg13g2_nor2_1 _21185_ (.A(_03564_),
    .B(_03655_),
    .Y(_03656_));
 sg13g2_o21ai_1 _21186_ (.B1(_03656_),
    .Y(_03657_),
    .A1(_03573_),
    .A2(_03580_));
 sg13g2_buf_2 _21187_ (.A(_03657_),
    .X(_03658_));
 sg13g2_mux2_1 _21188_ (.A0(net1023),
    .A1(_03654_),
    .S(_03658_),
    .X(_03659_));
 sg13g2_a21o_1 _21189_ (.A2(_03659_),
    .A1(net1124),
    .B1(net214),
    .X(_03660_));
 sg13g2_a221oi_1 _21190_ (.B2(_03653_),
    .C1(_03660_),
    .B1(_03652_),
    .A1(_11266_),
    .Y(_03661_),
    .A2(_03648_));
 sg13g2_nand2_1 _21191_ (.Y(_03662_),
    .A(net613),
    .B(net625));
 sg13g2_o21ai_1 _21192_ (.B1(net568),
    .Y(_03663_),
    .A1(\cpu.ex.r_mult[21] ),
    .A2(_11381_));
 sg13g2_a22oi_1 _21193_ (.Y(_00964_),
    .B1(_03662_),
    .B2(_03663_),
    .A2(_03661_),
    .A1(_03645_));
 sg13g2_xnor2_1 _21194_ (.Y(_03664_),
    .A(_11499_),
    .B(_11266_));
 sg13g2_nand4_1 _21195_ (.B(_11293_),
    .C(_03641_),
    .A(_11256_),
    .Y(_03665_),
    .D(_03664_));
 sg13g2_inv_1 _21196_ (.Y(_03666_),
    .A(_10660_));
 sg13g2_a21oi_1 _21197_ (.A1(_11286_),
    .A2(_11292_),
    .Y(_03667_),
    .B1(net231));
 sg13g2_a21oi_1 _21198_ (.A1(_11256_),
    .A2(_11317_),
    .Y(_03668_),
    .B1(_03667_));
 sg13g2_a21oi_1 _21199_ (.A1(net281),
    .A2(_03668_),
    .Y(_03669_),
    .B1(net216));
 sg13g2_a21oi_1 _21200_ (.A1(net1023),
    .A2(_11499_),
    .Y(_03670_),
    .B1(_11272_));
 sg13g2_o21ai_1 _21201_ (.B1(_03670_),
    .Y(_03671_),
    .A1(net281),
    .A2(_03668_));
 sg13g2_o21ai_1 _21202_ (.B1(_03671_),
    .Y(_03672_),
    .A1(_11261_),
    .A2(_03669_));
 sg13g2_a22oi_1 _21203_ (.Y(_03673_),
    .B1(_03672_),
    .B2(_11316_),
    .A2(_03668_),
    .A1(_03666_));
 sg13g2_o21ai_1 _21204_ (.B1(_03673_),
    .Y(_03674_),
    .A1(_03599_),
    .A2(_03665_));
 sg13g2_xnor2_1 _21205_ (.Y(_03675_),
    .A(net230),
    .B(_03674_));
 sg13g2_a21oi_1 _21206_ (.A1(_03651_),
    .A2(_03675_),
    .Y(_03676_),
    .B1(net79));
 sg13g2_o21ai_1 _21207_ (.B1(_11263_),
    .Y(_03677_),
    .A1(_03648_),
    .A2(_03676_));
 sg13g2_and2_1 _21208_ (.A(_11264_),
    .B(_03675_),
    .X(_03678_));
 sg13g2_nor3_1 _21209_ (.A(net1023),
    .B(_03593_),
    .C(_03655_),
    .Y(_03679_));
 sg13g2_xnor2_1 _21210_ (.Y(_03680_),
    .A(_11258_),
    .B(_03679_));
 sg13g2_a21o_1 _21211_ (.A2(net271),
    .A1(\cpu.ex.r_mult[22] ),
    .B1(net691),
    .X(_03681_));
 sg13g2_a221oi_1 _21212_ (.B2(_03613_),
    .C1(_03681_),
    .B1(_03680_),
    .A1(_11366_),
    .Y(_03682_),
    .A2(_03678_));
 sg13g2_a22oi_1 _21213_ (.Y(_00965_),
    .B1(_03677_),
    .B2(_03682_),
    .A2(net542),
    .A1(net675));
 sg13g2_nand3b_1 _21214_ (.B(net568),
    .C(_11700_),
    .Y(_03683_),
    .A_N(\cpu.ex.r_mult[23] ));
 sg13g2_o21ai_1 _21215_ (.B1(_03683_),
    .Y(_03684_),
    .A1(net1057),
    .A2(net568));
 sg13g2_or4_1 _21216_ (.A(_11258_),
    .B(net1023),
    .C(_03593_),
    .D(_03655_),
    .X(_03685_));
 sg13g2_buf_2 _21217_ (.A(_03685_),
    .X(_03686_));
 sg13g2_xor2_1 _21218_ (.B(_03686_),
    .A(net1110),
    .X(_03687_));
 sg13g2_a21o_1 _21219_ (.A2(_11260_),
    .A1(net216),
    .B1(_11270_),
    .X(_03688_));
 sg13g2_a21o_1 _21220_ (.A2(_11265_),
    .A1(_11262_),
    .B1(_03688_),
    .X(_03689_));
 sg13g2_nand2_1 _21221_ (.Y(_03690_),
    .A(net216),
    .B(_03639_));
 sg13g2_inv_1 _21222_ (.Y(_03691_),
    .A(_03639_));
 sg13g2_a221oi_1 _21223_ (.B2(_11499_),
    .C1(_11261_),
    .B1(_03691_),
    .A1(_11258_),
    .Y(_03692_),
    .A2(net230));
 sg13g2_a21oi_1 _21224_ (.A1(net230),
    .A2(_03690_),
    .Y(_03693_),
    .B1(_11258_));
 sg13g2_o21ai_1 _21225_ (.B1(_11316_),
    .Y(_03694_),
    .A1(_03692_),
    .A2(_03693_));
 sg13g2_o21ai_1 _21226_ (.B1(_03694_),
    .Y(_03695_),
    .A1(net230),
    .A2(_03690_));
 sg13g2_a21oi_1 _21227_ (.A1(_03689_),
    .A2(_03642_),
    .Y(_03696_),
    .B1(_03695_));
 sg13g2_xnor2_1 _21228_ (.Y(_03697_),
    .A(net242),
    .B(_03696_));
 sg13g2_nor2b_1 _21229_ (.A(_11277_),
    .B_N(_03697_),
    .Y(_03698_));
 sg13g2_a221oi_1 _21230_ (.B2(_11366_),
    .C1(net214),
    .B1(_03698_),
    .A1(net224),
    .Y(_03699_),
    .A2(_03687_));
 sg13g2_a21oi_1 _21231_ (.A1(_03651_),
    .A2(_03697_),
    .Y(_03700_),
    .B1(net79));
 sg13g2_nor3_1 _21232_ (.A(net1110),
    .B(net450),
    .C(_03684_),
    .Y(_03701_));
 sg13g2_o21ai_1 _21233_ (.B1(_03701_),
    .Y(_03702_),
    .A1(_03648_),
    .A2(_03700_));
 sg13g2_o21ai_1 _21234_ (.B1(_03702_),
    .Y(_00966_),
    .A1(_03684_),
    .A2(_03699_));
 sg13g2_buf_1 _21235_ (.A(_11297_),
    .X(_03703_));
 sg13g2_nand2_1 _21236_ (.Y(_03704_),
    .A(net74),
    .B(net97));
 sg13g2_xnor2_1 _21237_ (.Y(_03705_),
    .A(net192),
    .B(_03704_));
 sg13g2_nand2_1 _21238_ (.Y(_03706_),
    .A(_03651_),
    .B(_03705_));
 sg13g2_nor2_1 _21239_ (.A(net79),
    .B(_10750_),
    .Y(_03707_));
 sg13g2_o21ai_1 _21240_ (.B1(_03707_),
    .Y(_03708_),
    .A1(_03648_),
    .A2(_03706_));
 sg13g2_or3_1 _21241_ (.A(net1110),
    .B(_11258_),
    .C(net1023),
    .X(_03709_));
 sg13g2_buf_1 _21242_ (.A(_03709_),
    .X(_03710_));
 sg13g2_nor2_1 _21243_ (.A(_03658_),
    .B(_03710_),
    .Y(_03711_));
 sg13g2_xnor2_1 _21244_ (.Y(_03712_),
    .A(_10737_),
    .B(_03711_));
 sg13g2_and2_1 _21245_ (.A(_10750_),
    .B(_03705_),
    .X(_03713_));
 sg13g2_a21o_1 _21246_ (.A2(net271),
    .A1(\cpu.ex.r_mult[24] ),
    .B1(net691),
    .X(_03714_));
 sg13g2_a221oi_1 _21247_ (.B2(_11366_),
    .C1(_03714_),
    .B1(_03713_),
    .A1(net224),
    .Y(_03715_),
    .A2(_03712_));
 sg13g2_a22oi_1 _21248_ (.Y(_00967_),
    .B1(_03708_),
    .B2(_03715_),
    .A2(net542),
    .A1(net749));
 sg13g2_nor3_1 _21249_ (.A(_10737_),
    .B(net1110),
    .C(_03686_),
    .Y(_03716_));
 sg13g2_xnor2_1 _21250_ (.Y(_03717_),
    .A(_10725_),
    .B(_03716_));
 sg13g2_a221oi_1 _21251_ (.B2(_03717_),
    .C1(net625),
    .B1(net224),
    .A1(\cpu.ex.r_mult[25] ),
    .Y(_03718_),
    .A2(net271));
 sg13g2_inv_1 _21252_ (.Y(_03719_),
    .A(net446));
 sg13g2_a21oi_1 _21253_ (.A1(_03703_),
    .A2(_11336_),
    .Y(_03720_),
    .B1(_10750_));
 sg13g2_nand3_1 _21254_ (.B(_03703_),
    .C(_11336_),
    .A(_10750_),
    .Y(_03721_));
 sg13g2_o21ai_1 _21255_ (.B1(_03721_),
    .Y(_03722_),
    .A1(net191),
    .A2(_03720_));
 sg13g2_xnor2_1 _21256_ (.Y(_03723_),
    .A(net212),
    .B(_03722_));
 sg13g2_nand3_1 _21257_ (.B(_11362_),
    .C(_03723_),
    .A(_03719_),
    .Y(_03724_));
 sg13g2_o21ai_1 _21258_ (.B1(_03724_),
    .Y(_03725_),
    .A1(_03719_),
    .A2(_03723_));
 sg13g2_nor3_1 _21259_ (.A(net79),
    .B(net446),
    .C(_03646_),
    .Y(_03726_));
 sg13g2_nor3_1 _21260_ (.A(net79),
    .B(_03719_),
    .C(_03555_),
    .Y(_03727_));
 sg13g2_a221oi_1 _21261_ (.B2(_03723_),
    .C1(_03727_),
    .B1(_03726_),
    .A1(net75),
    .Y(_03728_),
    .A2(_03725_));
 sg13g2_a22oi_1 _21262_ (.Y(_00968_),
    .B1(_03718_),
    .B2(_03728_),
    .A2(net542),
    .A1(net748));
 sg13g2_buf_1 _21263_ (.A(_10762_),
    .X(_03729_));
 sg13g2_nand3b_1 _21264_ (.B(_10749_),
    .C(net445),
    .Y(_03730_),
    .A_N(_10725_));
 sg13g2_buf_1 _21265_ (.A(_03730_),
    .X(_03731_));
 sg13g2_nor3_1 _21266_ (.A(net1110),
    .B(_03686_),
    .C(_03731_),
    .Y(_03732_));
 sg13g2_xnor2_1 _21267_ (.Y(_03733_),
    .A(_10740_),
    .B(_03732_));
 sg13g2_a21o_1 _21268_ (.A2(net271),
    .A1(\cpu.ex.r_mult[26] ),
    .B1(net691),
    .X(_03734_));
 sg13g2_a221oi_1 _21269_ (.B2(net224),
    .C1(_03734_),
    .B1(_03733_),
    .A1(net392),
    .Y(_03735_),
    .A2(_03584_));
 sg13g2_nor2_1 _21270_ (.A(net212),
    .B(net446),
    .Y(_03736_));
 sg13g2_nand2_1 _21271_ (.Y(_03737_),
    .A(net212),
    .B(net446));
 sg13g2_o21ai_1 _21272_ (.B1(_03737_),
    .Y(_03738_),
    .A1(_03722_),
    .A2(_03736_));
 sg13g2_xnor2_1 _21273_ (.Y(_03739_),
    .A(net285),
    .B(_03738_));
 sg13g2_nor3_1 _21274_ (.A(net392),
    .B(net28),
    .C(_03739_),
    .Y(_03740_));
 sg13g2_and2_1 _21275_ (.A(net392),
    .B(_03739_),
    .X(_03741_));
 sg13g2_o21ai_1 _21276_ (.B1(net75),
    .Y(_03742_),
    .A1(_03740_),
    .A2(_03741_));
 sg13g2_a22oi_1 _21277_ (.Y(_00969_),
    .B1(_03735_),
    .B2(_03742_),
    .A2(net542),
    .A1(net747));
 sg13g2_nor4_1 _21278_ (.A(_10740_),
    .B(net1110),
    .C(_03686_),
    .D(_03731_),
    .Y(_03743_));
 sg13g2_xnor2_1 _21279_ (.Y(_03744_),
    .A(_10731_),
    .B(_03743_));
 sg13g2_a21oi_1 _21280_ (.A1(net224),
    .A2(_03744_),
    .Y(_03745_),
    .B1(net214));
 sg13g2_nor3_1 _21281_ (.A(net446),
    .B(_10756_),
    .C(net392),
    .Y(_03746_));
 sg13g2_nand3_1 _21282_ (.B(net97),
    .C(_03746_),
    .A(net74),
    .Y(_03747_));
 sg13g2_nor3_1 _21283_ (.A(net212),
    .B(_10756_),
    .C(net392),
    .Y(_03748_));
 sg13g2_nand3_1 _21284_ (.B(net97),
    .C(_03748_),
    .A(net74),
    .Y(_03749_));
 sg13g2_nand2_1 _21285_ (.Y(_03750_),
    .A(_03719_),
    .B(_10743_));
 sg13g2_nor2_1 _21286_ (.A(net191),
    .B(_03750_),
    .Y(_03751_));
 sg13g2_nand3_1 _21287_ (.B(net97),
    .C(_03751_),
    .A(net74),
    .Y(_03752_));
 sg13g2_nor3_1 _21288_ (.A(net212),
    .B(net191),
    .C(net392),
    .Y(_03753_));
 sg13g2_nand3_1 _21289_ (.B(net97),
    .C(_03753_),
    .A(net74),
    .Y(_03754_));
 sg13g2_nand4_1 _21290_ (.B(_03749_),
    .C(_03752_),
    .A(_03747_),
    .Y(_03755_),
    .D(_03754_));
 sg13g2_o21ai_1 _21291_ (.B1(net192),
    .Y(_03756_),
    .A1(_03746_),
    .A2(_03748_));
 sg13g2_o21ai_1 _21292_ (.B1(_03756_),
    .Y(_03757_),
    .A1(net212),
    .A2(_03750_));
 sg13g2_nand3_1 _21293_ (.B(_10756_),
    .C(net392),
    .A(_10727_),
    .Y(_03758_));
 sg13g2_nand3_1 _21294_ (.B(_10756_),
    .C(net392),
    .A(net243),
    .Y(_03759_));
 sg13g2_a22oi_1 _21295_ (.Y(_03760_),
    .B1(_03758_),
    .B2(_03759_),
    .A2(net97),
    .A1(net74));
 sg13g2_nand2_1 _21296_ (.Y(_03761_),
    .A(net446),
    .B(_03729_));
 sg13g2_nand2_1 _21297_ (.Y(_03762_),
    .A(net212),
    .B(_03729_));
 sg13g2_a221oi_1 _21298_ (.B2(_03762_),
    .C1(net192),
    .B1(_03761_),
    .A1(net74),
    .Y(_03763_),
    .A2(net97));
 sg13g2_a21oi_1 _21299_ (.A1(_03758_),
    .A2(_03759_),
    .Y(_03764_),
    .B1(net192));
 sg13g2_or2_1 _21300_ (.X(_03765_),
    .B(_03761_),
    .A(net228));
 sg13g2_nand2b_1 _21301_ (.Y(_03766_),
    .B(_03765_),
    .A_N(_03764_));
 sg13g2_nor4_1 _21302_ (.A(net285),
    .B(_03760_),
    .C(_03763_),
    .D(_03766_),
    .Y(_03767_));
 sg13g2_nor3_1 _21303_ (.A(_03755_),
    .B(_03757_),
    .C(_03767_),
    .Y(_03768_));
 sg13g2_xnor2_1 _21304_ (.Y(_03769_),
    .A(net280),
    .B(_03768_));
 sg13g2_o21ai_1 _21305_ (.B1(_10733_),
    .Y(_03770_),
    .A1(net28),
    .A2(_03769_));
 sg13g2_or3_1 _21306_ (.A(_10733_),
    .B(net28),
    .C(_03769_),
    .X(_03771_));
 sg13g2_a21o_1 _21307_ (.A2(_03771_),
    .A1(_03770_),
    .B1(_10724_),
    .X(_03772_));
 sg13g2_nor3_1 _21308_ (.A(\cpu.ex.r_mult[27] ),
    .B(net625),
    .C(_11381_),
    .Y(_03773_));
 sg13g2_a221oi_1 _21309_ (.B2(_03772_),
    .C1(_03773_),
    .B1(_03745_),
    .A1(_11032_),
    .Y(_00970_),
    .A2(net625));
 sg13g2_nor3_1 _21310_ (.A(_10773_),
    .B(_11312_),
    .C(_11318_),
    .Y(_03774_));
 sg13g2_a21oi_1 _21311_ (.A1(net74),
    .A2(_03774_),
    .Y(_03775_),
    .B1(_10774_));
 sg13g2_xnor2_1 _21312_ (.Y(_03776_),
    .A(net194),
    .B(_03775_));
 sg13g2_and3_1 _21313_ (.X(_03777_),
    .A(net85),
    .B(_11324_),
    .C(_03776_));
 sg13g2_nand2_1 _21314_ (.Y(_03778_),
    .A(net85),
    .B(_11337_));
 sg13g2_nor2_1 _21315_ (.A(_11362_),
    .B(_03778_),
    .Y(_03779_));
 sg13g2_mux2_1 _21316_ (.A0(_03777_),
    .A1(_03779_),
    .S(_03646_),
    .X(_03780_));
 sg13g2_or3_1 _21317_ (.A(_10731_),
    .B(_10740_),
    .C(_03731_),
    .X(_03781_));
 sg13g2_nor3_1 _21318_ (.A(_03658_),
    .B(_03710_),
    .C(_03781_),
    .Y(_03782_));
 sg13g2_xor2_1 _21319_ (.B(_03782_),
    .A(_11322_),
    .X(_03783_));
 sg13g2_nor2_1 _21320_ (.A(_03776_),
    .B(_03778_),
    .Y(_03784_));
 sg13g2_a221oi_1 _21321_ (.B2(_11362_),
    .C1(_03784_),
    .B1(_03777_),
    .A1(\cpu.ex.r_mult[28] ),
    .Y(_03785_),
    .A2(_11700_));
 sg13g2_o21ai_1 _21322_ (.B1(_03785_),
    .Y(_03786_),
    .A1(_03591_),
    .A2(_03783_));
 sg13g2_nor3_1 _21323_ (.A(net625),
    .B(_03780_),
    .C(_03786_),
    .Y(_03787_));
 sg13g2_a21oi_1 _21324_ (.A1(_09576_),
    .A2(net542),
    .Y(_00971_),
    .B1(_03787_));
 sg13g2_and3_1 _21325_ (.X(_03788_),
    .A(_11339_),
    .B(_11340_),
    .C(_11341_));
 sg13g2_buf_1 _21326_ (.A(_03788_),
    .X(_03789_));
 sg13g2_xnor2_1 _21327_ (.Y(_03790_),
    .A(net211),
    .B(_03789_));
 sg13g2_nand2_1 _21328_ (.Y(_03791_),
    .A(_03555_),
    .B(_03790_));
 sg13g2_xnor2_1 _21329_ (.Y(_03792_),
    .A(_11326_),
    .B(_03791_));
 sg13g2_or2_1 _21330_ (.X(_03793_),
    .B(_03781_),
    .A(_11322_));
 sg13g2_nor3_1 _21331_ (.A(_03658_),
    .B(_03710_),
    .C(_03793_),
    .Y(_03794_));
 sg13g2_xnor2_1 _21332_ (.Y(_03795_),
    .A(_11321_),
    .B(_03794_));
 sg13g2_a22oi_1 _21333_ (.Y(_03796_),
    .B1(net224),
    .B2(_03795_),
    .A2(net271),
    .A1(\cpu.ex.r_mult[29] ));
 sg13g2_nor2_1 _21334_ (.A(net696),
    .B(net568),
    .Y(_03797_));
 sg13g2_a21oi_1 _21335_ (.A1(net568),
    .A2(_03796_),
    .Y(_03798_),
    .B1(_03797_));
 sg13g2_a21o_1 _21336_ (.A2(_03792_),
    .A1(_11532_),
    .B1(_03798_),
    .X(_00972_));
 sg13g2_nand2_1 _21337_ (.Y(_03799_),
    .A(_11334_),
    .B(_11343_));
 sg13g2_xnor2_1 _21338_ (.Y(_03800_),
    .A(net142),
    .B(_03799_));
 sg13g2_nand2_1 _21339_ (.Y(_03801_),
    .A(net1109),
    .B(net210));
 sg13g2_nand3_1 _21340_ (.B(net500),
    .C(net75),
    .A(_11346_),
    .Y(_03802_));
 sg13g2_a21o_1 _21341_ (.A2(_03801_),
    .A1(_03800_),
    .B1(_03802_),
    .X(_03803_));
 sg13g2_nand2_1 _21342_ (.Y(_03804_),
    .A(net500),
    .B(net85));
 sg13g2_nor4_1 _21343_ (.A(net1109),
    .B(_11346_),
    .C(net210),
    .D(_03804_),
    .Y(_03805_));
 sg13g2_a22oi_1 _21344_ (.Y(_03806_),
    .B1(_03800_),
    .B2(_03805_),
    .A2(net271),
    .A1(\cpu.ex.r_mult[30] ));
 sg13g2_or4_1 _21345_ (.A(_11321_),
    .B(_03658_),
    .C(_03710_),
    .D(_03793_),
    .X(_03807_));
 sg13g2_buf_1 _21346_ (.A(_03807_),
    .X(_03808_));
 sg13g2_xnor2_1 _21347_ (.Y(_03809_),
    .A(_11346_),
    .B(_03808_));
 sg13g2_nand2_1 _21348_ (.Y(_03810_),
    .A(net224),
    .B(_03809_));
 sg13g2_and4_1 _21349_ (.A(net568),
    .B(_03803_),
    .C(_03806_),
    .D(_03810_),
    .X(_03811_));
 sg13g2_a21oi_1 _21350_ (.A1(_03537_),
    .A2(net542),
    .Y(_00973_),
    .B1(_03811_));
 sg13g2_a21oi_1 _21351_ (.A1(net142),
    .A2(_11347_),
    .Y(_03812_),
    .B1(_11343_));
 sg13g2_nor2_1 _21352_ (.A(net142),
    .B(_11347_),
    .Y(_03813_));
 sg13g2_o21ai_1 _21353_ (.B1(net235),
    .Y(_03814_),
    .A1(_03812_),
    .A2(_03813_));
 sg13g2_nand3_1 _21354_ (.B(_11346_),
    .C(_03603_),
    .A(net1109),
    .Y(_03815_));
 sg13g2_nand2b_1 _21355_ (.Y(_03816_),
    .B(_03603_),
    .A_N(net1109));
 sg13g2_mux2_1 _21356_ (.A0(_03815_),
    .A1(_03816_),
    .S(_03808_),
    .X(_03817_));
 sg13g2_nor2_1 _21357_ (.A(net1109),
    .B(_11346_),
    .Y(_03818_));
 sg13g2_a22oi_1 _21358_ (.Y(_03819_),
    .B1(_03603_),
    .B2(_03818_),
    .A2(_11700_),
    .A1(\cpu.ex.r_mult[31] ));
 sg13g2_nand3_1 _21359_ (.B(_03817_),
    .C(_03819_),
    .A(net568),
    .Y(_03820_));
 sg13g2_nor2_1 _21360_ (.A(_11321_),
    .B(net210),
    .Y(_03821_));
 sg13g2_o21ai_1 _21361_ (.B1(_03821_),
    .Y(_03822_),
    .A1(_11346_),
    .A2(net141));
 sg13g2_a21oi_1 _21362_ (.A1(net141),
    .A2(_03789_),
    .Y(_03823_),
    .B1(net500));
 sg13g2_a21oi_1 _21363_ (.A1(net500),
    .A2(_03789_),
    .Y(_03824_),
    .B1(net217));
 sg13g2_nor3_1 _21364_ (.A(_03822_),
    .B(_03823_),
    .C(_03824_),
    .Y(_03825_));
 sg13g2_nor3_1 _21365_ (.A(net28),
    .B(_03820_),
    .C(_03825_),
    .Y(_03826_));
 sg13g2_nor2_1 _21366_ (.A(net1109),
    .B(_03804_),
    .Y(_03827_));
 sg13g2_nand2_1 _21367_ (.Y(_03828_),
    .A(_09426_),
    .B(net691));
 sg13g2_o21ai_1 _21368_ (.B1(_03828_),
    .Y(_03829_),
    .A1(_03827_),
    .A2(_03820_));
 sg13g2_a21oi_1 _21369_ (.A1(_03814_),
    .A2(_03826_),
    .Y(_00974_),
    .B1(_03829_));
 sg13g2_inv_1 _21370_ (.Y(_03830_),
    .A(_00238_));
 sg13g2_nand2_1 _21371_ (.Y(_03831_),
    .A(_08331_),
    .B(_03830_));
 sg13g2_mux2_1 _21372_ (.A0(_03831_),
    .A1(net1132),
    .S(_11796_),
    .X(_03832_));
 sg13g2_and2_1 _21373_ (.A(_11159_),
    .B(_11160_),
    .X(_03833_));
 sg13g2_buf_2 _21374_ (.A(_03833_),
    .X(_03834_));
 sg13g2_nand3b_1 _21375_ (.B(_03834_),
    .C(net710),
    .Y(_03835_),
    .A_N(_03832_));
 sg13g2_buf_1 _21376_ (.A(_03835_),
    .X(_03836_));
 sg13g2_buf_1 _21377_ (.A(_03836_),
    .X(_03837_));
 sg13g2_buf_1 _21378_ (.A(_11389_),
    .X(_03838_));
 sg13g2_buf_1 _21379_ (.A(net239),
    .X(_03839_));
 sg13g2_nand2b_1 _21380_ (.Y(_03840_),
    .B(net201),
    .A_N(_10959_));
 sg13g2_o21ai_1 _21381_ (.B1(_03840_),
    .Y(_03841_),
    .A1(_10392_),
    .A2(net201));
 sg13g2_buf_2 _21382_ (.A(_03841_),
    .X(_03842_));
 sg13g2_buf_1 _21383_ (.A(_03842_),
    .X(_03843_));
 sg13g2_nor2_1 _21384_ (.A(net234),
    .B(net115),
    .Y(_03844_));
 sg13g2_nor2_1 _21385_ (.A(net202),
    .B(net237),
    .Y(_03845_));
 sg13g2_nand2_1 _21386_ (.Y(_03846_),
    .A(net232),
    .B(net283));
 sg13g2_buf_1 _21387_ (.A(_03846_),
    .X(_03847_));
 sg13g2_nor4_1 _21388_ (.A(net277),
    .B(_03844_),
    .C(_03845_),
    .D(net183),
    .Y(_03848_));
 sg13g2_nand2b_1 _21389_ (.Y(_03849_),
    .B(net239),
    .A_N(_11090_));
 sg13g2_o21ai_1 _21390_ (.B1(_03849_),
    .Y(_03850_),
    .A1(_10457_),
    .A2(_10796_));
 sg13g2_buf_1 _21391_ (.A(_03850_),
    .X(_03851_));
 sg13g2_buf_1 _21392_ (.A(_03851_),
    .X(_03852_));
 sg13g2_buf_1 _21393_ (.A(net139),
    .X(_03853_));
 sg13g2_nand2_2 _21394_ (.Y(_03854_),
    .A(_03558_),
    .B(net282));
 sg13g2_nor3_1 _21395_ (.A(net232),
    .B(net278),
    .C(_03854_),
    .Y(_03855_));
 sg13g2_buf_1 _21396_ (.A(_03855_),
    .X(_03856_));
 sg13g2_buf_1 _21397_ (.A(net182),
    .X(_03857_));
 sg13g2_nand2_1 _21398_ (.Y(_03858_),
    .A(net359),
    .B(net236));
 sg13g2_buf_1 _21399_ (.A(_03858_),
    .X(_03859_));
 sg13g2_nor3_1 _21400_ (.A(net213),
    .B(net278),
    .C(_03859_),
    .Y(_03860_));
 sg13g2_buf_1 _21401_ (.A(_03860_),
    .X(_03861_));
 sg13g2_buf_1 _21402_ (.A(_03861_),
    .X(_03862_));
 sg13g2_nand2b_1 _21403_ (.Y(_03863_),
    .B(net201),
    .A_N(_11071_));
 sg13g2_o21ai_1 _21404_ (.B1(_03863_),
    .Y(_03864_),
    .A1(_10330_),
    .A2(_03839_));
 sg13g2_buf_2 _21405_ (.A(_03864_),
    .X(_03865_));
 sg13g2_buf_1 _21406_ (.A(_03865_),
    .X(_03866_));
 sg13g2_a22oi_1 _21407_ (.Y(_03867_),
    .B1(net113),
    .B2(net112),
    .A2(net165),
    .A1(net114));
 sg13g2_nand2_2 _21408_ (.Y(_03868_),
    .A(net272),
    .B(net236));
 sg13g2_o21ai_1 _21409_ (.B1(_11253_),
    .Y(_03869_),
    .A1(_10487_),
    .A2(_10514_));
 sg13g2_buf_2 _21410_ (.A(_03869_),
    .X(_03870_));
 sg13g2_nor2_1 _21411_ (.A(_03868_),
    .B(_03870_),
    .Y(_03871_));
 sg13g2_buf_1 _21412_ (.A(_03871_),
    .X(_03872_));
 sg13g2_nor2_2 _21413_ (.A(net183),
    .B(_03859_),
    .Y(_03873_));
 sg13g2_a22oi_1 _21414_ (.Y(_03874_),
    .B1(_03873_),
    .B2(net238),
    .A2(net164),
    .A1(net215));
 sg13g2_nand2_1 _21415_ (.Y(_03875_),
    .A(_03867_),
    .B(_03874_));
 sg13g2_nand2_1 _21416_ (.Y(_03876_),
    .A(net1130),
    .B(net237));
 sg13g2_buf_1 _21417_ (.A(_03876_),
    .X(_03877_));
 sg13g2_nand2_2 _21418_ (.Y(_03878_),
    .A(net359),
    .B(net234));
 sg13g2_nor3_1 _21419_ (.A(net183),
    .B(net181),
    .C(_03878_),
    .Y(_03879_));
 sg13g2_mux2_1 _21420_ (.A0(_10486_),
    .A1(_11235_),
    .S(net239),
    .X(_03880_));
 sg13g2_buf_1 _21421_ (.A(_03880_),
    .X(_03881_));
 sg13g2_nor2_1 _21422_ (.A(_10567_),
    .B(net236),
    .Y(_03882_));
 sg13g2_nand2_1 _21423_ (.Y(_03883_),
    .A(_10549_),
    .B(_03882_));
 sg13g2_nor2_1 _21424_ (.A(net180),
    .B(_03883_),
    .Y(_03884_));
 sg13g2_buf_1 _21425_ (.A(_11133_),
    .X(_03885_));
 sg13g2_nand3_1 _21426_ (.B(net283),
    .C(_10602_),
    .A(_11290_),
    .Y(_03886_));
 sg13g2_buf_1 _21427_ (.A(_03886_),
    .X(_03887_));
 sg13g2_nor2_1 _21428_ (.A(net179),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_nor3_1 _21429_ (.A(_03879_),
    .B(_03884_),
    .C(_03888_),
    .Y(_03889_));
 sg13g2_buf_1 _21430_ (.A(_11048_),
    .X(_03890_));
 sg13g2_buf_1 _21431_ (.A(net178),
    .X(_03891_));
 sg13g2_nor2_1 _21432_ (.A(_03854_),
    .B(_03870_),
    .Y(_03892_));
 sg13g2_buf_1 _21433_ (.A(_03892_),
    .X(_03893_));
 sg13g2_nor2_1 _21434_ (.A(_03859_),
    .B(_03870_),
    .Y(_03894_));
 sg13g2_buf_1 _21435_ (.A(_03894_),
    .X(_03895_));
 sg13g2_buf_1 _21436_ (.A(_11008_),
    .X(_03896_));
 sg13g2_inv_1 _21437_ (.Y(_03897_),
    .A(net177));
 sg13g2_a22oi_1 _21438_ (.Y(_03898_),
    .B1(_03895_),
    .B2(net161),
    .A2(net162),
    .A1(net163));
 sg13g2_buf_1 _21439_ (.A(net193),
    .X(_03899_));
 sg13g2_nor2_1 _21440_ (.A(_03870_),
    .B(_03878_),
    .Y(_03900_));
 sg13g2_buf_2 _21441_ (.A(_03900_),
    .X(_03901_));
 sg13g2_buf_1 _21442_ (.A(_10989_),
    .X(_03902_));
 sg13g2_nor2_1 _21443_ (.A(net272),
    .B(net236),
    .Y(_03903_));
 sg13g2_nand3_1 _21444_ (.B(net233),
    .C(_03903_),
    .A(net231),
    .Y(_03904_));
 sg13g2_buf_1 _21445_ (.A(_03904_),
    .X(_03905_));
 sg13g2_nor2_1 _21446_ (.A(_03902_),
    .B(_03905_),
    .Y(_03906_));
 sg13g2_a21oi_1 _21447_ (.A1(net160),
    .A2(_03901_),
    .Y(_03907_),
    .B1(_03906_));
 sg13g2_nand3_1 _21448_ (.B(_03898_),
    .C(_03907_),
    .A(_03889_),
    .Y(_03908_));
 sg13g2_buf_8 _21449_ (.A(_11113_),
    .X(_03909_));
 sg13g2_buf_1 _21450_ (.A(net175),
    .X(_03910_));
 sg13g2_o21ai_1 _21451_ (.B1(net277),
    .Y(_03911_),
    .A1(net202),
    .A2(net159));
 sg13g2_inv_1 _21452_ (.Y(_03912_),
    .A(net1130));
 sg13g2_mux2_1 _21453_ (.A0(_00176_),
    .A1(_11793_),
    .S(_03839_),
    .X(_03913_));
 sg13g2_buf_1 _21454_ (.A(_03913_),
    .X(_03914_));
 sg13g2_nor2_1 _21455_ (.A(_03912_),
    .B(_03914_),
    .Y(_03915_));
 sg13g2_nand2_1 _21456_ (.Y(_03916_),
    .A(net202),
    .B(_03915_));
 sg13g2_or3_1 _21457_ (.A(_10487_),
    .B(_10514_),
    .C(net283),
    .X(_03917_));
 sg13g2_buf_2 _21458_ (.A(_03917_),
    .X(_03918_));
 sg13g2_a21oi_1 _21459_ (.A1(_03911_),
    .A2(_03916_),
    .Y(_03919_),
    .B1(_03918_));
 sg13g2_nor4_1 _21460_ (.A(_03848_),
    .B(_03875_),
    .C(_03908_),
    .D(_03919_),
    .Y(_03920_));
 sg13g2_buf_1 _21461_ (.A(_11157_),
    .X(_03921_));
 sg13g2_nor2_1 _21462_ (.A(net272),
    .B(net282),
    .Y(_03922_));
 sg13g2_nand2_1 _21463_ (.Y(_03923_),
    .A(_10549_),
    .B(_03922_));
 sg13g2_buf_1 _21464_ (.A(_03923_),
    .X(_03924_));
 sg13g2_or2_1 _21465_ (.X(_03925_),
    .B(_09831_),
    .A(net1130));
 sg13g2_buf_1 _21466_ (.A(_03925_),
    .X(_03926_));
 sg13g2_o21ai_1 _21467_ (.B1(_03926_),
    .Y(_03927_),
    .A1(net174),
    .A2(net158));
 sg13g2_a21oi_2 _21468_ (.B1(_11161_),
    .Y(_03928_),
    .A2(_11160_),
    .A1(_11159_));
 sg13g2_a21o_1 _21469_ (.A2(_11185_),
    .A1(net459),
    .B1(_11186_),
    .X(_03929_));
 sg13g2_buf_1 _21470_ (.A(_03929_),
    .X(_03930_));
 sg13g2_nor2_2 _21471_ (.A(_03928_),
    .B(_03930_),
    .Y(_03931_));
 sg13g2_nand2b_1 _21472_ (.Y(_03932_),
    .B(_10791_),
    .A_N(_10596_));
 sg13g2_a21o_1 _21473_ (.A2(_10790_),
    .A1(net459),
    .B1(_03932_),
    .X(_03933_));
 sg13g2_buf_1 _21474_ (.A(_03933_),
    .X(_03934_));
 sg13g2_nor4_2 _21475_ (.A(_08330_),
    .B(_10789_),
    .C(_11191_),
    .Y(_03935_),
    .D(_11211_));
 sg13g2_nor3_1 _21476_ (.A(_10791_),
    .B(_11191_),
    .C(_11211_),
    .Y(_03936_));
 sg13g2_a21oi_2 _21477_ (.B1(_03936_),
    .Y(_03937_),
    .A2(_03935_),
    .A1(net459));
 sg13g2_nand3_1 _21478_ (.B(_03934_),
    .C(_03937_),
    .A(net282),
    .Y(_03938_));
 sg13g2_a21oi_2 _21479_ (.B1(_03932_),
    .Y(_03939_),
    .A2(_10790_),
    .A1(net459));
 sg13g2_a21o_1 _21480_ (.A2(_03935_),
    .A1(_08402_),
    .B1(_03936_),
    .X(_03940_));
 sg13g2_buf_1 _21481_ (.A(_03940_),
    .X(_03941_));
 sg13g2_o21ai_1 _21482_ (.B1(_11243_),
    .Y(_03942_),
    .A1(_03939_),
    .A2(_03941_));
 sg13g2_inv_1 _21483_ (.Y(_03943_),
    .A(net1077));
 sg13g2_nor2_1 _21484_ (.A(_03943_),
    .B(_03931_),
    .Y(_03944_));
 sg13g2_a221oi_1 _21485_ (.B2(_03942_),
    .C1(_03944_),
    .B1(_03938_),
    .A1(_09069_),
    .Y(_03945_),
    .A2(_03931_));
 sg13g2_o21ai_1 _21486_ (.B1(net277),
    .Y(_03946_),
    .A1(_09069_),
    .A2(_03931_));
 sg13g2_nor3_1 _21487_ (.A(net236),
    .B(_03939_),
    .C(_03941_),
    .Y(_03947_));
 sg13g2_a21oi_1 _21488_ (.A1(_03934_),
    .A2(_03937_),
    .Y(_03948_),
    .B1(net282));
 sg13g2_nor2_1 _21489_ (.A(_03947_),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_a22oi_1 _21490_ (.Y(_03950_),
    .B1(_03946_),
    .B2(_03949_),
    .A2(_03945_),
    .A1(net277));
 sg13g2_nand2_1 _21491_ (.Y(_03951_),
    .A(_03931_),
    .B(_03949_));
 sg13g2_a21o_1 _21492_ (.A2(_03951_),
    .A1(_09069_),
    .B1(net1077),
    .X(_03952_));
 sg13g2_nor2_1 _21493_ (.A(net1130),
    .B(_09831_),
    .Y(_03953_));
 sg13g2_buf_2 _21494_ (.A(_03953_),
    .X(_03954_));
 sg13g2_nor2_2 _21495_ (.A(_09069_),
    .B(_09078_),
    .Y(_03955_));
 sg13g2_nor2_1 _21496_ (.A(_08279_),
    .B(_09073_),
    .Y(_03956_));
 sg13g2_nor4_1 _21497_ (.A(_09048_),
    .B(_09834_),
    .C(net1121),
    .D(_09850_),
    .Y(_03957_));
 sg13g2_nand4_1 _21498_ (.B(_03955_),
    .C(_03956_),
    .A(_03954_),
    .Y(_03958_),
    .D(_03957_));
 sg13g2_buf_1 _21499_ (.A(_03958_),
    .X(_03959_));
 sg13g2_nand2b_1 _21500_ (.Y(_03960_),
    .B(_03959_),
    .A_N(_09078_));
 sg13g2_o21ai_1 _21501_ (.B1(_10566_),
    .Y(_03961_),
    .A1(_03928_),
    .A2(_03930_));
 sg13g2_xor2_1 _21502_ (.B(_03961_),
    .A(_03949_),
    .X(_03962_));
 sg13g2_nor3_1 _21503_ (.A(net282),
    .B(_03939_),
    .C(_03941_),
    .Y(_03963_));
 sg13g2_a21oi_1 _21504_ (.A1(_03934_),
    .A2(_03937_),
    .Y(_03964_),
    .B1(_11243_));
 sg13g2_mux2_1 _21505_ (.A0(_09073_),
    .A1(net1121),
    .S(_03964_),
    .X(_03965_));
 sg13g2_nor2_1 _21506_ (.A(_09834_),
    .B(_03965_),
    .Y(_03966_));
 sg13g2_nor2_1 _21507_ (.A(_03918_),
    .B(_03859_),
    .Y(_03967_));
 sg13g2_buf_1 _21508_ (.A(_03967_),
    .X(_03968_));
 sg13g2_inv_1 _21509_ (.Y(_03969_),
    .A(_09850_));
 sg13g2_nor2_1 _21510_ (.A(net979),
    .B(_03931_),
    .Y(_03970_));
 sg13g2_nor2b_1 _21511_ (.A(_11379_),
    .B_N(_11387_),
    .Y(_03971_));
 sg13g2_buf_1 _21512_ (.A(_03971_),
    .X(_03972_));
 sg13g2_a221oi_1 _21513_ (.B2(_03970_),
    .C1(_03972_),
    .B1(net137),
    .A1(_09048_),
    .Y(_03973_),
    .A2(net228));
 sg13g2_o21ai_1 _21514_ (.B1(_03973_),
    .Y(_03974_),
    .A1(_03963_),
    .A2(_03966_));
 sg13g2_a221oi_1 _21515_ (.B2(_03962_),
    .C1(_03974_),
    .B1(_03960_),
    .A1(_03950_),
    .Y(_03975_),
    .A2(_03952_));
 sg13g2_o21ai_1 _21516_ (.B1(_03975_),
    .Y(_03976_),
    .A1(_03920_),
    .A2(_03927_));
 sg13g2_o21ai_1 _21517_ (.B1(_03976_),
    .Y(_03977_),
    .A1(net166),
    .A2(\cpu.ex.c_mult[1] ));
 sg13g2_and3_1 _21518_ (.X(_03978_),
    .A(_03834_),
    .B(_11396_),
    .C(_11797_));
 sg13g2_buf_1 _21519_ (.A(_03978_),
    .X(_03979_));
 sg13g2_nand2_1 _21520_ (.Y(_03980_),
    .A(_11159_),
    .B(_11160_));
 sg13g2_buf_1 _21521_ (.A(_03980_),
    .X(_03981_));
 sg13g2_nor3_2 _21522_ (.A(_11395_),
    .B(net352),
    .C(_03832_),
    .Y(_03982_));
 sg13g2_inv_1 _21523_ (.Y(_03983_),
    .A(_09087_));
 sg13g2_nor3_1 _21524_ (.A(_03983_),
    .B(_08404_),
    .C(_09263_),
    .Y(_03984_));
 sg13g2_a21oi_1 _21525_ (.A1(net288),
    .A2(_09263_),
    .Y(_03985_),
    .B1(_03984_));
 sg13g2_nor2_1 _21526_ (.A(_08341_),
    .B(_03985_),
    .Y(_03986_));
 sg13g2_nor2_1 _21527_ (.A(_09087_),
    .B(_08404_),
    .Y(_03987_));
 sg13g2_nand3_1 _21528_ (.B(_09135_),
    .C(_11396_),
    .A(_03987_),
    .Y(_03988_));
 sg13g2_nand2_1 _21529_ (.Y(_03989_),
    .A(_09081_),
    .B(_03988_));
 sg13g2_nor4_1 _21530_ (.A(_03982_),
    .B(net94),
    .C(_03986_),
    .D(_03989_),
    .Y(_03990_));
 sg13g2_buf_1 _21531_ (.A(_03990_),
    .X(_03991_));
 sg13g2_buf_1 _21532_ (.A(_03991_),
    .X(_03992_));
 sg13g2_a22oi_1 _21533_ (.Y(_03993_),
    .B1(net35),
    .B2(net803),
    .A2(net94),
    .A1(_10596_));
 sg13g2_o21ai_1 _21534_ (.B1(_03993_),
    .Y(_00975_),
    .A1(net84),
    .A2(_03977_));
 sg13g2_mux2_1 _21535_ (.A0(_10330_),
    .A1(_11071_),
    .S(_10796_),
    .X(_03994_));
 sg13g2_buf_2 _21536_ (.A(_03994_),
    .X(_03995_));
 sg13g2_nand2_1 _21537_ (.Y(_03996_),
    .A(net286),
    .B(_03995_));
 sg13g2_nand2_1 _21538_ (.Y(_03997_),
    .A(_11290_),
    .B(_03881_));
 sg13g2_nand2_1 _21539_ (.Y(_03998_),
    .A(net241),
    .B(net179));
 sg13g2_nand3_1 _21540_ (.B(_03997_),
    .C(_03998_),
    .A(_03625_),
    .Y(_03999_));
 sg13g2_nand3_1 _21541_ (.B(_03997_),
    .C(_03998_),
    .A(net175),
    .Y(_04000_));
 sg13g2_nand2b_1 _21542_ (.Y(_04001_),
    .B(net239),
    .A_N(_11235_));
 sg13g2_o21ai_1 _21543_ (.B1(_04001_),
    .Y(_04002_),
    .A1(_10486_),
    .A2(net201));
 sg13g2_buf_1 _21544_ (.A(_04002_),
    .X(_04003_));
 sg13g2_a21o_1 _21545_ (.A2(_11153_),
    .A1(net619),
    .B1(_11154_),
    .X(_04004_));
 sg13g2_mux2_1 _21546_ (.A0(_00271_),
    .A1(_04004_),
    .S(net239),
    .X(_04005_));
 sg13g2_buf_2 _21547_ (.A(_04005_),
    .X(_04006_));
 sg13g2_nand2_1 _21548_ (.Y(_04007_),
    .A(net278),
    .B(_04006_));
 sg13g2_o21ai_1 _21549_ (.B1(_10601_),
    .Y(_04008_),
    .A1(_03939_),
    .A2(_03941_));
 sg13g2_o21ai_1 _21550_ (.B1(_04008_),
    .Y(_04009_),
    .A1(_03961_),
    .A2(_03963_));
 sg13g2_buf_1 _21551_ (.A(_04009_),
    .X(_04010_));
 sg13g2_nor2_1 _21552_ (.A(net278),
    .B(_04006_),
    .Y(_04011_));
 sg13g2_a221oi_1 _21553_ (.B2(_04010_),
    .C1(_04011_),
    .B1(_04007_),
    .A1(net232),
    .Y(_04012_),
    .A2(_04003_));
 sg13g2_buf_1 _21554_ (.A(_04012_),
    .X(_04013_));
 sg13g2_a21o_1 _21555_ (.A2(_04000_),
    .A1(_03999_),
    .B1(_04013_),
    .X(_04014_));
 sg13g2_nand2_1 _21556_ (.Y(_04015_),
    .A(_03625_),
    .B(net175));
 sg13g2_and2_1 _21557_ (.A(net241),
    .B(net179),
    .X(_04016_));
 sg13g2_or2_1 _21558_ (.X(_04017_),
    .B(net179),
    .A(net241));
 sg13g2_buf_2 _21559_ (.A(_04017_),
    .X(_04018_));
 sg13g2_o21ai_1 _21560_ (.B1(_04018_),
    .Y(_04019_),
    .A1(_04015_),
    .A2(_04016_));
 sg13g2_buf_1 _21561_ (.A(_04019_),
    .X(_04020_));
 sg13g2_inv_1 _21562_ (.Y(_04021_),
    .A(_04020_));
 sg13g2_nand2_1 _21563_ (.Y(_04022_),
    .A(net276),
    .B(_03865_));
 sg13g2_nand3_1 _21564_ (.B(_04021_),
    .C(_04022_),
    .A(_04014_),
    .Y(_04023_));
 sg13g2_mux2_1 _21565_ (.A0(_10457_),
    .A1(_11090_),
    .S(net201),
    .X(_04024_));
 sg13g2_buf_1 _21566_ (.A(_04024_),
    .X(_04025_));
 sg13g2_xnor2_1 _21567_ (.Y(_04026_),
    .A(net242),
    .B(_04025_));
 sg13g2_inv_1 _21568_ (.Y(_04027_),
    .A(_04026_));
 sg13g2_a21oi_1 _21569_ (.A1(_03996_),
    .A2(_04023_),
    .Y(_04028_),
    .B1(_04027_));
 sg13g2_nand3_1 _21570_ (.B(_04023_),
    .C(_04027_),
    .A(_03996_),
    .Y(_04029_));
 sg13g2_nand3b_1 _21571_ (.B(_04029_),
    .C(_09069_),
    .Y(_04030_),
    .A_N(_04028_));
 sg13g2_buf_1 _21572_ (.A(_04030_),
    .X(_04031_));
 sg13g2_nand2_1 _21573_ (.Y(_04032_),
    .A(_03959_),
    .B(_04031_));
 sg13g2_buf_1 _21574_ (.A(_09834_),
    .X(_04033_));
 sg13g2_and2_1 _21575_ (.A(net240),
    .B(net178),
    .X(_04034_));
 sg13g2_mux2_1 _21576_ (.A0(net1060),
    .A1(net1048),
    .S(_04034_),
    .X(_04035_));
 sg13g2_or2_1 _21577_ (.X(_04036_),
    .B(net178),
    .A(net240));
 sg13g2_buf_1 _21578_ (.A(_04036_),
    .X(_04037_));
 sg13g2_o21ai_1 _21579_ (.B1(_04037_),
    .Y(_04038_),
    .A1(_04033_),
    .A2(_04035_));
 sg13g2_buf_1 _21580_ (.A(_03972_),
    .X(_04039_));
 sg13g2_a21oi_1 _21581_ (.A1(_09049_),
    .A2(net213),
    .Y(_04040_),
    .B1(_04039_));
 sg13g2_nand2b_1 _21582_ (.Y(_04041_),
    .B(net201),
    .A_N(_10987_));
 sg13g2_o21ai_1 _21583_ (.B1(_04041_),
    .Y(_04042_),
    .A1(_10427_),
    .A2(net201));
 sg13g2_buf_1 _21584_ (.A(_04042_),
    .X(_04043_));
 sg13g2_nor2_1 _21585_ (.A(_03918_),
    .B(_03878_),
    .Y(_04044_));
 sg13g2_buf_1 _21586_ (.A(_04044_),
    .X(_04045_));
 sg13g2_buf_1 _21587_ (.A(_04045_),
    .X(_04046_));
 sg13g2_a21oi_1 _21588_ (.A1(_04043_),
    .A2(_04046_),
    .Y(_04047_),
    .B1(_03968_));
 sg13g2_nand2_1 _21589_ (.Y(_04048_),
    .A(_03934_),
    .B(_03937_));
 sg13g2_buf_1 _21590_ (.A(_04048_),
    .X(_04049_));
 sg13g2_buf_1 _21591_ (.A(_04049_),
    .X(_04050_));
 sg13g2_a22oi_1 _21592_ (.Y(_04051_),
    .B1(_03893_),
    .B2(_04050_),
    .A2(net113),
    .A1(net112));
 sg13g2_nand2_1 _21593_ (.Y(_04052_),
    .A(_04047_),
    .B(_04051_));
 sg13g2_buf_1 _21594_ (.A(_04003_),
    .X(_04053_));
 sg13g2_buf_1 _21595_ (.A(_11189_),
    .X(_04054_));
 sg13g2_a22oi_1 _21596_ (.Y(_04055_),
    .B1(_03901_),
    .B2(net223),
    .A2(net134),
    .A1(_03872_));
 sg13g2_nor3_2 _21597_ (.A(net213),
    .B(net278),
    .C(_03878_),
    .Y(_04056_));
 sg13g2_buf_1 _21598_ (.A(_04056_),
    .X(_04057_));
 sg13g2_nand2_1 _21599_ (.Y(_04058_),
    .A(_03910_),
    .B(_04057_));
 sg13g2_nor3_1 _21600_ (.A(net232),
    .B(net278),
    .C(_03868_),
    .Y(_04059_));
 sg13g2_buf_2 _21601_ (.A(_04059_),
    .X(_04060_));
 sg13g2_buf_1 _21602_ (.A(_04060_),
    .X(_04061_));
 sg13g2_a22oi_1 _21603_ (.Y(_04062_),
    .B1(net138),
    .B2(net174),
    .A2(_04061_),
    .A1(_03853_));
 sg13g2_inv_2 _21604_ (.Y(_04063_),
    .A(net179));
 sg13g2_mux2_1 _21605_ (.A0(_10293_),
    .A1(_11027_),
    .S(net201),
    .X(_04064_));
 sg13g2_buf_1 _21606_ (.A(_04064_),
    .X(_04065_));
 sg13g2_nor2_1 _21607_ (.A(net154),
    .B(_03883_),
    .Y(_04066_));
 sg13g2_a21oi_1 _21608_ (.A1(_04063_),
    .A2(net165),
    .Y(_04067_),
    .B1(_04066_));
 sg13g2_nand4_1 _21609_ (.B(_04058_),
    .C(_04062_),
    .A(_04055_),
    .Y(_04068_),
    .D(_04067_));
 sg13g2_buf_1 _21610_ (.A(net137),
    .X(_04069_));
 sg13g2_buf_1 _21611_ (.A(net111),
    .X(_04070_));
 sg13g2_a21oi_1 _21612_ (.A1(net177),
    .A2(_04070_),
    .Y(_04071_),
    .B1(net979));
 sg13g2_o21ai_1 _21613_ (.B1(_04071_),
    .Y(_04072_),
    .A1(_04052_),
    .A2(_04068_));
 sg13g2_nand2b_1 _21614_ (.Y(_04073_),
    .B(_04070_),
    .A_N(net160));
 sg13g2_nand2_1 _21615_ (.Y(_04074_),
    .A(_09831_),
    .B(net237));
 sg13g2_nor3_1 _21616_ (.A(_03918_),
    .B(net202),
    .C(_03842_),
    .Y(_04075_));
 sg13g2_a21oi_1 _21617_ (.A1(net202),
    .A2(net181),
    .Y(_04076_),
    .B1(_04075_));
 sg13g2_a21oi_1 _21618_ (.A1(_08402_),
    .A2(_10790_),
    .Y(_04077_),
    .B1(_10792_));
 sg13g2_nor2_1 _21619_ (.A(_04077_),
    .B(_11790_),
    .Y(_04078_));
 sg13g2_a21oi_1 _21620_ (.A1(_10248_),
    .A2(_04077_),
    .Y(_04079_),
    .B1(_04078_));
 sg13g2_buf_1 _21621_ (.A(_04079_),
    .X(_04080_));
 sg13g2_a221oi_1 _21622_ (.B2(net222),
    .C1(_03954_),
    .B1(net135),
    .A1(_03918_),
    .Y(_04081_),
    .A2(net181));
 sg13g2_o21ai_1 _21623_ (.B1(_04081_),
    .Y(_04082_),
    .A1(net277),
    .A2(_04076_));
 sg13g2_o21ai_1 _21624_ (.B1(_04082_),
    .Y(_04083_),
    .A1(_03887_),
    .A2(_04074_));
 sg13g2_nand2_1 _21625_ (.Y(_04084_),
    .A(_04073_),
    .B(_04083_));
 sg13g2_nand4_1 _21626_ (.B(_04040_),
    .C(_04072_),
    .A(_04038_),
    .Y(_04085_),
    .D(_04084_));
 sg13g2_nor2_1 _21627_ (.A(_04032_),
    .B(_04085_),
    .Y(_04086_));
 sg13g2_nand2b_1 _21628_ (.Y(_04087_),
    .B(_10717_),
    .A_N(net178));
 sg13g2_buf_1 _21629_ (.A(_04087_),
    .X(_04088_));
 sg13g2_nand2_2 _21630_ (.Y(_04089_),
    .A(net280),
    .B(net178));
 sg13g2_nand2_1 _21631_ (.Y(_04090_),
    .A(_04088_),
    .B(_04089_));
 sg13g2_nor2_1 _21632_ (.A(_10658_),
    .B(net175),
    .Y(_04091_));
 sg13g2_buf_2 _21633_ (.A(_04091_),
    .X(_04092_));
 sg13g2_nor2_1 _21634_ (.A(_11252_),
    .B(_11157_),
    .Y(_04093_));
 sg13g2_nand3_1 _21635_ (.B(_11162_),
    .C(_11187_),
    .A(_10566_),
    .Y(_04094_));
 sg13g2_a221oi_1 _21636_ (.B2(_04094_),
    .C1(_03948_),
    .B1(_03938_),
    .A1(_11252_),
    .Y(_04095_),
    .A2(_11157_));
 sg13g2_buf_1 _21637_ (.A(_04095_),
    .X(_04096_));
 sg13g2_nand2b_1 _21638_ (.Y(_04097_),
    .B(net241),
    .A_N(net180));
 sg13g2_nor4_1 _21639_ (.A(_04092_),
    .B(_04093_),
    .C(_04096_),
    .D(_04097_),
    .Y(_04098_));
 sg13g2_nand2_1 _21640_ (.Y(_04099_),
    .A(_11290_),
    .B(_10634_));
 sg13g2_nor4_1 _21641_ (.A(_04092_),
    .B(_04093_),
    .C(_04096_),
    .D(_04099_),
    .Y(_04100_));
 sg13g2_nor3_1 _21642_ (.A(_11451_),
    .B(_04092_),
    .C(_04097_),
    .Y(_04101_));
 sg13g2_and2_1 _21643_ (.A(_10658_),
    .B(net175),
    .X(_04102_));
 sg13g2_buf_1 _21644_ (.A(_04102_),
    .X(_04103_));
 sg13g2_and2_1 _21645_ (.A(_10634_),
    .B(_04103_),
    .X(_04104_));
 sg13g2_nor4_1 _21646_ (.A(_04098_),
    .B(_04100_),
    .C(_04101_),
    .D(_04104_),
    .Y(_04105_));
 sg13g2_nor2_1 _21647_ (.A(net283),
    .B(_04006_),
    .Y(_04106_));
 sg13g2_nor3_1 _21648_ (.A(_03558_),
    .B(_03928_),
    .C(_03930_),
    .Y(_04107_));
 sg13g2_a21oi_1 _21649_ (.A1(_03942_),
    .A2(_04107_),
    .Y(_04108_),
    .B1(_03947_));
 sg13g2_a21oi_1 _21650_ (.A1(net283),
    .A2(_04006_),
    .Y(_04109_),
    .B1(net232));
 sg13g2_a221oi_1 _21651_ (.B2(_04109_),
    .C1(_04003_),
    .B1(_04108_),
    .A1(_11290_),
    .Y(_04110_),
    .A2(_04106_));
 sg13g2_nand2_1 _21652_ (.Y(_04111_),
    .A(_11451_),
    .B(_04096_));
 sg13g2_nor3_1 _21653_ (.A(_11290_),
    .B(net278),
    .C(_11157_),
    .Y(_04112_));
 sg13g2_nor3_1 _21654_ (.A(net179),
    .B(_04092_),
    .C(_04112_),
    .Y(_04113_));
 sg13g2_nand3b_1 _21655_ (.B(_04111_),
    .C(_04113_),
    .Y(_04114_),
    .A_N(_04110_));
 sg13g2_nor2_1 _21656_ (.A(net276),
    .B(_03995_),
    .Y(_04115_));
 sg13g2_a21o_1 _21657_ (.A2(_04115_),
    .A1(_03851_),
    .B1(net242),
    .X(_04116_));
 sg13g2_o21ai_1 _21658_ (.B1(_04116_),
    .Y(_04117_),
    .A1(net139),
    .A2(_04115_));
 sg13g2_o21ai_1 _21659_ (.B1(net155),
    .Y(_04118_),
    .A1(net216),
    .A2(_04103_));
 sg13g2_nand4_1 _21660_ (.B(_04114_),
    .C(_04117_),
    .A(_04105_),
    .Y(_04119_),
    .D(_04118_));
 sg13g2_buf_2 _21661_ (.A(_04119_),
    .X(_04120_));
 sg13g2_nand2_1 _21662_ (.Y(_04121_),
    .A(net276),
    .B(_03995_));
 sg13g2_inv_1 _21663_ (.Y(_04122_),
    .A(_04121_));
 sg13g2_nor2_1 _21664_ (.A(net242),
    .B(net139),
    .Y(_04123_));
 sg13g2_a21oi_2 _21665_ (.B1(_04123_),
    .Y(_04124_),
    .A2(_04122_),
    .A1(_04117_));
 sg13g2_nand2_1 _21666_ (.Y(_04125_),
    .A(_10989_),
    .B(net154));
 sg13g2_nand2_1 _21667_ (.Y(_04126_),
    .A(net228),
    .B(_10989_));
 sg13g2_nor2_1 _21668_ (.A(_11608_),
    .B(net177),
    .Y(_04127_));
 sg13g2_buf_1 _21669_ (.A(_04127_),
    .X(_04128_));
 sg13g2_a221oi_1 _21670_ (.B2(_04126_),
    .C1(_04128_),
    .B1(_04125_),
    .A1(_04120_),
    .Y(_04129_),
    .A2(_04124_));
 sg13g2_buf_2 _21671_ (.A(_04129_),
    .X(_04130_));
 sg13g2_nand2_1 _21672_ (.Y(_04131_),
    .A(_11535_),
    .B(net154));
 sg13g2_a221oi_1 _21673_ (.B2(_11597_),
    .C1(_04128_),
    .B1(_04131_),
    .A1(_04120_),
    .Y(_04132_),
    .A2(_04124_));
 sg13g2_buf_2 _21674_ (.A(_04132_),
    .X(_04133_));
 sg13g2_nand2_1 _21675_ (.Y(_04134_),
    .A(net228),
    .B(net154));
 sg13g2_nor2_1 _21676_ (.A(_04128_),
    .B(_04131_),
    .Y(_04135_));
 sg13g2_nand2_1 _21677_ (.Y(_04136_),
    .A(net192),
    .B(_10989_));
 sg13g2_nor2_1 _21678_ (.A(_04128_),
    .B(_04136_),
    .Y(_04137_));
 sg13g2_a22oi_1 _21679_ (.Y(_04138_),
    .B1(_04137_),
    .B2(net228),
    .A2(_04135_),
    .A1(_10989_));
 sg13g2_o21ai_1 _21680_ (.B1(_04138_),
    .Y(_04139_),
    .A1(_04128_),
    .A2(_04134_));
 sg13g2_buf_1 _21681_ (.A(_04139_),
    .X(_04140_));
 sg13g2_nor2_1 _21682_ (.A(net285),
    .B(net161),
    .Y(_04141_));
 sg13g2_nor4_2 _21683_ (.A(_04130_),
    .B(_04133_),
    .C(_04140_),
    .Y(_04142_),
    .D(_04141_));
 sg13g2_xnor2_1 _21684_ (.Y(_04143_),
    .A(_04090_),
    .B(_04142_));
 sg13g2_nand2_1 _21685_ (.Y(_04144_),
    .A(_08281_),
    .B(_04143_));
 sg13g2_or2_1 _21686_ (.X(_04145_),
    .B(net175),
    .A(_03625_));
 sg13g2_buf_1 _21687_ (.A(_04145_),
    .X(_04146_));
 sg13g2_nor2_1 _21688_ (.A(net232),
    .B(_04003_),
    .Y(_04147_));
 sg13g2_o21ai_1 _21689_ (.B1(_04015_),
    .Y(_04148_),
    .A1(_04147_),
    .A2(_04013_));
 sg13g2_nand2_1 _21690_ (.Y(_04149_),
    .A(net229),
    .B(net139));
 sg13g2_buf_1 _21691_ (.A(_04149_),
    .X(_04150_));
 sg13g2_nand3_1 _21692_ (.B(_04018_),
    .C(_04150_),
    .A(_03995_),
    .Y(_04151_));
 sg13g2_nand3_1 _21693_ (.B(_04018_),
    .C(_04150_),
    .A(net286),
    .Y(_04152_));
 sg13g2_a22oi_1 _21694_ (.Y(_04153_),
    .B1(_04151_),
    .B2(_04152_),
    .A2(_04148_),
    .A1(_04146_));
 sg13g2_nor2_1 _21695_ (.A(net230),
    .B(_03865_),
    .Y(_04154_));
 sg13g2_a221oi_1 _21696_ (.B2(net229),
    .C1(_03998_),
    .B1(net139),
    .A1(net230),
    .Y(_04155_),
    .A2(_03865_));
 sg13g2_a21o_1 _21697_ (.A2(_04150_),
    .A1(_04154_),
    .B1(_04155_),
    .X(_04156_));
 sg13g2_nor2_1 _21698_ (.A(_11522_),
    .B(net139),
    .Y(_04157_));
 sg13g2_nor3_2 _21699_ (.A(_04153_),
    .B(_04156_),
    .C(_04157_),
    .Y(_04158_));
 sg13g2_or2_1 _21700_ (.X(_04159_),
    .B(net177),
    .A(net285));
 sg13g2_buf_1 _21701_ (.A(_04159_),
    .X(_04160_));
 sg13g2_nand2_1 _21702_ (.Y(_04161_),
    .A(net154),
    .B(_04160_));
 sg13g2_nand2_1 _21703_ (.Y(_04162_),
    .A(_11562_),
    .B(_04160_));
 sg13g2_a21oi_1 _21704_ (.A1(_03999_),
    .A2(_04000_),
    .Y(_04163_),
    .B1(_04013_));
 sg13g2_nand3_1 _21705_ (.B(_03995_),
    .C(_04150_),
    .A(_10989_),
    .Y(_04164_));
 sg13g2_nor3_1 _21706_ (.A(_04163_),
    .B(_04020_),
    .C(_04164_),
    .Y(_04165_));
 sg13g2_nand3_1 _21707_ (.B(_10989_),
    .C(_04150_),
    .A(net286),
    .Y(_04166_));
 sg13g2_nor3_1 _21708_ (.A(_04163_),
    .B(_04020_),
    .C(_04166_),
    .Y(_04167_));
 sg13g2_nand2_1 _21709_ (.Y(_04168_),
    .A(net176),
    .B(_04157_));
 sg13g2_o21ai_1 _21710_ (.B1(_04168_),
    .Y(_04169_),
    .A1(net230),
    .A2(_04164_));
 sg13g2_nor4_1 _21711_ (.A(net191),
    .B(_04165_),
    .C(_04167_),
    .D(_04169_),
    .Y(_04170_));
 sg13g2_a221oi_1 _21712_ (.B2(_04162_),
    .C1(_04170_),
    .B1(_04161_),
    .A1(net136),
    .Y(_04171_),
    .A2(_04158_));
 sg13g2_nand2_1 _21713_ (.Y(_04172_),
    .A(_10390_),
    .B(net177));
 sg13g2_nand2_1 _21714_ (.Y(_04173_),
    .A(net243),
    .B(net154));
 sg13g2_nor2_1 _21715_ (.A(_10390_),
    .B(net177),
    .Y(_04174_));
 sg13g2_a21oi_1 _21716_ (.A1(_04172_),
    .A2(_04173_),
    .Y(_04175_),
    .B1(_04174_));
 sg13g2_nor2_1 _21717_ (.A(_04171_),
    .B(_04175_),
    .Y(_04176_));
 sg13g2_xnor2_1 _21718_ (.Y(_04177_),
    .A(_04090_),
    .B(_04176_));
 sg13g2_nor2_1 _21719_ (.A(net157),
    .B(_03959_),
    .Y(_04178_));
 sg13g2_a22oi_1 _21720_ (.Y(_04179_),
    .B1(_04177_),
    .B2(_04178_),
    .A2(_04144_),
    .A1(_04086_));
 sg13g2_o21ai_1 _21721_ (.B1(_04179_),
    .Y(_04180_),
    .A1(net166),
    .A2(\cpu.ex.c_mult[11] ));
 sg13g2_nand2_2 _21722_ (.Y(_04181_),
    .A(net1062),
    .B(net716));
 sg13g2_nor2_2 _21723_ (.A(_08444_),
    .B(_04181_),
    .Y(_04182_));
 sg13g2_nand4_1 _21724_ (.B(_08624_),
    .C(_08633_),
    .A(_08667_),
    .Y(_04183_),
    .D(_04182_));
 sg13g2_nor2_1 _21725_ (.A(_08615_),
    .B(_04183_),
    .Y(_04184_));
 sg13g2_nand3_1 _21726_ (.B(_08652_),
    .C(_04184_),
    .A(_08680_),
    .Y(_04185_));
 sg13g2_xnor2_1 _21727_ (.Y(_04186_),
    .A(_11031_),
    .B(_04185_));
 sg13g2_buf_1 _21728_ (.A(_03979_),
    .X(_04187_));
 sg13g2_a22oi_1 _21729_ (.Y(_04188_),
    .B1(_04186_),
    .B2(_04187_),
    .A2(_03992_),
    .A1(\cpu.ex.pc[11] ));
 sg13g2_o21ai_1 _21730_ (.B1(_04188_),
    .Y(_00976_),
    .A1(net84),
    .A2(_04180_));
 sg13g2_buf_1 _21731_ (.A(net157),
    .X(_04189_));
 sg13g2_nand3_1 _21732_ (.B(_03956_),
    .C(_03957_),
    .A(_03954_),
    .Y(_04190_));
 sg13g2_buf_1 _21733_ (.A(_04190_),
    .X(_04191_));
 sg13g2_nor3_1 _21734_ (.A(_09069_),
    .B(_09078_),
    .C(_04191_),
    .Y(_04192_));
 sg13g2_buf_2 _21735_ (.A(_04192_),
    .X(_04193_));
 sg13g2_nand2b_1 _21736_ (.Y(_04194_),
    .B(net194),
    .A_N(net193));
 sg13g2_buf_1 _21737_ (.A(_04194_),
    .X(_04195_));
 sg13g2_nand2_1 _21738_ (.Y(_04196_),
    .A(_11300_),
    .B(net193));
 sg13g2_and2_1 _21739_ (.A(_04195_),
    .B(_04196_),
    .X(_04197_));
 sg13g2_buf_1 _21740_ (.A(_04197_),
    .X(_04198_));
 sg13g2_nor2_1 _21741_ (.A(net191),
    .B(_03902_),
    .Y(_04199_));
 sg13g2_o21ai_1 _21742_ (.B1(_04037_),
    .Y(_04200_),
    .A1(net192),
    .A2(net136));
 sg13g2_nor2_1 _21743_ (.A(_04175_),
    .B(_04200_),
    .Y(_04201_));
 sg13g2_o21ai_1 _21744_ (.B1(_04201_),
    .Y(_04202_),
    .A1(_04158_),
    .A2(_04199_));
 sg13g2_nand2_2 _21745_ (.Y(_04203_),
    .A(_10729_),
    .B(net215));
 sg13g2_nand2_1 _21746_ (.Y(_04204_),
    .A(_04203_),
    .B(_04160_));
 sg13g2_and2_1 _21747_ (.A(_04172_),
    .B(_04204_),
    .X(_04205_));
 sg13g2_o21ai_1 _21748_ (.B1(_04037_),
    .Y(_04206_),
    .A1(_04034_),
    .A2(_04205_));
 sg13g2_nand2_1 _21749_ (.Y(_04207_),
    .A(_04202_),
    .B(_04206_));
 sg13g2_xor2_1 _21750_ (.B(_04207_),
    .A(_04198_),
    .X(_04208_));
 sg13g2_a22oi_1 _21751_ (.Y(_04209_),
    .B1(_03901_),
    .B2(net200),
    .A2(_03862_),
    .A1(net114));
 sg13g2_a22oi_1 _21752_ (.Y(_04210_),
    .B1(net162),
    .B2(net174),
    .A2(net165),
    .A1(net112));
 sg13g2_nor2_1 _21753_ (.A(_03918_),
    .B(_03854_),
    .Y(_04211_));
 sg13g2_buf_1 _21754_ (.A(_04211_),
    .X(_04212_));
 sg13g2_buf_1 _21755_ (.A(_04212_),
    .X(_04213_));
 sg13g2_nor2_2 _21756_ (.A(_03868_),
    .B(_03847_),
    .Y(_04214_));
 sg13g2_a22oi_1 _21757_ (.Y(_04215_),
    .B1(_04214_),
    .B2(net223),
    .A2(net131),
    .A1(net161));
 sg13g2_a21oi_1 _21758_ (.A1(net215),
    .A2(_04045_),
    .Y(_04216_),
    .B1(_03967_));
 sg13g2_and4_1 _21759_ (.A(_04209_),
    .B(_04210_),
    .C(_04215_),
    .D(_04216_),
    .X(_04217_));
 sg13g2_a22oi_1 _21760_ (.Y(_04218_),
    .B1(net134),
    .B2(net138),
    .A2(net164),
    .A1(net159));
 sg13g2_a22oi_1 _21761_ (.Y(_04219_),
    .B1(net156),
    .B2(net155),
    .A2(net133),
    .A1(net136));
 sg13g2_and2_1 _21762_ (.A(_04218_),
    .B(_04219_),
    .X(_04220_));
 sg13g2_o21ai_1 _21763_ (.B1(_09850_),
    .Y(_04221_),
    .A1(net163),
    .A2(net158));
 sg13g2_a21oi_1 _21764_ (.A1(_04217_),
    .A2(_04220_),
    .Y(_04222_),
    .B1(_04221_));
 sg13g2_mux2_1 _21765_ (.A0(_04089_),
    .A1(_04088_),
    .S(_04198_),
    .X(_04223_));
 sg13g2_buf_1 _21766_ (.A(_03914_),
    .X(_04224_));
 sg13g2_nand2_1 _21767_ (.Y(_04225_),
    .A(_10549_),
    .B(_11421_));
 sg13g2_a22oi_1 _21768_ (.Y(_04226_),
    .B1(_04225_),
    .B2(net1130),
    .A2(net359),
    .A1(_10549_));
 sg13g2_o21ai_1 _21769_ (.B1(_03859_),
    .Y(_04227_),
    .A1(net222),
    .A2(_03854_));
 sg13g2_nand2_1 _21770_ (.Y(_04228_),
    .A(_10549_),
    .B(_04227_));
 sg13g2_o21ai_1 _21771_ (.B1(_04228_),
    .Y(_04229_),
    .A1(net130),
    .A2(_04226_));
 sg13g2_a21oi_1 _21772_ (.A1(_10961_),
    .A2(net111),
    .Y(_04230_),
    .B1(_03954_));
 sg13g2_nand2_1 _21773_ (.Y(_04231_),
    .A(_04229_),
    .B(_04230_));
 sg13g2_o21ai_1 _21774_ (.B1(_04231_),
    .Y(_04232_),
    .A1(_03943_),
    .A2(_04223_));
 sg13g2_inv_1 _21775_ (.Y(_04233_),
    .A(_09048_));
 sg13g2_nand2_1 _21776_ (.Y(_04234_),
    .A(net194),
    .B(net193));
 sg13g2_mux2_1 _21777_ (.A0(net1048),
    .A1(net1060),
    .S(_04234_),
    .X(_04235_));
 sg13g2_or2_1 _21778_ (.X(_04236_),
    .B(net193),
    .A(_10690_));
 sg13g2_buf_1 _21779_ (.A(_04236_),
    .X(_04237_));
 sg13g2_o21ai_1 _21780_ (.B1(_04237_),
    .Y(_04238_),
    .A1(net978),
    .A2(_04235_));
 sg13g2_o21ai_1 _21781_ (.B1(_04238_),
    .Y(_04239_),
    .A1(_04233_),
    .A2(_10659_));
 sg13g2_nor4_1 _21782_ (.A(_04032_),
    .B(_04222_),
    .C(_04232_),
    .D(_04239_),
    .Y(_04240_));
 sg13g2_nand3_1 _21783_ (.B(_04089_),
    .C(_04198_),
    .A(net1077),
    .Y(_04241_));
 sg13g2_nand3b_1 _21784_ (.B(net1077),
    .C(_04088_),
    .Y(_04242_),
    .A_N(_04198_));
 sg13g2_mux2_1 _21785_ (.A0(_04241_),
    .A1(_04242_),
    .S(_04142_),
    .X(_04243_));
 sg13g2_a221oi_1 _21786_ (.B2(_04243_),
    .C1(net132),
    .B1(_04240_),
    .A1(_04193_),
    .Y(_04244_),
    .A2(_04208_));
 sg13g2_a21oi_1 _21787_ (.A1(_04189_),
    .A2(\cpu.ex.c_mult[12] ),
    .Y(_04245_),
    .B1(_04244_));
 sg13g2_nor2_2 _21788_ (.A(_08643_),
    .B(_04185_),
    .Y(_04246_));
 sg13g2_xnor2_1 _21789_ (.Y(_04247_),
    .A(_10661_),
    .B(_04246_));
 sg13g2_a22oi_1 _21790_ (.Y(_04248_),
    .B1(_04247_),
    .B2(net83),
    .A2(net35),
    .A1(net727));
 sg13g2_o21ai_1 _21791_ (.B1(_04248_),
    .Y(_00977_),
    .A1(net84),
    .A2(_04245_));
 sg13g2_inv_1 _21792_ (.Y(_04249_),
    .A(_04141_));
 sg13g2_nand3_1 _21793_ (.B(_04249_),
    .C(_04195_),
    .A(net178),
    .Y(_04250_));
 sg13g2_nor4_2 _21794_ (.A(_04130_),
    .B(_04133_),
    .C(_04140_),
    .Y(_04251_),
    .D(_04250_));
 sg13g2_nand3_1 _21795_ (.B(_04249_),
    .C(_04195_),
    .A(_10761_),
    .Y(_04252_));
 sg13g2_nor4_2 _21796_ (.A(_04130_),
    .B(_04133_),
    .C(_04140_),
    .Y(_04253_),
    .D(_04252_));
 sg13g2_inv_1 _21797_ (.Y(_04254_),
    .A(_04195_));
 sg13g2_o21ai_1 _21798_ (.B1(_04196_),
    .Y(_04255_),
    .A1(_04089_),
    .A2(_04254_));
 sg13g2_nor3_2 _21799_ (.A(_04251_),
    .B(_04253_),
    .C(_04255_),
    .Y(_04256_));
 sg13g2_nor2_1 _21800_ (.A(net217),
    .B(net115),
    .Y(_04257_));
 sg13g2_nor2_1 _21801_ (.A(net211),
    .B(_10961_),
    .Y(_04258_));
 sg13g2_nor2_1 _21802_ (.A(_04257_),
    .B(_04258_),
    .Y(_04259_));
 sg13g2_xor2_1 _21803_ (.B(_04259_),
    .A(_04256_),
    .X(_04260_));
 sg13g2_nor2_1 _21804_ (.A(net130),
    .B(_03883_),
    .Y(_04261_));
 sg13g2_nor2_1 _21805_ (.A(net222),
    .B(net158),
    .Y(_04262_));
 sg13g2_o21ai_1 _21806_ (.B1(_09831_),
    .Y(_04263_),
    .A1(_04261_),
    .A2(_04262_));
 sg13g2_nand2_1 _21807_ (.Y(_04264_),
    .A(net222),
    .B(net93));
 sg13g2_a21oi_1 _21808_ (.A1(net130),
    .A2(net158),
    .Y(_04265_),
    .B1(_03912_));
 sg13g2_a22oi_1 _21809_ (.Y(_04266_),
    .B1(_04264_),
    .B2(_04265_),
    .A2(_11499_),
    .A1(net1061));
 sg13g2_nand2_1 _21810_ (.Y(_04267_),
    .A(net211),
    .B(net115));
 sg13g2_mux2_1 _21811_ (.A0(_09848_),
    .A1(_09074_),
    .S(_04267_),
    .X(_04268_));
 sg13g2_nand2_1 _21812_ (.Y(_04269_),
    .A(net217),
    .B(_10961_));
 sg13g2_o21ai_1 _21813_ (.B1(_04269_),
    .Y(_04270_),
    .A1(net978),
    .A2(_04268_));
 sg13g2_nand2_1 _21814_ (.Y(_04271_),
    .A(_10549_),
    .B(_03903_));
 sg13g2_o21ai_1 _21815_ (.B1(net158),
    .Y(_04272_),
    .A1(net177),
    .A2(_04271_));
 sg13g2_a221oi_1 _21816_ (.B2(_04214_),
    .C1(_04272_),
    .B1(net200),
    .A1(_03866_),
    .Y(_04273_),
    .A2(net156));
 sg13g2_a22oi_1 _21817_ (.Y(_04274_),
    .B1(net138),
    .B2(_03910_),
    .A2(_03873_),
    .A1(net223));
 sg13g2_nand3_1 _21818_ (.B(net283),
    .C(_03922_),
    .A(_11290_),
    .Y(_04275_));
 sg13g2_buf_1 _21819_ (.A(_04275_),
    .X(_04276_));
 sg13g2_nand2_1 _21820_ (.Y(_04277_),
    .A(net215),
    .B(_04060_));
 sg13g2_o21ai_1 _21821_ (.B1(_04277_),
    .Y(_04278_),
    .A1(net176),
    .A2(_04276_));
 sg13g2_a221oi_1 _21822_ (.B2(net163),
    .C1(_04278_),
    .B1(net131),
    .A1(_03853_),
    .Y(_04279_),
    .A2(net165));
 sg13g2_mux2_1 _21823_ (.A0(net155),
    .A1(net134),
    .S(net234),
    .X(_04280_));
 sg13g2_a22oi_1 _21824_ (.Y(_04281_),
    .B1(_04280_),
    .B2(net272),
    .A2(_03903_),
    .A1(net174));
 sg13g2_or2_1 _21825_ (.X(_04282_),
    .B(_04281_),
    .A(_03870_));
 sg13g2_nand4_1 _21826_ (.B(_04274_),
    .C(_04279_),
    .A(_04273_),
    .Y(_04283_),
    .D(_04282_));
 sg13g2_nand3_1 _21827_ (.B(_04073_),
    .C(_04283_),
    .A(_09850_),
    .Y(_04284_));
 sg13g2_nand4_1 _21828_ (.B(_04266_),
    .C(_04270_),
    .A(_04263_),
    .Y(_04285_),
    .D(_04284_));
 sg13g2_nor2_1 _21829_ (.A(_04032_),
    .B(_04285_),
    .Y(_04286_));
 sg13g2_o21ai_1 _21830_ (.B1(_04286_),
    .Y(_04287_),
    .A1(_03943_),
    .A2(_04260_));
 sg13g2_nand2_1 _21831_ (.Y(_04288_),
    .A(_03865_),
    .B(net139));
 sg13g2_nand2_1 _21832_ (.Y(_04289_),
    .A(_11497_),
    .B(net139));
 sg13g2_a22oi_1 _21833_ (.Y(_04290_),
    .B1(_04288_),
    .B2(_04289_),
    .A2(_04021_),
    .A1(_04014_));
 sg13g2_o21ai_1 _21834_ (.B1(_10483_),
    .Y(_04291_),
    .A1(_10364_),
    .A2(_04288_));
 sg13g2_or2_1 _21835_ (.X(_04292_),
    .B(_04291_),
    .A(_04290_));
 sg13g2_nor2_1 _21836_ (.A(_03865_),
    .B(_03852_),
    .Y(_04293_));
 sg13g2_nand2_1 _21837_ (.Y(_04294_),
    .A(_04018_),
    .B(_04293_));
 sg13g2_nor2_1 _21838_ (.A(_11497_),
    .B(_03852_),
    .Y(_04295_));
 sg13g2_nand2_1 _21839_ (.Y(_04296_),
    .A(_04018_),
    .B(_04295_));
 sg13g2_a22oi_1 _21840_ (.Y(_04297_),
    .B1(_04294_),
    .B2(_04296_),
    .A2(_04148_),
    .A1(_04146_));
 sg13g2_inv_1 _21841_ (.Y(_04298_),
    .A(_04293_));
 sg13g2_o21ai_1 _21842_ (.B1(_04016_),
    .Y(_04299_),
    .A1(_04293_),
    .A2(_04295_));
 sg13g2_o21ai_1 _21843_ (.B1(_04299_),
    .Y(_04300_),
    .A1(_11514_),
    .A2(_04298_));
 sg13g2_nand2_1 _21844_ (.Y(_04301_),
    .A(_04201_),
    .B(_04237_));
 sg13g2_nor3_1 _21845_ (.A(_04297_),
    .B(_04300_),
    .C(_04301_),
    .Y(_04302_));
 sg13g2_nand2_1 _21846_ (.Y(_04303_),
    .A(_04206_),
    .B(_04234_));
 sg13g2_and3_1 _21847_ (.X(_04304_),
    .A(_04199_),
    .B(_04201_),
    .C(_04237_));
 sg13g2_a221oi_1 _21848_ (.B2(_04237_),
    .C1(_04304_),
    .B1(_04303_),
    .A1(_04292_),
    .Y(_04305_),
    .A2(_04302_));
 sg13g2_xnor2_1 _21849_ (.Y(_04306_),
    .A(_04259_),
    .B(_04305_));
 sg13g2_a21oi_1 _21850_ (.A1(_04193_),
    .A2(_04306_),
    .Y(_04307_),
    .B1(_04189_));
 sg13g2_nor2_1 _21851_ (.A(net166),
    .B(_11679_),
    .Y(_04308_));
 sg13g2_a22oi_1 _21852_ (.Y(_04309_),
    .B1(_04308_),
    .B2(_11706_),
    .A2(_04307_),
    .A1(_04287_));
 sg13g2_nand2_1 _21853_ (.Y(_04310_),
    .A(net727),
    .B(_04246_));
 sg13g2_xor2_1 _21854_ (.B(_04310_),
    .A(_10392_),
    .X(_04311_));
 sg13g2_a22oi_1 _21855_ (.Y(_04312_),
    .B1(_04311_),
    .B2(net83),
    .A2(net35),
    .A1(net822));
 sg13g2_o21ai_1 _21856_ (.B1(_04312_),
    .Y(_00978_),
    .A1(net84),
    .A2(_04309_));
 sg13g2_xnor2_1 _21857_ (.Y(_04313_),
    .A(_10292_),
    .B(net222));
 sg13g2_nor2_1 _21858_ (.A(net211),
    .B(net115),
    .Y(_04314_));
 sg13g2_o21ai_1 _21859_ (.B1(_04267_),
    .Y(_04315_),
    .A1(_04314_),
    .A2(_04305_));
 sg13g2_xor2_1 _21860_ (.B(_04315_),
    .A(_04313_),
    .X(_04316_));
 sg13g2_nor2b_1 _21861_ (.A(_04257_),
    .B_N(_04313_),
    .Y(_04317_));
 sg13g2_nor2_1 _21862_ (.A(_04258_),
    .B(_04313_),
    .Y(_04318_));
 sg13g2_mux2_1 _21863_ (.A0(_04317_),
    .A1(_04318_),
    .S(_04256_),
    .X(_04319_));
 sg13g2_and2_1 _21864_ (.A(_11389_),
    .B(_04031_),
    .X(_04320_));
 sg13g2_buf_1 _21865_ (.A(_04320_),
    .X(_04321_));
 sg13g2_o21ai_1 _21866_ (.B1(net1060),
    .Y(_04322_),
    .A1(net141),
    .A2(_04080_));
 sg13g2_nor2_1 _21867_ (.A(_11709_),
    .B(net222),
    .Y(_04323_));
 sg13g2_nand2_1 _21868_ (.Y(_04324_),
    .A(net1048),
    .B(_04323_));
 sg13g2_nand3_1 _21869_ (.B(_04322_),
    .C(_04324_),
    .A(_09835_),
    .Y(_04325_));
 sg13g2_nand2_1 _21870_ (.Y(_04326_),
    .A(_11709_),
    .B(net222));
 sg13g2_mux2_1 _21871_ (.A0(_04257_),
    .A1(_04258_),
    .S(_04313_),
    .X(_04327_));
 sg13g2_nand2_1 _21872_ (.Y(_04328_),
    .A(net1061),
    .B(_11514_));
 sg13g2_o21ai_1 _21873_ (.B1(_04328_),
    .Y(_04329_),
    .A1(net158),
    .A2(_04074_));
 sg13g2_a221oi_1 _21874_ (.B2(net1077),
    .C1(_04329_),
    .B1(_04327_),
    .A1(_04325_),
    .Y(_04330_),
    .A2(_04326_));
 sg13g2_nand2_1 _21875_ (.Y(_04331_),
    .A(net213),
    .B(_11189_));
 sg13g2_o21ai_1 _21876_ (.B1(_04331_),
    .Y(_04332_),
    .A1(net213),
    .A2(net176));
 sg13g2_nand3_1 _21877_ (.B(_03882_),
    .C(_04332_),
    .A(net233),
    .Y(_04333_));
 sg13g2_a22oi_1 _21878_ (.Y(_04334_),
    .B1(net200),
    .B2(_03873_),
    .A2(net162),
    .A1(net159));
 sg13g2_a22oi_1 _21879_ (.Y(_04335_),
    .B1(net134),
    .B2(_03901_),
    .A2(net164),
    .A1(net112));
 sg13g2_nand3_1 _21880_ (.B(_04334_),
    .C(_04335_),
    .A(_04333_),
    .Y(_04336_));
 sg13g2_a21oi_1 _21881_ (.A1(net163),
    .A2(net135),
    .Y(_04337_),
    .B1(net111));
 sg13g2_nor2_1 _21882_ (.A(net154),
    .B(_04276_),
    .Y(_04338_));
 sg13g2_a21oi_1 _21883_ (.A1(net160),
    .A2(net131),
    .Y(_04339_),
    .B1(_04338_));
 sg13g2_nor2_1 _21884_ (.A(_04025_),
    .B(_03905_),
    .Y(_04340_));
 sg13g2_a21oi_1 _21885_ (.A1(net174),
    .A2(_04214_),
    .Y(_04341_),
    .B1(_04340_));
 sg13g2_nor2_1 _21886_ (.A(net177),
    .B(_03887_),
    .Y(_04342_));
 sg13g2_a21oi_1 _21887_ (.A1(net155),
    .A2(net138),
    .Y(_04343_),
    .B1(_04342_));
 sg13g2_nand4_1 _21888_ (.B(_04339_),
    .C(_04341_),
    .A(_04337_),
    .Y(_04344_),
    .D(_04343_));
 sg13g2_a21oi_1 _21889_ (.A1(_10961_),
    .A2(net93),
    .Y(_04345_),
    .B1(_03969_));
 sg13g2_o21ai_1 _21890_ (.B1(_04345_),
    .Y(_04346_),
    .A1(_04336_),
    .A2(_04344_));
 sg13g2_nand4_1 _21891_ (.B(_04321_),
    .C(_04330_),
    .A(net181),
    .Y(_04347_),
    .D(_04346_));
 sg13g2_a221oi_1 _21892_ (.B2(net935),
    .C1(_04347_),
    .B1(_04319_),
    .A1(_04193_),
    .Y(_04348_),
    .A2(_04316_));
 sg13g2_inv_1 _21893_ (.Y(_04349_),
    .A(_11743_));
 sg13g2_nor3_1 _21894_ (.A(net166),
    .B(_11742_),
    .C(_04349_),
    .Y(_04350_));
 sg13g2_nor3_1 _21895_ (.A(_03836_),
    .B(_04348_),
    .C(_04350_),
    .Y(_04351_));
 sg13g2_nand3_1 _21896_ (.B(net822),
    .C(_04246_),
    .A(net727),
    .Y(_04352_));
 sg13g2_xnor2_1 _21897_ (.Y(_04353_),
    .A(_00177_),
    .B(_04352_));
 sg13g2_inv_1 _21898_ (.Y(_04354_),
    .A(_04353_));
 sg13g2_a22oi_1 _21899_ (.Y(_04355_),
    .B1(_04354_),
    .B2(net83),
    .A2(net35),
    .A1(net820));
 sg13g2_nand2b_1 _21900_ (.Y(_00979_),
    .B(_04355_),
    .A_N(_04351_));
 sg13g2_xnor2_1 _21901_ (.Y(_04356_),
    .A(net210),
    .B(net130));
 sg13g2_nor2_1 _21902_ (.A(_03959_),
    .B(_04356_),
    .Y(_04357_));
 sg13g2_and2_1 _21903_ (.A(_04193_),
    .B(_04356_),
    .X(_04358_));
 sg13g2_a21oi_1 _21904_ (.A1(_04315_),
    .A2(_04326_),
    .Y(_04359_),
    .B1(_04323_));
 sg13g2_mux2_1 _21905_ (.A0(_04357_),
    .A1(_04358_),
    .S(_04359_),
    .X(_04360_));
 sg13g2_a22oi_1 _21906_ (.Y(_04361_),
    .B1(_03901_),
    .B2(net159),
    .A2(net164),
    .A1(net114));
 sg13g2_a22oi_1 _21907_ (.Y(_04362_),
    .B1(net133),
    .B2(net163),
    .A2(_04213_),
    .A1(net115));
 sg13g2_nand2_1 _21908_ (.Y(_04363_),
    .A(net234),
    .B(_11189_));
 sg13g2_nand2_1 _21909_ (.Y(_04364_),
    .A(net202),
    .B(net134));
 sg13g2_nor2_1 _21910_ (.A(net359),
    .B(_03964_),
    .Y(_04365_));
 sg13g2_a221oi_1 _21911_ (.B2(_04365_),
    .C1(net183),
    .B1(_04364_),
    .A1(net359),
    .Y(_04366_),
    .A2(_04363_));
 sg13g2_a22oi_1 _21912_ (.Y(_04367_),
    .B1(net113),
    .B2(net161),
    .A2(net182),
    .A1(net215));
 sg13g2_a22oi_1 _21913_ (.Y(_04368_),
    .B1(_03894_),
    .B2(net112),
    .A2(net162),
    .A1(net155));
 sg13g2_a21oi_1 _21914_ (.A1(net193),
    .A2(_04045_),
    .Y(_04369_),
    .B1(_03967_));
 sg13g2_a21oi_1 _21915_ (.A1(_11157_),
    .A2(_03873_),
    .Y(_04370_),
    .B1(_03906_));
 sg13g2_nand4_1 _21916_ (.B(_04368_),
    .C(_04369_),
    .A(_04367_),
    .Y(_04371_),
    .D(_04370_));
 sg13g2_nor2_1 _21917_ (.A(_04366_),
    .B(_04371_),
    .Y(_04372_));
 sg13g2_nand3_1 _21918_ (.B(_04362_),
    .C(_04372_),
    .A(_04361_),
    .Y(_04373_));
 sg13g2_nand3_1 _21919_ (.B(_04264_),
    .C(_04373_),
    .A(_09850_),
    .Y(_04374_));
 sg13g2_nor2_1 _21920_ (.A(_11707_),
    .B(_04080_),
    .Y(_04375_));
 sg13g2_and2_1 _21921_ (.A(net1077),
    .B(_04356_),
    .X(_04376_));
 sg13g2_o21ai_1 _21922_ (.B1(_09073_),
    .Y(_04377_),
    .A1(net235),
    .A2(_04224_));
 sg13g2_nand3_1 _21923_ (.B(_11763_),
    .C(net237),
    .A(_09847_),
    .Y(_04378_));
 sg13g2_and3_1 _21924_ (.X(_04379_),
    .A(_09835_),
    .B(_04377_),
    .C(_04378_));
 sg13g2_a21oi_1 _21925_ (.A1(_11359_),
    .A2(_04224_),
    .Y(_04380_),
    .B1(_04379_));
 sg13g2_a221oi_1 _21926_ (.B2(_04376_),
    .C1(_04380_),
    .B1(_04375_),
    .A1(net1061),
    .Y(_04381_),
    .A2(_11522_));
 sg13g2_and4_1 _21927_ (.A(_03877_),
    .B(_04321_),
    .C(_04374_),
    .D(_04381_),
    .X(_04382_));
 sg13g2_nand2_1 _21928_ (.Y(_04383_),
    .A(net935),
    .B(_04356_));
 sg13g2_nand2_1 _21929_ (.Y(_04384_),
    .A(net168),
    .B(_04079_));
 sg13g2_o21ai_1 _21930_ (.B1(_10961_),
    .Y(_04385_),
    .A1(_11695_),
    .A2(_04196_));
 sg13g2_nand4_1 _21931_ (.B(_04088_),
    .C(_04195_),
    .A(_10426_),
    .Y(_04386_),
    .D(_04384_));
 sg13g2_nor2_1 _21932_ (.A(_04141_),
    .B(_04386_),
    .Y(_04387_));
 sg13g2_nor3_1 _21933_ (.A(_04130_),
    .B(_04133_),
    .C(_04140_),
    .Y(_04388_));
 sg13g2_nor2_1 _21934_ (.A(_04089_),
    .B(_04386_),
    .Y(_04389_));
 sg13g2_a221oi_1 _21935_ (.B2(_04388_),
    .C1(_04389_),
    .B1(_04387_),
    .A1(_04384_),
    .Y(_04390_),
    .A2(_04385_));
 sg13g2_nor4_1 _21936_ (.A(_10426_),
    .B(_04251_),
    .C(_04253_),
    .D(_04255_),
    .Y(_04391_));
 sg13g2_or3_1 _21937_ (.A(_04383_),
    .B(_04390_),
    .C(_04391_),
    .X(_04392_));
 sg13g2_nor3_1 _21938_ (.A(_03943_),
    .B(_04375_),
    .C(_04356_),
    .Y(_04393_));
 sg13g2_o21ai_1 _21939_ (.B1(_04393_),
    .Y(_04394_),
    .A1(_04390_),
    .A2(_04391_));
 sg13g2_nand3_1 _21940_ (.B(_04392_),
    .C(_04394_),
    .A(_04382_),
    .Y(_04395_));
 sg13g2_nand2_1 _21941_ (.Y(_04396_),
    .A(net132),
    .B(_11774_));
 sg13g2_o21ai_1 _21942_ (.B1(_04396_),
    .Y(_04397_),
    .A1(_04360_),
    .A2(_04395_));
 sg13g2_nand4_1 _21943_ (.B(net822),
    .C(net820),
    .A(net727),
    .Y(_04398_),
    .D(_04246_));
 sg13g2_xnor2_1 _21944_ (.Y(_04399_),
    .A(_10915_),
    .B(_04398_));
 sg13g2_a22oi_1 _21945_ (.Y(_04400_),
    .B1(_04399_),
    .B2(net83),
    .A2(net35),
    .A1(_08363_));
 sg13g2_o21ai_1 _21946_ (.B1(_04400_),
    .Y(_00980_),
    .A1(_03837_),
    .A2(_04397_));
 sg13g2_buf_1 _21947_ (.A(_11159_),
    .X(_04401_));
 sg13g2_nand4_1 _21948_ (.B(_09087_),
    .C(net391),
    .A(_08399_),
    .Y(_04402_),
    .D(_09265_));
 sg13g2_a21oi_1 _21949_ (.A1(_08868_),
    .A2(net94),
    .Y(_04403_),
    .B1(_03991_));
 sg13g2_nand2b_1 _21950_ (.Y(_04404_),
    .B(net724),
    .A_N(_04403_));
 sg13g2_nand3_1 _21951_ (.B(net803),
    .C(net94),
    .A(net717),
    .Y(_04405_));
 sg13g2_nor2_1 _21952_ (.A(net278),
    .B(net277),
    .Y(_04406_));
 sg13g2_a21oi_1 _21953_ (.A1(net272),
    .A2(net181),
    .Y(_04407_),
    .B1(net233));
 sg13g2_a21oi_1 _21954_ (.A1(_03866_),
    .A2(_04406_),
    .Y(_04408_),
    .B1(_04407_));
 sg13g2_nor3_1 _21955_ (.A(_11452_),
    .B(net234),
    .C(_04408_),
    .Y(_04409_));
 sg13g2_nor2_1 _21956_ (.A(net202),
    .B(net181),
    .Y(_04410_));
 sg13g2_nand2_1 _21957_ (.Y(_04411_),
    .A(_10567_),
    .B(_03914_));
 sg13g2_o21ai_1 _21958_ (.B1(_04411_),
    .Y(_04412_),
    .A1(net359),
    .A2(net238));
 sg13g2_nor2_1 _21959_ (.A(net234),
    .B(_04412_),
    .Y(_04413_));
 sg13g2_nor2_1 _21960_ (.A(_04410_),
    .B(_04413_),
    .Y(_04414_));
 sg13g2_nand2_1 _21961_ (.Y(_04415_),
    .A(net115),
    .B(_03901_));
 sg13g2_a22oi_1 _21962_ (.Y(_04416_),
    .B1(net156),
    .B2(net215),
    .A2(net138),
    .A1(_03891_));
 sg13g2_a22oi_1 _21963_ (.Y(_04417_),
    .B1(_04046_),
    .B2(net155),
    .A2(_04213_),
    .A1(net175));
 sg13g2_a22oi_1 _21964_ (.Y(_04418_),
    .B1(_03893_),
    .B2(net160),
    .A2(_03871_),
    .A1(net161));
 sg13g2_nand4_1 _21965_ (.B(_04416_),
    .C(_04417_),
    .A(_04415_),
    .Y(_04419_),
    .D(_04418_));
 sg13g2_a221oi_1 _21966_ (.B2(net114),
    .C1(_04419_),
    .B1(net113),
    .A1(net136),
    .Y(_04420_),
    .A2(_03857_));
 sg13g2_o21ai_1 _21967_ (.B1(_04420_),
    .Y(_04421_),
    .A1(net183),
    .A2(_04414_));
 sg13g2_a21oi_1 _21968_ (.A1(net180),
    .A2(net93),
    .Y(_04422_),
    .B1(_03954_));
 sg13g2_o21ai_1 _21969_ (.B1(_04422_),
    .Y(_04423_),
    .A1(_04409_),
    .A2(_04421_));
 sg13g2_or2_1 _21970_ (.X(_04424_),
    .B(_04093_),
    .A(_04106_));
 sg13g2_buf_1 _21971_ (.A(_04424_),
    .X(_04425_));
 sg13g2_xnor2_1 _21972_ (.Y(_04426_),
    .A(_04108_),
    .B(_04425_));
 sg13g2_nand2_2 _21973_ (.Y(_04427_),
    .A(_03955_),
    .B(_04191_));
 sg13g2_xor2_1 _21974_ (.B(_04425_),
    .A(_04010_),
    .X(_04428_));
 sg13g2_nor2b_1 _21975_ (.A(_04011_),
    .B_N(net1060),
    .Y(_04429_));
 sg13g2_o21ai_1 _21976_ (.B1(_04007_),
    .Y(_04430_),
    .A1(net978),
    .A2(_04429_));
 sg13g2_a221oi_1 _21977_ (.B2(net1048),
    .C1(_03972_),
    .B1(_04011_),
    .A1(_09048_),
    .Y(_04431_),
    .A2(_11609_));
 sg13g2_a22oi_1 _21978_ (.Y(_04432_),
    .B1(net111),
    .B2(net200),
    .A2(net131),
    .A1(net223));
 sg13g2_nand2b_1 _21979_ (.Y(_04433_),
    .B(_09850_),
    .A_N(_04432_));
 sg13g2_nand3_1 _21980_ (.B(_04431_),
    .C(_04433_),
    .A(_04430_),
    .Y(_04434_));
 sg13g2_a221oi_1 _21981_ (.B2(_04428_),
    .C1(_04434_),
    .B1(_04427_),
    .A1(net935),
    .Y(_04435_),
    .A2(_04426_));
 sg13g2_a22oi_1 _21982_ (.Y(_04436_),
    .B1(_04423_),
    .B2(_04435_),
    .A2(_11445_),
    .A1(net157));
 sg13g2_nand2_1 _21983_ (.Y(_04437_),
    .A(_03982_),
    .B(_04436_));
 sg13g2_nand4_1 _21984_ (.B(_04404_),
    .C(_04405_),
    .A(_04402_),
    .Y(_00981_),
    .D(_04437_));
 sg13g2_a21oi_1 _21985_ (.A1(_04007_),
    .A2(_04010_),
    .Y(_04438_),
    .B1(_04011_));
 sg13g2_xnor2_1 _21986_ (.Y(_04439_),
    .A(net231),
    .B(net180));
 sg13g2_xor2_1 _21987_ (.B(_04439_),
    .A(_04438_),
    .X(_04440_));
 sg13g2_a221oi_1 _21988_ (.B2(_04107_),
    .C1(_03947_),
    .B1(_03942_),
    .A1(_10547_),
    .Y(_04441_),
    .A2(_04006_));
 sg13g2_nor2_1 _21989_ (.A(_04106_),
    .B(_04441_),
    .Y(_04442_));
 sg13g2_xnor2_1 _21990_ (.Y(_04443_),
    .A(_04442_),
    .B(_04439_));
 sg13g2_nor2_1 _21991_ (.A(net231),
    .B(net180),
    .Y(_04444_));
 sg13g2_mux2_1 _21992_ (.A0(net1060),
    .A1(net1048),
    .S(_04444_),
    .X(_04445_));
 sg13g2_o21ai_1 _21993_ (.B1(_03997_),
    .Y(_04446_),
    .A1(net978),
    .A2(_04445_));
 sg13g2_a21oi_1 _21994_ (.A1(net1061),
    .A2(_10717_),
    .Y(_04447_),
    .B1(_04039_));
 sg13g2_nand2_1 _21995_ (.Y(_04448_),
    .A(_03585_),
    .B(net174));
 sg13g2_and3_1 _21996_ (.X(_04449_),
    .A(_11367_),
    .B(_04363_),
    .C(_04448_));
 sg13g2_or4_1 _21997_ (.A(net979),
    .B(_03918_),
    .C(_04365_),
    .D(_04449_),
    .X(_04450_));
 sg13g2_a22oi_1 _21998_ (.Y(_04451_),
    .B1(net156),
    .B2(net161),
    .A2(_03901_),
    .A1(net238));
 sg13g2_a22oi_1 _21999_ (.Y(_04452_),
    .B1(_03862_),
    .B2(net136),
    .A2(net182),
    .A1(net215));
 sg13g2_a22oi_1 _22000_ (.Y(_04453_),
    .B1(_03895_),
    .B2(net160),
    .A2(_03872_),
    .A1(_03891_));
 sg13g2_nor2_1 _22001_ (.A(net179),
    .B(_03883_),
    .Y(_04454_));
 sg13g2_a21oi_1 _22002_ (.A1(net237),
    .A2(_04214_),
    .Y(_04455_),
    .B1(_04454_));
 sg13g2_and4_1 _22003_ (.A(_04451_),
    .B(_04452_),
    .C(_04453_),
    .D(_04455_),
    .X(_04456_));
 sg13g2_a21oi_1 _22004_ (.A1(net112),
    .A2(net135),
    .Y(_04457_),
    .B1(net137));
 sg13g2_o21ai_1 _22005_ (.B1(_10604_),
    .Y(_04458_),
    .A1(_10602_),
    .A2(net183));
 sg13g2_nand2_1 _22006_ (.Y(_04459_),
    .A(_03915_),
    .B(_04458_));
 sg13g2_a22oi_1 _22007_ (.Y(_04460_),
    .B1(net162),
    .B2(net115),
    .A2(net133),
    .A1(net114));
 sg13g2_nand4_1 _22008_ (.B(_04457_),
    .C(_04459_),
    .A(_04456_),
    .Y(_04461_),
    .D(_04460_));
 sg13g2_nand2b_1 _22009_ (.Y(_04462_),
    .B(net111),
    .A_N(net159));
 sg13g2_nand3_1 _22010_ (.B(_04461_),
    .C(_04462_),
    .A(_03926_),
    .Y(_04463_));
 sg13g2_nand4_1 _22011_ (.B(_04447_),
    .C(_04450_),
    .A(_04446_),
    .Y(_04464_),
    .D(_04463_));
 sg13g2_a221oi_1 _22012_ (.B2(net935),
    .C1(_04464_),
    .B1(_04443_),
    .A1(_04427_),
    .Y(_04465_),
    .A2(_04440_));
 sg13g2_a21o_1 _22013_ (.A2(_11468_),
    .A1(net132),
    .B1(_04465_),
    .X(_04466_));
 sg13g2_nand2_1 _22014_ (.Y(_04467_),
    .A(net724),
    .B(net803));
 sg13g2_a21o_1 _22015_ (.A2(_04467_),
    .A1(net94),
    .B1(_03991_),
    .X(_04468_));
 sg13g2_nor2_1 _22016_ (.A(net642),
    .B(_04467_),
    .Y(_04469_));
 sg13g2_o21ai_1 _22017_ (.B1(_03988_),
    .Y(_04470_),
    .A1(_00255_),
    .A2(_04402_));
 sg13g2_a221oi_1 _22018_ (.B2(net94),
    .C1(_04470_),
    .B1(_04469_),
    .A1(net642),
    .Y(_04471_),
    .A2(_04468_));
 sg13g2_o21ai_1 _22019_ (.B1(_04471_),
    .Y(_00982_),
    .A1(net84),
    .A2(_04466_));
 sg13g2_nor3_1 _22020_ (.A(_03914_),
    .B(_03870_),
    .C(_03878_),
    .Y(_04472_));
 sg13g2_a21o_1 _22021_ (.A2(net162),
    .A1(net238),
    .B1(_04472_),
    .X(_04473_));
 sg13g2_a221oi_1 _22022_ (.B2(_10879_),
    .C1(_04473_),
    .B1(_03871_),
    .A1(net161),
    .Y(_04474_),
    .A2(net182));
 sg13g2_nor2_1 _22023_ (.A(_04025_),
    .B(_04271_),
    .Y(_04475_));
 sg13g2_a221oi_1 _22024_ (.B2(_03842_),
    .C1(_04475_),
    .B1(_03894_),
    .A1(net136),
    .Y(_04476_),
    .A2(_04060_));
 sg13g2_a21oi_1 _22025_ (.A1(net112),
    .A2(_04212_),
    .Y(_04477_),
    .B1(net137));
 sg13g2_nand2_1 _22026_ (.Y(_04478_),
    .A(_10604_),
    .B(net183));
 sg13g2_a221oi_1 _22027_ (.B2(_03915_),
    .C1(_04338_),
    .B1(_04478_),
    .A1(net178),
    .Y(_04479_),
    .A2(_04056_));
 sg13g2_nand4_1 _22028_ (.B(_04476_),
    .C(_04477_),
    .A(_04474_),
    .Y(_04480_),
    .D(_04479_));
 sg13g2_a21oi_1 _22029_ (.A1(_03885_),
    .A2(net137),
    .Y(_04481_),
    .B1(_03954_));
 sg13g2_o21ai_1 _22030_ (.B1(net180),
    .Y(_04482_),
    .A1(net233),
    .A2(_04006_));
 sg13g2_o21ai_1 _22031_ (.B1(_11454_),
    .Y(_04483_),
    .A1(_04441_),
    .A2(_04482_));
 sg13g2_o21ai_1 _22032_ (.B1(_04483_),
    .Y(_04484_),
    .A1(net180),
    .A2(_04442_));
 sg13g2_nor2_1 _22033_ (.A(_04103_),
    .B(_04092_),
    .Y(_04485_));
 sg13g2_xor2_1 _22034_ (.B(_04485_),
    .A(_04484_),
    .X(_04486_));
 sg13g2_nor3_1 _22035_ (.A(_03918_),
    .B(_04006_),
    .C(_03854_),
    .Y(_04487_));
 sg13g2_a21oi_1 _22036_ (.A1(_04049_),
    .A2(_04045_),
    .Y(_04488_),
    .B1(_04487_));
 sg13g2_a21oi_1 _22037_ (.A1(_11189_),
    .A2(_04060_),
    .Y(_04489_),
    .B1(_03967_));
 sg13g2_a221oi_1 _22038_ (.B2(_04489_),
    .C1(net979),
    .B1(_04488_),
    .A1(net180),
    .Y(_04490_),
    .A2(net137));
 sg13g2_a21oi_1 _22039_ (.A1(_09048_),
    .A2(_10690_),
    .Y(_04491_),
    .B1(_04193_));
 sg13g2_mux2_1 _22040_ (.A0(net1121),
    .A1(_09073_),
    .S(_04015_),
    .X(_04492_));
 sg13g2_o21ai_1 _22041_ (.B1(_04146_),
    .Y(_04493_),
    .A1(_09834_),
    .A2(_04492_));
 sg13g2_nand3b_1 _22042_ (.B(_04491_),
    .C(_04493_),
    .Y(_04494_),
    .A_N(_04490_));
 sg13g2_a221oi_1 _22043_ (.B2(net1077),
    .C1(_04494_),
    .B1(_04486_),
    .A1(_04480_),
    .Y(_04495_),
    .A2(_04481_));
 sg13g2_nor2_1 _22044_ (.A(_04147_),
    .B(_04013_),
    .Y(_04496_));
 sg13g2_xor2_1 _22045_ (.B(_04485_),
    .A(_04496_),
    .X(_04497_));
 sg13g2_a21oi_1 _22046_ (.A1(_03955_),
    .A2(_04495_),
    .Y(_04498_),
    .B1(_04497_));
 sg13g2_nor2_1 _22047_ (.A(_04193_),
    .B(_04495_),
    .Y(_04499_));
 sg13g2_nor3_1 _22048_ (.A(net157),
    .B(_04498_),
    .C(_04499_),
    .Y(_04500_));
 sg13g2_a21o_1 _22049_ (.A2(_11479_),
    .A1(net157),
    .B1(_04500_),
    .X(_04501_));
 sg13g2_nor2_1 _22050_ (.A(_08442_),
    .B(_04181_),
    .Y(_04502_));
 sg13g2_nor3_1 _22051_ (.A(_08341_),
    .B(net916),
    .C(_11393_),
    .Y(_04503_));
 sg13g2_a21oi_1 _22052_ (.A1(net94),
    .A2(_04181_),
    .Y(_04504_),
    .B1(_03991_));
 sg13g2_nor2_1 _22053_ (.A(_08444_),
    .B(_04504_),
    .Y(_04505_));
 sg13g2_a221oi_1 _22054_ (.B2(net288),
    .C1(_04505_),
    .B1(_04503_),
    .A1(net94),
    .Y(_04506_),
    .A2(_04502_));
 sg13g2_o21ai_1 _22055_ (.B1(_04506_),
    .Y(_00983_),
    .A1(net84),
    .A2(_04501_));
 sg13g2_nand2_1 _22056_ (.Y(_04507_),
    .A(_04146_),
    .B(_04148_));
 sg13g2_xnor2_1 _22057_ (.Y(_04508_),
    .A(net216),
    .B(net179));
 sg13g2_xor2_1 _22058_ (.B(_04508_),
    .A(_04507_),
    .X(_04509_));
 sg13g2_nand2_1 _22059_ (.Y(_04510_),
    .A(_04427_),
    .B(_04509_));
 sg13g2_inv_1 _22060_ (.Y(_04511_),
    .A(_04092_));
 sg13g2_a21oi_1 _22061_ (.A1(_04511_),
    .A2(_04484_),
    .Y(_04512_),
    .B1(_04103_));
 sg13g2_xnor2_1 _22062_ (.Y(_04513_),
    .A(_04512_),
    .B(_04508_));
 sg13g2_o21ai_1 _22063_ (.B1(_04277_),
    .Y(_04514_),
    .A1(_03896_),
    .A2(_04276_));
 sg13g2_a221oi_1 _22064_ (.B2(net160),
    .C1(_04514_),
    .B1(_04057_),
    .A1(net163),
    .Y(_04515_),
    .A2(net165));
 sg13g2_o21ai_1 _22065_ (.B1(_11452_),
    .Y(_04516_),
    .A1(_11432_),
    .A2(net234));
 sg13g2_a21o_1 _22066_ (.A2(_04516_),
    .A1(_10604_),
    .B1(net181),
    .X(_04517_));
 sg13g2_and2_1 _22067_ (.A(net238),
    .B(net138),
    .X(_04518_));
 sg13g2_a21o_1 _22068_ (.A2(net164),
    .A1(_03843_),
    .B1(_04518_),
    .X(_04519_));
 sg13g2_a221oi_1 _22069_ (.B2(net237),
    .C1(_04519_),
    .B1(net162),
    .A1(net114),
    .Y(_04520_),
    .A2(net131));
 sg13g2_nand4_1 _22070_ (.B(_04515_),
    .C(_04517_),
    .A(_04047_),
    .Y(_04521_),
    .D(_04520_));
 sg13g2_a21oi_1 _22071_ (.A1(_03995_),
    .A2(net93),
    .Y(_04522_),
    .B1(_03954_));
 sg13g2_a221oi_1 _22072_ (.B2(net174),
    .C1(_03884_),
    .B1(net135),
    .A1(_04054_),
    .Y(_04523_),
    .A2(net113));
 sg13g2_a21oi_1 _22073_ (.A1(net133),
    .A2(net200),
    .Y(_04524_),
    .B1(net111));
 sg13g2_nand2_1 _22074_ (.Y(_04525_),
    .A(_04523_),
    .B(_04524_));
 sg13g2_nand3_1 _22075_ (.B(_04462_),
    .C(_04525_),
    .A(_09850_),
    .Y(_04526_));
 sg13g2_mux2_1 _22076_ (.A0(net1048),
    .A1(_09074_),
    .S(_04018_),
    .X(_04527_));
 sg13g2_o21ai_1 _22077_ (.B1(_03998_),
    .Y(_04528_),
    .A1(net978),
    .A2(_04527_));
 sg13g2_a21oi_1 _22078_ (.A1(net1061),
    .A2(_11695_),
    .Y(_04529_),
    .B1(net157));
 sg13g2_nand3_1 _22079_ (.B(_04528_),
    .C(_04529_),
    .A(_04526_),
    .Y(_04530_));
 sg13g2_a221oi_1 _22080_ (.B2(_04522_),
    .C1(_04530_),
    .B1(_04521_),
    .A1(_08281_),
    .Y(_04531_),
    .A2(_04513_));
 sg13g2_a22oi_1 _22081_ (.Y(_04532_),
    .B1(_04510_),
    .B2(_04531_),
    .A2(_11494_),
    .A1(net132));
 sg13g2_nand2_1 _22082_ (.Y(_04533_),
    .A(_03982_),
    .B(_04532_));
 sg13g2_buf_1 _22083_ (.A(_08667_),
    .X(_04534_));
 sg13g2_xnor2_1 _22084_ (.Y(_04535_),
    .A(_10629_),
    .B(_04182_));
 sg13g2_a22oi_1 _22085_ (.Y(_04536_),
    .B1(_04535_),
    .B2(net83),
    .A2(net35),
    .A1(net977));
 sg13g2_nand2_1 _22086_ (.Y(_00984_),
    .A(_04533_),
    .B(_04536_));
 sg13g2_nand3_1 _22087_ (.B(_04114_),
    .C(_04118_),
    .A(_04105_),
    .Y(_04537_));
 sg13g2_nand2b_1 _22088_ (.Y(_04538_),
    .B(_04121_),
    .A_N(_04115_));
 sg13g2_xnor2_1 _22089_ (.Y(_04539_),
    .A(_04537_),
    .B(_04538_));
 sg13g2_nor2_1 _22090_ (.A(_04163_),
    .B(_04020_),
    .Y(_04540_));
 sg13g2_xnor2_1 _22091_ (.Y(_04541_),
    .A(_04540_),
    .B(_04538_));
 sg13g2_mux2_1 _22092_ (.A0(net1121),
    .A1(_09073_),
    .S(_04022_),
    .X(_04542_));
 sg13g2_o21ai_1 _22093_ (.B1(_03996_),
    .Y(_04543_),
    .A1(_09834_),
    .A2(_04542_));
 sg13g2_a22oi_1 _22094_ (.Y(_04544_),
    .B1(_04045_),
    .B2(net134),
    .A2(_04212_),
    .A1(net175));
 sg13g2_a22oi_1 _22095_ (.Y(_04545_),
    .B1(_04060_),
    .B2(_11157_),
    .A2(net182),
    .A1(_11189_));
 sg13g2_a21oi_1 _22096_ (.A1(_03861_),
    .A2(_04049_),
    .Y(_04546_),
    .B1(_03968_));
 sg13g2_nand3_1 _22097_ (.B(_04545_),
    .C(_04546_),
    .A(_04544_),
    .Y(_04547_));
 sg13g2_a21oi_1 _22098_ (.A1(_03885_),
    .A2(net137),
    .Y(_04548_),
    .B1(net979));
 sg13g2_a221oi_1 _22099_ (.B2(_04548_),
    .C1(_03972_),
    .B1(_04547_),
    .A1(_09048_),
    .Y(_04549_),
    .A2(_10292_));
 sg13g2_nand2_1 _22100_ (.Y(_04550_),
    .A(_04543_),
    .B(_04549_));
 sg13g2_nand2_1 _22101_ (.Y(_04551_),
    .A(net237),
    .B(_03894_));
 sg13g2_nand2_1 _22102_ (.Y(_04552_),
    .A(_04043_),
    .B(_04212_));
 sg13g2_a22oi_1 _22103_ (.Y(_04553_),
    .B1(_04056_),
    .B2(_03842_),
    .A2(_03871_),
    .A1(net238));
 sg13g2_nand4_1 _22104_ (.B(_04551_),
    .C(_04552_),
    .A(_04216_),
    .Y(_04554_),
    .D(_04553_));
 sg13g2_a22oi_1 _22105_ (.Y(_04555_),
    .B1(_03861_),
    .B2(net178),
    .A2(_03856_),
    .A1(net193));
 sg13g2_nand2b_1 _22106_ (.Y(_04556_),
    .B(_04555_),
    .A_N(_04342_));
 sg13g2_o21ai_1 _22107_ (.B1(_03926_),
    .Y(_04557_),
    .A1(_04554_),
    .A2(_04556_));
 sg13g2_a22oi_1 _22108_ (.Y(_04558_),
    .B1(_04517_),
    .B2(_04557_),
    .A2(net111),
    .A1(_04025_));
 sg13g2_or2_1 _22109_ (.X(_04559_),
    .B(_04558_),
    .A(_04550_));
 sg13g2_a221oi_1 _22110_ (.B2(_04427_),
    .C1(_04559_),
    .B1(_04541_),
    .A1(net1077),
    .Y(_04560_),
    .A2(_04539_));
 sg13g2_a21o_1 _22111_ (.A2(_11518_),
    .A1(net157),
    .B1(_04560_),
    .X(_04561_));
 sg13g2_buf_1 _22112_ (.A(_08624_),
    .X(_04562_));
 sg13g2_nand2_1 _22113_ (.Y(_04563_),
    .A(_08667_),
    .B(_04182_));
 sg13g2_xor2_1 _22114_ (.B(_04563_),
    .A(_10330_),
    .X(_04564_));
 sg13g2_a22oi_1 _22115_ (.Y(_04565_),
    .B1(_04564_),
    .B2(net83),
    .A2(net35),
    .A1(net976));
 sg13g2_o21ai_1 _22116_ (.B1(_04565_),
    .Y(_00985_),
    .A1(_03837_),
    .A2(_04561_));
 sg13g2_a22oi_1 _22117_ (.Y(_04566_),
    .B1(_03861_),
    .B2(_03899_),
    .A2(_03856_),
    .A1(_03842_));
 sg13g2_a221oi_1 _22118_ (.B2(net238),
    .C1(_04066_),
    .B1(_04056_),
    .A1(_03890_),
    .Y(_04567_),
    .A2(net133));
 sg13g2_nand3b_1 _22119_ (.B(_04566_),
    .C(_04567_),
    .Y(_04568_),
    .A_N(_04272_));
 sg13g2_nor3_1 _22120_ (.A(_03868_),
    .B(net130),
    .C(_03870_),
    .Y(_04569_));
 sg13g2_o21ai_1 _22121_ (.B1(_09831_),
    .Y(_04570_),
    .A1(_04568_),
    .A2(_04569_));
 sg13g2_a21oi_1 _22122_ (.A1(_11454_),
    .A2(_10604_),
    .Y(_04571_),
    .B1(net130));
 sg13g2_o21ai_1 _22123_ (.B1(net1130),
    .Y(_04572_),
    .A1(_04568_),
    .A2(_04571_));
 sg13g2_a22oi_1 _22124_ (.Y(_04573_),
    .B1(_04570_),
    .B2(_04572_),
    .A2(net93),
    .A1(net176));
 sg13g2_a221oi_1 _22125_ (.B2(net165),
    .C1(_04454_),
    .B1(_04050_),
    .A1(_04053_),
    .Y(_04574_),
    .A2(net133));
 sg13g2_o21ai_1 _22126_ (.B1(net158),
    .Y(_04575_),
    .A1(_04006_),
    .A2(_04276_));
 sg13g2_a221oi_1 _22127_ (.B2(net159),
    .C1(_04575_),
    .B1(net135),
    .A1(_04054_),
    .Y(_04576_),
    .A2(net156));
 sg13g2_a221oi_1 _22128_ (.B2(_04576_),
    .C1(_03969_),
    .B1(_04574_),
    .A1(_03995_),
    .Y(_04577_),
    .A2(net93));
 sg13g2_mux2_1 _22129_ (.A0(_09848_),
    .A1(net1060),
    .S(_04150_),
    .X(_04578_));
 sg13g2_nor2_1 _22130_ (.A(net978),
    .B(_04578_),
    .Y(_04579_));
 sg13g2_a21oi_1 _22131_ (.A1(_09049_),
    .A2(_11763_),
    .Y(_04580_),
    .B1(net157));
 sg13g2_o21ai_1 _22132_ (.B1(_04580_),
    .Y(_04581_),
    .A1(_04157_),
    .A2(_04579_));
 sg13g2_nor3_1 _22133_ (.A(_04573_),
    .B(_04577_),
    .C(_04581_),
    .Y(_04582_));
 sg13g2_nor2b_1 _22134_ (.A(_04028_),
    .B_N(_04029_),
    .Y(_04583_));
 sg13g2_a21oi_1 _22135_ (.A1(_04537_),
    .A2(_04121_),
    .Y(_04584_),
    .B1(_04115_));
 sg13g2_xnor2_1 _22136_ (.Y(_04585_),
    .A(_04026_),
    .B(_04584_));
 sg13g2_a22oi_1 _22137_ (.Y(_04586_),
    .B1(_04585_),
    .B2(net935),
    .A2(_04427_),
    .A1(_04583_));
 sg13g2_nand2_1 _22138_ (.Y(_04587_),
    .A(_04582_),
    .B(_04586_));
 sg13g2_o21ai_1 _22139_ (.B1(_04587_),
    .Y(_04588_),
    .A1(net166),
    .A2(\cpu.ex.c_mult[7] ));
 sg13g2_buf_1 _22140_ (.A(_08633_),
    .X(_04589_));
 sg13g2_nand3_1 _22141_ (.B(_08624_),
    .C(_04182_),
    .A(_08667_),
    .Y(_04590_));
 sg13g2_xor2_1 _22142_ (.B(_04590_),
    .A(_10457_),
    .X(_04591_));
 sg13g2_a22oi_1 _22143_ (.Y(_04592_),
    .B1(_04591_),
    .B2(net83),
    .A2(net35),
    .A1(net975));
 sg13g2_o21ai_1 _22144_ (.B1(_04592_),
    .Y(_00986_),
    .A1(net84),
    .A2(_04588_));
 sg13g2_nand3b_1 _22145_ (.B(_11561_),
    .C(net132),
    .Y(_04593_),
    .A_N(_11559_));
 sg13g2_and2_1 _22146_ (.A(_04120_),
    .B(_04124_),
    .X(_04594_));
 sg13g2_nor2_1 _22147_ (.A(net192),
    .B(net176),
    .Y(_04595_));
 sg13g2_inv_1 _22148_ (.Y(_04596_),
    .A(_04136_));
 sg13g2_nor2_1 _22149_ (.A(_04595_),
    .B(_04596_),
    .Y(_04597_));
 sg13g2_xor2_1 _22150_ (.B(_04597_),
    .A(_04594_),
    .X(_04598_));
 sg13g2_nand2_1 _22151_ (.Y(_04599_),
    .A(net1130),
    .B(_04571_));
 sg13g2_a22oi_1 _22152_ (.Y(_04600_),
    .B1(_04061_),
    .B2(net160),
    .A2(net113),
    .A1(_03843_));
 sg13g2_nor2_1 _22153_ (.A(net130),
    .B(_03905_),
    .Y(_04601_));
 sg13g2_a221oi_1 _22154_ (.B2(net161),
    .C1(_04601_),
    .B1(net131),
    .A1(_10914_),
    .Y(_04602_),
    .A2(net165));
 sg13g2_nand4_1 _22155_ (.B(_04599_),
    .C(_04600_),
    .A(_04337_),
    .Y(_04603_),
    .D(_04602_));
 sg13g2_a21oi_1 _22156_ (.A1(_04065_),
    .A2(net93),
    .Y(_04604_),
    .B1(_03954_));
 sg13g2_mux2_1 _22157_ (.A0(_09073_),
    .A1(net1121),
    .S(_04199_),
    .X(_04605_));
 sg13g2_nand2_1 _22158_ (.Y(_04606_),
    .A(_11600_),
    .B(net176));
 sg13g2_o21ai_1 _22159_ (.B1(_04606_),
    .Y(_04607_),
    .A1(_04033_),
    .A2(_04605_));
 sg13g2_a22oi_1 _22160_ (.Y(_04608_),
    .B1(net135),
    .B2(net155),
    .A2(net133),
    .A1(_03909_));
 sg13g2_a22oi_1 _22161_ (.Y(_04609_),
    .B1(net113),
    .B2(net134),
    .A2(net182),
    .A1(net174));
 sg13g2_a22oi_1 _22162_ (.Y(_04610_),
    .B1(net156),
    .B2(_04049_),
    .A2(net164),
    .A1(_11189_));
 sg13g2_nand4_1 _22163_ (.B(_04608_),
    .C(_04609_),
    .A(_04477_),
    .Y(_04611_),
    .D(_04610_));
 sg13g2_a21oi_1 _22164_ (.A1(_04025_),
    .A2(net111),
    .Y(_04612_),
    .B1(net979));
 sg13g2_nand2_1 _22165_ (.Y(_04613_),
    .A(_04611_),
    .B(_04612_));
 sg13g2_nand2_1 _22166_ (.Y(_04614_),
    .A(net1061),
    .B(_11367_));
 sg13g2_nand3_1 _22167_ (.B(_04613_),
    .C(_04614_),
    .A(_04607_),
    .Y(_04615_));
 sg13g2_a221oi_1 _22168_ (.B2(_04604_),
    .C1(_04615_),
    .B1(_04603_),
    .A1(_08280_),
    .Y(_04616_),
    .A2(_04598_));
 sg13g2_nor2b_1 _22169_ (.A(_04032_),
    .B_N(_04616_),
    .Y(_04617_));
 sg13g2_xnor2_1 _22170_ (.Y(_04618_),
    .A(_04158_),
    .B(_04597_));
 sg13g2_nor2_1 _22171_ (.A(_03959_),
    .B(_04618_),
    .Y(_04619_));
 sg13g2_o21ai_1 _22172_ (.B1(net166),
    .Y(_04620_),
    .A1(_04617_),
    .A2(_04619_));
 sg13g2_nand2_1 _22173_ (.Y(_04621_),
    .A(_04593_),
    .B(_04620_));
 sg13g2_xor2_1 _22174_ (.B(_04183_),
    .A(_10427_),
    .X(_04622_));
 sg13g2_a22oi_1 _22175_ (.Y(_04623_),
    .B1(_04622_),
    .B2(net83),
    .A2(_03991_),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_o21ai_1 _22176_ (.B1(_04623_),
    .Y(_00987_),
    .A1(net84),
    .A2(_04621_));
 sg13g2_nor4_1 _22177_ (.A(_03838_),
    .B(_11573_),
    .C(_11578_),
    .D(_11582_),
    .Y(_04624_));
 sg13g2_a21oi_1 _22178_ (.A1(net136),
    .A2(_04158_),
    .Y(_04625_),
    .B1(_04170_));
 sg13g2_xnor2_1 _22179_ (.Y(_04626_),
    .A(net228),
    .B(net154));
 sg13g2_xnor2_1 _22180_ (.Y(_04627_),
    .A(_04625_),
    .B(_04626_));
 sg13g2_a21oi_1 _22181_ (.A1(_04594_),
    .A2(_04136_),
    .Y(_04628_),
    .B1(_04595_));
 sg13g2_xor2_1 _22182_ (.B(_04626_),
    .A(_04628_),
    .X(_04629_));
 sg13g2_a22oi_1 _22183_ (.Y(_04630_),
    .B1(net156),
    .B2(_03921_),
    .A2(net138),
    .A1(net223));
 sg13g2_a22oi_1 _22184_ (.Y(_04631_),
    .B1(_04053_),
    .B2(net165),
    .A2(net113),
    .A1(net159));
 sg13g2_a221oi_1 _22185_ (.B2(net164),
    .C1(_03888_),
    .B1(net200),
    .A1(net114),
    .Y(_04632_),
    .A2(net131));
 sg13g2_nand4_1 _22186_ (.B(_04630_),
    .C(_04631_),
    .A(_04457_),
    .Y(_04633_),
    .D(_04632_));
 sg13g2_a21oi_1 _22187_ (.A1(net176),
    .A2(_04069_),
    .Y(_04634_),
    .B1(net979));
 sg13g2_a22oi_1 _22188_ (.Y(_04635_),
    .B1(_04212_),
    .B2(_03890_),
    .A2(_03861_),
    .A1(net238));
 sg13g2_a22oi_1 _22189_ (.Y(_04636_),
    .B1(_04060_),
    .B2(_03842_),
    .A2(net182),
    .A1(_10937_));
 sg13g2_nand3_1 _22190_ (.B(_04635_),
    .C(_04636_),
    .A(_04369_),
    .Y(_04637_));
 sg13g2_a21o_1 _22191_ (.A2(_04637_),
    .A1(_09831_),
    .B1(_09066_),
    .X(_04638_));
 sg13g2_nor3_1 _22192_ (.A(_04571_),
    .B(_04601_),
    .C(_04637_),
    .Y(_04639_));
 sg13g2_a21oi_1 _22193_ (.A1(_03896_),
    .A2(_04069_),
    .Y(_04640_),
    .B1(_04639_));
 sg13g2_mux2_1 _22194_ (.A0(net1121),
    .A1(_09073_),
    .S(_04203_),
    .X(_04641_));
 sg13g2_o21ai_1 _22195_ (.B1(_04173_),
    .Y(_04642_),
    .A1(_09834_),
    .A2(_04641_));
 sg13g2_o21ai_1 _22196_ (.B1(_04642_),
    .Y(_04643_),
    .A1(_04233_),
    .A2(net202));
 sg13g2_a221oi_1 _22197_ (.B2(_04640_),
    .C1(_04643_),
    .B1(_04638_),
    .A1(_04633_),
    .Y(_04644_),
    .A2(_04634_));
 sg13g2_nand3_1 _22198_ (.B(_04031_),
    .C(_04644_),
    .A(_03838_),
    .Y(_04645_));
 sg13g2_a221oi_1 _22199_ (.B2(net935),
    .C1(_04645_),
    .B1(_04629_),
    .A1(_04193_),
    .Y(_04646_),
    .A2(_04627_));
 sg13g2_or2_1 _22200_ (.X(_04647_),
    .B(_04646_),
    .A(_04624_));
 sg13g2_buf_1 _22201_ (.A(_08680_),
    .X(_04648_));
 sg13g2_xnor2_1 _22202_ (.Y(_04649_),
    .A(_10293_),
    .B(_04184_));
 sg13g2_a22oi_1 _22203_ (.Y(_04650_),
    .B1(_04649_),
    .B2(_03979_),
    .A2(_03991_),
    .A1(net974));
 sg13g2_o21ai_1 _22204_ (.B1(_04650_),
    .Y(_00988_),
    .A1(_03836_),
    .A2(_04647_));
 sg13g2_or2_1 _22205_ (.X(_04651_),
    .B(_04141_),
    .A(_04128_));
 sg13g2_buf_1 _22206_ (.A(_04651_),
    .X(_04652_));
 sg13g2_nand3_1 _22207_ (.B(_04203_),
    .C(_04652_),
    .A(_04625_),
    .Y(_04653_));
 sg13g2_nor2b_1 _22208_ (.A(_04652_),
    .B_N(_04173_),
    .Y(_04654_));
 sg13g2_nand2b_1 _22209_ (.Y(_04655_),
    .B(_04654_),
    .A_N(_04625_));
 sg13g2_a21o_1 _22210_ (.A2(_04655_),
    .A1(_04653_),
    .B1(_03959_),
    .X(_04656_));
 sg13g2_nand2b_1 _22211_ (.Y(_04657_),
    .B(_04652_),
    .A_N(_04173_));
 sg13g2_o21ai_1 _22212_ (.B1(_04657_),
    .Y(_04658_),
    .A1(_04203_),
    .A2(_04652_));
 sg13g2_a21oi_1 _22213_ (.A1(net155),
    .A2(_03861_),
    .Y(_04659_),
    .B1(net137));
 sg13g2_a22oi_1 _22214_ (.Y(_04660_),
    .B1(net133),
    .B2(net112),
    .A2(net164),
    .A1(_03921_));
 sg13g2_nand2_1 _22215_ (.Y(_04661_),
    .A(_04659_),
    .B(_04660_));
 sg13g2_a221oi_1 _22216_ (.B2(net114),
    .C1(_04661_),
    .B1(net135),
    .A1(net159),
    .Y(_04662_),
    .A2(_03857_));
 sg13g2_a22oi_1 _22217_ (.Y(_04663_),
    .B1(net200),
    .B2(net138),
    .A2(net156),
    .A1(net134));
 sg13g2_nand2_1 _22218_ (.Y(_04664_),
    .A(net223),
    .B(net162));
 sg13g2_nand4_1 _22219_ (.B(_04662_),
    .C(_04663_),
    .A(_04552_),
    .Y(_04665_),
    .D(_04664_));
 sg13g2_a21oi_1 _22220_ (.A1(_04065_),
    .A2(net93),
    .Y(_04666_),
    .B1(net979));
 sg13g2_o21ai_1 _22221_ (.B1(_03926_),
    .Y(_04667_),
    .A1(net163),
    .A2(_03924_));
 sg13g2_o21ai_1 _22222_ (.B1(_03924_),
    .Y(_04668_),
    .A1(net130),
    .A2(_04276_));
 sg13g2_a221oi_1 _22223_ (.B2(net115),
    .C1(_04668_),
    .B1(net135),
    .A1(net160),
    .Y(_04669_),
    .A2(net131));
 sg13g2_o21ai_1 _22224_ (.B1(_04669_),
    .Y(_04670_),
    .A1(net222),
    .A2(_03887_));
 sg13g2_nand2b_1 _22225_ (.Y(_04671_),
    .B(_04670_),
    .A_N(_04667_));
 sg13g2_o21ai_1 _22226_ (.B1(_11432_),
    .Y(_04672_),
    .A1(net1061),
    .A2(_04410_));
 sg13g2_mux2_1 _22227_ (.A0(net1060),
    .A1(net1048),
    .S(_04174_),
    .X(_04673_));
 sg13g2_o21ai_1 _22228_ (.B1(_04172_),
    .Y(_04674_),
    .A1(net978),
    .A2(_04673_));
 sg13g2_nand4_1 _22229_ (.B(_04671_),
    .C(_04672_),
    .A(_04599_),
    .Y(_04675_),
    .D(_04674_));
 sg13g2_a221oi_1 _22230_ (.B2(_04666_),
    .C1(_04675_),
    .B1(_04665_),
    .A1(_04193_),
    .Y(_04676_),
    .A2(_04658_));
 sg13g2_a22oi_1 _22231_ (.Y(_04677_),
    .B1(_04125_),
    .B2(_04126_),
    .A2(_04124_),
    .A1(_04120_));
 sg13g2_a22oi_1 _22232_ (.Y(_04678_),
    .B1(_04131_),
    .B2(_11597_),
    .A2(_04124_),
    .A1(_04120_));
 sg13g2_inv_1 _22233_ (.Y(_04679_),
    .A(_04131_));
 sg13g2_a22oi_1 _22234_ (.Y(_04680_),
    .B1(_04679_),
    .B2(net176),
    .A2(_04596_),
    .A1(net228));
 sg13g2_nand2_1 _22235_ (.Y(_04681_),
    .A(_04134_),
    .B(_04680_));
 sg13g2_nor3_1 _22236_ (.A(_04677_),
    .B(_04678_),
    .C(_04681_),
    .Y(_04682_));
 sg13g2_xnor2_1 _22237_ (.Y(_04683_),
    .A(_04682_),
    .B(_04652_));
 sg13g2_nand2_1 _22238_ (.Y(_04684_),
    .A(net935),
    .B(_04683_));
 sg13g2_nand4_1 _22239_ (.B(_04656_),
    .C(_04676_),
    .A(_04321_),
    .Y(_04685_),
    .D(_04684_));
 sg13g2_nand3_1 _22240_ (.B(_11617_),
    .C(_11619_),
    .A(net132),
    .Y(_04686_));
 sg13g2_nand3_1 _22241_ (.B(_04685_),
    .C(_04686_),
    .A(_03982_),
    .Y(_04687_));
 sg13g2_buf_1 _22242_ (.A(_08652_),
    .X(_04688_));
 sg13g2_nand2_1 _22243_ (.Y(_04689_),
    .A(_08680_),
    .B(_04184_));
 sg13g2_xor2_1 _22244_ (.B(_04689_),
    .A(_10365_),
    .X(_04690_));
 sg13g2_a22oi_1 _22245_ (.Y(_04691_),
    .B1(_04690_),
    .B2(_04187_),
    .A2(_03992_),
    .A1(net973));
 sg13g2_nand2_1 _22246_ (.Y(_00989_),
    .A(_04687_),
    .B(_04691_));
 sg13g2_buf_1 _22247_ (.A(_00236_),
    .X(_04692_));
 sg13g2_nor4_1 _22248_ (.A(net1117),
    .B(_10140_),
    .C(_04692_),
    .D(_03457_),
    .Y(_04693_));
 sg13g2_buf_2 _22249_ (.A(_04693_),
    .X(_04694_));
 sg13g2_buf_1 _22250_ (.A(_04694_),
    .X(_04695_));
 sg13g2_mux2_1 _22251_ (.A0(_10589_),
    .A1(net552),
    .S(net541),
    .X(_00992_));
 sg13g2_mux2_1 _22252_ (.A0(_10697_),
    .A1(net852),
    .S(net541),
    .X(_00993_));
 sg13g2_buf_1 _22253_ (.A(net611),
    .X(_04696_));
 sg13g2_mux2_1 _22254_ (.A0(_10664_),
    .A1(_04696_),
    .S(net541),
    .X(_00994_));
 sg13g2_mux2_1 _22255_ (.A0(_10394_),
    .A1(net547),
    .S(_04695_),
    .X(_00995_));
 sg13g2_mux2_1 _22256_ (.A0(_10278_),
    .A1(net674),
    .S(_04695_),
    .X(_00996_));
 sg13g2_mux2_1 _22257_ (.A0(_10200_),
    .A1(net744),
    .S(net541),
    .X(_00997_));
 sg13g2_mux2_1 _22258_ (.A0(_10524_),
    .A1(net434),
    .S(net541),
    .X(_00998_));
 sg13g2_mux2_1 _22259_ (.A0(_10492_),
    .A1(net435),
    .S(net541),
    .X(_00999_));
 sg13g2_mux2_1 _22260_ (.A0(_10644_),
    .A1(net477),
    .S(net541),
    .X(_01000_));
 sg13g2_mux2_1 _22261_ (.A0(_10622_),
    .A1(net556),
    .S(net541),
    .X(_01001_));
 sg13g2_mux2_1 _22262_ (.A0(_10354_),
    .A1(net743),
    .S(_04694_),
    .X(_01002_));
 sg13g2_mux2_1 _22263_ (.A0(_10460_),
    .A1(net742),
    .S(_04694_),
    .X(_01003_));
 sg13g2_mux2_1 _22264_ (.A0(_10449_),
    .A1(net850),
    .S(_04694_),
    .X(_01004_));
 sg13g2_mux2_1 _22265_ (.A0(_10310_),
    .A1(net849),
    .S(_04694_),
    .X(_01005_));
 sg13g2_mux2_1 _22266_ (.A0(_10376_),
    .A1(net851),
    .S(_04694_),
    .X(_01006_));
 sg13g2_or2_1 _22267_ (.X(_04697_),
    .B(_03457_),
    .A(_10141_));
 sg13g2_buf_1 _22268_ (.A(_04697_),
    .X(_04698_));
 sg13g2_buf_1 _22269_ (.A(_04698_),
    .X(_04699_));
 sg13g2_nor2_1 _22270_ (.A(_08428_),
    .B(_04692_),
    .Y(_04700_));
 sg13g2_nand2_1 _22271_ (.Y(_04701_),
    .A(_03455_),
    .B(_04700_));
 sg13g2_nor2_1 _22272_ (.A(net819),
    .B(_11374_),
    .Y(_04702_));
 sg13g2_a21oi_1 _22273_ (.A1(_11374_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_or4_1 _22274_ (.A(net1117),
    .B(_04692_),
    .C(_03457_),
    .D(_04703_),
    .X(_04704_));
 sg13g2_buf_1 _22275_ (.A(_04704_),
    .X(_04705_));
 sg13g2_buf_1 _22276_ (.A(net476),
    .X(_04706_));
 sg13g2_nand2_1 _22277_ (.Y(_04707_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net433));
 sg13g2_o21ai_1 _22278_ (.B1(_04707_),
    .Y(_01007_),
    .A1(net539),
    .A2(_04701_));
 sg13g2_buf_1 _22279_ (.A(net476),
    .X(_04708_));
 sg13g2_buf_1 _22280_ (.A(net598),
    .X(_04709_));
 sg13g2_nor2_1 _22281_ (.A(_02931_),
    .B(_04709_),
    .Y(_04710_));
 sg13g2_a21oi_1 _22282_ (.A1(_10376_),
    .A2(net539),
    .Y(_04711_),
    .B1(_04710_));
 sg13g2_nand2_1 _22283_ (.Y(_04712_),
    .A(\cpu.ex.r_stmp[10] ),
    .B(net433));
 sg13g2_o21ai_1 _22284_ (.B1(_04712_),
    .Y(_01008_),
    .A1(net432),
    .A2(_04711_));
 sg13g2_mux2_1 _22285_ (.A0(_10693_),
    .A1(_10697_),
    .S(net538),
    .X(_04713_));
 sg13g2_mux2_1 _22286_ (.A0(_04713_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net433),
    .X(_01009_));
 sg13g2_mux2_1 _22287_ (.A0(net695),
    .A1(_10664_),
    .S(net538),
    .X(_04714_));
 sg13g2_mux2_1 _22288_ (.A0(_04714_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net433),
    .X(_01010_));
 sg13g2_mux2_1 _22289_ (.A0(net696),
    .A1(_10394_),
    .S(net538),
    .X(_04715_));
 sg13g2_mux2_1 _22290_ (.A0(_04715_),
    .A1(\cpu.ex.r_stmp[13] ),
    .S(net433),
    .X(_01011_));
 sg13g2_nor2_1 _22291_ (.A(_03536_),
    .B(net538),
    .Y(_04716_));
 sg13g2_a21oi_1 _22292_ (.A1(_10278_),
    .A2(_04699_),
    .Y(_04717_),
    .B1(_04716_));
 sg13g2_nand2_1 _22293_ (.Y(_04718_),
    .A(\cpu.ex.r_stmp[14] ),
    .B(net433));
 sg13g2_o21ai_1 _22294_ (.B1(_04718_),
    .Y(_01012_),
    .A1(_04708_),
    .A2(_04717_));
 sg13g2_nor2_1 _22295_ (.A(net630),
    .B(net538),
    .Y(_04719_));
 sg13g2_a21oi_1 _22296_ (.A1(_10200_),
    .A2(_04699_),
    .Y(_04720_),
    .B1(_04719_));
 sg13g2_nand2_1 _22297_ (.Y(_04721_),
    .A(\cpu.ex.r_stmp[15] ),
    .B(net433));
 sg13g2_o21ai_1 _22298_ (.B1(_04721_),
    .Y(_01013_),
    .A1(_04708_),
    .A2(_04720_));
 sg13g2_nor2_1 _22299_ (.A(net601),
    .B(net538),
    .Y(_04722_));
 sg13g2_a21oi_1 _22300_ (.A1(_10589_),
    .A2(net539),
    .Y(_04723_),
    .B1(_04722_));
 sg13g2_nand2_1 _22301_ (.Y(_04724_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net433));
 sg13g2_o21ai_1 _22302_ (.B1(_04724_),
    .Y(_01014_),
    .A1(net432),
    .A2(_04723_));
 sg13g2_nor2_1 _22303_ (.A(_03541_),
    .B(net598),
    .Y(_04725_));
 sg13g2_a21oi_1 _22304_ (.A1(_10524_),
    .A2(net539),
    .Y(_04726_),
    .B1(_04725_));
 sg13g2_nand2_1 _22305_ (.Y(_04727_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net476));
 sg13g2_o21ai_1 _22306_ (.B1(_04727_),
    .Y(_01015_),
    .A1(net432),
    .A2(_04726_));
 sg13g2_nor2_1 _22307_ (.A(net679),
    .B(net598),
    .Y(_04728_));
 sg13g2_a21oi_1 _22308_ (.A1(_10492_),
    .A2(net539),
    .Y(_04729_),
    .B1(_04728_));
 sg13g2_nand2_1 _22309_ (.Y(_04730_),
    .A(\cpu.ex.r_stmp[3] ),
    .B(net476));
 sg13g2_o21ai_1 _22310_ (.B1(_04730_),
    .Y(_01016_),
    .A1(net432),
    .A2(_04729_));
 sg13g2_nor2_1 _22311_ (.A(net599),
    .B(net598),
    .Y(_04731_));
 sg13g2_a21oi_1 _22312_ (.A1(_10644_),
    .A2(net539),
    .Y(_04732_),
    .B1(_04731_));
 sg13g2_nand2_1 _22313_ (.Y(_04733_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(net476));
 sg13g2_o21ai_1 _22314_ (.B1(_04733_),
    .Y(_01017_),
    .A1(net432),
    .A2(_04732_));
 sg13g2_buf_2 _22315_ (.A(net757),
    .X(_04734_));
 sg13g2_mux2_1 _22316_ (.A0(net668),
    .A1(_10622_),
    .S(net538),
    .X(_04735_));
 sg13g2_mux2_1 _22317_ (.A0(_04735_),
    .A1(\cpu.ex.r_stmp[5] ),
    .S(_04706_),
    .X(_01018_));
 sg13g2_nor2_1 _22318_ (.A(_02918_),
    .B(net598),
    .Y(_04736_));
 sg13g2_a21oi_1 _22319_ (.A1(_10354_),
    .A2(net539),
    .Y(_04737_),
    .B1(_04736_));
 sg13g2_nand2_1 _22320_ (.Y(_04738_),
    .A(\cpu.ex.r_stmp[6] ),
    .B(net476));
 sg13g2_o21ai_1 _22321_ (.B1(_04738_),
    .Y(_01019_),
    .A1(net432),
    .A2(_04737_));
 sg13g2_nor2_1 _22322_ (.A(net864),
    .B(net598),
    .Y(_04739_));
 sg13g2_a21oi_1 _22323_ (.A1(_10460_),
    .A2(net539),
    .Y(_04740_),
    .B1(_04739_));
 sg13g2_nand2_1 _22324_ (.Y(_04741_),
    .A(\cpu.ex.r_stmp[7] ),
    .B(net476));
 sg13g2_o21ai_1 _22325_ (.B1(_04741_),
    .Y(_01020_),
    .A1(net432),
    .A2(_04740_));
 sg13g2_nor2_1 _22326_ (.A(_09153_),
    .B(net598),
    .Y(_04742_));
 sg13g2_a21oi_1 _22327_ (.A1(_10449_),
    .A2(net538),
    .Y(_04743_),
    .B1(_04742_));
 sg13g2_nand2_1 _22328_ (.Y(_04744_),
    .A(\cpu.ex.r_stmp[8] ),
    .B(_04705_));
 sg13g2_o21ai_1 _22329_ (.B1(_04744_),
    .Y(_01021_),
    .A1(net432),
    .A2(_04743_));
 sg13g2_nor2_1 _22330_ (.A(_11012_),
    .B(net598),
    .Y(_04745_));
 sg13g2_a21oi_1 _22331_ (.A1(_10310_),
    .A2(_04709_),
    .Y(_04746_),
    .B1(_04745_));
 sg13g2_nand2_1 _22332_ (.Y(_04747_),
    .A(\cpu.ex.r_stmp[9] ),
    .B(net476));
 sg13g2_o21ai_1 _22333_ (.B1(_04747_),
    .Y(_01022_),
    .A1(_04706_),
    .A2(_04746_));
 sg13g2_nor2_1 _22334_ (.A(_08399_),
    .B(_11410_),
    .Y(_04748_));
 sg13g2_buf_1 _22335_ (.A(_04748_),
    .X(_04749_));
 sg13g2_buf_1 _22336_ (.A(_04749_),
    .X(_04750_));
 sg13g2_nand4_1 _22337_ (.B(_09146_),
    .C(net1132),
    .A(_11784_),
    .Y(_04751_),
    .D(_09769_));
 sg13g2_buf_1 _22338_ (.A(_04751_),
    .X(_04752_));
 sg13g2_buf_1 _22339_ (.A(_04752_),
    .X(_04753_));
 sg13g2_nand2_1 _22340_ (.Y(_04754_),
    .A(\cpu.dcache.r_data[1][0] ),
    .B(net484));
 sg13g2_buf_1 _22341_ (.A(net615),
    .X(_04755_));
 sg13g2_a22oi_1 _22342_ (.Y(_04756_),
    .B1(_04755_),
    .B2(\cpu.dcache.r_data[5][0] ),
    .A2(net482),
    .A1(\cpu.dcache.r_data[3][0] ));
 sg13g2_buf_1 _22343_ (.A(net632),
    .X(_04757_));
 sg13g2_buf_1 _22344_ (.A(net536),
    .X(_04758_));
 sg13g2_a22oi_1 _22345_ (.Y(_04759_),
    .B1(net483),
    .B2(\cpu.dcache.r_data[2][0] ),
    .A2(net475),
    .A1(\cpu.dcache.r_data[0][0] ));
 sg13g2_mux2_1 _22346_ (.A0(\cpu.dcache.r_data[4][0] ),
    .A1(\cpu.dcache.r_data[6][0] ),
    .S(net575),
    .X(_04760_));
 sg13g2_a22oi_1 _22347_ (.Y(_04761_),
    .B1(_04760_),
    .B2(net782),
    .A2(net693),
    .A1(\cpu.dcache.r_data[7][0] ));
 sg13g2_nand2b_1 _22348_ (.Y(_04762_),
    .B(net779),
    .A_N(_04761_));
 sg13g2_nand4_1 _22349_ (.B(_04756_),
    .C(_04759_),
    .A(_04754_),
    .Y(_04763_),
    .D(_04762_));
 sg13g2_nand2_1 _22350_ (.Y(_04764_),
    .A(\cpu.dcache.r_data[1][16] ),
    .B(net484));
 sg13g2_a22oi_1 _22351_ (.Y(_04765_),
    .B1(net537),
    .B2(\cpu.dcache.r_data[5][16] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[3][16] ));
 sg13g2_buf_1 _22352_ (.A(net563),
    .X(_04766_));
 sg13g2_a22oi_1 _22353_ (.Y(_04767_),
    .B1(net474),
    .B2(\cpu.dcache.r_data[2][16] ),
    .A2(net536),
    .A1(\cpu.dcache.r_data[0][16] ));
 sg13g2_mux2_1 _22354_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(\cpu.dcache.r_data[6][16] ),
    .S(net575),
    .X(_04768_));
 sg13g2_a22oi_1 _22355_ (.Y(_04769_),
    .B1(_04768_),
    .B2(net782),
    .A2(net693),
    .A1(\cpu.dcache.r_data[7][16] ));
 sg13g2_nand2b_1 _22356_ (.Y(_04770_),
    .B(net779),
    .A_N(_04769_));
 sg13g2_nand4_1 _22357_ (.B(_04765_),
    .C(_04767_),
    .A(_04764_),
    .Y(_04771_),
    .D(_04770_));
 sg13g2_buf_1 _22358_ (.A(_04771_),
    .X(_04772_));
 sg13g2_mux2_1 _22359_ (.A0(_04763_),
    .A1(_04772_),
    .S(net609),
    .X(_04773_));
 sg13g2_nand2_1 _22360_ (.Y(_04774_),
    .A(net1132),
    .B(_08322_));
 sg13g2_or2_1 _22361_ (.X(_04775_),
    .B(_04774_),
    .A(_08333_));
 sg13g2_buf_1 _22362_ (.A(_04775_),
    .X(_04776_));
 sg13g2_buf_1 _22363_ (.A(net667),
    .X(_04777_));
 sg13g2_buf_1 _22364_ (.A(_11898_),
    .X(_04778_));
 sg13g2_mux2_1 _22365_ (.A0(\cpu.dcache.r_data[5][24] ),
    .A1(\cpu.dcache.r_data[7][24] ),
    .S(_09165_),
    .X(_04779_));
 sg13g2_a22oi_1 _22366_ (.Y(_04780_),
    .B1(_04779_),
    .B2(net574),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][24] ));
 sg13g2_nor2_1 _22367_ (.A(net758),
    .B(_04780_),
    .Y(_04781_));
 sg13g2_buf_1 _22368_ (.A(_09364_),
    .X(_04782_));
 sg13g2_a22oi_1 _22369_ (.Y(_04783_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][24] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][24] ));
 sg13g2_o21ai_1 _22370_ (.B1(_04783_),
    .Y(_04784_),
    .A1(_00295_),
    .A2(net535));
 sg13g2_a221oi_1 _22371_ (.B2(\cpu.dcache.r_data[2][24] ),
    .C1(_04784_),
    .B1(net474),
    .A1(\cpu.dcache.r_data[3][24] ),
    .Y(_04785_),
    .A2(net562));
 sg13g2_nor2b_1 _22372_ (.A(_04781_),
    .B_N(_04785_),
    .Y(_04786_));
 sg13g2_buf_1 _22373_ (.A(net575),
    .X(_04787_));
 sg13g2_mux2_1 _22374_ (.A0(\cpu.dcache.r_data[4][8] ),
    .A1(\cpu.dcache.r_data[6][8] ),
    .S(net473),
    .X(_04788_));
 sg13g2_a22oi_1 _22375_ (.Y(_04789_),
    .B1(_04788_),
    .B2(net669),
    .A2(net693),
    .A1(\cpu.dcache.r_data[7][8] ));
 sg13g2_a22oi_1 _22376_ (.Y(_04790_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][8] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][8] ));
 sg13g2_o21ai_1 _22377_ (.B1(_04790_),
    .Y(_04791_),
    .A1(_00296_),
    .A2(net535));
 sg13g2_a221oi_1 _22378_ (.B2(\cpu.dcache.r_data[5][8] ),
    .C1(_04791_),
    .B1(net537),
    .A1(\cpu.dcache.r_data[2][8] ),
    .Y(_04792_),
    .A2(net483));
 sg13g2_o21ai_1 _22379_ (.B1(_04792_),
    .Y(_04793_),
    .A1(net680),
    .A2(_04789_));
 sg13g2_nand2_1 _22380_ (.Y(_04794_),
    .A(net780),
    .B(_04793_));
 sg13g2_o21ai_1 _22381_ (.B1(_04794_),
    .Y(_04795_),
    .A1(net972),
    .A2(_04786_));
 sg13g2_nor2_2 _22382_ (.A(net780),
    .B(_11898_),
    .Y(_04796_));
 sg13g2_a22oi_1 _22383_ (.Y(_04797_),
    .B1(_04772_),
    .B2(_04796_),
    .A2(_04763_),
    .A1(_11898_));
 sg13g2_nand2_1 _22384_ (.Y(_04798_),
    .A(net667),
    .B(_04797_));
 sg13g2_o21ai_1 _22385_ (.B1(_04798_),
    .Y(_04799_),
    .A1(_04777_),
    .A2(_04795_));
 sg13g2_nand2_1 _22386_ (.Y(_04800_),
    .A(_04799_),
    .B(_04753_));
 sg13g2_o21ai_1 _22387_ (.B1(_04800_),
    .Y(_04801_),
    .A1(net597),
    .A2(_04773_));
 sg13g2_nand2_1 _22388_ (.Y(_04802_),
    .A(_09153_),
    .B(net1057));
 sg13g2_nor2_1 _22389_ (.A(net1058),
    .B(_04802_),
    .Y(_04803_));
 sg13g2_buf_2 _22390_ (.A(_04803_),
    .X(_04804_));
 sg13g2_nand2_1 _22391_ (.Y(_04805_),
    .A(net714),
    .B(_09900_));
 sg13g2_buf_1 _22392_ (.A(_04805_),
    .X(_04806_));
 sg13g2_nor3_1 _22393_ (.A(net1120),
    .B(net781),
    .C(net534),
    .Y(_04807_));
 sg13g2_buf_2 _22394_ (.A(_04807_),
    .X(_04808_));
 sg13g2_nand2_1 _22395_ (.Y(_04809_),
    .A(net910),
    .B(net634));
 sg13g2_nor3_1 _22396_ (.A(net782),
    .B(_09740_),
    .C(_04809_),
    .Y(_04810_));
 sg13g2_buf_2 _22397_ (.A(_04810_),
    .X(_04811_));
 sg13g2_buf_2 _22398_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04812_));
 sg13g2_buf_2 _22399_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04813_));
 sg13g2_mux2_1 _22400_ (.A0(_04812_),
    .A1(_04813_),
    .S(net673),
    .X(_04814_));
 sg13g2_a22oi_1 _22401_ (.Y(_04815_),
    .B1(_04811_),
    .B2(_04814_),
    .A2(_04808_),
    .A1(_09107_));
 sg13g2_buf_2 _22402_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04816_));
 sg13g2_buf_1 _22403_ (.A(_09740_),
    .X(_04817_));
 sg13g2_nor3_2 _22404_ (.A(net971),
    .B(net781),
    .C(net534),
    .Y(_04818_));
 sg13g2_nand2_2 _22405_ (.Y(_04819_),
    .A(_09142_),
    .B(net1128));
 sg13g2_nor2_1 _22406_ (.A(net781),
    .B(_04819_),
    .Y(_04820_));
 sg13g2_buf_1 _22407_ (.A(_04820_),
    .X(_04821_));
 sg13g2_and2_1 _22408_ (.A(net1016),
    .B(net472),
    .X(_04822_));
 sg13g2_buf_1 _22409_ (.A(_04822_),
    .X(_04823_));
 sg13g2_buf_2 _22410_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04824_));
 sg13g2_a22oi_1 _22411_ (.Y(_04825_),
    .B1(_04823_),
    .B2(_04824_),
    .A2(_04818_),
    .A1(_04816_));
 sg13g2_buf_2 _22412_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04826_));
 sg13g2_nand2_2 _22413_ (.Y(_04827_),
    .A(net915),
    .B(net615));
 sg13g2_nor2_1 _22414_ (.A(_09741_),
    .B(_04827_),
    .Y(_04828_));
 sg13g2_nor3_2 _22415_ (.A(net1120),
    .B(net1128),
    .C(_09400_),
    .Y(_04829_));
 sg13g2_buf_2 _22416_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04830_));
 sg13g2_a22oi_1 _22417_ (.Y(_04831_),
    .B1(_04829_),
    .B2(_04830_),
    .A2(_04828_),
    .A1(_04826_));
 sg13g2_o21ai_1 _22418_ (.B1(_09740_),
    .Y(_04832_),
    .A1(net1128),
    .A2(_09903_));
 sg13g2_nor2_1 _22419_ (.A(net1120),
    .B(net713),
    .Y(_04833_));
 sg13g2_and2_1 _22420_ (.A(net1120),
    .B(_09164_),
    .X(_04834_));
 sg13g2_a21oi_1 _22421_ (.A1(_04832_),
    .A2(_04833_),
    .Y(_04835_),
    .B1(_04834_));
 sg13g2_nand2_1 _22422_ (.Y(_04836_),
    .A(net903),
    .B(_09741_));
 sg13g2_o21ai_1 _22423_ (.B1(_04836_),
    .Y(_04837_),
    .A1(net679),
    .A2(_09741_));
 sg13g2_nand2_1 _22424_ (.Y(_04838_),
    .A(net910),
    .B(_09740_));
 sg13g2_o21ai_1 _22425_ (.B1(_04836_),
    .Y(_04839_),
    .A1(_04806_),
    .A2(_04838_));
 sg13g2_a22oi_1 _22426_ (.Y(_04840_),
    .B1(_09741_),
    .B2(_04833_),
    .A2(net634),
    .A1(net903));
 sg13g2_nor2_1 _22427_ (.A(_09900_),
    .B(_04840_),
    .Y(_04841_));
 sg13g2_a221oi_1 _22428_ (.B2(net1120),
    .C1(_04841_),
    .B1(_04839_),
    .A1(net633),
    .Y(_04842_),
    .A2(_04837_));
 sg13g2_o21ai_1 _22429_ (.B1(_04842_),
    .Y(_04843_),
    .A1(net633),
    .A2(_04835_));
 sg13g2_buf_2 _22430_ (.A(_04843_),
    .X(_04844_));
 sg13g2_nor2_1 _22431_ (.A(net903),
    .B(net789),
    .Y(_04845_));
 sg13g2_and2_1 _22432_ (.A(_09144_),
    .B(_04845_),
    .X(_04846_));
 sg13g2_buf_2 _22433_ (.A(_04846_),
    .X(_04847_));
 sg13g2_nor2b_1 _22434_ (.A(_11833_),
    .B_N(_04847_),
    .Y(_04848_));
 sg13g2_buf_1 _22435_ (.A(_04848_),
    .X(_04849_));
 sg13g2_a21oi_1 _22436_ (.A1(_09107_),
    .A2(_04844_),
    .Y(_04850_),
    .B1(net390));
 sg13g2_nand2b_1 _22437_ (.Y(_04851_),
    .B(\cpu.gpio.r_enable_in[0] ),
    .A_N(_04850_));
 sg13g2_nand4_1 _22438_ (.B(_04825_),
    .C(_04831_),
    .A(_04815_),
    .Y(_04852_),
    .D(_04851_));
 sg13g2_buf_1 _22439_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04853_));
 sg13g2_nor2_1 _22440_ (.A(_09142_),
    .B(_09900_),
    .Y(_04854_));
 sg13g2_nand2_2 _22441_ (.Y(_04855_),
    .A(_04845_),
    .B(_04854_));
 sg13g2_nor2_1 _22442_ (.A(_04817_),
    .B(_04855_),
    .Y(_04856_));
 sg13g2_buf_2 _22443_ (.A(_04856_),
    .X(_04857_));
 sg13g2_nand2_1 _22444_ (.Y(_04858_),
    .A(_09164_),
    .B(_04836_));
 sg13g2_nand2_1 _22445_ (.Y(_04859_),
    .A(net789),
    .B(_09086_));
 sg13g2_o21ai_1 _22446_ (.B1(_04859_),
    .Y(_04860_),
    .A1(net633),
    .A2(_04838_));
 sg13g2_nor2_1 _22447_ (.A(_09333_),
    .B(_09511_),
    .Y(_04861_));
 sg13g2_nor2_1 _22448_ (.A(_09143_),
    .B(_04861_),
    .Y(_04862_));
 sg13g2_a221oi_1 _22449_ (.B2(net1052),
    .C1(_04862_),
    .B1(_04860_),
    .A1(_09537_),
    .Y(_04863_),
    .A2(_04858_));
 sg13g2_nor2_1 _22450_ (.A(net1120),
    .B(_04855_),
    .Y(_04864_));
 sg13g2_nor3_1 _22451_ (.A(_04829_),
    .B(_04863_),
    .C(_04864_),
    .Y(_04865_));
 sg13g2_buf_2 _22452_ (.A(_04865_),
    .X(_04866_));
 sg13g2_nor2_1 _22453_ (.A(net1052),
    .B(_09400_),
    .Y(_04867_));
 sg13g2_buf_1 _22454_ (.A(_04867_),
    .X(_04868_));
 sg13g2_nand2b_1 _22455_ (.Y(_04869_),
    .B(_04847_),
    .A_N(_00205_));
 sg13g2_o21ai_1 _22456_ (.B1(_04869_),
    .Y(_04870_),
    .A1(_00298_),
    .A2(_04855_));
 sg13g2_a21oi_1 _22457_ (.A1(\cpu.spi.r_mode[1][0] ),
    .A2(_04868_),
    .Y(_04871_),
    .B1(_04870_));
 sg13g2_a22oi_1 _22458_ (.Y(_04872_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net507),
    .A2(_09085_),
    .A1(_09121_));
 sg13g2_nand2b_1 _22459_ (.Y(_04873_),
    .B(net915),
    .A_N(_04872_));
 sg13g2_nand3_1 _22460_ (.B(net679),
    .C(\cpu.spi.r_ready ),
    .A(net901),
    .Y(_04874_));
 sg13g2_a21oi_1 _22461_ (.A1(_04873_),
    .A2(_04874_),
    .Y(_04875_),
    .B1(net669));
 sg13g2_nand3_1 _22462_ (.B(_09740_),
    .C(net631),
    .A(net1052),
    .Y(_04876_));
 sg13g2_buf_2 _22463_ (.A(_04876_),
    .X(_04877_));
 sg13g2_nand3_1 _22464_ (.B(\cpu.spi.r_mode[2][0] ),
    .C(_04847_),
    .A(net1016),
    .Y(_04878_));
 sg13g2_o21ai_1 _22465_ (.B1(_04878_),
    .Y(_04879_),
    .A1(_00297_),
    .A2(_04877_));
 sg13g2_nor2_1 _22466_ (.A(_04875_),
    .B(_04879_),
    .Y(_04880_));
 sg13g2_o21ai_1 _22467_ (.B1(_04880_),
    .Y(_04881_),
    .A1(net874),
    .A2(_04871_));
 sg13g2_a221oi_1 _22468_ (.B2(_09189_),
    .C1(_04881_),
    .B1(_04866_),
    .A1(_04853_),
    .Y(_04882_),
    .A2(_04857_));
 sg13g2_and2_1 _22469_ (.A(net1058),
    .B(_09908_),
    .X(_04883_));
 sg13g2_buf_1 _22470_ (.A(_04883_),
    .X(_04884_));
 sg13g2_buf_1 _22471_ (.A(net797),
    .X(_04885_));
 sg13g2_a22oi_1 _22472_ (.Y(_04886_),
    .B1(net559),
    .B2(\cpu.intr.r_timer_reload[16] ),
    .A2(net442),
    .A1(_09933_));
 sg13g2_a221oi_1 _22473_ (.B2(_10052_),
    .C1(net797),
    .B1(net503),
    .A1(\cpu.intr.r_clock_cmp[0] ),
    .Y(_04887_),
    .A2(net561));
 sg13g2_a21o_1 _22474_ (.A2(_04886_),
    .A1(net666),
    .B1(_04887_),
    .X(_04888_));
 sg13g2_nor2_1 _22475_ (.A(net781),
    .B(net534),
    .Y(_04889_));
 sg13g2_buf_1 _22476_ (.A(_04889_),
    .X(_04890_));
 sg13g2_buf_1 _22477_ (.A(_04890_),
    .X(_04891_));
 sg13g2_nand2_1 _22478_ (.Y(_04892_),
    .A(_09537_),
    .B(net1128));
 sg13g2_buf_1 _22479_ (.A(_04892_),
    .X(_04893_));
 sg13g2_nor3_1 _22480_ (.A(net910),
    .B(net634),
    .C(net595),
    .Y(_04894_));
 sg13g2_buf_1 _22481_ (.A(_04894_),
    .X(_04895_));
 sg13g2_buf_1 _22482_ (.A(_04895_),
    .X(_04896_));
 sg13g2_buf_1 _22483_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04897_));
 sg13g2_nor3_1 _22484_ (.A(net797),
    .B(_00266_),
    .C(_09400_),
    .Y(_04898_));
 sg13g2_a221oi_1 _22485_ (.B2(_04897_),
    .C1(_04898_),
    .B1(net431),
    .A1(_09129_),
    .Y(_04899_),
    .A2(net389));
 sg13g2_nor2_1 _22486_ (.A(_09900_),
    .B(_09395_),
    .Y(_04900_));
 sg13g2_buf_1 _22487_ (.A(_04900_),
    .X(_04901_));
 sg13g2_nor2_1 _22488_ (.A(net915),
    .B(_09906_),
    .Y(_04902_));
 sg13g2_a22oi_1 _22489_ (.Y(_04903_),
    .B1(_04902_),
    .B2(\cpu.intr.r_timer_reload[0] ),
    .A2(_04901_),
    .A1(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_a21oi_1 _22490_ (.A1(net534),
    .A2(net595),
    .Y(_04904_),
    .B1(net634));
 sg13g2_nor2_1 _22491_ (.A(net779),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_buf_1 _22492_ (.A(_04905_),
    .X(_04906_));
 sg13g2_nor2_1 _22493_ (.A(net781),
    .B(net595),
    .Y(_04907_));
 sg13g2_buf_1 _22494_ (.A(_04907_),
    .X(_04908_));
 sg13g2_buf_1 _22495_ (.A(_04908_),
    .X(_04909_));
 sg13g2_a21o_1 _22496_ (.A2(net388),
    .A1(_09129_),
    .B1(net430),
    .X(_04910_));
 sg13g2_o21ai_1 _22497_ (.B1(_04910_),
    .Y(_04911_),
    .A1(_09127_),
    .A2(_09128_));
 sg13g2_nand4_1 _22498_ (.B(_04899_),
    .C(_04903_),
    .A(_04888_),
    .Y(_04912_),
    .D(_04911_));
 sg13g2_nand2_1 _22499_ (.Y(_04913_),
    .A(_04802_),
    .B(_09910_));
 sg13g2_buf_1 _22500_ (.A(_04913_),
    .X(_04914_));
 sg13g2_o21ai_1 _22501_ (.B1(net758),
    .Y(_04915_),
    .A1(net706),
    .A2(_09641_));
 sg13g2_buf_2 _22502_ (.A(_04915_),
    .X(_04916_));
 sg13g2_nor2_1 _22503_ (.A(_04809_),
    .B(net595),
    .Y(_04917_));
 sg13g2_buf_2 _22504_ (.A(_04917_),
    .X(_04918_));
 sg13g2_a22oi_1 _22505_ (.Y(_04919_),
    .B1(_04918_),
    .B2(\cpu.uart.r_div_value[8] ),
    .A2(_04847_),
    .A1(\cpu.uart.r_div_value[0] ));
 sg13g2_a22oi_1 _22506_ (.Y(_04920_),
    .B1(net472),
    .B2(\cpu.uart.r_x_invert ),
    .A2(_04890_),
    .A1(_09127_));
 sg13g2_nand2_1 _22507_ (.Y(_04921_),
    .A(_04919_),
    .B(_04920_));
 sg13g2_a21oi_1 _22508_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04916_),
    .Y(_04922_),
    .B1(_04921_));
 sg13g2_o21ai_1 _22509_ (.B1(_08321_),
    .Y(_04923_),
    .A1(net533),
    .A2(_04922_));
 sg13g2_a21oi_1 _22510_ (.A1(_04884_),
    .A2(_04912_),
    .Y(_04924_),
    .B1(_04923_));
 sg13g2_o21ai_1 _22511_ (.B1(_04924_),
    .Y(_04925_),
    .A1(net800),
    .A2(_04882_));
 sg13g2_a21oi_1 _22512_ (.A1(_04804_),
    .A2(_04852_),
    .Y(_04926_),
    .B1(_04925_));
 sg13g2_a21oi_1 _22513_ (.A1(net902),
    .A2(_04801_),
    .Y(_04927_),
    .B1(_04926_));
 sg13g2_nand2_1 _22514_ (.Y(_04928_),
    .A(net73),
    .B(_04927_));
 sg13g2_o21ai_1 _22515_ (.B1(_04928_),
    .Y(_04929_),
    .A1(_03552_),
    .A2(_04750_));
 sg13g2_nand2_1 _22516_ (.Y(_04930_),
    .A(_11384_),
    .B(_03972_));
 sg13g2_nor2b_1 _22517_ (.A(_04930_),
    .B_N(_11371_),
    .Y(_04931_));
 sg13g2_nand3_1 _22518_ (.B(_03956_),
    .C(_04191_),
    .A(_03955_),
    .Y(_04932_));
 sg13g2_o21ai_1 _22519_ (.B1(net223),
    .Y(_04933_),
    .A1(net978),
    .A2(_04932_));
 sg13g2_or2_1 _22520_ (.X(_04934_),
    .B(_03961_),
    .A(net1121));
 sg13g2_o21ai_1 _22521_ (.B1(_04934_),
    .Y(_04935_),
    .A1(net223),
    .A2(_04932_));
 sg13g2_a22oi_1 _22522_ (.Y(_04936_),
    .B1(_04935_),
    .B2(_09835_),
    .A2(_04933_),
    .A1(_03559_));
 sg13g2_o21ai_1 _22523_ (.B1(net166),
    .Y(_04937_),
    .A1(_04233_),
    .A2(_11600_));
 sg13g2_nor2_1 _22524_ (.A(_04936_),
    .B(_04937_),
    .Y(_04938_));
 sg13g2_a21oi_1 _22525_ (.A1(_03842_),
    .A2(_03873_),
    .Y(_04939_),
    .B1(_04340_));
 sg13g2_a22oi_1 _22526_ (.Y(_04940_),
    .B1(_04214_),
    .B2(_03899_),
    .A2(_03901_),
    .A1(net163));
 sg13g2_nor3_1 _22527_ (.A(net236),
    .B(net183),
    .C(_04412_),
    .Y(_04941_));
 sg13g2_a22oi_1 _22528_ (.Y(_04942_),
    .B1(_04045_),
    .B2(_04003_),
    .A2(_04060_),
    .A1(_03909_));
 sg13g2_a21oi_1 _22529_ (.A1(_03865_),
    .A2(net182),
    .Y(_04943_),
    .B1(_04487_));
 sg13g2_nand2_1 _22530_ (.Y(_04944_),
    .A(_04942_),
    .B(_04943_));
 sg13g2_nor2_1 _22531_ (.A(_04941_),
    .B(_04944_),
    .Y(_04945_));
 sg13g2_nand4_1 _22532_ (.B(_04939_),
    .C(_04940_),
    .A(_04659_),
    .Y(_04946_),
    .D(_04945_));
 sg13g2_mux2_1 _22533_ (.A0(net136),
    .A1(_03897_),
    .S(net234),
    .X(_04947_));
 sg13g2_a22oi_1 _22534_ (.Y(_04948_),
    .B1(_04947_),
    .B2(_03559_),
    .A2(_03922_),
    .A1(_11030_));
 sg13g2_nor2_1 _22535_ (.A(_03870_),
    .B(_04948_),
    .Y(_04949_));
 sg13g2_o21ai_1 _22536_ (.B1(_03926_),
    .Y(_04950_),
    .A1(_04946_),
    .A2(_04949_));
 sg13g2_o21ai_1 _22537_ (.B1(_04950_),
    .Y(_04951_),
    .A1(_10604_),
    .A2(net181));
 sg13g2_o21ai_1 _22538_ (.B1(_04951_),
    .Y(_04952_),
    .A1(net158),
    .A2(net200));
 sg13g2_nor2_1 _22539_ (.A(net85),
    .B(_04930_),
    .Y(_04953_));
 sg13g2_nor3_1 _22540_ (.A(_11373_),
    .B(net618),
    .C(net166),
    .Y(_04954_));
 sg13g2_a21o_1 _22541_ (.A2(_04953_),
    .A1(_11371_),
    .B1(_04954_),
    .X(_04955_));
 sg13g2_a221oi_1 _22542_ (.B2(_04952_),
    .C1(_04955_),
    .B1(_04938_),
    .A1(net28),
    .Y(_04956_),
    .A2(_04931_));
 sg13g2_buf_1 _22543_ (.A(_04956_),
    .X(_04957_));
 sg13g2_buf_1 _22544_ (.A(_11399_),
    .X(_04958_));
 sg13g2_nand2_1 _22545_ (.Y(_04959_),
    .A(_03834_),
    .B(net665));
 sg13g2_mux2_1 _22546_ (.A0(_04957_),
    .A1(net982),
    .S(_04959_),
    .X(_04960_));
 sg13g2_buf_1 _22547_ (.A(net86),
    .X(_04961_));
 sg13g2_mux2_1 _22548_ (.A0(_04929_),
    .A1(_04960_),
    .S(net72),
    .X(_01023_));
 sg13g2_nand3_1 _22549_ (.B(_04685_),
    .C(_04686_),
    .A(_04958_),
    .Y(_04962_));
 sg13g2_a21oi_1 _22550_ (.A1(_00238_),
    .A2(_11397_),
    .Y(_04963_),
    .B1(_11784_));
 sg13g2_buf_1 _22551_ (.A(_04963_),
    .X(_04964_));
 sg13g2_buf_1 _22552_ (.A(net740),
    .X(_04965_));
 sg13g2_nand2_1 _22553_ (.Y(_04966_),
    .A(_03834_),
    .B(_11405_));
 sg13g2_buf_1 _22554_ (.A(_04966_),
    .X(_04967_));
 sg13g2_a21oi_1 _22555_ (.A1(net664),
    .A2(_04690_),
    .Y(_04968_),
    .B1(_04967_));
 sg13g2_nand2_2 _22556_ (.Y(_04969_),
    .A(net352),
    .B(_11405_));
 sg13g2_nor2_1 _22557_ (.A(_11405_),
    .B(_04749_),
    .Y(_04970_));
 sg13g2_buf_1 _22558_ (.A(_04970_),
    .X(_04971_));
 sg13g2_nor3_1 _22559_ (.A(net902),
    .B(_09910_),
    .C(_04906_),
    .Y(_04972_));
 sg13g2_buf_2 _22560_ (.A(_04972_),
    .X(_04973_));
 sg13g2_buf_1 _22561_ (.A(_04902_),
    .X(_04974_));
 sg13g2_nor2_1 _22562_ (.A(net1128),
    .B(_09395_),
    .Y(_04975_));
 sg13g2_buf_1 _22563_ (.A(_04975_),
    .X(_04976_));
 sg13g2_buf_1 _22564_ (.A(_04976_),
    .X(_04977_));
 sg13g2_a22oi_1 _22565_ (.Y(_04978_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net429),
    .A1(\cpu.intr.r_timer_reload[10] ));
 sg13g2_buf_1 _22566_ (.A(_04901_),
    .X(_04979_));
 sg13g2_a22oi_1 _22567_ (.Y(_04980_),
    .B1(net593),
    .B2(\cpu.intr.r_clock_cmp[26] ),
    .A2(net447),
    .A1(_10101_));
 sg13g2_buf_1 _22568_ (.A(_04868_),
    .X(_04981_));
 sg13g2_buf_1 _22569_ (.A(_04896_),
    .X(_04982_));
 sg13g2_buf_2 _22570_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_04983_));
 sg13g2_a22oi_1 _22571_ (.Y(_04984_),
    .B1(net387),
    .B2(_04983_),
    .A2(net532),
    .A1(\cpu.intr.r_timer_count[10] ));
 sg13g2_nand3_1 _22572_ (.B(_04980_),
    .C(_04984_),
    .A(_04978_),
    .Y(_04985_));
 sg13g2_a22oi_1 _22573_ (.Y(_04986_),
    .B1(net559),
    .B2(\cpu.dcache.r_data[7][26] ),
    .A2(net503),
    .A1(\cpu.dcache.r_data[4][26] ));
 sg13g2_a22oi_1 _22574_ (.Y(_04987_),
    .B1(_02900_),
    .B2(\cpu.dcache.r_data[5][26] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[2][26] ));
 sg13g2_inv_1 _22575_ (.Y(_04988_),
    .A(_00310_));
 sg13g2_a22oi_1 _22576_ (.Y(_04989_),
    .B1(_02904_),
    .B2(\cpu.dcache.r_data[6][26] ),
    .A2(net475),
    .A1(_04988_));
 sg13g2_a22oi_1 _22577_ (.Y(_04990_),
    .B1(_02889_),
    .B2(\cpu.dcache.r_data[1][26] ),
    .A2(net482),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_nand4_1 _22578_ (.B(_04987_),
    .C(_04989_),
    .A(_04986_),
    .Y(_04991_),
    .D(_04990_));
 sg13g2_mux2_1 _22579_ (.A0(\cpu.dcache.r_data[1][10] ),
    .A1(\cpu.dcache.r_data[3][10] ),
    .S(net507),
    .X(_04992_));
 sg13g2_a22oi_1 _22580_ (.Y(_04993_),
    .B1(_04992_),
    .B2(net574),
    .A2(net706),
    .A1(\cpu.dcache.r_data[2][10] ));
 sg13g2_inv_1 _22581_ (.Y(_04994_),
    .A(_00091_));
 sg13g2_mux2_1 _22582_ (.A0(\cpu.dcache.r_data[5][10] ),
    .A1(\cpu.dcache.r_data[7][10] ),
    .S(net473),
    .X(_04995_));
 sg13g2_a22oi_1 _22583_ (.Y(_04996_),
    .B1(_04995_),
    .B2(net574),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][10] ));
 sg13g2_nor2_1 _22584_ (.A(net680),
    .B(_04996_),
    .Y(_04997_));
 sg13g2_a221oi_1 _22585_ (.B2(\cpu.dcache.r_data[6][10] ),
    .C1(_04997_),
    .B1(_02904_),
    .A1(_04994_),
    .Y(_04998_),
    .A2(net475));
 sg13g2_o21ai_1 _22586_ (.B1(_04998_),
    .Y(_04999_),
    .A1(_09310_),
    .A2(_04993_));
 sg13g2_mux2_1 _22587_ (.A0(_04991_),
    .A1(_04999_),
    .S(net672),
    .X(_05000_));
 sg13g2_nor3_2 _22588_ (.A(net1133),
    .B(_08331_),
    .C(_04774_),
    .Y(_05001_));
 sg13g2_buf_1 _22589_ (.A(_05001_),
    .X(_05002_));
 sg13g2_a22oi_1 _22590_ (.Y(_05003_),
    .B1(_05000_),
    .B2(net663),
    .A2(_04985_),
    .A1(_04973_));
 sg13g2_nor2_1 _22591_ (.A(net692),
    .B(net388),
    .Y(_05004_));
 sg13g2_mux2_1 _22592_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(\cpu.intr.r_timer_reload[23] ),
    .S(net1052),
    .X(_05005_));
 sg13g2_mux2_1 _22593_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(\cpu.intr.r_clock_cmp[23] ),
    .S(net1052),
    .X(_05006_));
 sg13g2_a22oi_1 _22594_ (.Y(_05007_),
    .B1(_05006_),
    .B2(net700),
    .A2(_05005_),
    .A1(net697));
 sg13g2_buf_2 _22595_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05008_));
 sg13g2_mux2_1 _22596_ (.A0(\cpu.intr.r_timer_count[7] ),
    .A1(_09930_),
    .S(net1052),
    .X(_05009_));
 sg13g2_a22oi_1 _22597_ (.Y(_05010_),
    .B1(_05009_),
    .B2(net560),
    .A2(_04895_),
    .A1(_05008_));
 sg13g2_nand2_1 _22598_ (.Y(_05011_),
    .A(_10083_),
    .B(_10043_));
 sg13g2_nand3_1 _22599_ (.B(_05010_),
    .C(_05011_),
    .A(_05007_),
    .Y(_05012_));
 sg13g2_inv_1 _22600_ (.Y(_05013_),
    .A(_00144_));
 sg13g2_nand2_1 _22601_ (.Y(_05014_),
    .A(net1016),
    .B(_04821_));
 sg13g2_buf_1 _22602_ (.A(_05014_),
    .X(_05015_));
 sg13g2_nor2_1 _22603_ (.A(_00143_),
    .B(net386),
    .Y(_05016_));
 sg13g2_a221oi_1 _22604_ (.B2(_05013_),
    .C1(_05016_),
    .B1(_04818_),
    .A1(_09109_),
    .Y(_05017_),
    .A2(_04808_));
 sg13g2_buf_1 _22605_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05018_));
 sg13g2_nand2_1 _22606_ (.Y(_05019_),
    .A(_09900_),
    .B(_05018_));
 sg13g2_o21ai_1 _22607_ (.B1(_05019_),
    .Y(_05020_),
    .A1(_09900_),
    .A2(_00142_));
 sg13g2_a22oi_1 _22608_ (.Y(_05021_),
    .B1(_05020_),
    .B2(_04811_),
    .A2(_04864_),
    .A1(_09095_));
 sg13g2_nand2_1 _22609_ (.Y(_05022_),
    .A(net1016),
    .B(_04908_));
 sg13g2_nor2_1 _22610_ (.A(_00145_),
    .B(_05022_),
    .Y(_05023_));
 sg13g2_a21oi_1 _22611_ (.A1(_09108_),
    .A2(net390),
    .Y(_05024_),
    .B1(_05023_));
 sg13g2_and2_1 _22612_ (.A(_09108_),
    .B(_09109_),
    .X(_05025_));
 sg13g2_inv_1 _22613_ (.Y(_05026_),
    .A(_00146_));
 sg13g2_a22oi_1 _22614_ (.Y(_05027_),
    .B1(_04976_),
    .B2(net11),
    .A2(_04901_),
    .A1(_05026_));
 sg13g2_a22oi_1 _22615_ (.Y(_05028_),
    .B1(_04895_),
    .B2(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A2(_10043_),
    .A1(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_a21oi_1 _22616_ (.A1(_09095_),
    .A2(_04908_),
    .Y(_05029_),
    .B1(net472));
 sg13g2_nand2b_1 _22617_ (.Y(_05030_),
    .B(_09096_),
    .A_N(_05029_));
 sg13g2_nand3_1 _22618_ (.B(_05028_),
    .C(_05030_),
    .A(_05027_),
    .Y(_05031_));
 sg13g2_a22oi_1 _22619_ (.Y(_05032_),
    .B1(_05031_),
    .B2(net971),
    .A2(_04844_),
    .A1(_05025_));
 sg13g2_nand4_1 _22620_ (.B(_05021_),
    .C(_05024_),
    .A(_05017_),
    .Y(_05033_),
    .D(_05032_));
 sg13g2_buf_1 _22621_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05034_));
 sg13g2_buf_1 _22622_ (.A(_04864_),
    .X(_05035_));
 sg13g2_inv_1 _22623_ (.Y(_05036_),
    .A(_00141_));
 sg13g2_nor2_1 _22624_ (.A(net679),
    .B(_04819_),
    .Y(_05037_));
 sg13g2_buf_2 _22625_ (.A(_05037_),
    .X(_05038_));
 sg13g2_nand2_1 _22626_ (.Y(_05039_),
    .A(\cpu.spi.r_timeout[7] ),
    .B(_05038_));
 sg13g2_o21ai_1 _22627_ (.B1(_05039_),
    .Y(_05040_),
    .A1(_00140_),
    .A2(_04877_));
 sg13g2_a221oi_1 _22628_ (.B2(_05036_),
    .C1(_05040_),
    .B1(net428),
    .A1(_05034_),
    .Y(_05041_),
    .A2(_04857_));
 sg13g2_nand2b_1 _22629_ (.Y(_05042_),
    .B(_04866_),
    .A_N(_00202_));
 sg13g2_a21oi_1 _22630_ (.A1(_05041_),
    .A2(_05042_),
    .Y(_05043_),
    .B1(net800));
 sg13g2_a221oi_1 _22631_ (.B2(_04804_),
    .C1(_05043_),
    .B1(_05033_),
    .A1(_05004_),
    .Y(_05044_),
    .A2(_05012_));
 sg13g2_a221oi_1 _22632_ (.B2(\cpu.uart.r_in[7] ),
    .C1(_04913_),
    .B1(_04916_),
    .A1(\cpu.uart.r_div_value[7] ),
    .Y(_05045_),
    .A2(_04847_));
 sg13g2_a21oi_1 _22633_ (.A1(net533),
    .A2(_05044_),
    .Y(_05046_),
    .B1(_05045_));
 sg13g2_and2_1 _22634_ (.A(net634),
    .B(\cpu.dcache.r_data[6][23] ),
    .X(_05047_));
 sg13g2_a21oi_1 _22635_ (.A1(net679),
    .A2(\cpu.dcache.r_data[4][23] ),
    .Y(_05048_),
    .B1(_05047_));
 sg13g2_nand2_1 _22636_ (.Y(_05049_),
    .A(\cpu.dcache.r_data[7][23] ),
    .B(net693));
 sg13g2_o21ai_1 _22637_ (.B1(_05049_),
    .Y(_05050_),
    .A1(net633),
    .A2(_05048_));
 sg13g2_nand2b_1 _22638_ (.Y(_05051_),
    .B(net536),
    .A_N(_00137_));
 sg13g2_a22oi_1 _22639_ (.Y(_05052_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][23] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_a22oi_1 _22640_ (.Y(_05053_),
    .B1(net700),
    .B2(\cpu.dcache.r_data[5][23] ),
    .A2(net563),
    .A1(\cpu.dcache.r_data[2][23] ));
 sg13g2_nand3_1 _22641_ (.B(_05052_),
    .C(_05053_),
    .A(_05051_),
    .Y(_05054_));
 sg13g2_a21oi_2 _22642_ (.B1(_05054_),
    .Y(_05055_),
    .A2(_05050_),
    .A1(net779));
 sg13g2_nor2_1 _22643_ (.A(net901),
    .B(_05055_),
    .Y(_05056_));
 sg13g2_a22oi_1 _22644_ (.Y(_05057_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][31] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_a22oi_1 _22645_ (.Y(_05058_),
    .B1(net628),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(net563),
    .A1(\cpu.dcache.r_data[2][31] ));
 sg13g2_mux2_1 _22646_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(\cpu.dcache.r_data[7][31] ),
    .S(net713),
    .X(_05059_));
 sg13g2_a22oi_1 _22647_ (.Y(_05060_),
    .B1(_05059_),
    .B2(net633),
    .A2(net706),
    .A1(\cpu.dcache.r_data[6][31] ));
 sg13g2_nand2b_1 _22648_ (.Y(_05061_),
    .B(net779),
    .A_N(_05060_));
 sg13g2_and4_1 _22649_ (.A(_09364_),
    .B(_05057_),
    .C(_05058_),
    .D(_05061_),
    .X(_05062_));
 sg13g2_a21oi_2 _22650_ (.B1(_05062_),
    .Y(_05063_),
    .A2(_04757_),
    .A1(_00138_));
 sg13g2_nor2b_1 _22651_ (.A(net667),
    .B_N(_05063_),
    .Y(_05064_));
 sg13g2_a21oi_1 _22652_ (.A1(net667),
    .A2(_05056_),
    .Y(_05065_),
    .B1(_05064_));
 sg13g2_nor2_1 _22653_ (.A(_11898_),
    .B(_05065_),
    .Y(_05066_));
 sg13g2_a22oi_1 _22654_ (.Y(_05067_),
    .B1(net698),
    .B2(\cpu.dcache.r_data[3][7] ),
    .A2(net631),
    .A1(\cpu.dcache.r_data[6][7] ));
 sg13g2_a22oi_1 _22655_ (.Y(_05068_),
    .B1(net697),
    .B2(\cpu.dcache.r_data[7][7] ),
    .A2(net700),
    .A1(\cpu.dcache.r_data[5][7] ));
 sg13g2_a22oi_1 _22656_ (.Y(_05069_),
    .B1(net628),
    .B2(\cpu.dcache.r_data[4][7] ),
    .A2(net629),
    .A1(\cpu.dcache.r_data[2][7] ));
 sg13g2_nand3_1 _22657_ (.B(_05068_),
    .C(_05069_),
    .A(_05067_),
    .Y(_05070_));
 sg13g2_nand2_1 _22658_ (.Y(_05071_),
    .A(_00136_),
    .B(_09362_));
 sg13g2_o21ai_1 _22659_ (.B1(_05071_),
    .Y(_05072_),
    .A1(_09362_),
    .A2(_05070_));
 sg13g2_nor3_1 _22660_ (.A(\cpu.dcache.r_data[1][7] ),
    .B(net572),
    .C(_05070_),
    .Y(_05073_));
 sg13g2_a21o_1 _22661_ (.A2(_05072_),
    .A1(net572),
    .B1(_05073_),
    .X(_05074_));
 sg13g2_buf_1 _22662_ (.A(_05074_),
    .X(_05075_));
 sg13g2_nand2_1 _22663_ (.Y(_05076_),
    .A(_11898_),
    .B(net667));
 sg13g2_mux2_1 _22664_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(\cpu.dcache.r_data[6][15] ),
    .S(net634),
    .X(_05077_));
 sg13g2_a22oi_1 _22665_ (.Y(_05078_),
    .B1(_05077_),
    .B2(net782),
    .A2(_09641_),
    .A1(\cpu.dcache.r_data[5][15] ));
 sg13g2_a22oi_1 _22666_ (.Y(_05079_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][15] ),
    .A2(_02891_),
    .A1(\cpu.dcache.r_data[2][15] ));
 sg13g2_o21ai_1 _22667_ (.B1(_05079_),
    .Y(_05080_),
    .A1(_00139_),
    .A2(_09364_));
 sg13g2_a221oi_1 _22668_ (.B2(\cpu.dcache.r_data[7][15] ),
    .C1(_05080_),
    .B1(_09484_),
    .A1(\cpu.dcache.r_data[3][15] ),
    .Y(_05081_),
    .A2(net616));
 sg13g2_o21ai_1 _22669_ (.B1(_05081_),
    .Y(_05082_),
    .A1(net910),
    .A2(_05078_));
 sg13g2_nor2_1 _22670_ (.A(_09244_),
    .B(net667),
    .Y(_05083_));
 sg13g2_nand2_1 _22671_ (.Y(_05084_),
    .A(_05082_),
    .B(_05083_));
 sg13g2_o21ai_1 _22672_ (.B1(_05084_),
    .Y(_05085_),
    .A1(_05075_),
    .A2(_05076_));
 sg13g2_nor3_1 _22673_ (.A(_05001_),
    .B(_05066_),
    .C(_05085_),
    .Y(_05086_));
 sg13g2_nor2_1 _22674_ (.A(_09244_),
    .B(_05075_),
    .Y(_05087_));
 sg13g2_nor3_1 _22675_ (.A(_04752_),
    .B(_05056_),
    .C(_05087_),
    .Y(_05088_));
 sg13g2_nor3_1 _22676_ (.A(_08321_),
    .B(_05086_),
    .C(_05088_),
    .Y(_05089_));
 sg13g2_a21oi_2 _22677_ (.B1(_05089_),
    .Y(_05090_),
    .A2(_05046_),
    .A1(_08321_));
 sg13g2_inv_1 _22678_ (.Y(_05091_),
    .A(_05090_));
 sg13g2_a21oi_1 _22679_ (.A1(net1133),
    .A2(_05091_),
    .Y(_05092_),
    .B1(_11405_));
 sg13g2_buf_2 _22680_ (.A(_05092_),
    .X(_05093_));
 sg13g2_o21ai_1 _22681_ (.B1(_05093_),
    .Y(_05094_),
    .A1(net983),
    .A2(_05003_));
 sg13g2_nor2_1 _22682_ (.A(net34),
    .B(_05094_),
    .Y(_05095_));
 sg13g2_a21oi_1 _22683_ (.A1(_02932_),
    .A2(net34),
    .Y(_05096_),
    .B1(_05095_));
 sg13g2_o21ai_1 _22684_ (.B1(_05096_),
    .Y(_05097_),
    .A1(net973),
    .A2(_04969_));
 sg13g2_a21oi_1 _22685_ (.A1(_04962_),
    .A2(_04968_),
    .Y(_01024_),
    .B1(_05097_));
 sg13g2_nor2_1 _22686_ (.A(net664),
    .B(_04967_),
    .Y(_05098_));
 sg13g2_nor2_1 _22687_ (.A(_04958_),
    .B(_04186_),
    .Y(_05099_));
 sg13g2_nand2_1 _22688_ (.Y(_05100_),
    .A(_09082_),
    .B(_11403_));
 sg13g2_buf_2 _22689_ (.A(_05100_),
    .X(_05101_));
 sg13g2_nor2_1 _22690_ (.A(net352),
    .B(_05101_),
    .Y(_05102_));
 sg13g2_a22oi_1 _22691_ (.Y(_05103_),
    .B1(net429),
    .B2(\cpu.intr.r_timer_reload[11] ),
    .A2(net532),
    .A1(_09915_));
 sg13g2_a22oi_1 _22692_ (.Y(_05104_),
    .B1(net593),
    .B2(\cpu.intr.r_clock_cmp[27] ),
    .A2(net447),
    .A1(_10106_));
 sg13g2_buf_1 _22693_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05105_));
 sg13g2_a22oi_1 _22694_ (.Y(_05106_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net387),
    .A1(_05105_));
 sg13g2_nand3_1 _22695_ (.B(_05104_),
    .C(_05106_),
    .A(_05103_),
    .Y(_05107_));
 sg13g2_mux2_1 _22696_ (.A0(\cpu.dcache.r_data[1][27] ),
    .A1(\cpu.dcache.r_data[3][27] ),
    .S(net507),
    .X(_05108_));
 sg13g2_a22oi_1 _22697_ (.Y(_05109_),
    .B1(_05108_),
    .B2(net574),
    .A2(_09314_),
    .A1(\cpu.dcache.r_data[2][27] ));
 sg13g2_inv_1 _22698_ (.Y(_05110_),
    .A(_00100_));
 sg13g2_mux2_1 _22699_ (.A0(\cpu.dcache.r_data[5][27] ),
    .A1(\cpu.dcache.r_data[7][27] ),
    .S(_09165_),
    .X(_05111_));
 sg13g2_a22oi_1 _22700_ (.Y(_05112_),
    .B1(_05111_),
    .B2(_09242_),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][27] ));
 sg13g2_nor2_1 _22701_ (.A(net758),
    .B(_05112_),
    .Y(_05113_));
 sg13g2_a221oi_1 _22702_ (.B2(\cpu.dcache.r_data[6][27] ),
    .C1(_05113_),
    .B1(net481),
    .A1(_05110_),
    .Y(_05114_),
    .A2(_04758_));
 sg13g2_o21ai_1 _22703_ (.B1(_05114_),
    .Y(_05115_),
    .A1(_09310_),
    .A2(_05109_));
 sg13g2_nand2_1 _22704_ (.Y(_05116_),
    .A(net673),
    .B(_05115_));
 sg13g2_nand2_1 _22705_ (.Y(_05117_),
    .A(\cpu.dcache.r_data[3][11] ),
    .B(net562));
 sg13g2_a22oi_1 _22706_ (.Y(_05118_),
    .B1(net563),
    .B2(\cpu.dcache.r_data[2][11] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][11] ));
 sg13g2_a22oi_1 _22707_ (.Y(_05119_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][11] ),
    .A2(net615),
    .A1(\cpu.dcache.r_data[5][11] ));
 sg13g2_a22oi_1 _22708_ (.Y(_05120_),
    .B1(_02906_),
    .B2(\cpu.dcache.r_data[7][11] ),
    .A2(_10035_),
    .A1(\cpu.dcache.r_data[4][11] ));
 sg13g2_nand4_1 _22709_ (.B(_05118_),
    .C(_05119_),
    .A(_05117_),
    .Y(_05121_),
    .D(_05120_));
 sg13g2_nor2_1 _22710_ (.A(net475),
    .B(_05121_),
    .Y(_05122_));
 sg13g2_a21oi_1 _22711_ (.A1(_00101_),
    .A2(net475),
    .Y(_05123_),
    .B1(_05122_));
 sg13g2_nand2_1 _22712_ (.Y(_05124_),
    .A(net780),
    .B(_05123_));
 sg13g2_nand2_1 _22713_ (.Y(_05125_),
    .A(_05116_),
    .B(_05124_));
 sg13g2_a22oi_1 _22714_ (.Y(_05126_),
    .B1(_05125_),
    .B2(net663),
    .A2(_05107_),
    .A1(_04973_));
 sg13g2_o21ai_1 _22715_ (.B1(_05093_),
    .Y(_05127_),
    .A1(net983),
    .A2(_05126_));
 sg13g2_mux2_1 _22716_ (.A0(_05127_),
    .A1(_10693_),
    .S(net34),
    .X(_05128_));
 sg13g2_o21ai_1 _22717_ (.B1(_05128_),
    .Y(_05129_),
    .A1(\cpu.ex.pc[11] ),
    .A2(_04969_));
 sg13g2_a221oi_1 _22718_ (.B2(_05102_),
    .C1(_05129_),
    .B1(_05099_),
    .A1(_04180_),
    .Y(_01025_),
    .A2(_05098_));
 sg13g2_a221oi_1 _22719_ (.B2(net132),
    .C1(_04244_),
    .B1(\cpu.ex.c_mult[12] ),
    .A1(_03011_),
    .Y(_05130_),
    .A2(_11398_));
 sg13g2_a22oi_1 _22720_ (.Y(_05131_),
    .B1(net429),
    .B2(\cpu.intr.r_timer_reload[12] ),
    .A2(_04901_),
    .A1(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_a22oi_1 _22721_ (.Y(_05132_),
    .B1(net532),
    .B2(\cpu.intr.r_timer_count[12] ),
    .A2(net502),
    .A1(_10114_));
 sg13g2_buf_2 _22722_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05133_));
 sg13g2_a22oi_1 _22723_ (.Y(_05134_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net431),
    .A1(_05133_));
 sg13g2_nand3_1 _22724_ (.B(_05132_),
    .C(_05134_),
    .A(_05131_),
    .Y(_05135_));
 sg13g2_mux2_1 _22725_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(\cpu.dcache.r_data[6][28] ),
    .S(net473),
    .X(_05136_));
 sg13g2_a22oi_1 _22726_ (.Y(_05137_),
    .B1(_05136_),
    .B2(net782),
    .A2(net693),
    .A1(\cpu.dcache.r_data[7][28] ));
 sg13g2_a22oi_1 _22727_ (.Y(_05138_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][28] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][28] ));
 sg13g2_o21ai_1 _22728_ (.B1(_05138_),
    .Y(_05139_),
    .A1(_00110_),
    .A2(net535));
 sg13g2_a221oi_1 _22729_ (.B2(\cpu.dcache.r_data[5][28] ),
    .C1(_05139_),
    .B1(net615),
    .A1(\cpu.dcache.r_data[2][28] ),
    .Y(_05140_),
    .A2(net474));
 sg13g2_o21ai_1 _22730_ (.B1(_05140_),
    .Y(_05141_),
    .A1(net758),
    .A2(_05137_));
 sg13g2_mux2_1 _22731_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(\cpu.dcache.r_data[6][12] ),
    .S(net473),
    .X(_05142_));
 sg13g2_a22oi_1 _22732_ (.Y(_05143_),
    .B1(_05142_),
    .B2(net669),
    .A2(_09904_),
    .A1(\cpu.dcache.r_data[7][12] ));
 sg13g2_a22oi_1 _22733_ (.Y(_05144_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][12] ),
    .A2(_02894_),
    .A1(\cpu.dcache.r_data[3][12] ));
 sg13g2_o21ai_1 _22734_ (.B1(_05144_),
    .Y(_05145_),
    .A1(_00111_),
    .A2(net535));
 sg13g2_a221oi_1 _22735_ (.B2(\cpu.dcache.r_data[5][12] ),
    .C1(_05145_),
    .B1(net537),
    .A1(\cpu.dcache.r_data[2][12] ),
    .Y(_05146_),
    .A2(_04766_));
 sg13g2_o21ai_1 _22736_ (.B1(_05146_),
    .Y(_05147_),
    .A1(net680),
    .A2(_05143_));
 sg13g2_mux2_1 _22737_ (.A0(_05141_),
    .A1(_05147_),
    .S(_09902_),
    .X(_05148_));
 sg13g2_a22oi_1 _22738_ (.Y(_05149_),
    .B1(_05148_),
    .B2(net663),
    .A2(_05135_),
    .A1(_04973_));
 sg13g2_o21ai_1 _22739_ (.B1(_05093_),
    .Y(_05150_),
    .A1(net1133),
    .A2(_05149_));
 sg13g2_mux2_1 _22740_ (.A0(_05150_),
    .A1(net695),
    .S(net34),
    .X(_05151_));
 sg13g2_o21ai_1 _22741_ (.B1(_05151_),
    .Y(_05152_),
    .A1(_08408_),
    .A2(_04969_));
 sg13g2_nor3_1 _22742_ (.A(net665),
    .B(_04247_),
    .C(_04967_),
    .Y(_05153_));
 sg13g2_or2_1 _22743_ (.X(_05154_),
    .B(_05153_),
    .A(_05152_));
 sg13g2_a21oi_1 _22744_ (.A1(_05102_),
    .A2(_05130_),
    .Y(_01026_),
    .B1(_05154_));
 sg13g2_buf_1 _22745_ (.A(_05101_),
    .X(_05155_));
 sg13g2_a22oi_1 _22746_ (.Y(_05156_),
    .B1(net429),
    .B2(\cpu.intr.r_timer_reload[13] ),
    .A2(net593),
    .A1(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_a22oi_1 _22747_ (.Y(_05157_),
    .B1(net532),
    .B2(\cpu.intr.r_timer_count[13] ),
    .A2(net447),
    .A1(_10120_));
 sg13g2_buf_1 _22748_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05158_));
 sg13g2_a22oi_1 _22749_ (.Y(_05159_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net387),
    .A1(_05158_));
 sg13g2_nand3_1 _22750_ (.B(_05157_),
    .C(_05159_),
    .A(_05156_),
    .Y(_05160_));
 sg13g2_mux2_1 _22751_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(\cpu.dcache.r_data[7][29] ),
    .S(net473),
    .X(_05161_));
 sg13g2_a22oi_1 _22752_ (.Y(_05162_),
    .B1(_05161_),
    .B2(net574),
    .A2(net706),
    .A1(\cpu.dcache.r_data[6][29] ));
 sg13g2_a22oi_1 _22753_ (.Y(_05163_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][29] ),
    .A2(net564),
    .A1(\cpu.dcache.r_data[1][29] ));
 sg13g2_o21ai_1 _22754_ (.B1(_05163_),
    .Y(_05164_),
    .A1(_00116_),
    .A2(_04782_));
 sg13g2_a221oi_1 _22755_ (.B2(\cpu.dcache.r_data[2][29] ),
    .C1(_05164_),
    .B1(net483),
    .A1(\cpu.dcache.r_data[3][29] ),
    .Y(_05165_),
    .A2(net482));
 sg13g2_o21ai_1 _22756_ (.B1(_05165_),
    .Y(_05166_),
    .A1(_11839_),
    .A2(_05162_));
 sg13g2_mux2_1 _22757_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(\cpu.dcache.r_data[6][13] ),
    .S(_04787_),
    .X(_05167_));
 sg13g2_a22oi_1 _22758_ (.Y(_05168_),
    .B1(_05167_),
    .B2(net669),
    .A2(_09904_),
    .A1(\cpu.dcache.r_data[7][13] ));
 sg13g2_a22oi_1 _22759_ (.Y(_05169_),
    .B1(_02888_),
    .B2(\cpu.dcache.r_data[1][13] ),
    .A2(_02895_),
    .A1(\cpu.dcache.r_data[3][13] ));
 sg13g2_o21ai_1 _22760_ (.B1(_05169_),
    .Y(_05170_),
    .A1(_00117_),
    .A2(net535));
 sg13g2_a221oi_1 _22761_ (.B2(\cpu.dcache.r_data[5][13] ),
    .C1(_05170_),
    .B1(_04755_),
    .A1(\cpu.dcache.r_data[2][13] ),
    .Y(_05171_),
    .A2(net483));
 sg13g2_o21ai_1 _22762_ (.B1(_05171_),
    .Y(_05172_),
    .A1(net680),
    .A2(_05168_));
 sg13g2_mux2_1 _22763_ (.A0(_05166_),
    .A1(_05172_),
    .S(net672),
    .X(_05173_));
 sg13g2_a22oi_1 _22764_ (.Y(_05174_),
    .B1(_05173_),
    .B2(net663),
    .A2(_05160_),
    .A1(_04973_));
 sg13g2_o21ai_1 _22765_ (.B1(_05093_),
    .Y(_05175_),
    .A1(net983),
    .A2(_05174_));
 sg13g2_buf_1 _22766_ (.A(_04749_),
    .X(_05176_));
 sg13g2_mux2_1 _22767_ (.A0(net696),
    .A1(_05175_),
    .S(net71),
    .X(_05177_));
 sg13g2_nand2_1 _22768_ (.Y(_05178_),
    .A(_08416_),
    .B(net352));
 sg13g2_o21ai_1 _22769_ (.B1(_03834_),
    .Y(_05179_),
    .A1(net665),
    .A2(_04311_));
 sg13g2_a21oi_1 _22770_ (.A1(_05178_),
    .A2(_05179_),
    .Y(_05180_),
    .B1(_05101_));
 sg13g2_a21oi_1 _22771_ (.A1(net82),
    .A2(_05177_),
    .Y(_05181_),
    .B1(_05180_));
 sg13g2_a21oi_1 _22772_ (.A1(_04309_),
    .A2(_05098_),
    .Y(_01027_),
    .B1(_05181_));
 sg13g2_a22oi_1 _22773_ (.Y(_05182_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[14] ),
    .A2(_04974_),
    .A1(\cpu.intr.r_timer_reload[14] ));
 sg13g2_a22oi_1 _22774_ (.Y(_05183_),
    .B1(net532),
    .B2(_09914_),
    .A2(net502),
    .A1(_10126_));
 sg13g2_buf_1 _22775_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05184_));
 sg13g2_a22oi_1 _22776_ (.Y(_05185_),
    .B1(net387),
    .B2(_05184_),
    .A2(net593),
    .A1(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_nand3_1 _22777_ (.B(_05183_),
    .C(_05185_),
    .A(_05182_),
    .Y(_05186_));
 sg13g2_mux2_1 _22778_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(\cpu.dcache.r_data[6][30] ),
    .S(net473),
    .X(_05187_));
 sg13g2_a22oi_1 _22779_ (.Y(_05188_),
    .B1(_05187_),
    .B2(net669),
    .A2(net693),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_a22oi_1 _22780_ (.Y(_05189_),
    .B1(_09678_),
    .B2(\cpu.dcache.r_data[1][30] ),
    .A2(_02894_),
    .A1(\cpu.dcache.r_data[3][30] ));
 sg13g2_o21ai_1 _22781_ (.B1(_05189_),
    .Y(_05190_),
    .A1(_00127_),
    .A2(net535));
 sg13g2_a221oi_1 _22782_ (.B2(\cpu.dcache.r_data[5][30] ),
    .C1(_05190_),
    .B1(_02899_),
    .A1(\cpu.dcache.r_data[2][30] ),
    .Y(_05191_),
    .A2(_04766_));
 sg13g2_o21ai_1 _22783_ (.B1(_05191_),
    .Y(_05192_),
    .A1(_11838_),
    .A2(_05188_));
 sg13g2_a22oi_1 _22784_ (.Y(_05193_),
    .B1(_02889_),
    .B2(\cpu.dcache.r_data[1][14] ),
    .A2(_02896_),
    .A1(\cpu.dcache.r_data[3][14] ));
 sg13g2_a22oi_1 _22785_ (.Y(_05194_),
    .B1(_10036_),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(_02892_),
    .A1(\cpu.dcache.r_data[2][14] ));
 sg13g2_mux2_1 _22786_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(\cpu.dcache.r_data[7][14] ),
    .S(_04787_),
    .X(_05195_));
 sg13g2_a22oi_1 _22787_ (.Y(_05196_),
    .B1(_05195_),
    .B2(net574),
    .A2(net706),
    .A1(\cpu.dcache.r_data[6][14] ));
 sg13g2_nand2b_1 _22788_ (.Y(_05197_),
    .B(net779),
    .A_N(_05196_));
 sg13g2_and4_1 _22789_ (.A(_04782_),
    .B(_05193_),
    .C(_05194_),
    .D(_05197_),
    .X(_05198_));
 sg13g2_a21oi_2 _22790_ (.B1(_05198_),
    .Y(_05199_),
    .A2(_04758_),
    .A1(_00128_));
 sg13g2_mux2_1 _22791_ (.A0(_05192_),
    .A1(_05199_),
    .S(net672),
    .X(_05200_));
 sg13g2_a22oi_1 _22792_ (.Y(_05201_),
    .B1(_05200_),
    .B2(_05002_),
    .A2(_05186_),
    .A1(_04973_));
 sg13g2_o21ai_1 _22793_ (.B1(_05093_),
    .Y(_05202_),
    .A1(net1133),
    .A2(_05201_));
 sg13g2_nand2_1 _22794_ (.Y(_05203_),
    .A(net71),
    .B(_05202_));
 sg13g2_o21ai_1 _22795_ (.B1(_05203_),
    .Y(_05204_),
    .A1(_03536_),
    .A2(net71));
 sg13g2_nand2_1 _22796_ (.Y(_05205_),
    .A(_05155_),
    .B(_05204_));
 sg13g2_buf_1 _22797_ (.A(_03834_),
    .X(_05206_));
 sg13g2_o21ai_1 _22798_ (.B1(net86),
    .Y(_05207_),
    .A1(_08424_),
    .A2(_05206_));
 sg13g2_or3_1 _22799_ (.A(net664),
    .B(_04348_),
    .C(_04350_),
    .X(_05208_));
 sg13g2_a21oi_1 _22800_ (.A1(net664),
    .A2(_04354_),
    .Y(_05209_),
    .B1(_04967_));
 sg13g2_a22oi_1 _22801_ (.Y(_01028_),
    .B1(_05208_),
    .B2(_05209_),
    .A2(_05207_),
    .A1(_05205_));
 sg13g2_a22oi_1 _22802_ (.Y(_05210_),
    .B1(_04902_),
    .B2(\cpu.intr.r_timer_reload[15] ),
    .A2(_04868_),
    .A1(_09913_));
 sg13g2_a22oi_1 _22803_ (.Y(_05211_),
    .B1(_04901_),
    .B2(\cpu.intr.r_clock_cmp[31] ),
    .A2(net502),
    .A1(_10131_));
 sg13g2_a22oi_1 _22804_ (.Y(_05212_),
    .B1(_04977_),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net431),
    .A1(\cpu.intr.r_clock_count[31] ));
 sg13g2_nand3_1 _22805_ (.B(_05211_),
    .C(_05212_),
    .A(_05210_),
    .Y(_05213_));
 sg13g2_mux2_1 _22806_ (.A0(_05082_),
    .A1(_05063_),
    .S(net666),
    .X(_05214_));
 sg13g2_a22oi_1 _22807_ (.Y(_05215_),
    .B1(_05214_),
    .B2(_05002_),
    .A2(_05213_),
    .A1(_04973_));
 sg13g2_o21ai_1 _22808_ (.B1(_05093_),
    .Y(_05216_),
    .A1(net1133),
    .A2(_05215_));
 sg13g2_nand2_1 _22809_ (.Y(_05217_),
    .A(_04749_),
    .B(_05216_));
 sg13g2_o21ai_1 _22810_ (.B1(_05217_),
    .Y(_05218_),
    .A1(_09426_),
    .A2(_05176_));
 sg13g2_nand2_1 _22811_ (.Y(_05219_),
    .A(net82),
    .B(_05218_));
 sg13g2_o21ai_1 _22812_ (.B1(_05216_),
    .Y(_05220_),
    .A1(_08363_),
    .A2(_03834_));
 sg13g2_or2_1 _22813_ (.X(_05221_),
    .B(_05220_),
    .A(_04971_));
 sg13g2_a21oi_1 _22814_ (.A1(net132),
    .A2(_11774_),
    .Y(_05222_),
    .B1(_04965_));
 sg13g2_o21ai_1 _22815_ (.B1(_05222_),
    .Y(_05223_),
    .A1(_04360_),
    .A2(_04395_));
 sg13g2_a221oi_1 _22816_ (.B2(_05101_),
    .C1(net352),
    .B1(_05218_),
    .A1(net664),
    .Y(_05224_),
    .A2(_04399_));
 sg13g2_a22oi_1 _22817_ (.Y(_01029_),
    .B1(_05223_),
    .B2(_05224_),
    .A2(_05221_),
    .A1(_05219_));
 sg13g2_nand2_1 _22818_ (.Y(_05225_),
    .A(_10596_),
    .B(_04963_));
 sg13g2_o21ai_1 _22819_ (.B1(_05225_),
    .Y(_05226_),
    .A1(net740),
    .A2(_03977_));
 sg13g2_mux2_1 _22820_ (.A0(net803),
    .A1(_05226_),
    .S(net270),
    .X(_05227_));
 sg13g2_mux2_1 _22821_ (.A0(\cpu.dcache.r_data[1][1] ),
    .A1(\cpu.dcache.r_data[3][1] ),
    .S(net473),
    .X(_05228_));
 sg13g2_a22oi_1 _22822_ (.Y(_05229_),
    .B1(_05228_),
    .B2(net574),
    .A2(net706),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_mux2_1 _22823_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(\cpu.dcache.r_data[7][1] ),
    .S(net575),
    .X(_05230_));
 sg13g2_a22oi_1 _22824_ (.Y(_05231_),
    .B1(_05230_),
    .B2(net633),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][1] ));
 sg13g2_nor2_1 _22825_ (.A(net758),
    .B(_05231_),
    .Y(_05232_));
 sg13g2_a221oi_1 _22826_ (.B2(\cpu.dcache.r_data[6][1] ),
    .C1(_05232_),
    .B1(_02903_),
    .A1(\cpu.dcache.r_data[0][1] ),
    .Y(_05233_),
    .A2(net475));
 sg13g2_o21ai_1 _22827_ (.B1(_05233_),
    .Y(_05234_),
    .A1(_09310_),
    .A2(_05229_));
 sg13g2_mux2_1 _22828_ (.A0(\cpu.dcache.r_data[1][17] ),
    .A1(\cpu.dcache.r_data[3][17] ),
    .S(net575),
    .X(_05235_));
 sg13g2_a22oi_1 _22829_ (.Y(_05236_),
    .B1(_05235_),
    .B2(net633),
    .A2(net706),
    .A1(\cpu.dcache.r_data[2][17] ));
 sg13g2_inv_1 _22830_ (.Y(_05237_),
    .A(_00299_));
 sg13g2_mux2_1 _22831_ (.A0(\cpu.dcache.r_data[5][17] ),
    .A1(\cpu.dcache.r_data[7][17] ),
    .S(net575),
    .X(_05238_));
 sg13g2_a22oi_1 _22832_ (.Y(_05239_),
    .B1(_05238_),
    .B2(net633),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][17] ));
 sg13g2_nor2_1 _22833_ (.A(net758),
    .B(_05239_),
    .Y(_05240_));
 sg13g2_a221oi_1 _22834_ (.B2(\cpu.dcache.r_data[6][17] ),
    .C1(_05240_),
    .B1(_02902_),
    .A1(_05237_),
    .Y(_05241_),
    .A2(net536));
 sg13g2_o21ai_1 _22835_ (.B1(_05241_),
    .Y(_05242_),
    .A1(_09310_),
    .A2(_05236_));
 sg13g2_mux2_1 _22836_ (.A0(_05234_),
    .A1(_05242_),
    .S(net609),
    .X(_05243_));
 sg13g2_mux2_1 _22837_ (.A0(\cpu.dcache.r_data[5][25] ),
    .A1(\cpu.dcache.r_data[7][25] ),
    .S(net575),
    .X(_05244_));
 sg13g2_a22oi_1 _22838_ (.Y(_05245_),
    .B1(_05244_),
    .B2(_09241_),
    .A2(_09314_),
    .A1(\cpu.dcache.r_data[6][25] ));
 sg13g2_nor2_1 _22839_ (.A(_11838_),
    .B(_05245_),
    .Y(_05246_));
 sg13g2_a22oi_1 _22840_ (.Y(_05247_),
    .B1(net628),
    .B2(\cpu.dcache.r_data[4][25] ),
    .A2(_09678_),
    .A1(\cpu.dcache.r_data[1][25] ));
 sg13g2_o21ai_1 _22841_ (.B1(_05247_),
    .Y(_05248_),
    .A1(_00300_),
    .A2(_09364_));
 sg13g2_a221oi_1 _22842_ (.B2(\cpu.dcache.r_data[2][25] ),
    .C1(_05248_),
    .B1(_02891_),
    .A1(\cpu.dcache.r_data[3][25] ),
    .Y(_05249_),
    .A2(net562));
 sg13g2_nor2b_1 _22843_ (.A(_05246_),
    .B_N(_05249_),
    .Y(_05250_));
 sg13g2_mux2_1 _22844_ (.A0(\cpu.dcache.r_data[5][9] ),
    .A1(\cpu.dcache.r_data[7][9] ),
    .S(net473),
    .X(_05251_));
 sg13g2_a22oi_1 _22845_ (.Y(_05252_),
    .B1(_05251_),
    .B2(net574),
    .A2(net705),
    .A1(\cpu.dcache.r_data[4][9] ));
 sg13g2_nor2_1 _22846_ (.A(net758),
    .B(_05252_),
    .Y(_05253_));
 sg13g2_a22oi_1 _22847_ (.Y(_05254_),
    .B1(_02888_),
    .B2(\cpu.dcache.r_data[1][9] ),
    .A2(_02902_),
    .A1(\cpu.dcache.r_data[6][9] ));
 sg13g2_o21ai_1 _22848_ (.B1(_05254_),
    .Y(_05255_),
    .A1(_00301_),
    .A2(net535));
 sg13g2_a221oi_1 _22849_ (.B2(\cpu.dcache.r_data[2][9] ),
    .C1(_05255_),
    .B1(_02892_),
    .A1(\cpu.dcache.r_data[3][9] ),
    .Y(_05256_),
    .A2(_02896_));
 sg13g2_nor2b_1 _22850_ (.A(_05253_),
    .B_N(_05256_),
    .Y(_05257_));
 sg13g2_or2_1 _22851_ (.X(_05258_),
    .B(_05257_),
    .A(net666));
 sg13g2_o21ai_1 _22852_ (.B1(_05258_),
    .Y(_05259_),
    .A1(net972),
    .A2(_05250_));
 sg13g2_a22oi_1 _22853_ (.Y(_05260_),
    .B1(_05242_),
    .B2(_04796_),
    .A2(_05234_),
    .A1(net972));
 sg13g2_nand2_1 _22854_ (.Y(_05261_),
    .A(net596),
    .B(_05260_));
 sg13g2_o21ai_1 _22855_ (.B1(_05261_),
    .Y(_05262_),
    .A1(net596),
    .A2(_05259_));
 sg13g2_nand2_1 _22856_ (.Y(_05263_),
    .A(net597),
    .B(_05262_));
 sg13g2_o21ai_1 _22857_ (.B1(_05263_),
    .Y(_05264_),
    .A1(net597),
    .A2(_05243_));
 sg13g2_nand2_2 _22858_ (.Y(_05265_),
    .A(_09741_),
    .B(_04890_));
 sg13g2_nand2_1 _22859_ (.Y(_05266_),
    .A(_09093_),
    .B(_04849_));
 sg13g2_o21ai_1 _22860_ (.B1(_05266_),
    .Y(_05267_),
    .A1(_00306_),
    .A2(_05265_));
 sg13g2_nor2_1 _22861_ (.A(net780),
    .B(_00304_),
    .Y(_05268_));
 sg13g2_buf_2 _22862_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05269_));
 sg13g2_nor2b_1 _22863_ (.A(net666),
    .B_N(_05269_),
    .Y(_05270_));
 sg13g2_o21ai_1 _22864_ (.B1(_04811_),
    .Y(_05271_),
    .A1(_05268_),
    .A2(_05270_));
 sg13g2_o21ai_1 _22865_ (.B1(_05271_),
    .Y(_05272_),
    .A1(_00305_),
    .A2(net386));
 sg13g2_nand2b_1 _22866_ (.Y(_05273_),
    .B(_04868_),
    .A_N(net874));
 sg13g2_buf_2 _22867_ (.A(_05273_),
    .X(_05274_));
 sg13g2_nand2b_1 _22868_ (.Y(_05275_),
    .B(_04828_),
    .A_N(_00308_));
 sg13g2_o21ai_1 _22869_ (.B1(_05275_),
    .Y(_05276_),
    .A1(_00307_),
    .A2(_05274_));
 sg13g2_a21oi_1 _22870_ (.A1(_09093_),
    .A2(_04844_),
    .Y(_05277_),
    .B1(_04808_));
 sg13g2_nor2b_1 _22871_ (.A(_05277_),
    .B_N(_09094_),
    .Y(_05278_));
 sg13g2_nor4_1 _22872_ (.A(_05267_),
    .B(_05272_),
    .C(_05276_),
    .D(_05278_),
    .Y(_05279_));
 sg13g2_nand2b_1 _22873_ (.Y(_05280_),
    .B(_04804_),
    .A_N(_05279_));
 sg13g2_buf_1 _22874_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05281_));
 sg13g2_inv_1 _22875_ (.Y(_05282_),
    .A(_00303_));
 sg13g2_a22oi_1 _22876_ (.Y(_05283_),
    .B1(net428),
    .B2(_05282_),
    .A2(_04857_),
    .A1(_05281_));
 sg13g2_mux2_1 _22877_ (.A0(_11825_),
    .A1(_11830_),
    .S(net1016),
    .X(_05284_));
 sg13g2_buf_1 _22878_ (.A(_04847_),
    .X(_05285_));
 sg13g2_a22oi_1 _22879_ (.Y(_05286_),
    .B1(_05284_),
    .B2(_05285_),
    .A2(_05038_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_or2_1 _22880_ (.X(_05287_),
    .B(_04877_),
    .A(_00302_));
 sg13g2_nand3_1 _22881_ (.B(_05286_),
    .C(_05287_),
    .A(_05283_),
    .Y(_05288_));
 sg13g2_a221oi_1 _22882_ (.B2(_09188_),
    .C1(_05288_),
    .B1(_04866_),
    .A1(_11826_),
    .Y(_05289_),
    .A2(_04829_));
 sg13g2_nor2_1 _22883_ (.A(_09157_),
    .B(_05289_),
    .Y(_05290_));
 sg13g2_a22oi_1 _22884_ (.Y(_05291_),
    .B1(net559),
    .B2(\cpu.intr.r_timer_reload[17] ),
    .A2(net442),
    .A1(_09932_));
 sg13g2_a221oi_1 _22885_ (.B2(\cpu.intr.r_clock_cmp[1] ),
    .C1(net673),
    .B1(net561),
    .A1(_09917_),
    .Y(_05292_),
    .A2(net442));
 sg13g2_a21oi_1 _22886_ (.A1(net673),
    .A2(_05291_),
    .Y(_05293_),
    .B1(_05292_));
 sg13g2_nand2_1 _22887_ (.Y(_05294_),
    .A(\cpu.intr.r_timer_reload[1] ),
    .B(net429));
 sg13g2_buf_2 _22888_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05295_));
 sg13g2_a22oi_1 _22889_ (.Y(_05296_),
    .B1(_04982_),
    .B2(_05295_),
    .A2(net389),
    .A1(_09124_));
 sg13g2_a22oi_1 _22890_ (.Y(_05297_),
    .B1(net593),
    .B2(\cpu.intr.r_clock_cmp[17] ),
    .A2(net502),
    .A1(_10053_));
 sg13g2_nand3_1 _22891_ (.B(_05296_),
    .C(_05297_),
    .A(_05294_),
    .Y(_05298_));
 sg13g2_nor2_1 _22892_ (.A(_05293_),
    .B(_05298_),
    .Y(_05299_));
 sg13g2_a21oi_1 _22893_ (.A1(_09124_),
    .A2(net388),
    .Y(_05300_),
    .B1(net430));
 sg13g2_nand2b_1 _22894_ (.Y(_05301_),
    .B(\cpu.intr.r_clock ),
    .A_N(_05300_));
 sg13g2_a21oi_1 _22895_ (.A1(_05299_),
    .A2(_05301_),
    .Y(_05302_),
    .B1(net692));
 sg13g2_a22oi_1 _22896_ (.Y(_05303_),
    .B1(_04918_),
    .B2(\cpu.uart.r_div_value[9] ),
    .A2(_04847_),
    .A1(\cpu.uart.r_div_value[1] ));
 sg13g2_a22oi_1 _22897_ (.Y(_05304_),
    .B1(net472),
    .B2(\cpu.uart.r_r_invert ),
    .A2(net389),
    .A1(_09128_));
 sg13g2_nand2_1 _22898_ (.Y(_05305_),
    .A(_05303_),
    .B(_05304_));
 sg13g2_a21oi_1 _22899_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04916_),
    .Y(_05306_),
    .B1(_05305_));
 sg13g2_o21ai_1 _22900_ (.B1(net987),
    .Y(_05307_),
    .A1(net533),
    .A2(_05306_));
 sg13g2_nor3_1 _22901_ (.A(_05290_),
    .B(_05302_),
    .C(_05307_),
    .Y(_05308_));
 sg13g2_a22oi_1 _22902_ (.Y(_05309_),
    .B1(_05280_),
    .B2(_05308_),
    .A2(_05264_),
    .A1(net902));
 sg13g2_mux2_1 _22903_ (.A0(net609),
    .A1(_05309_),
    .S(net73),
    .X(_05310_));
 sg13g2_mux2_1 _22904_ (.A0(_05227_),
    .A1(_05310_),
    .S(net82),
    .X(_01030_));
 sg13g2_o21ai_1 _22905_ (.B1(net270),
    .Y(_05311_),
    .A1(net803),
    .A2(net665));
 sg13g2_nand3_1 _22906_ (.B(net803),
    .C(net740),
    .A(net724),
    .Y(_05312_));
 sg13g2_o21ai_1 _22907_ (.B1(_05312_),
    .Y(_05313_),
    .A1(net740),
    .A2(_04436_));
 sg13g2_a22oi_1 _22908_ (.Y(_05314_),
    .B1(_05313_),
    .B2(net270),
    .A2(_05311_),
    .A1(net717));
 sg13g2_a22oi_1 _22909_ (.Y(_05315_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[5][2] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][2] ));
 sg13g2_a22oi_1 _22910_ (.Y(_05316_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][2] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[3][2] ));
 sg13g2_a22oi_1 _22911_ (.Y(_05317_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][2] ),
    .A2(net563),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_nand3_1 _22912_ (.B(_05316_),
    .C(_05317_),
    .A(_05315_),
    .Y(_05318_));
 sg13g2_mux2_1 _22913_ (.A0(\cpu.dcache.r_data[0][2] ),
    .A1(_05318_),
    .S(net781),
    .X(_05319_));
 sg13g2_or3_1 _22914_ (.A(\cpu.dcache.r_data[1][2] ),
    .B(net572),
    .C(_05318_),
    .X(_05320_));
 sg13g2_o21ai_1 _22915_ (.B1(_05320_),
    .Y(_05321_),
    .A1(net484),
    .A2(_05319_));
 sg13g2_a22oi_1 _22916_ (.Y(_05322_),
    .B1(net700),
    .B2(\cpu.dcache.r_data[5][18] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][18] ));
 sg13g2_a22oi_1 _22917_ (.Y(_05323_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][18] ),
    .A2(net563),
    .A1(\cpu.dcache.r_data[2][18] ));
 sg13g2_a22oi_1 _22918_ (.Y(_05324_),
    .B1(net628),
    .B2(\cpu.dcache.r_data[4][18] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][18] ));
 sg13g2_nand3_1 _22919_ (.B(_05323_),
    .C(_05324_),
    .A(_05322_),
    .Y(_05325_));
 sg13g2_nand2_1 _22920_ (.Y(_05326_),
    .A(_00309_),
    .B(_09362_));
 sg13g2_o21ai_1 _22921_ (.B1(_05326_),
    .Y(_05327_),
    .A1(_09362_),
    .A2(_05325_));
 sg13g2_nor3_1 _22922_ (.A(\cpu.dcache.r_data[1][18] ),
    .B(net572),
    .C(_05325_),
    .Y(_05328_));
 sg13g2_a21o_1 _22923_ (.A2(_05327_),
    .A1(net572),
    .B1(_05328_),
    .X(_05329_));
 sg13g2_nand2b_1 _22924_ (.Y(_05330_),
    .B(net666),
    .A_N(_05329_));
 sg13g2_o21ai_1 _22925_ (.B1(_05330_),
    .Y(_05331_),
    .A1(net609),
    .A2(_05321_));
 sg13g2_nand2_1 _22926_ (.Y(_05332_),
    .A(net663),
    .B(_05331_));
 sg13g2_mux2_1 _22927_ (.A0(_05321_),
    .A1(_05330_),
    .S(net1012),
    .X(_05333_));
 sg13g2_a221oi_1 _22928_ (.B2(net672),
    .C1(_04777_),
    .B1(_04999_),
    .A1(net1012),
    .Y(_05334_),
    .A2(_04991_));
 sg13g2_a21oi_1 _22929_ (.A1(net596),
    .A2(_05333_),
    .Y(_05335_),
    .B1(_05334_));
 sg13g2_nand2_1 _22930_ (.Y(_05336_),
    .A(net597),
    .B(_05335_));
 sg13g2_nand3_1 _22931_ (.B(_05332_),
    .C(_05336_),
    .A(net902),
    .Y(_05337_));
 sg13g2_buf_1 _22932_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05338_));
 sg13g2_inv_1 _22933_ (.Y(_05339_),
    .A(_00093_));
 sg13g2_nand2_1 _22934_ (.Y(_05340_),
    .A(net1016),
    .B(_11811_));
 sg13g2_o21ai_1 _22935_ (.B1(_05340_),
    .Y(_05341_),
    .A1(net1016),
    .A2(_00263_));
 sg13g2_a22oi_1 _22936_ (.Y(_05342_),
    .B1(_05341_),
    .B2(_04847_),
    .A2(_05038_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _22937_ (.B1(_05342_),
    .Y(_05343_),
    .A1(_00092_),
    .A2(_04877_));
 sg13g2_a221oi_1 _22938_ (.B2(_05339_),
    .C1(_05343_),
    .B1(net428),
    .A1(_05338_),
    .Y(_05344_),
    .A2(_04857_));
 sg13g2_o21ai_1 _22939_ (.B1(_05344_),
    .Y(_05345_),
    .A1(_00264_),
    .A2(_05274_));
 sg13g2_a21oi_1 _22940_ (.A1(_09192_),
    .A2(_04866_),
    .Y(_05346_),
    .B1(_05345_));
 sg13g2_nand3_1 _22941_ (.B(_09089_),
    .C(_04844_),
    .A(_09088_),
    .Y(_05347_));
 sg13g2_nand2b_1 _22942_ (.Y(_05348_),
    .B(_04829_),
    .A_N(_00097_));
 sg13g2_inv_1 _22943_ (.Y(_05349_),
    .A(_00095_));
 sg13g2_nand2_1 _22944_ (.Y(_05350_),
    .A(net797),
    .B(_04811_));
 sg13g2_buf_1 _22945_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05351_));
 sg13g2_and2_1 _22946_ (.A(net901),
    .B(_04811_),
    .X(_05352_));
 sg13g2_buf_1 _22947_ (.A(_05352_),
    .X(_05353_));
 sg13g2_nand2_1 _22948_ (.Y(_05354_),
    .A(_05351_),
    .B(_05353_));
 sg13g2_o21ai_1 _22949_ (.B1(_05354_),
    .Y(_05355_),
    .A1(_00094_),
    .A2(_05350_));
 sg13g2_a221oi_1 _22950_ (.B2(_05349_),
    .C1(_05355_),
    .B1(_04823_),
    .A1(_09089_),
    .Y(_05356_),
    .A2(_04808_));
 sg13g2_inv_1 _22951_ (.Y(_05357_),
    .A(_00098_));
 sg13g2_nor2_1 _22952_ (.A(_00096_),
    .B(_05265_),
    .Y(_05358_));
 sg13g2_a221oi_1 _22953_ (.B2(_09088_),
    .C1(_05358_),
    .B1(net390),
    .A1(_05357_),
    .Y(_05359_),
    .A2(_04828_));
 sg13g2_nand4_1 _22954_ (.B(_05348_),
    .C(_05356_),
    .A(_05347_),
    .Y(_05360_),
    .D(_05359_));
 sg13g2_nand2_1 _22955_ (.Y(_05361_),
    .A(\cpu.intr.r_timer_count[2] ),
    .B(net532));
 sg13g2_a22oi_1 _22956_ (.Y(_05362_),
    .B1(net593),
    .B2(\cpu.intr.r_clock_cmp[18] ),
    .A2(net447),
    .A1(_10058_));
 sg13g2_inv_1 _22957_ (.Y(_05363_),
    .A(\cpu.intr.r_timer_reload[18] ));
 sg13g2_nor2_1 _22958_ (.A(net901),
    .B(_05363_),
    .Y(_05364_));
 sg13g2_a21oi_1 _22959_ (.A1(net780),
    .A2(\cpu.intr.r_timer_reload[2] ),
    .Y(_05365_),
    .B1(_05364_));
 sg13g2_buf_2 _22960_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05366_));
 sg13g2_a22oi_1 _22961_ (.Y(_05367_),
    .B1(net431),
    .B2(_05366_),
    .A2(net389),
    .A1(_09125_));
 sg13g2_o21ai_1 _22962_ (.B1(_05367_),
    .Y(_05368_),
    .A1(_09906_),
    .A2(_05365_));
 sg13g2_nand2_1 _22963_ (.Y(_05369_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(net561));
 sg13g2_nand3_1 _22964_ (.B(_09935_),
    .C(net442),
    .A(net666),
    .Y(_05370_));
 sg13g2_o21ai_1 _22965_ (.B1(_05370_),
    .Y(_05371_),
    .A1(net666),
    .A2(_05369_));
 sg13g2_nor2_1 _22966_ (.A(_05368_),
    .B(_05371_),
    .Y(_05372_));
 sg13g2_a21oi_1 _22967_ (.A1(_09125_),
    .A2(_04906_),
    .Y(_05373_),
    .B1(net430));
 sg13g2_nand2b_1 _22968_ (.Y(_05374_),
    .B(\cpu.intr.r_timer ),
    .A_N(_05373_));
 sg13g2_nand4_1 _22969_ (.B(_05362_),
    .C(_05372_),
    .A(_05361_),
    .Y(_05375_),
    .D(_05374_));
 sg13g2_and2_1 _22970_ (.A(\cpu.uart.r_in[2] ),
    .B(_04916_),
    .X(_05376_));
 sg13g2_a221oi_1 _22971_ (.B2(_09891_),
    .C1(_05376_),
    .B1(_04918_),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05377_),
    .A2(net427));
 sg13g2_o21ai_1 _22972_ (.B1(_08321_),
    .Y(_05378_),
    .A1(_04914_),
    .A2(_05377_));
 sg13g2_a221oi_1 _22973_ (.B2(_04884_),
    .C1(_05378_),
    .B1(_05375_),
    .A1(_04804_),
    .Y(_05379_),
    .A2(_05360_));
 sg13g2_o21ai_1 _22974_ (.B1(_05379_),
    .Y(_05380_),
    .A1(net800),
    .A2(_05346_));
 sg13g2_nand3_1 _22975_ (.B(_05337_),
    .C(_05380_),
    .A(net71),
    .Y(_05381_));
 sg13g2_o21ai_1 _22976_ (.B1(_05381_),
    .Y(_05382_),
    .A1(_03541_),
    .A2(net73));
 sg13g2_mux2_1 _22977_ (.A0(_05314_),
    .A1(_05382_),
    .S(net82),
    .X(_01031_));
 sg13g2_nor2_1 _22978_ (.A(_05101_),
    .B(_04959_),
    .Y(_05383_));
 sg13g2_a21oi_1 _22979_ (.A1(net740),
    .A2(_04467_),
    .Y(_05384_),
    .B1(_03981_));
 sg13g2_nor2_1 _22980_ (.A(_08441_),
    .B(_04467_),
    .Y(_05385_));
 sg13g2_nand3_1 _22981_ (.B(net740),
    .C(_05385_),
    .A(net270),
    .Y(_05386_));
 sg13g2_o21ai_1 _22982_ (.B1(_05386_),
    .Y(_05387_),
    .A1(net642),
    .A2(_05384_));
 sg13g2_nand3_1 _22983_ (.B(_09112_),
    .C(_04844_),
    .A(_09111_),
    .Y(_05388_));
 sg13g2_buf_1 _22984_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05389_));
 sg13g2_nand2_1 _22985_ (.Y(_05390_),
    .A(net672),
    .B(_05389_));
 sg13g2_o21ai_1 _22986_ (.B1(_05390_),
    .Y(_05391_),
    .A1(net672),
    .A2(_00104_));
 sg13g2_a22oi_1 _22987_ (.Y(_05392_),
    .B1(_05391_),
    .B2(_04811_),
    .A2(net390),
    .A1(_09111_));
 sg13g2_nand2_1 _22988_ (.Y(_05393_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(_10044_));
 sg13g2_o21ai_1 _22989_ (.B1(_05393_),
    .Y(_05394_),
    .A1(_00107_),
    .A2(_04827_));
 sg13g2_inv_1 _22990_ (.Y(_05395_),
    .A(_00106_));
 sg13g2_a22oi_1 _22991_ (.Y(_05396_),
    .B1(_04818_),
    .B2(_05395_),
    .A2(_04808_),
    .A1(_09112_));
 sg13g2_o21ai_1 _22992_ (.B1(_05396_),
    .Y(_05397_),
    .A1(_00105_),
    .A2(net386));
 sg13g2_a21oi_1 _22993_ (.A1(net971),
    .A2(_05394_),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nand3_1 _22994_ (.B(_05392_),
    .C(_05398_),
    .A(_05388_),
    .Y(_05399_));
 sg13g2_nand2_1 _22995_ (.Y(_05400_),
    .A(_04804_),
    .B(_05399_));
 sg13g2_buf_1 _22996_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05401_));
 sg13g2_inv_1 _22997_ (.Y(_05402_),
    .A(_00103_));
 sg13g2_nand2_1 _22998_ (.Y(_05403_),
    .A(\cpu.spi.r_timeout[3] ),
    .B(_05038_));
 sg13g2_o21ai_1 _22999_ (.B1(_05403_),
    .Y(_05404_),
    .A1(_00102_),
    .A2(_04877_));
 sg13g2_a221oi_1 _23000_ (.B2(_05402_),
    .C1(_05404_),
    .B1(net428),
    .A1(_05401_),
    .Y(_05405_),
    .A2(_04857_));
 sg13g2_nand2_1 _23001_ (.Y(_05406_),
    .A(_09186_),
    .B(_04866_));
 sg13g2_a21oi_1 _23002_ (.A1(_05405_),
    .A2(_05406_),
    .Y(_05407_),
    .B1(net800));
 sg13g2_a22oi_1 _23003_ (.Y(_05408_),
    .B1(net559),
    .B2(\cpu.intr.r_timer_reload[19] ),
    .A2(net442),
    .A1(_09934_));
 sg13g2_a221oi_1 _23004_ (.B2(\cpu.intr.r_timer_reload[3] ),
    .C1(net666),
    .B1(net559),
    .A1(\cpu.intr.r_clock_cmp[3] ),
    .Y(_05409_),
    .A2(net561));
 sg13g2_a21oi_1 _23005_ (.A1(net673),
    .A2(_05408_),
    .Y(_05410_),
    .B1(_05409_));
 sg13g2_buf_1 _23006_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05411_));
 sg13g2_a22oi_1 _23007_ (.Y(_05412_),
    .B1(net430),
    .B2(_09120_),
    .A2(net431),
    .A1(_05411_));
 sg13g2_nand2_1 _23008_ (.Y(_05413_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_04979_));
 sg13g2_a22oi_1 _23009_ (.Y(_05414_),
    .B1(_04981_),
    .B2(\cpu.intr.r_timer_count[3] ),
    .A2(net502),
    .A1(_10063_));
 sg13g2_nand3_1 _23010_ (.B(_05413_),
    .C(_05414_),
    .A(_05412_),
    .Y(_05415_));
 sg13g2_nor2_1 _23011_ (.A(_05410_),
    .B(_05415_),
    .Y(_05416_));
 sg13g2_a21oi_1 _23012_ (.A1(_09120_),
    .A2(net388),
    .Y(_05417_),
    .B1(net389));
 sg13g2_nand2b_1 _23013_ (.Y(_05418_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05417_));
 sg13g2_a21oi_1 _23014_ (.A1(_05416_),
    .A2(_05418_),
    .Y(_05419_),
    .B1(net692));
 sg13g2_nand2_1 _23015_ (.Y(_05420_),
    .A(\cpu.uart.r_div_value[11] ),
    .B(_04918_));
 sg13g2_a22oi_1 _23016_ (.Y(_05421_),
    .B1(_04916_),
    .B2(\cpu.uart.r_in[3] ),
    .A2(net427),
    .A1(\cpu.uart.r_div_value[3] ));
 sg13g2_a21oi_1 _23017_ (.A1(_05420_),
    .A2(_05421_),
    .Y(_05422_),
    .B1(net533));
 sg13g2_nor4_1 _23018_ (.A(net902),
    .B(_05407_),
    .C(_05419_),
    .D(_05422_),
    .Y(_05423_));
 sg13g2_a22oi_1 _23019_ (.Y(_05424_),
    .B1(net561),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[2][19] ));
 sg13g2_a22oi_1 _23020_ (.Y(_05425_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][19] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[6][19] ));
 sg13g2_a22oi_1 _23021_ (.Y(_05426_),
    .B1(_02907_),
    .B2(\cpu.dcache.r_data[7][19] ),
    .A2(net482),
    .A1(\cpu.dcache.r_data[3][19] ));
 sg13g2_inv_1 _23022_ (.Y(_05427_),
    .A(_00099_));
 sg13g2_a22oi_1 _23023_ (.Y(_05428_),
    .B1(net503),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net475),
    .A1(_05427_));
 sg13g2_and4_1 _23024_ (.A(_05424_),
    .B(_05425_),
    .C(_05426_),
    .D(_05428_),
    .X(_05429_));
 sg13g2_nand2b_1 _23025_ (.Y(_05430_),
    .B(_04885_),
    .A_N(_05429_));
 sg13g2_nand2_1 _23026_ (.Y(_05431_),
    .A(\cpu.dcache.r_data[3][3] ),
    .B(net482));
 sg13g2_a22oi_1 _23027_ (.Y(_05432_),
    .B1(net474),
    .B2(\cpu.dcache.r_data[2][3] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_a22oi_1 _23028_ (.Y(_05433_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][3] ),
    .A2(net615),
    .A1(\cpu.dcache.r_data[5][3] ));
 sg13g2_a22oi_1 _23029_ (.Y(_05434_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][3] ),
    .A2(net571),
    .A1(\cpu.dcache.r_data[4][3] ));
 sg13g2_nand4_1 _23030_ (.B(_05432_),
    .C(_05433_),
    .A(_05431_),
    .Y(_05435_),
    .D(_05434_));
 sg13g2_mux2_1 _23031_ (.A0(\cpu.dcache.r_data[0][3] ),
    .A1(_05435_),
    .S(net535),
    .X(_05436_));
 sg13g2_nand2_1 _23032_ (.Y(_05437_),
    .A(net601),
    .B(_05436_));
 sg13g2_a21oi_1 _23033_ (.A1(_05430_),
    .A2(_05437_),
    .Y(_05438_),
    .B1(net597));
 sg13g2_nand2_1 _23034_ (.Y(_05439_),
    .A(net972),
    .B(_05436_));
 sg13g2_o21ai_1 _23035_ (.B1(_05439_),
    .Y(_05440_),
    .A1(net972),
    .A2(_05430_));
 sg13g2_nand2_1 _23036_ (.Y(_05441_),
    .A(net1012),
    .B(_05115_));
 sg13g2_a21oi_1 _23037_ (.A1(_05124_),
    .A2(_05441_),
    .Y(_05442_),
    .B1(net596));
 sg13g2_a21oi_1 _23038_ (.A1(net596),
    .A2(_05440_),
    .Y(_05443_),
    .B1(_05442_));
 sg13g2_nor2_1 _23039_ (.A(net663),
    .B(_05443_),
    .Y(_05444_));
 sg13g2_nor3_1 _23040_ (.A(net987),
    .B(_05438_),
    .C(_05444_),
    .Y(_05445_));
 sg13g2_a21oi_1 _23041_ (.A1(_05400_),
    .A2(_05423_),
    .Y(_05446_),
    .B1(_05445_));
 sg13g2_nor2_1 _23042_ (.A(net679),
    .B(net71),
    .Y(_05447_));
 sg13g2_a221oi_1 _23043_ (.B2(_05446_),
    .C1(_05447_),
    .B1(net73),
    .A1(_09083_),
    .Y(_05448_),
    .A2(_11403_));
 sg13g2_a221oi_1 _23044_ (.B2(_04961_),
    .C1(_05448_),
    .B1(_05387_),
    .A1(_04466_),
    .Y(_01032_),
    .A2(_05383_));
 sg13g2_o21ai_1 _23045_ (.B1(net270),
    .Y(_05449_),
    .A1(net665),
    .A2(_05385_));
 sg13g2_mux2_1 _23046_ (.A0(_04182_),
    .A1(_04501_),
    .S(net665),
    .X(_05450_));
 sg13g2_a22oi_1 _23047_ (.Y(_05451_),
    .B1(_05450_),
    .B2(net270),
    .A2(_05449_),
    .A1(_08444_));
 sg13g2_a22oi_1 _23048_ (.Y(_05452_),
    .B1(net537),
    .B2(\cpu.dcache.r_data[5][4] ),
    .A2(net474),
    .A1(\cpu.dcache.r_data[2][4] ));
 sg13g2_a22oi_1 _23049_ (.Y(_05453_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][4] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[6][4] ));
 sg13g2_a22oi_1 _23050_ (.Y(_05454_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][4] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_inv_1 _23051_ (.Y(_05455_),
    .A(_00108_));
 sg13g2_a22oi_1 _23052_ (.Y(_05456_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][4] ),
    .A2(_04757_),
    .A1(_05455_));
 sg13g2_nand4_1 _23053_ (.B(_05453_),
    .C(_05454_),
    .A(_05452_),
    .Y(_05457_),
    .D(_05456_));
 sg13g2_buf_1 _23054_ (.A(_05457_),
    .X(_05458_));
 sg13g2_a22oi_1 _23055_ (.Y(_05459_),
    .B1(net537),
    .B2(\cpu.dcache.r_data[5][20] ),
    .A2(net474),
    .A1(\cpu.dcache.r_data[2][20] ));
 sg13g2_a22oi_1 _23056_ (.Y(_05460_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][20] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[6][20] ));
 sg13g2_a22oi_1 _23057_ (.Y(_05461_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][20] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[3][20] ));
 sg13g2_inv_1 _23058_ (.Y(_05462_),
    .A(_00109_));
 sg13g2_a22oi_1 _23059_ (.Y(_05463_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][20] ),
    .A2(net536),
    .A1(_05462_));
 sg13g2_nand4_1 _23060_ (.B(_05460_),
    .C(_05461_),
    .A(_05459_),
    .Y(_05464_),
    .D(_05463_));
 sg13g2_buf_1 _23061_ (.A(_05464_),
    .X(_05465_));
 sg13g2_a22oi_1 _23062_ (.Y(_05466_),
    .B1(_05465_),
    .B2(_04796_),
    .A2(_05458_),
    .A1(net972));
 sg13g2_a221oi_1 _23063_ (.B2(net672),
    .C1(net596),
    .B1(_05147_),
    .A1(net1012),
    .Y(_05467_),
    .A2(_05141_));
 sg13g2_a21oi_1 _23064_ (.A1(net596),
    .A2(_05466_),
    .Y(_05468_),
    .B1(_05467_));
 sg13g2_nand2_1 _23065_ (.Y(_05469_),
    .A(_03471_),
    .B(_05465_));
 sg13g2_nand2_1 _23066_ (.Y(_05470_),
    .A(_03526_),
    .B(_05458_));
 sg13g2_a21oi_1 _23067_ (.A1(_05469_),
    .A2(_05470_),
    .Y(_05471_),
    .B1(_04752_));
 sg13g2_a21oi_1 _23068_ (.A1(net597),
    .A2(_05468_),
    .Y(_05472_),
    .B1(_05471_));
 sg13g2_a221oi_1 _23069_ (.B2(\cpu.uart.r_in[4] ),
    .C1(net533),
    .B1(_04916_),
    .A1(\cpu.uart.r_div_value[4] ),
    .Y(_05473_),
    .A2(net427));
 sg13g2_and2_1 _23070_ (.A(net915),
    .B(\cpu.intr.r_timer_count[20] ),
    .X(_05474_));
 sg13g2_nor2b_1 _23071_ (.A(net915),
    .B_N(_10068_),
    .Y(_05475_));
 sg13g2_a22oi_1 _23072_ (.Y(_05476_),
    .B1(_05475_),
    .B2(net503),
    .A2(_05474_),
    .A1(net481));
 sg13g2_buf_1 _23073_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05477_));
 sg13g2_inv_1 _23074_ (.Y(_05478_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_nor2_1 _23075_ (.A(net901),
    .B(_05478_),
    .Y(_05479_));
 sg13g2_a21oi_1 _23076_ (.A1(net901),
    .A2(\cpu.intr.r_timer_reload[4] ),
    .Y(_05480_),
    .B1(_05479_));
 sg13g2_nor2_1 _23077_ (.A(_09906_),
    .B(_05480_),
    .Y(_05481_));
 sg13g2_a221oi_1 _23078_ (.B2(_05477_),
    .C1(_05481_),
    .B1(net431),
    .A1(_09118_),
    .Y(_05482_),
    .A2(_04890_));
 sg13g2_a22oi_1 _23079_ (.Y(_05483_),
    .B1(_04976_),
    .B2(\cpu.intr.r_clock_cmp[4] ),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[4] ));
 sg13g2_a21oi_1 _23080_ (.A1(\cpu.intr.r_clock_cmp[20] ),
    .A2(_04901_),
    .Y(_05484_),
    .B1(net388));
 sg13g2_and4_1 _23081_ (.A(_05476_),
    .B(_05482_),
    .C(_05483_),
    .D(_05484_),
    .X(_05485_));
 sg13g2_nand2_1 _23082_ (.Y(_05486_),
    .A(_09362_),
    .B(_04854_));
 sg13g2_a221oi_1 _23083_ (.B2(_05486_),
    .C1(net692),
    .B1(_05485_),
    .A1(_10777_),
    .Y(_05487_),
    .A2(net388));
 sg13g2_nor2_1 _23084_ (.A(_09098_),
    .B(_09117_),
    .Y(_05488_));
 sg13g2_o21ai_1 _23085_ (.B1(_05488_),
    .Y(_05489_),
    .A1(net388),
    .A2(_05485_));
 sg13g2_buf_1 _23086_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05490_));
 sg13g2_inv_1 _23087_ (.Y(_05491_),
    .A(_00113_));
 sg13g2_nand2_1 _23088_ (.Y(_05492_),
    .A(\cpu.spi.r_timeout[4] ),
    .B(_05038_));
 sg13g2_o21ai_1 _23089_ (.B1(_05492_),
    .Y(_05493_),
    .A1(_00112_),
    .A2(_04877_));
 sg13g2_a221oi_1 _23090_ (.B2(_05491_),
    .C1(_05493_),
    .B1(net428),
    .A1(_05490_),
    .Y(_05494_),
    .A2(_04857_));
 sg13g2_nand2_1 _23091_ (.Y(_05495_),
    .A(_09194_),
    .B(_04866_));
 sg13g2_a21oi_1 _23092_ (.A1(_05494_),
    .A2(_05495_),
    .Y(_05496_),
    .B1(net800));
 sg13g2_a21oi_1 _23093_ (.A1(_05487_),
    .A2(_05489_),
    .Y(_05497_),
    .B1(_05496_));
 sg13g2_buf_2 _23094_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05498_));
 sg13g2_nand3_1 _23095_ (.B(_05498_),
    .C(_04909_),
    .A(_11834_),
    .Y(_05499_));
 sg13g2_buf_2 _23096_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05500_));
 sg13g2_a22oi_1 _23097_ (.Y(_05501_),
    .B1(_04823_),
    .B2(_05500_),
    .A2(_04808_),
    .A1(_09091_));
 sg13g2_a22oi_1 _23098_ (.Y(_05502_),
    .B1(net428),
    .B2(_09103_),
    .A2(net390),
    .A1(_09090_));
 sg13g2_buf_2 _23099_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05503_));
 sg13g2_buf_2 _23100_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05504_));
 sg13g2_buf_2 _23101_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05505_));
 sg13g2_mux2_1 _23102_ (.A0(_05504_),
    .A1(_05505_),
    .S(_09245_),
    .X(_05506_));
 sg13g2_a22oi_1 _23103_ (.Y(_05507_),
    .B1(_05506_),
    .B2(_04811_),
    .A2(_04818_),
    .A1(_05503_));
 sg13g2_nand4_1 _23104_ (.B(_05501_),
    .C(_05502_),
    .A(_05499_),
    .Y(_05508_),
    .D(_05507_));
 sg13g2_a21o_1 _23105_ (.A2(net430),
    .A1(_09103_),
    .B1(net472),
    .X(_05509_));
 sg13g2_a22oi_1 _23106_ (.Y(_05510_),
    .B1(net503),
    .B2(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A2(net537),
    .A1(net8));
 sg13g2_buf_2 _23107_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05511_));
 sg13g2_a21oi_1 _23108_ (.A1(_05511_),
    .A2(net561),
    .Y(_05512_),
    .B1(net901));
 sg13g2_a21oi_1 _23109_ (.A1(net780),
    .A2(_05510_),
    .Y(_05513_),
    .B1(_05512_));
 sg13g2_a221oi_1 _23110_ (.B2(_09104_),
    .C1(_05513_),
    .B1(_05509_),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .Y(_05514_),
    .A2(_04896_));
 sg13g2_nand3_1 _23111_ (.B(_09091_),
    .C(_04844_),
    .A(_09090_),
    .Y(_05515_));
 sg13g2_o21ai_1 _23112_ (.B1(_05515_),
    .Y(_05516_),
    .A1(_09741_),
    .A2(_05514_));
 sg13g2_o21ai_1 _23113_ (.B1(_04804_),
    .Y(_05517_),
    .A1(_05508_),
    .A2(_05516_));
 sg13g2_nand3_1 _23114_ (.B(_05497_),
    .C(_05517_),
    .A(net533),
    .Y(_05518_));
 sg13g2_nand3b_1 _23115_ (.B(net987),
    .C(_05518_),
    .Y(_05519_),
    .A_N(_05473_));
 sg13g2_o21ai_1 _23116_ (.B1(_05519_),
    .Y(_05520_),
    .A1(net987),
    .A2(_05472_));
 sg13g2_nand2_1 _23117_ (.Y(_05521_),
    .A(net73),
    .B(_05520_));
 sg13g2_o21ai_1 _23118_ (.B1(_05521_),
    .Y(_05522_),
    .A1(net599),
    .A2(net73));
 sg13g2_mux2_1 _23119_ (.A0(_05451_),
    .A1(_05522_),
    .S(net82),
    .X(_01033_));
 sg13g2_a22oi_1 _23120_ (.Y(_05523_),
    .B1(net559),
    .B2(\cpu.intr.r_timer_reload[21] ),
    .A2(net442),
    .A1(_09929_));
 sg13g2_a221oi_1 _23121_ (.B2(_10073_),
    .C1(net673),
    .B1(net503),
    .A1(\cpu.intr.r_clock_cmp[5] ),
    .Y(_05524_),
    .A2(net561));
 sg13g2_a21o_1 _23122_ (.A2(_05523_),
    .A1(net673),
    .B1(_05524_),
    .X(_05525_));
 sg13g2_buf_2 _23123_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05526_));
 sg13g2_and2_1 _23124_ (.A(_09122_),
    .B(net389),
    .X(_05527_));
 sg13g2_a221oi_1 _23125_ (.B2(\cpu.intr.r_timer_reload[5] ),
    .C1(_05527_),
    .B1(net429),
    .A1(_05526_),
    .Y(_05528_),
    .A2(_04982_));
 sg13g2_a22oi_1 _23126_ (.Y(_05529_),
    .B1(_04981_),
    .B2(\cpu.intr.r_timer_count[5] ),
    .A2(_04979_),
    .A1(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_a21oi_1 _23127_ (.A1(_09122_),
    .A2(net388),
    .Y(_05530_),
    .B1(net430));
 sg13g2_nand2b_1 _23128_ (.Y(_05531_),
    .B(_09121_),
    .A_N(_05530_));
 sg13g2_nand4_1 _23129_ (.B(_05528_),
    .C(_05529_),
    .A(_05525_),
    .Y(_05532_),
    .D(_05531_));
 sg13g2_nor2_1 _23130_ (.A(_00122_),
    .B(_05265_),
    .Y(_05533_));
 sg13g2_nor2_1 _23131_ (.A(_00121_),
    .B(net386),
    .Y(_05534_));
 sg13g2_nand2_1 _23132_ (.Y(_05535_),
    .A(_09114_),
    .B(_04808_));
 sg13g2_o21ai_1 _23133_ (.B1(_05535_),
    .Y(_05536_),
    .A1(_00120_),
    .A2(_05350_));
 sg13g2_nor3_1 _23134_ (.A(_05533_),
    .B(_05534_),
    .C(_05536_),
    .Y(_05537_));
 sg13g2_buf_2 _23135_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05538_));
 sg13g2_nand2_1 _23136_ (.Y(_05539_),
    .A(_05538_),
    .B(_05353_));
 sg13g2_o21ai_1 _23137_ (.B1(_05539_),
    .Y(_05540_),
    .A1(_00123_),
    .A2(_05022_));
 sg13g2_a221oi_1 _23138_ (.B2(_09105_),
    .C1(_05540_),
    .B1(_05035_),
    .A1(_09113_),
    .Y(_05541_),
    .A2(net390));
 sg13g2_inv_1 _23139_ (.Y(_05542_),
    .A(net3));
 sg13g2_a21oi_1 _23140_ (.A1(_09105_),
    .A2(_04909_),
    .Y(_05543_),
    .B1(net472));
 sg13g2_nand2b_1 _23141_ (.Y(_05544_),
    .B(net915),
    .A_N(_00124_));
 sg13g2_nand2_1 _23142_ (.Y(_05545_),
    .A(net901),
    .B(net9));
 sg13g2_a21oi_1 _23143_ (.A1(_05544_),
    .A2(_05545_),
    .Y(_05546_),
    .B1(_09395_));
 sg13g2_a221oi_1 _23144_ (.B2(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .C1(_05546_),
    .B1(net431),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .Y(_05547_),
    .A2(net502));
 sg13g2_o21ai_1 _23145_ (.B1(_05547_),
    .Y(_05548_),
    .A1(_05542_),
    .A2(_05543_));
 sg13g2_nand2_1 _23146_ (.Y(_05549_),
    .A(net971),
    .B(_05548_));
 sg13g2_nand3_1 _23147_ (.B(_09114_),
    .C(_04844_),
    .A(_09113_),
    .Y(_05550_));
 sg13g2_nand4_1 _23148_ (.B(_05541_),
    .C(_05549_),
    .A(_05537_),
    .Y(_05551_),
    .D(_05550_));
 sg13g2_a22oi_1 _23149_ (.Y(_05552_),
    .B1(_04916_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net427),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_buf_1 _23150_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05553_));
 sg13g2_inv_1 _23151_ (.Y(_05554_),
    .A(_00119_));
 sg13g2_nand2_1 _23152_ (.Y(_05555_),
    .A(\cpu.spi.r_timeout[5] ),
    .B(_05038_));
 sg13g2_o21ai_1 _23153_ (.B1(_05555_),
    .Y(_05556_),
    .A1(_00118_),
    .A2(_04877_));
 sg13g2_a221oi_1 _23154_ (.B2(_05554_),
    .C1(_05556_),
    .B1(net428),
    .A1(_05553_),
    .Y(_05557_),
    .A2(_04857_));
 sg13g2_nand2_1 _23155_ (.Y(_05558_),
    .A(_09193_),
    .B(_04866_));
 sg13g2_a21o_1 _23156_ (.A2(_05558_),
    .A1(_05557_),
    .B1(net800),
    .X(_05559_));
 sg13g2_o21ai_1 _23157_ (.B1(_05559_),
    .Y(_05560_),
    .A1(net533),
    .A2(_05552_));
 sg13g2_a221oi_1 _23158_ (.B2(_04804_),
    .C1(_05560_),
    .B1(_05551_),
    .A1(_04884_),
    .Y(_05561_),
    .A2(_05532_));
 sg13g2_a22oi_1 _23159_ (.Y(_05562_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][5] ),
    .A2(net571),
    .A1(\cpu.dcache.r_data[4][5] ));
 sg13g2_a22oi_1 _23160_ (.Y(_05563_),
    .B1(net537),
    .B2(\cpu.dcache.r_data[5][5] ),
    .A2(net474),
    .A1(\cpu.dcache.r_data[2][5] ));
 sg13g2_inv_1 _23161_ (.Y(_05564_),
    .A(_00114_));
 sg13g2_a22oi_1 _23162_ (.Y(_05565_),
    .B1(net481),
    .B2(\cpu.dcache.r_data[6][5] ),
    .A2(net536),
    .A1(_05564_));
 sg13g2_a22oi_1 _23163_ (.Y(_05566_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(net482),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_nand4_1 _23164_ (.B(_05563_),
    .C(_05565_),
    .A(_05562_),
    .Y(_05567_),
    .D(_05566_));
 sg13g2_buf_1 _23165_ (.A(_05567_),
    .X(_05568_));
 sg13g2_a22oi_1 _23166_ (.Y(_05569_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[5][21] ),
    .A2(net616),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_a22oi_1 _23167_ (.Y(_05570_),
    .B1(net563),
    .B2(\cpu.dcache.r_data[2][21] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][21] ));
 sg13g2_a22oi_1 _23168_ (.Y(_05571_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][21] ),
    .A2(net628),
    .A1(\cpu.dcache.r_data[4][21] ));
 sg13g2_inv_1 _23169_ (.Y(_05572_),
    .A(_00115_));
 sg13g2_a22oi_1 _23170_ (.Y(_05573_),
    .B1(net627),
    .B2(\cpu.dcache.r_data[1][21] ),
    .A2(net536),
    .A1(_05572_));
 sg13g2_nand4_1 _23171_ (.B(_05570_),
    .C(_05571_),
    .A(_05569_),
    .Y(_05574_),
    .D(_05573_));
 sg13g2_and2_1 _23172_ (.A(_03471_),
    .B(_05574_),
    .X(_05575_));
 sg13g2_a21oi_1 _23173_ (.A1(net601),
    .A2(_05568_),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_a22oi_1 _23174_ (.Y(_05577_),
    .B1(_05574_),
    .B2(_04796_),
    .A2(_05568_),
    .A1(net972));
 sg13g2_a221oi_1 _23175_ (.B2(_09902_),
    .C1(net667),
    .B1(_05172_),
    .A1(net1012),
    .Y(_05578_),
    .A2(_05166_));
 sg13g2_a21oi_1 _23176_ (.A1(net596),
    .A2(_05577_),
    .Y(_05579_),
    .B1(_05578_));
 sg13g2_nand2_1 _23177_ (.Y(_05580_),
    .A(_04752_),
    .B(_05579_));
 sg13g2_o21ai_1 _23178_ (.B1(_05580_),
    .Y(_05581_),
    .A1(net597),
    .A2(_05576_));
 sg13g2_nor2_1 _23179_ (.A(net987),
    .B(_05581_),
    .Y(_05582_));
 sg13g2_a21oi_1 _23180_ (.A1(net987),
    .A2(_05561_),
    .Y(_05583_),
    .B1(_05582_));
 sg13g2_nor2b_1 _23181_ (.A(_05176_),
    .B_N(_02909_),
    .Y(_05584_));
 sg13g2_a21oi_1 _23182_ (.A1(net73),
    .A2(_05583_),
    .Y(_05585_),
    .B1(_05584_));
 sg13g2_and2_1 _23183_ (.A(net740),
    .B(_04535_),
    .X(_05586_));
 sg13g2_a21oi_1 _23184_ (.A1(net665),
    .A2(_04532_),
    .Y(_05587_),
    .B1(_05586_));
 sg13g2_nor3_1 _23185_ (.A(net977),
    .B(_05206_),
    .C(_05101_),
    .Y(_05588_));
 sg13g2_a221oi_1 _23186_ (.B2(_05102_),
    .C1(_05588_),
    .B1(_05587_),
    .A1(net82),
    .Y(_01034_),
    .A2(_05585_));
 sg13g2_nand2_1 _23187_ (.Y(_05589_),
    .A(_04964_),
    .B(_04564_));
 sg13g2_o21ai_1 _23188_ (.B1(_05589_),
    .Y(_05590_),
    .A1(_04964_),
    .A2(_04561_));
 sg13g2_mux2_1 _23189_ (.A0(net976),
    .A1(_05590_),
    .S(net270),
    .X(_05591_));
 sg13g2_a22oi_1 _23190_ (.Y(_05592_),
    .B1(net615),
    .B2(\cpu.dcache.r_data[5][22] ),
    .A2(net474),
    .A1(\cpu.dcache.r_data[2][22] ));
 sg13g2_a22oi_1 _23191_ (.Y(_05593_),
    .B1(net564),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net560),
    .A1(\cpu.dcache.r_data[6][22] ));
 sg13g2_a22oi_1 _23192_ (.Y(_05594_),
    .B1(net614),
    .B2(\cpu.dcache.r_data[7][22] ),
    .A2(net562),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_inv_1 _23193_ (.Y(_05595_),
    .A(_00126_));
 sg13g2_a22oi_1 _23194_ (.Y(_05596_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][22] ),
    .A2(net536),
    .A1(_05595_));
 sg13g2_and4_1 _23195_ (.A(_05592_),
    .B(_05593_),
    .C(_05594_),
    .D(_05596_),
    .X(_05597_));
 sg13g2_buf_1 _23196_ (.A(_05597_),
    .X(_05598_));
 sg13g2_a22oi_1 _23197_ (.Y(_05599_),
    .B1(net537),
    .B2(\cpu.dcache.r_data[5][6] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_a22oi_1 _23198_ (.Y(_05600_),
    .B1(net484),
    .B2(\cpu.dcache.r_data[1][6] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[6][6] ));
 sg13g2_a22oi_1 _23199_ (.Y(_05601_),
    .B1(net559),
    .B2(\cpu.dcache.r_data[7][6] ),
    .A2(net482),
    .A1(\cpu.dcache.r_data[3][6] ));
 sg13g2_inv_1 _23200_ (.Y(_05602_),
    .A(_00125_));
 sg13g2_a22oi_1 _23201_ (.Y(_05603_),
    .B1(net571),
    .B2(\cpu.dcache.r_data[4][6] ),
    .A2(net475),
    .A1(_05602_));
 sg13g2_and4_1 _23202_ (.A(_05599_),
    .B(_05600_),
    .C(_05601_),
    .D(_05603_),
    .X(_05604_));
 sg13g2_buf_1 _23203_ (.A(_05604_),
    .X(_05605_));
 sg13g2_and2_1 _23204_ (.A(_03526_),
    .B(_05605_),
    .X(_05606_));
 sg13g2_a21oi_1 _23205_ (.A1(net609),
    .A2(_05598_),
    .Y(_05607_),
    .B1(_05606_));
 sg13g2_nand2_1 _23206_ (.Y(_05608_),
    .A(_04885_),
    .B(net667));
 sg13g2_nand2b_1 _23207_ (.Y(_05609_),
    .B(_05192_),
    .A_N(_04776_));
 sg13g2_o21ai_1 _23208_ (.B1(_05609_),
    .Y(_05610_),
    .A1(_05608_),
    .A2(_05598_));
 sg13g2_nor2_1 _23209_ (.A(_05076_),
    .B(_05605_),
    .Y(_05611_));
 sg13g2_a221oi_1 _23210_ (.B2(net1012),
    .C1(_05611_),
    .B1(_05610_),
    .A1(_05083_),
    .Y(_05612_),
    .A2(_05199_));
 sg13g2_nand2_1 _23211_ (.Y(_05613_),
    .A(net597),
    .B(_05612_));
 sg13g2_o21ai_1 _23212_ (.B1(_05613_),
    .Y(_05614_),
    .A1(_04753_),
    .A2(_05607_));
 sg13g2_buf_2 _23213_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05615_));
 sg13g2_mux2_1 _23214_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .S(net915),
    .X(_05616_));
 sg13g2_a22oi_1 _23215_ (.Y(_05617_),
    .B1(_05616_),
    .B2(net559),
    .A2(net431),
    .A1(_05615_));
 sg13g2_nand2_1 _23216_ (.Y(_05618_),
    .A(_10079_),
    .B(net502));
 sg13g2_a22oi_1 _23217_ (.Y(_05619_),
    .B1(net561),
    .B2(\cpu.intr.r_clock_cmp[22] ),
    .A2(net442),
    .A1(_09931_));
 sg13g2_nand2b_1 _23218_ (.Y(_05620_),
    .B(net797),
    .A_N(_05619_));
 sg13g2_a22oi_1 _23219_ (.Y(_05621_),
    .B1(_04976_),
    .B2(\cpu.intr.r_clock_cmp[6] ),
    .A2(_04868_),
    .A1(\cpu.intr.r_timer_count[6] ));
 sg13g2_nand4_1 _23220_ (.B(_05618_),
    .C(_05620_),
    .A(_05617_),
    .Y(_05622_),
    .D(_05621_));
 sg13g2_a22oi_1 _23221_ (.Y(_05623_),
    .B1(_04895_),
    .B2(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A2(net472),
    .A1(_09101_));
 sg13g2_o21ai_1 _23222_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_00135_),
    .A2(_04827_));
 sg13g2_a221oi_1 _23223_ (.B2(net10),
    .C1(_05624_),
    .B1(_04976_),
    .A1(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .Y(_05625_),
    .A2(_10044_));
 sg13g2_nand2b_1 _23224_ (.Y(_05626_),
    .B(net971),
    .A_N(_05625_));
 sg13g2_nand3_1 _23225_ (.B(net971),
    .C(_04908_),
    .A(_09101_),
    .Y(_05627_));
 sg13g2_nand2b_1 _23226_ (.Y(_05628_),
    .B(_05627_),
    .A_N(_05035_));
 sg13g2_nor2_1 _23227_ (.A(_09901_),
    .B(_00131_),
    .Y(_05629_));
 sg13g2_buf_1 _23228_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05630_));
 sg13g2_nor2b_1 _23229_ (.A(_09245_),
    .B_N(_05630_),
    .Y(_05631_));
 sg13g2_o21ai_1 _23230_ (.B1(_04811_),
    .Y(_05632_),
    .A1(_05629_),
    .A2(_05631_));
 sg13g2_o21ai_1 _23231_ (.B1(_05632_),
    .Y(_05633_),
    .A1(_00134_),
    .A2(_05022_));
 sg13g2_a21oi_1 _23232_ (.A1(\cpu.gpio.r_enable_io[6] ),
    .A2(_05628_),
    .Y(_05634_),
    .B1(_05633_));
 sg13g2_inv_1 _23233_ (.Y(_05635_),
    .A(_00132_));
 sg13g2_nand2_1 _23234_ (.Y(_05636_),
    .A(_09100_),
    .B(_04808_));
 sg13g2_o21ai_1 _23235_ (.B1(_05636_),
    .Y(_05637_),
    .A1(_00133_),
    .A2(_05265_));
 sg13g2_a221oi_1 _23236_ (.B2(_09099_),
    .C1(_05637_),
    .B1(net390),
    .A1(_05635_),
    .Y(_05638_),
    .A2(_04823_));
 sg13g2_nand3_1 _23237_ (.B(_09100_),
    .C(_04844_),
    .A(_09099_),
    .Y(_05639_));
 sg13g2_nand4_1 _23238_ (.B(_05634_),
    .C(_05638_),
    .A(_05626_),
    .Y(_05640_),
    .D(_05639_));
 sg13g2_buf_1 _23239_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05641_));
 sg13g2_inv_1 _23240_ (.Y(_05642_),
    .A(_00130_));
 sg13g2_nand2_1 _23241_ (.Y(_05643_),
    .A(\cpu.spi.r_timeout[6] ),
    .B(_05038_));
 sg13g2_o21ai_1 _23242_ (.B1(_05643_),
    .Y(_05644_),
    .A1(_00129_),
    .A2(_04877_));
 sg13g2_a221oi_1 _23243_ (.B2(_05642_),
    .C1(_05644_),
    .B1(net428),
    .A1(_05641_),
    .Y(_05645_),
    .A2(_04857_));
 sg13g2_nand2_1 _23244_ (.Y(_05646_),
    .A(_09187_),
    .B(_04866_));
 sg13g2_a21oi_1 _23245_ (.A1(_05645_),
    .A2(_05646_),
    .Y(_05647_),
    .B1(net800));
 sg13g2_a221oi_1 _23246_ (.B2(_04804_),
    .C1(_05647_),
    .B1(_05640_),
    .A1(_05004_),
    .Y(_05648_),
    .A2(_05622_));
 sg13g2_a221oi_1 _23247_ (.B2(\cpu.uart.r_in[6] ),
    .C1(net533),
    .B1(_04916_),
    .A1(\cpu.uart.r_div_value[6] ),
    .Y(_05649_),
    .A2(net427));
 sg13g2_a21oi_1 _23248_ (.A1(_04914_),
    .A2(_05648_),
    .Y(_05650_),
    .B1(_05649_));
 sg13g2_nand2_1 _23249_ (.Y(_05651_),
    .A(net987),
    .B(_05650_));
 sg13g2_o21ai_1 _23250_ (.B1(_05651_),
    .Y(_05652_),
    .A1(net987),
    .A2(_05614_));
 sg13g2_nand2_1 _23251_ (.Y(_05653_),
    .A(net71),
    .B(_05652_));
 sg13g2_o21ai_1 _23252_ (.B1(_05653_),
    .Y(_05654_),
    .A1(_02919_),
    .A2(net73));
 sg13g2_mux2_1 _23253_ (.A0(_05591_),
    .A1(_05654_),
    .S(net82),
    .X(_01035_));
 sg13g2_nand2_1 _23254_ (.Y(_05655_),
    .A(net664),
    .B(_04591_));
 sg13g2_o21ai_1 _23255_ (.B1(_05655_),
    .Y(_05656_),
    .A1(net664),
    .A2(_04588_));
 sg13g2_nand2_1 _23256_ (.Y(_05657_),
    .A(net71),
    .B(_05090_));
 sg13g2_o21ai_1 _23257_ (.B1(_05657_),
    .Y(_05658_),
    .A1(_09155_),
    .A2(net71));
 sg13g2_nand3_1 _23258_ (.B(net352),
    .C(net86),
    .A(net975),
    .Y(_05659_));
 sg13g2_o21ai_1 _23259_ (.B1(_05659_),
    .Y(_05660_),
    .A1(net86),
    .A2(_05658_));
 sg13g2_a21o_1 _23260_ (.A2(_05656_),
    .A1(_05102_),
    .B1(_05660_),
    .X(_01036_));
 sg13g2_nand3_1 _23261_ (.B(_04593_),
    .C(_04620_),
    .A(net665),
    .Y(_05661_));
 sg13g2_a21oi_1 _23262_ (.A1(_04965_),
    .A2(_04622_),
    .Y(_05662_),
    .B1(_04967_));
 sg13g2_a22oi_1 _23263_ (.Y(_05663_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(net429),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_a22oi_1 _23264_ (.Y(_05664_),
    .B1(net532),
    .B2(_09916_),
    .A2(net447),
    .A1(_10088_));
 sg13g2_buf_2 _23265_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05665_));
 sg13g2_a22oi_1 _23266_ (.Y(_05666_),
    .B1(net387),
    .B2(_05665_),
    .A2(net593),
    .A1(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_nand3_1 _23267_ (.B(_05664_),
    .C(_05666_),
    .A(_05663_),
    .Y(_05667_));
 sg13g2_o21ai_1 _23268_ (.B1(_04794_),
    .Y(_05668_),
    .A1(net601),
    .A2(_04786_));
 sg13g2_a22oi_1 _23269_ (.Y(_05669_),
    .B1(_05668_),
    .B2(net663),
    .A2(_05667_),
    .A1(_04973_));
 sg13g2_o21ai_1 _23270_ (.B1(_05093_),
    .Y(_05670_),
    .A1(net983),
    .A2(_05669_));
 sg13g2_nor2_1 _23271_ (.A(net34),
    .B(_05670_),
    .Y(_05671_));
 sg13g2_a21oi_1 _23272_ (.A1(_02925_),
    .A2(net34),
    .Y(_05672_),
    .B1(_05671_));
 sg13g2_o21ai_1 _23273_ (.B1(_05672_),
    .Y(_05673_),
    .A1(\cpu.ex.pc[8] ),
    .A2(_04969_));
 sg13g2_a21oi_1 _23274_ (.A1(_05661_),
    .A2(_05662_),
    .Y(_01037_),
    .B1(_05673_));
 sg13g2_a22oi_1 _23275_ (.Y(_05674_),
    .B1(net429),
    .B2(\cpu.intr.r_timer_reload[9] ),
    .A2(net532),
    .A1(\cpu.intr.r_timer_count[9] ));
 sg13g2_a22oi_1 _23276_ (.Y(_05675_),
    .B1(net593),
    .B2(\cpu.intr.r_clock_cmp[25] ),
    .A2(net447),
    .A1(_10095_));
 sg13g2_buf_2 _23277_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05676_));
 sg13g2_a22oi_1 _23278_ (.Y(_05677_),
    .B1(net594),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(net387),
    .A1(_05676_));
 sg13g2_nand3_1 _23279_ (.B(_05675_),
    .C(_05677_),
    .A(_05674_),
    .Y(_05678_));
 sg13g2_o21ai_1 _23280_ (.B1(_05258_),
    .Y(_05679_),
    .A1(net601),
    .A2(_05250_));
 sg13g2_a22oi_1 _23281_ (.Y(_05680_),
    .B1(_05679_),
    .B2(net663),
    .A2(_05678_),
    .A1(_04973_));
 sg13g2_o21ai_1 _23282_ (.B1(_05093_),
    .Y(_05681_),
    .A1(net983),
    .A2(_05680_));
 sg13g2_nor2_1 _23283_ (.A(net34),
    .B(_05681_),
    .Y(_05682_));
 sg13g2_a21oi_1 _23284_ (.A1(_02928_),
    .A2(net34),
    .Y(_05683_),
    .B1(_05682_));
 sg13g2_o21ai_1 _23285_ (.B1(_05683_),
    .Y(_05684_),
    .A1(net974),
    .A2(_04969_));
 sg13g2_a21oi_1 _23286_ (.A1(net740),
    .A2(_04649_),
    .Y(_05685_),
    .B1(_04967_));
 sg13g2_o21ai_1 _23287_ (.B1(_05685_),
    .Y(_05686_),
    .A1(net664),
    .A2(_04647_));
 sg13g2_nor2b_1 _23288_ (.A(_05684_),
    .B_N(_05686_),
    .Y(_01038_));
 sg13g2_nand2b_1 _23289_ (.Y(_05687_),
    .B(\cpu.dec.r_rd[0] ),
    .A_N(_03416_));
 sg13g2_a21oi_1 _23290_ (.A1(net270),
    .A2(_05687_),
    .Y(_05688_),
    .B1(_05101_));
 sg13g2_a21o_1 _23291_ (.A2(net82),
    .A1(_10144_),
    .B1(_05688_),
    .X(_01039_));
 sg13g2_buf_1 _23292_ (.A(net86),
    .X(_05689_));
 sg13g2_nor2b_1 _23293_ (.A(_03416_),
    .B_N(\cpu.dec.r_rd[1] ),
    .Y(_05690_));
 sg13g2_buf_1 _23294_ (.A(net86),
    .X(_05691_));
 sg13g2_o21ai_1 _23295_ (.B1(_05691_),
    .Y(_05692_),
    .A1(net352),
    .A2(_05690_));
 sg13g2_o21ai_1 _23296_ (.B1(_05692_),
    .Y(_01040_),
    .A1(_03490_),
    .A2(net70));
 sg13g2_nor3_1 _23297_ (.A(_03416_),
    .B(_09231_),
    .C(_03981_),
    .Y(_05693_));
 sg13g2_nand3_1 _23298_ (.B(_11406_),
    .C(_05693_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05694_));
 sg13g2_o21ai_1 _23299_ (.B1(_05694_),
    .Y(_01041_),
    .A1(_11374_),
    .A2(_05689_));
 sg13g2_nand3_1 _23300_ (.B(_11406_),
    .C(_05693_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05695_));
 sg13g2_o21ai_1 _23301_ (.B1(_05695_),
    .Y(_01042_),
    .A1(_10139_),
    .A2(_05689_));
 sg13g2_mux2_1 _23302_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05155_),
    .X(_01043_));
 sg13g2_buf_1 _23303_ (.A(net570),
    .X(_05696_));
 sg13g2_a22oi_1 _23304_ (.Y(_05697_),
    .B1(net501),
    .B2(_10564_),
    .A2(net471),
    .A1(_03455_));
 sg13g2_nor2_1 _23305_ (.A(net865),
    .B(net69),
    .Y(_05698_));
 sg13g2_a21oi_1 _23306_ (.A1(_05697_),
    .A2(net70),
    .Y(_01044_),
    .B1(_05698_));
 sg13g2_a221oi_1 _23307_ (.B2(_10385_),
    .C1(net983),
    .B1(net501),
    .A1(_10368_),
    .Y(_05699_),
    .A2(net471));
 sg13g2_a21oi_1 _23308_ (.A1(net854),
    .A2(_10538_),
    .Y(_05700_),
    .B1(_05699_));
 sg13g2_mux2_1 _23309_ (.A0(_10099_),
    .A1(_05700_),
    .S(net72),
    .X(_01045_));
 sg13g2_a22oi_1 _23310_ (.Y(_05701_),
    .B1(net501),
    .B2(_10512_),
    .A2(net471),
    .A1(_09166_));
 sg13g2_a221oi_1 _23311_ (.B2(_10712_),
    .C1(_03010_),
    .B1(_10251_),
    .A1(_10693_),
    .Y(_05702_),
    .A2(net471));
 sg13g2_a21oi_1 _23312_ (.A1(net854),
    .A2(_05701_),
    .Y(_05703_),
    .B1(_05702_));
 sg13g2_mux2_1 _23313_ (.A0(_10105_),
    .A1(_05703_),
    .S(net72),
    .X(_01046_));
 sg13g2_a21oi_2 _23314_ (.B1(_10653_),
    .Y(_05704_),
    .A2(net471),
    .A1(net551));
 sg13g2_a221oi_1 _23315_ (.B2(_10684_),
    .C1(net983),
    .B1(_10251_),
    .A1(net695),
    .Y(_05705_),
    .A2(_05696_));
 sg13g2_a21oi_1 _23316_ (.A1(net854),
    .A2(_05704_),
    .Y(_05706_),
    .B1(_05705_));
 sg13g2_mux2_1 _23317_ (.A0(_10113_),
    .A1(_05706_),
    .S(net72),
    .X(_01047_));
 sg13g2_a22oi_1 _23318_ (.Y(_05707_),
    .B1(net501),
    .B2(_10625_),
    .A2(net471),
    .A1(_02909_));
 sg13g2_nand2_1 _23319_ (.Y(_05708_),
    .A(_11784_),
    .B(_10420_));
 sg13g2_o21ai_1 _23320_ (.B1(_05708_),
    .Y(_05709_),
    .A1(_11784_),
    .A2(_05707_));
 sg13g2_mux2_1 _23321_ (.A0(_10119_),
    .A1(_05709_),
    .S(net72),
    .X(_01048_));
 sg13g2_a22oi_1 _23322_ (.Y(_05710_),
    .B1(net501),
    .B2(_10359_),
    .A2(net471),
    .A1(_09151_));
 sg13g2_nand2b_1 _23323_ (.Y(_05711_),
    .B(net854),
    .A_N(_05710_));
 sg13g2_o21ai_1 _23324_ (.B1(_05711_),
    .Y(_05712_),
    .A1(net854),
    .A2(_10287_));
 sg13g2_mux2_1 _23325_ (.A0(_10125_),
    .A1(_05712_),
    .S(net72),
    .X(_01049_));
 sg13g2_mux2_1 _23326_ (.A0(_10240_),
    .A1(_10478_),
    .S(net854),
    .X(_05713_));
 sg13g2_mux2_1 _23327_ (.A0(_10130_),
    .A1(_05713_),
    .S(_04961_),
    .X(_01050_));
 sg13g2_nand2_1 _23328_ (.Y(_05714_),
    .A(_03472_),
    .B(net471));
 sg13g2_and2_1 _23329_ (.A(_10594_),
    .B(_05714_),
    .X(_05715_));
 sg13g2_nor2_1 _23330_ (.A(net1040),
    .B(net69),
    .Y(_05716_));
 sg13g2_a21oi_1 _23331_ (.A1(_05715_),
    .A2(net70),
    .Y(_01051_),
    .B1(_05716_));
 sg13g2_nor2_1 _23332_ (.A(net898),
    .B(net69),
    .Y(_05717_));
 sg13g2_a21oi_1 _23333_ (.A1(_10538_),
    .A2(net70),
    .Y(_01052_),
    .B1(_05717_));
 sg13g2_nor2_1 _23334_ (.A(_10062_),
    .B(net69),
    .Y(_05718_));
 sg13g2_a21oi_1 _23335_ (.A1(_05701_),
    .A2(net70),
    .Y(_01053_),
    .B1(_05718_));
 sg13g2_nor2_1 _23336_ (.A(net1043),
    .B(net69),
    .Y(_05719_));
 sg13g2_a21oi_1 _23337_ (.A1(_05704_),
    .A2(net70),
    .Y(_01054_),
    .B1(_05719_));
 sg13g2_nor2_1 _23338_ (.A(net1042),
    .B(net69),
    .Y(_05720_));
 sg13g2_a21oi_1 _23339_ (.A1(_05707_),
    .A2(net70),
    .Y(_01055_),
    .B1(_05720_));
 sg13g2_nor2_1 _23340_ (.A(_10078_),
    .B(net69),
    .Y(_05721_));
 sg13g2_a21oi_1 _23341_ (.A1(_05710_),
    .A2(net70),
    .Y(_01056_),
    .B1(_05721_));
 sg13g2_nand2_1 _23342_ (.Y(_05722_),
    .A(_10478_),
    .B(net69));
 sg13g2_o21ai_1 _23343_ (.B1(_05722_),
    .Y(_01057_),
    .A1(_12648_),
    .A2(net72));
 sg13g2_o21ai_1 _23344_ (.B1(_11784_),
    .Y(_05723_),
    .A1(_10452_),
    .A2(_10453_));
 sg13g2_o21ai_1 _23345_ (.B1(_05723_),
    .Y(_05724_),
    .A1(_11784_),
    .A2(_05697_));
 sg13g2_mux2_1 _23346_ (.A0(_10087_),
    .A1(_05724_),
    .S(net72),
    .X(_01058_));
 sg13g2_a221oi_1 _23347_ (.B2(_10323_),
    .C1(net983),
    .B1(net501),
    .A1(_10297_),
    .Y(_05725_),
    .A2(_05696_));
 sg13g2_a21oi_1 _23348_ (.A1(net854),
    .A2(_05715_),
    .Y(_05726_),
    .B1(_05725_));
 sg13g2_mux2_1 _23349_ (.A0(_10094_),
    .A1(_05726_),
    .S(_05691_),
    .X(_01059_));
 sg13g2_mux2_1 _23350_ (.A0(net695),
    .A1(_08408_),
    .S(_08398_),
    .X(_05727_));
 sg13g2_nor3_1 _23351_ (.A(_10550_),
    .B(_10542_),
    .C(_10488_),
    .Y(_05728_));
 sg13g2_inv_1 _23352_ (.Y(_05729_),
    .A(_05728_));
 sg13g2_o21ai_1 _23353_ (.B1(_03312_),
    .Y(_05730_),
    .A1(_10597_),
    .A2(_05729_));
 sg13g2_buf_2 _23354_ (.A(_05730_),
    .X(_05731_));
 sg13g2_nor4_1 _23355_ (.A(_08286_),
    .B(_04692_),
    .C(_10141_),
    .D(_03491_),
    .Y(_05732_));
 sg13g2_buf_2 _23356_ (.A(_05732_),
    .X(_05733_));
 sg13g2_buf_1 _23357_ (.A(_00269_),
    .X(_05734_));
 sg13g2_nand2b_1 _23358_ (.Y(_05735_),
    .B(net981),
    .A_N(net1086));
 sg13g2_o21ai_1 _23359_ (.B1(_05735_),
    .Y(_05736_),
    .A1(net981),
    .A2(net695));
 sg13g2_nand3_1 _23360_ (.B(_05733_),
    .C(_05736_),
    .A(_05731_),
    .Y(_05737_));
 sg13g2_mux2_1 _23361_ (.A0(_05727_),
    .A1(_05737_),
    .S(net391),
    .X(_05738_));
 sg13g2_nor2_1 _23362_ (.A(net796),
    .B(_05738_),
    .Y(_05739_));
 sg13g2_buf_1 _23363_ (.A(_10676_),
    .X(_05740_));
 sg13g2_nand2_2 _23364_ (.Y(_05741_),
    .A(_05731_),
    .B(_05733_));
 sg13g2_a21oi_2 _23365_ (.B1(_09231_),
    .Y(_05742_),
    .A2(_05741_),
    .A1(net391));
 sg13g2_nor2_1 _23366_ (.A(net970),
    .B(_05742_),
    .Y(_05743_));
 sg13g2_nor2_1 _23367_ (.A(_05739_),
    .B(_05743_),
    .Y(_01062_));
 sg13g2_mux2_1 _23368_ (.A0(_09563_),
    .A1(_08416_),
    .S(_08398_),
    .X(_05744_));
 sg13g2_and2_1 _23369_ (.A(_10676_),
    .B(_10401_),
    .X(_05745_));
 sg13g2_buf_2 _23370_ (.A(_05745_),
    .X(_05746_));
 sg13g2_buf_1 _23371_ (.A(_10401_),
    .X(_05747_));
 sg13g2_nor2_2 _23372_ (.A(_05740_),
    .B(_05747_),
    .Y(_05748_));
 sg13g2_o21ai_1 _23373_ (.B1(net981),
    .Y(_05749_),
    .A1(_05746_),
    .A2(_05748_));
 sg13g2_o21ai_1 _23374_ (.B1(_05749_),
    .Y(_05750_),
    .A1(net981),
    .A2(_09563_));
 sg13g2_nand3_1 _23375_ (.B(_05733_),
    .C(_05750_),
    .A(_05731_),
    .Y(_05751_));
 sg13g2_mux2_1 _23376_ (.A0(_05744_),
    .A1(_05751_),
    .S(net391),
    .X(_05752_));
 sg13g2_nor2_1 _23377_ (.A(net796),
    .B(_05752_),
    .Y(_05753_));
 sg13g2_nor2_1 _23378_ (.A(net969),
    .B(_05742_),
    .Y(_05754_));
 sg13g2_nor2_1 _23379_ (.A(_05753_),
    .B(_05754_),
    .Y(_01063_));
 sg13g2_buf_1 _23380_ (.A(_10275_),
    .X(_05755_));
 sg13g2_inv_1 _23381_ (.Y(_05756_),
    .A(net968));
 sg13g2_nand2_1 _23382_ (.Y(_05757_),
    .A(_10676_),
    .B(_10401_));
 sg13g2_buf_2 _23383_ (.A(_05757_),
    .X(_05758_));
 sg13g2_nor2_2 _23384_ (.A(net848),
    .B(_05758_),
    .Y(_05759_));
 sg13g2_buf_1 _23385_ (.A(net968),
    .X(_05760_));
 sg13g2_nor2_1 _23386_ (.A(net847),
    .B(_05746_),
    .Y(_05761_));
 sg13g2_o21ai_1 _23387_ (.B1(_03454_),
    .Y(_05762_),
    .A1(_05759_),
    .A2(_05761_));
 sg13g2_o21ai_1 _23388_ (.B1(_05762_),
    .Y(_05763_),
    .A1(_03454_),
    .A2(net783));
 sg13g2_nand2b_1 _23389_ (.Y(_05764_),
    .B(_05763_),
    .A_N(_05741_));
 sg13g2_nand2_1 _23390_ (.Y(_05765_),
    .A(_08424_),
    .B(_08398_));
 sg13g2_o21ai_1 _23391_ (.B1(_05765_),
    .Y(_05766_),
    .A1(net600),
    .A2(_08398_));
 sg13g2_mux2_1 _23392_ (.A0(_05764_),
    .A1(_05766_),
    .S(_08405_),
    .X(_05767_));
 sg13g2_nor2_1 _23393_ (.A(net796),
    .B(_05767_),
    .Y(_05768_));
 sg13g2_nor2_1 _23394_ (.A(net847),
    .B(_05742_),
    .Y(_05769_));
 sg13g2_nor2_1 _23395_ (.A(_05768_),
    .B(_05769_),
    .Y(_01064_));
 sg13g2_nor2_1 _23396_ (.A(net904),
    .B(_08398_),
    .Y(_05770_));
 sg13g2_a21oi_1 _23397_ (.A1(_08422_),
    .A2(_08398_),
    .Y(_05771_),
    .B1(_05770_));
 sg13g2_buf_1 _23398_ (.A(_10192_),
    .X(_05772_));
 sg13g2_xnor2_1 _23399_ (.Y(_05773_),
    .A(_05772_),
    .B(_05759_));
 sg13g2_nand2_1 _23400_ (.Y(_05774_),
    .A(net981),
    .B(_05773_));
 sg13g2_o21ai_1 _23401_ (.B1(_05774_),
    .Y(_05775_),
    .A1(net981),
    .A2(net904));
 sg13g2_nand4_1 _23402_ (.B(_05731_),
    .C(_05733_),
    .A(net391),
    .Y(_05776_),
    .D(_05775_));
 sg13g2_o21ai_1 _23403_ (.B1(_05776_),
    .Y(_05777_),
    .A1(net391),
    .A2(_05771_));
 sg13g2_nor2_1 _23404_ (.A(net967),
    .B(_05742_),
    .Y(_05778_));
 sg13g2_a21oi_1 _23405_ (.A1(_09084_),
    .A2(_05777_),
    .Y(_01065_),
    .B1(_05778_));
 sg13g2_buf_1 _23406_ (.A(net551),
    .X(_05779_));
 sg13g2_buf_2 _23407_ (.A(_00170_),
    .X(_05780_));
 sg13g2_nor2_1 _23408_ (.A(net1113),
    .B(_10192_),
    .Y(_05781_));
 sg13g2_buf_2 _23409_ (.A(_05781_),
    .X(_05782_));
 sg13g2_nand2_1 _23410_ (.Y(_05783_),
    .A(_05780_),
    .B(_05782_));
 sg13g2_nand3b_1 _23411_ (.B(_05733_),
    .C(_08332_),
    .Y(_05784_),
    .A_N(_10505_));
 sg13g2_buf_1 _23412_ (.A(_05784_),
    .X(_05785_));
 sg13g2_or3_1 _23413_ (.A(net970),
    .B(net969),
    .C(_05785_),
    .X(_05786_));
 sg13g2_buf_1 _23414_ (.A(_05786_),
    .X(_05787_));
 sg13g2_nor2_1 _23415_ (.A(_05783_),
    .B(_05787_),
    .Y(_05788_));
 sg13g2_buf_1 _23416_ (.A(_05788_),
    .X(_05789_));
 sg13g2_buf_1 _23417_ (.A(_05789_),
    .X(_05790_));
 sg13g2_mux2_1 _23418_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(net470),
    .S(net269),
    .X(_01133_));
 sg13g2_mux2_1 _23419_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(_03469_),
    .S(net269),
    .X(_01134_));
 sg13g2_buf_1 _23420_ (.A(net904),
    .X(_05791_));
 sg13g2_mux2_1 _23421_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(_05791_),
    .S(net269),
    .X(_01135_));
 sg13g2_buf_1 _23422_ (.A(net668),
    .X(_05792_));
 sg13g2_mux2_1 _23423_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net592),
    .S(net269),
    .X(_01136_));
 sg13g2_mux2_1 _23424_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(net743),
    .S(net269),
    .X(_01137_));
 sg13g2_mux2_1 _23425_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net742),
    .S(_05790_),
    .X(_01138_));
 sg13g2_mux2_1 _23426_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net850),
    .S(_05790_),
    .X(_01139_));
 sg13g2_mux2_1 _23427_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net849),
    .S(net269),
    .X(_01140_));
 sg13g2_mux2_1 _23428_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net851),
    .S(net269),
    .X(_01141_));
 sg13g2_mux2_1 _23429_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net852),
    .S(net269),
    .X(_01142_));
 sg13g2_mux2_1 _23430_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(net540),
    .S(_05789_),
    .X(_01143_));
 sg13g2_mux2_1 _23431_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net547),
    .S(_05789_),
    .X(_01144_));
 sg13g2_buf_1 _23432_ (.A(_05785_),
    .X(_05793_));
 sg13g2_nand2b_1 _23433_ (.Y(_05794_),
    .B(_05747_),
    .A_N(_10676_));
 sg13g2_buf_1 _23434_ (.A(_05794_),
    .X(_05795_));
 sg13g2_inv_1 _23435_ (.Y(_05796_),
    .A(net1113));
 sg13g2_nand2_1 _23436_ (.Y(_05797_),
    .A(_05796_),
    .B(_05772_));
 sg13g2_buf_2 _23437_ (.A(_05797_),
    .X(_05798_));
 sg13g2_nor3_2 _23438_ (.A(net968),
    .B(net738),
    .C(_05798_),
    .Y(_05799_));
 sg13g2_nor2b_1 _23439_ (.A(net469),
    .B_N(_05799_),
    .Y(_05800_));
 sg13g2_buf_1 _23440_ (.A(_05800_),
    .X(_05801_));
 sg13g2_buf_1 _23441_ (.A(_05801_),
    .X(_05802_));
 sg13g2_mux2_1 _23442_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net470),
    .S(net351),
    .X(_01145_));
 sg13g2_buf_1 _23443_ (.A(net783),
    .X(_05803_));
 sg13g2_mux2_1 _23444_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net662),
    .S(net351),
    .X(_01146_));
 sg13g2_mux2_1 _23445_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net739),
    .S(net351),
    .X(_01147_));
 sg13g2_mux2_1 _23446_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net592),
    .S(net351),
    .X(_01148_));
 sg13g2_mux2_1 _23447_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net743),
    .S(net351),
    .X(_01149_));
 sg13g2_mux2_1 _23448_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net742),
    .S(_05802_),
    .X(_01150_));
 sg13g2_mux2_1 _23449_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net850),
    .S(_05802_),
    .X(_01151_));
 sg13g2_mux2_1 _23450_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net849),
    .S(net351),
    .X(_01152_));
 sg13g2_mux2_1 _23451_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net851),
    .S(net351),
    .X(_01153_));
 sg13g2_mux2_1 _23452_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(_03495_),
    .S(net351),
    .X(_01154_));
 sg13g2_mux2_1 _23453_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net540),
    .S(_05801_),
    .X(_01155_));
 sg13g2_mux2_1 _23454_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net547),
    .S(_05801_),
    .X(_01156_));
 sg13g2_nor3_1 _23455_ (.A(_05755_),
    .B(_05758_),
    .C(_05798_),
    .Y(_05804_));
 sg13g2_buf_2 _23456_ (.A(_05804_),
    .X(_05805_));
 sg13g2_nor2b_1 _23457_ (.A(net469),
    .B_N(_05805_),
    .Y(_05806_));
 sg13g2_buf_1 _23458_ (.A(_05806_),
    .X(_05807_));
 sg13g2_buf_1 _23459_ (.A(_05807_),
    .X(_05808_));
 sg13g2_mux2_1 _23460_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net470),
    .S(net350),
    .X(_01157_));
 sg13g2_mux2_1 _23461_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(net662),
    .S(net350),
    .X(_01158_));
 sg13g2_mux2_1 _23462_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net739),
    .S(net350),
    .X(_01159_));
 sg13g2_mux2_1 _23463_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net592),
    .S(net350),
    .X(_01160_));
 sg13g2_mux2_1 _23464_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(_03506_),
    .S(net350),
    .X(_01161_));
 sg13g2_mux2_1 _23465_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(_03507_),
    .S(_05808_),
    .X(_01162_));
 sg13g2_mux2_1 _23466_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(_03508_),
    .S(_05808_),
    .X(_01163_));
 sg13g2_mux2_1 _23467_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(_03509_),
    .S(net350),
    .X(_01164_));
 sg13g2_mux2_1 _23468_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(_03502_),
    .S(net350),
    .X(_01165_));
 sg13g2_mux2_1 _23469_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(_03495_),
    .S(net350),
    .X(_01166_));
 sg13g2_mux2_1 _23470_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(_04696_),
    .S(_05807_),
    .X(_01167_));
 sg13g2_mux2_1 _23471_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net547),
    .S(_05807_),
    .X(_01168_));
 sg13g2_nor2b_2 _23472_ (.A(net1113),
    .B_N(net967),
    .Y(_05809_));
 sg13g2_nand2b_1 _23473_ (.Y(_05810_),
    .B(_05809_),
    .A_N(_05780_));
 sg13g2_buf_1 _23474_ (.A(_05810_),
    .X(_05811_));
 sg13g2_nor2_1 _23475_ (.A(_05787_),
    .B(_05811_),
    .Y(_05812_));
 sg13g2_buf_1 _23476_ (.A(_05812_),
    .X(_05813_));
 sg13g2_buf_1 _23477_ (.A(_05813_),
    .X(_05814_));
 sg13g2_mux2_1 _23478_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net470),
    .S(net268),
    .X(_01169_));
 sg13g2_mux2_1 _23479_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net662),
    .S(net268),
    .X(_01170_));
 sg13g2_mux2_1 _23480_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net739),
    .S(net268),
    .X(_01171_));
 sg13g2_mux2_1 _23481_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(net592),
    .S(net268),
    .X(_01172_));
 sg13g2_mux2_1 _23482_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(_03506_),
    .S(_05814_),
    .X(_01173_));
 sg13g2_mux2_1 _23483_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(_03507_),
    .S(_05814_),
    .X(_01174_));
 sg13g2_mux2_1 _23484_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(_03508_),
    .S(net268),
    .X(_01175_));
 sg13g2_mux2_1 _23485_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(_03509_),
    .S(net268),
    .X(_01176_));
 sg13g2_mux2_1 _23486_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(_03502_),
    .S(net268),
    .X(_01177_));
 sg13g2_buf_1 _23487_ (.A(_02955_),
    .X(_05815_));
 sg13g2_mux2_1 _23488_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net846),
    .S(net268),
    .X(_01178_));
 sg13g2_mux2_1 _23489_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net540),
    .S(_05813_),
    .X(_01179_));
 sg13g2_mux2_1 _23490_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net547),
    .S(_05813_),
    .X(_01180_));
 sg13g2_nand2b_1 _23491_ (.Y(_05816_),
    .B(net970),
    .A_N(net969));
 sg13g2_buf_1 _23492_ (.A(_05816_),
    .X(_05817_));
 sg13g2_or2_1 _23493_ (.X(_05818_),
    .B(_05785_),
    .A(_05817_));
 sg13g2_buf_2 _23494_ (.A(_05818_),
    .X(_05819_));
 sg13g2_nor2_1 _23495_ (.A(_05811_),
    .B(_05819_),
    .Y(_05820_));
 sg13g2_buf_1 _23496_ (.A(_05820_),
    .X(_05821_));
 sg13g2_buf_1 _23497_ (.A(_05821_),
    .X(_05822_));
 sg13g2_mux2_1 _23498_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net470),
    .S(net267),
    .X(_01181_));
 sg13g2_mux2_1 _23499_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net662),
    .S(net267),
    .X(_01182_));
 sg13g2_mux2_1 _23500_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net739),
    .S(net267),
    .X(_01183_));
 sg13g2_mux2_1 _23501_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(net592),
    .S(net267),
    .X(_01184_));
 sg13g2_buf_1 _23502_ (.A(_09151_),
    .X(_05823_));
 sg13g2_mux2_1 _23503_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net845),
    .S(_05822_),
    .X(_01185_));
 sg13g2_buf_1 _23504_ (.A(_09155_),
    .X(_05824_));
 sg13g2_mux2_1 _23505_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net844),
    .S(_05822_),
    .X(_01186_));
 sg13g2_buf_1 _23506_ (.A(_09152_),
    .X(_05825_));
 sg13g2_mux2_1 _23507_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(net966),
    .S(net267),
    .X(_01187_));
 sg13g2_buf_1 _23508_ (.A(_10297_),
    .X(_05826_));
 sg13g2_mux2_1 _23509_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(net965),
    .S(net267),
    .X(_01188_));
 sg13g2_buf_1 _23510_ (.A(_10368_),
    .X(_05827_));
 sg13g2_mux2_1 _23511_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net964),
    .S(net267),
    .X(_01189_));
 sg13g2_mux2_1 _23512_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net846),
    .S(net267),
    .X(_01190_));
 sg13g2_mux2_1 _23513_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net540),
    .S(_05821_),
    .X(_01191_));
 sg13g2_mux2_1 _23514_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net547),
    .S(_05821_),
    .X(_01192_));
 sg13g2_buf_1 _23515_ (.A(_05785_),
    .X(_05828_));
 sg13g2_nor3_1 _23516_ (.A(net738),
    .B(_05828_),
    .C(_05811_),
    .Y(_05829_));
 sg13g2_buf_1 _23517_ (.A(_05829_),
    .X(_05830_));
 sg13g2_buf_1 _23518_ (.A(_05830_),
    .X(_05831_));
 sg13g2_mux2_1 _23519_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(net470),
    .S(net349),
    .X(_01193_));
 sg13g2_mux2_1 _23520_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net662),
    .S(net349),
    .X(_01194_));
 sg13g2_mux2_1 _23521_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(_05791_),
    .S(net349),
    .X(_01195_));
 sg13g2_mux2_1 _23522_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(net592),
    .S(net349),
    .X(_01196_));
 sg13g2_mux2_1 _23523_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(net845),
    .S(_05831_),
    .X(_01197_));
 sg13g2_mux2_1 _23524_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net844),
    .S(net349),
    .X(_01198_));
 sg13g2_mux2_1 _23525_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(net966),
    .S(_05831_),
    .X(_01199_));
 sg13g2_mux2_1 _23526_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net965),
    .S(net349),
    .X(_01200_));
 sg13g2_mux2_1 _23527_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(net964),
    .S(net349),
    .X(_01201_));
 sg13g2_mux2_1 _23528_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(_05815_),
    .S(net349),
    .X(_01202_));
 sg13g2_mux2_1 _23529_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(net540),
    .S(_05830_),
    .X(_01203_));
 sg13g2_mux2_1 _23530_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03520_),
    .S(_05830_),
    .X(_01204_));
 sg13g2_nor3_1 _23531_ (.A(_05758_),
    .B(_05828_),
    .C(_05811_),
    .Y(_05832_));
 sg13g2_buf_1 _23532_ (.A(_05832_),
    .X(_05833_));
 sg13g2_buf_1 _23533_ (.A(_05833_),
    .X(_05834_));
 sg13g2_mux2_1 _23534_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(net470),
    .S(net348),
    .X(_01205_));
 sg13g2_mux2_1 _23535_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net662),
    .S(net348),
    .X(_01206_));
 sg13g2_mux2_1 _23536_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(net739),
    .S(net348),
    .X(_01207_));
 sg13g2_mux2_1 _23537_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(net592),
    .S(net348),
    .X(_01208_));
 sg13g2_mux2_1 _23538_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(net845),
    .S(_05834_),
    .X(_01209_));
 sg13g2_mux2_1 _23539_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(net844),
    .S(net348),
    .X(_01210_));
 sg13g2_mux2_1 _23540_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(net966),
    .S(_05834_),
    .X(_01211_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(_05826_),
    .S(net348),
    .X(_01212_));
 sg13g2_mux2_1 _23542_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net964),
    .S(net348),
    .X(_01213_));
 sg13g2_mux2_1 _23543_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(_05815_),
    .S(net348),
    .X(_01214_));
 sg13g2_mux2_1 _23544_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(net540),
    .S(_05833_),
    .X(_01215_));
 sg13g2_mux2_1 _23545_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03520_),
    .S(_05833_),
    .X(_01216_));
 sg13g2_nand2b_1 _23546_ (.Y(_05835_),
    .B(net1113),
    .A_N(net967));
 sg13g2_buf_2 _23547_ (.A(_05835_),
    .X(_05836_));
 sg13g2_nand2_2 _23548_ (.Y(_05837_),
    .A(net848),
    .B(_05748_));
 sg13g2_nor3_1 _23549_ (.A(net468),
    .B(_05836_),
    .C(_05837_),
    .Y(_05838_));
 sg13g2_buf_1 _23550_ (.A(_05838_),
    .X(_05839_));
 sg13g2_buf_1 _23551_ (.A(_05839_),
    .X(_05840_));
 sg13g2_mux2_1 _23552_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(_05779_),
    .S(net347),
    .X(_01217_));
 sg13g2_mux2_1 _23553_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net662),
    .S(net347),
    .X(_01218_));
 sg13g2_mux2_1 _23554_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net739),
    .S(net347),
    .X(_01219_));
 sg13g2_mux2_1 _23555_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(_05792_),
    .S(net347),
    .X(_01220_));
 sg13g2_mux2_1 _23556_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net845),
    .S(_05840_),
    .X(_01221_));
 sg13g2_mux2_1 _23557_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(net844),
    .S(_05840_),
    .X(_01222_));
 sg13g2_mux2_1 _23558_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(_05825_),
    .S(net347),
    .X(_01223_));
 sg13g2_mux2_1 _23559_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net965),
    .S(net347),
    .X(_01224_));
 sg13g2_mux2_1 _23560_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net964),
    .S(net347),
    .X(_01225_));
 sg13g2_mux2_1 _23561_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net846),
    .S(net347),
    .X(_01226_));
 sg13g2_mux2_1 _23562_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net540),
    .S(_05839_),
    .X(_01227_));
 sg13g2_buf_1 _23563_ (.A(net696),
    .X(_05841_));
 sg13g2_mux2_1 _23564_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net591),
    .S(_05839_),
    .X(_01228_));
 sg13g2_nor3_1 _23565_ (.A(net847),
    .B(_05819_),
    .C(_05836_),
    .Y(_05842_));
 sg13g2_buf_1 _23566_ (.A(_05842_),
    .X(_05843_));
 sg13g2_buf_1 _23567_ (.A(_05843_),
    .X(_05844_));
 sg13g2_mux2_1 _23568_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net470),
    .S(net266),
    .X(_01229_));
 sg13g2_mux2_1 _23569_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net662),
    .S(net266),
    .X(_01230_));
 sg13g2_mux2_1 _23570_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net739),
    .S(net266),
    .X(_01231_));
 sg13g2_mux2_1 _23571_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net592),
    .S(net266),
    .X(_01232_));
 sg13g2_mux2_1 _23572_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net845),
    .S(_05844_),
    .X(_01233_));
 sg13g2_mux2_1 _23573_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net844),
    .S(_05844_),
    .X(_01234_));
 sg13g2_mux2_1 _23574_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net966),
    .S(net266),
    .X(_01235_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net965),
    .S(net266),
    .X(_01236_));
 sg13g2_mux2_1 _23576_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net964),
    .S(net266),
    .X(_01237_));
 sg13g2_mux2_1 _23577_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(net846),
    .S(net266),
    .X(_01238_));
 sg13g2_mux2_1 _23578_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net540),
    .S(_05843_),
    .X(_01239_));
 sg13g2_mux2_1 _23579_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net591),
    .S(_05843_),
    .X(_01240_));
 sg13g2_nor2_1 _23580_ (.A(_05796_),
    .B(net970),
    .Y(_05845_));
 sg13g2_and3_1 _23581_ (.X(_05846_),
    .A(net969),
    .B(net848),
    .C(_05845_));
 sg13g2_nor2b_1 _23582_ (.A(net967),
    .B_N(_05846_),
    .Y(_05847_));
 sg13g2_buf_1 _23583_ (.A(_05847_),
    .X(_05848_));
 sg13g2_nor2b_1 _23584_ (.A(net469),
    .B_N(_05848_),
    .Y(_05849_));
 sg13g2_buf_1 _23585_ (.A(_05849_),
    .X(_05850_));
 sg13g2_buf_1 _23586_ (.A(_05850_),
    .X(_05851_));
 sg13g2_mux2_1 _23587_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(_05779_),
    .S(net346),
    .X(_01241_));
 sg13g2_mux2_1 _23588_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(_05803_),
    .S(net346),
    .X(_01242_));
 sg13g2_mux2_1 _23589_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(net739),
    .S(net346),
    .X(_01243_));
 sg13g2_mux2_1 _23590_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(_05792_),
    .S(net346),
    .X(_01244_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(net845),
    .S(_05851_),
    .X(_01245_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(net844),
    .S(_05851_),
    .X(_01246_));
 sg13g2_mux2_1 _23593_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net966),
    .S(net346),
    .X(_01247_));
 sg13g2_mux2_1 _23594_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(net965),
    .S(net346),
    .X(_01248_));
 sg13g2_mux2_1 _23595_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net964),
    .S(net346),
    .X(_01249_));
 sg13g2_mux2_1 _23596_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net846),
    .S(net346),
    .X(_01250_));
 sg13g2_buf_1 _23597_ (.A(_09575_),
    .X(_05852_));
 sg13g2_mux2_1 _23598_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net590),
    .S(_05850_),
    .X(_01251_));
 sg13g2_mux2_1 _23599_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net591),
    .S(_05850_),
    .X(_01252_));
 sg13g2_buf_1 _23600_ (.A(net551),
    .X(_05853_));
 sg13g2_nor3_1 _23601_ (.A(net968),
    .B(_05758_),
    .C(_05836_),
    .Y(_05854_));
 sg13g2_buf_2 _23602_ (.A(_05854_),
    .X(_05855_));
 sg13g2_nor2b_1 _23603_ (.A(net469),
    .B_N(_05855_),
    .Y(_05856_));
 sg13g2_buf_1 _23604_ (.A(_05856_),
    .X(_05857_));
 sg13g2_buf_1 _23605_ (.A(_05857_),
    .X(_05858_));
 sg13g2_mux2_1 _23606_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(_05853_),
    .S(net345),
    .X(_01253_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(_05803_),
    .S(net345),
    .X(_01254_));
 sg13g2_buf_1 _23608_ (.A(net904),
    .X(_05859_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(_05859_),
    .S(net345),
    .X(_01255_));
 sg13g2_buf_1 _23610_ (.A(_04734_),
    .X(_05860_));
 sg13g2_mux2_1 _23611_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net589),
    .S(net345),
    .X(_01256_));
 sg13g2_mux2_1 _23612_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(net845),
    .S(_05858_),
    .X(_01257_));
 sg13g2_mux2_1 _23613_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(_05824_),
    .S(_05858_),
    .X(_01258_));
 sg13g2_mux2_1 _23614_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net966),
    .S(net345),
    .X(_01259_));
 sg13g2_mux2_1 _23615_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net965),
    .S(net345),
    .X(_01260_));
 sg13g2_mux2_1 _23616_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(net964),
    .S(net345),
    .X(_01261_));
 sg13g2_mux2_1 _23617_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(net846),
    .S(net345),
    .X(_01262_));
 sg13g2_mux2_1 _23618_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net590),
    .S(_05857_),
    .X(_01263_));
 sg13g2_mux2_1 _23619_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net591),
    .S(_05857_),
    .X(_01264_));
 sg13g2_nor2_1 _23620_ (.A(_05783_),
    .B(_05819_),
    .Y(_05861_));
 sg13g2_buf_1 _23621_ (.A(_05861_),
    .X(_05862_));
 sg13g2_buf_1 _23622_ (.A(_05862_),
    .X(_05863_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(net467),
    .S(net265),
    .X(_01265_));
 sg13g2_buf_1 _23624_ (.A(net783),
    .X(_05864_));
 sg13g2_mux2_1 _23625_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(net661),
    .S(net265),
    .X(_01266_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05859_),
    .S(net265),
    .X(_01267_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(net589),
    .S(_05863_),
    .X(_01268_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(net845),
    .S(net265),
    .X(_01269_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(net844),
    .S(net265),
    .X(_01270_));
 sg13g2_mux2_1 _23630_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(net966),
    .S(_05863_),
    .X(_01271_));
 sg13g2_mux2_1 _23631_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05826_),
    .S(net265),
    .X(_01272_));
 sg13g2_mux2_1 _23632_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(net964),
    .S(net265),
    .X(_01273_));
 sg13g2_mux2_1 _23633_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(net846),
    .S(net265),
    .X(_01274_));
 sg13g2_mux2_1 _23634_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net590),
    .S(_05862_),
    .X(_01275_));
 sg13g2_mux2_1 _23635_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(net591),
    .S(_05862_),
    .X(_01276_));
 sg13g2_or2_1 _23636_ (.X(_05865_),
    .B(_05836_),
    .A(_05780_));
 sg13g2_buf_1 _23637_ (.A(_05865_),
    .X(_05866_));
 sg13g2_nor2_1 _23638_ (.A(_05787_),
    .B(_05866_),
    .Y(_05867_));
 sg13g2_buf_1 _23639_ (.A(_05867_),
    .X(_05868_));
 sg13g2_buf_2 _23640_ (.A(_05868_),
    .X(_05869_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net467),
    .S(net264),
    .X(_01277_));
 sg13g2_mux2_1 _23642_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net661),
    .S(net264),
    .X(_01278_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net737),
    .S(net264),
    .X(_01279_));
 sg13g2_mux2_1 _23644_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net589),
    .S(_05869_),
    .X(_01280_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(_05823_),
    .S(_05869_),
    .X(_01281_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net844),
    .S(net264),
    .X(_01282_));
 sg13g2_mux2_1 _23647_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(_05825_),
    .S(net264),
    .X(_01283_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net965),
    .S(net264),
    .X(_01284_));
 sg13g2_mux2_1 _23649_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(_05827_),
    .S(net264),
    .X(_01285_));
 sg13g2_mux2_1 _23650_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net846),
    .S(net264),
    .X(_01286_));
 sg13g2_mux2_1 _23651_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net590),
    .S(_05868_),
    .X(_01287_));
 sg13g2_mux2_1 _23652_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net591),
    .S(_05868_),
    .X(_01288_));
 sg13g2_nor2_1 _23653_ (.A(_05819_),
    .B(_05866_),
    .Y(_05870_));
 sg13g2_buf_1 _23654_ (.A(_05870_),
    .X(_05871_));
 sg13g2_buf_2 _23655_ (.A(_05871_),
    .X(_05872_));
 sg13g2_mux2_1 _23656_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net467),
    .S(net263),
    .X(_01289_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net661),
    .S(net263),
    .X(_01290_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net737),
    .S(net263),
    .X(_01291_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net589),
    .S(_05872_),
    .X(_01292_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(_05823_),
    .S(_05872_),
    .X(_01293_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(_05824_),
    .S(net263),
    .X(_01294_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net966),
    .S(net263),
    .X(_01295_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net965),
    .S(net263),
    .X(_01296_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(_05827_),
    .S(net263),
    .X(_01297_));
 sg13g2_buf_1 _23665_ (.A(_02955_),
    .X(_05873_));
 sg13g2_mux2_1 _23666_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net843),
    .S(net263),
    .X(_01298_));
 sg13g2_mux2_1 _23667_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net590),
    .S(_05871_),
    .X(_01299_));
 sg13g2_mux2_1 _23668_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net591),
    .S(_05871_),
    .X(_01300_));
 sg13g2_nor3_1 _23669_ (.A(net738),
    .B(net468),
    .C(_05866_),
    .Y(_05874_));
 sg13g2_buf_1 _23670_ (.A(_05874_),
    .X(_05875_));
 sg13g2_buf_2 _23671_ (.A(_05875_),
    .X(_05876_));
 sg13g2_mux2_1 _23672_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net467),
    .S(net344),
    .X(_01301_));
 sg13g2_mux2_1 _23673_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net661),
    .S(net344),
    .X(_01302_));
 sg13g2_mux2_1 _23674_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net737),
    .S(net344),
    .X(_01303_));
 sg13g2_mux2_1 _23675_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(_05860_),
    .S(_05876_),
    .X(_01304_));
 sg13g2_buf_1 _23676_ (.A(net1058),
    .X(_05877_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(_05877_),
    .S(_05876_),
    .X(_01305_));
 sg13g2_buf_1 _23678_ (.A(net1057),
    .X(_05878_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net841),
    .S(net344),
    .X(_01306_));
 sg13g2_buf_1 _23680_ (.A(_09152_),
    .X(_05879_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(_05879_),
    .S(net344),
    .X(_01307_));
 sg13g2_buf_1 _23682_ (.A(_10297_),
    .X(_05880_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net962),
    .S(net344),
    .X(_01308_));
 sg13g2_buf_1 _23684_ (.A(_10368_),
    .X(_05881_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net961),
    .S(net344),
    .X(_01309_));
 sg13g2_mux2_1 _23686_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net843),
    .S(net344),
    .X(_01310_));
 sg13g2_mux2_1 _23687_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(_05852_),
    .S(_05875_),
    .X(_01311_));
 sg13g2_mux2_1 _23688_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(_05841_),
    .S(_05875_),
    .X(_01312_));
 sg13g2_nor3_1 _23689_ (.A(_05758_),
    .B(net468),
    .C(_05866_),
    .Y(_05882_));
 sg13g2_buf_1 _23690_ (.A(_05882_),
    .X(_05883_));
 sg13g2_buf_2 _23691_ (.A(_05883_),
    .X(_05884_));
 sg13g2_mux2_1 _23692_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net467),
    .S(net343),
    .X(_01313_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net661),
    .S(net343),
    .X(_01314_));
 sg13g2_mux2_1 _23694_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net737),
    .S(net343),
    .X(_01315_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(_05860_),
    .S(_05884_),
    .X(_01316_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(_05877_),
    .S(_05884_),
    .X(_01317_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net841),
    .S(net343),
    .X(_01318_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(_05879_),
    .S(net343),
    .X(_01319_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net962),
    .S(net343),
    .X(_01320_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net961),
    .S(net343),
    .X(_01321_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(_05873_),
    .S(net343),
    .X(_01322_));
 sg13g2_mux2_1 _23702_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(_05852_),
    .S(_05883_),
    .X(_01323_));
 sg13g2_mux2_1 _23703_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(_05841_),
    .S(_05883_),
    .X(_01324_));
 sg13g2_nand2_1 _23704_ (.Y(_05885_),
    .A(net1113),
    .B(_10192_));
 sg13g2_buf_2 _23705_ (.A(_05885_),
    .X(_05886_));
 sg13g2_nor3_1 _23706_ (.A(net468),
    .B(_05837_),
    .C(_05886_),
    .Y(_05887_));
 sg13g2_buf_1 _23707_ (.A(_05887_),
    .X(_05888_));
 sg13g2_buf_1 _23708_ (.A(_05888_),
    .X(_05889_));
 sg13g2_mux2_1 _23709_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(_05853_),
    .S(net342),
    .X(_01325_));
 sg13g2_mux2_1 _23710_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net661),
    .S(net342),
    .X(_01326_));
 sg13g2_mux2_1 _23711_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net737),
    .S(net342),
    .X(_01327_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net589),
    .S(net342),
    .X(_01328_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(net842),
    .S(_05889_),
    .X(_01329_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net841),
    .S(_05889_),
    .X(_01330_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net963),
    .S(net342),
    .X(_01331_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net962),
    .S(net342),
    .X(_01332_));
 sg13g2_mux2_1 _23717_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net961),
    .S(net342),
    .X(_01333_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net843),
    .S(net342),
    .X(_01334_));
 sg13g2_mux2_1 _23719_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(net590),
    .S(_05888_),
    .X(_01335_));
 sg13g2_mux2_1 _23720_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(net591),
    .S(_05888_),
    .X(_01336_));
 sg13g2_nor3_1 _23721_ (.A(_05760_),
    .B(_05819_),
    .C(_05886_),
    .Y(_05890_));
 sg13g2_buf_1 _23722_ (.A(_05890_),
    .X(_05891_));
 sg13g2_buf_1 _23723_ (.A(_05891_),
    .X(_05892_));
 sg13g2_mux2_1 _23724_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net467),
    .S(net262),
    .X(_01337_));
 sg13g2_mux2_1 _23725_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(net661),
    .S(net262),
    .X(_01338_));
 sg13g2_mux2_1 _23726_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net737),
    .S(net262),
    .X(_01339_));
 sg13g2_mux2_1 _23727_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net589),
    .S(net262),
    .X(_01340_));
 sg13g2_mux2_1 _23728_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(net842),
    .S(_05892_),
    .X(_01341_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net841),
    .S(_05892_),
    .X(_01342_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net963),
    .S(net262),
    .X(_01343_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net962),
    .S(net262),
    .X(_01344_));
 sg13g2_mux2_1 _23732_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net961),
    .S(net262),
    .X(_01345_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(net843),
    .S(net262),
    .X(_01346_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(net590),
    .S(_05891_),
    .X(_01347_));
 sg13g2_buf_1 _23735_ (.A(net696),
    .X(_05893_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net588),
    .S(_05891_),
    .X(_01348_));
 sg13g2_and2_1 _23737_ (.A(net967),
    .B(_05846_),
    .X(_05894_));
 sg13g2_buf_1 _23738_ (.A(_05894_),
    .X(_05895_));
 sg13g2_nor2b_1 _23739_ (.A(net469),
    .B_N(_05895_),
    .Y(_05896_));
 sg13g2_buf_1 _23740_ (.A(_05896_),
    .X(_05897_));
 sg13g2_buf_1 _23741_ (.A(_05897_),
    .X(_05898_));
 sg13g2_mux2_1 _23742_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(net467),
    .S(net341),
    .X(_01349_));
 sg13g2_mux2_1 _23743_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(_05864_),
    .S(net341),
    .X(_01350_));
 sg13g2_mux2_1 _23744_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net737),
    .S(net341),
    .X(_01351_));
 sg13g2_mux2_1 _23745_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net589),
    .S(net341),
    .X(_01352_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net842),
    .S(_05898_),
    .X(_01353_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net841),
    .S(_05898_),
    .X(_01354_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net963),
    .S(net341),
    .X(_01355_));
 sg13g2_mux2_1 _23749_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net962),
    .S(net341),
    .X(_01356_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net961),
    .S(net341),
    .X(_01357_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(net843),
    .S(net341),
    .X(_01358_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net590),
    .S(_05897_),
    .X(_01359_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net588),
    .S(_05897_),
    .X(_01360_));
 sg13g2_nor3_1 _23754_ (.A(net968),
    .B(_05758_),
    .C(_05886_),
    .Y(_05899_));
 sg13g2_buf_2 _23755_ (.A(_05899_),
    .X(_05900_));
 sg13g2_nor2b_1 _23756_ (.A(net469),
    .B_N(_05900_),
    .Y(_05901_));
 sg13g2_buf_1 _23757_ (.A(_05901_),
    .X(_05902_));
 sg13g2_buf_1 _23758_ (.A(_05902_),
    .X(_05903_));
 sg13g2_mux2_1 _23759_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(net467),
    .S(net340),
    .X(_01361_));
 sg13g2_mux2_1 _23760_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(_05864_),
    .S(net340),
    .X(_01362_));
 sg13g2_mux2_1 _23761_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net737),
    .S(net340),
    .X(_01363_));
 sg13g2_mux2_1 _23762_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net589),
    .S(net340),
    .X(_01364_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net842),
    .S(_05903_),
    .X(_01365_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net841),
    .S(_05903_),
    .X(_01366_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net963),
    .S(net340),
    .X(_01367_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net962),
    .S(net340),
    .X(_01368_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net961),
    .S(net340),
    .X(_01369_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(_05873_),
    .S(net340),
    .X(_01370_));
 sg13g2_buf_1 _23769_ (.A(_09575_),
    .X(_05904_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net587),
    .S(_05902_),
    .X(_01371_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net588),
    .S(_05902_),
    .X(_01372_));
 sg13g2_buf_1 _23772_ (.A(net551),
    .X(_05905_));
 sg13g2_or2_1 _23773_ (.X(_05906_),
    .B(_05886_),
    .A(_05780_));
 sg13g2_buf_1 _23774_ (.A(_05906_),
    .X(_05907_));
 sg13g2_nor2_1 _23775_ (.A(_05787_),
    .B(_05907_),
    .Y(_05908_));
 sg13g2_buf_1 _23776_ (.A(_05908_),
    .X(_05909_));
 sg13g2_buf_1 _23777_ (.A(_05909_),
    .X(_05910_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net466),
    .S(net261),
    .X(_01373_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net661),
    .S(net261),
    .X(_01374_));
 sg13g2_buf_1 _23780_ (.A(net904),
    .X(_05911_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net736),
    .S(net261),
    .X(_01375_));
 sg13g2_buf_1 _23782_ (.A(_04734_),
    .X(_05912_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net586),
    .S(net261),
    .X(_01376_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net842),
    .S(_05910_),
    .X(_01377_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net841),
    .S(_05910_),
    .X(_01378_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net963),
    .S(net261),
    .X(_01379_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net962),
    .S(net261),
    .X(_01380_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net961),
    .S(net261),
    .X(_01381_));
 sg13g2_mux2_1 _23789_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net843),
    .S(net261),
    .X(_01382_));
 sg13g2_mux2_1 _23790_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net587),
    .S(_05909_),
    .X(_01383_));
 sg13g2_mux2_1 _23791_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net588),
    .S(_05909_),
    .X(_01384_));
 sg13g2_nor2_1 _23792_ (.A(_05819_),
    .B(_05907_),
    .Y(_05913_));
 sg13g2_buf_1 _23793_ (.A(_05913_),
    .X(_05914_));
 sg13g2_buf_1 _23794_ (.A(_05914_),
    .X(_05915_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net466),
    .S(net260),
    .X(_01385_));
 sg13g2_buf_1 _23796_ (.A(_09492_),
    .X(_05916_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net660),
    .S(net260),
    .X(_01386_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net736),
    .S(net260),
    .X(_01387_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net586),
    .S(net260),
    .X(_01388_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net842),
    .S(_05915_),
    .X(_01389_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(_05878_),
    .S(_05915_),
    .X(_01390_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net963),
    .S(net260),
    .X(_01391_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net962),
    .S(net260),
    .X(_01392_));
 sg13g2_mux2_1 _23804_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net961),
    .S(net260),
    .X(_01393_));
 sg13g2_mux2_1 _23805_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net843),
    .S(net260),
    .X(_01394_));
 sg13g2_mux2_1 _23806_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net587),
    .S(_05914_),
    .X(_01395_));
 sg13g2_mux2_1 _23807_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net588),
    .S(_05914_),
    .X(_01396_));
 sg13g2_nor3_1 _23808_ (.A(net738),
    .B(_05783_),
    .C(net469),
    .Y(_05917_));
 sg13g2_buf_1 _23809_ (.A(_05917_),
    .X(_05918_));
 sg13g2_buf_1 _23810_ (.A(_05918_),
    .X(_05919_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net466),
    .S(net339),
    .X(_01397_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net660),
    .S(net339),
    .X(_01398_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(net736),
    .S(net339),
    .X(_01399_));
 sg13g2_mux2_1 _23814_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(net586),
    .S(net339),
    .X(_01400_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net842),
    .S(net339),
    .X(_01401_));
 sg13g2_mux2_1 _23816_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(net841),
    .S(_05919_),
    .X(_01402_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(net963),
    .S(_05919_),
    .X(_01403_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(_05880_),
    .S(net339),
    .X(_01404_));
 sg13g2_mux2_1 _23819_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(_05881_),
    .S(net339),
    .X(_01405_));
 sg13g2_mux2_1 _23820_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net843),
    .S(net339),
    .X(_01406_));
 sg13g2_mux2_1 _23821_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(_05904_),
    .S(_05918_),
    .X(_01407_));
 sg13g2_mux2_1 _23822_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net588),
    .S(_05918_),
    .X(_01408_));
 sg13g2_nor3_1 _23823_ (.A(_05795_),
    .B(net468),
    .C(_05907_),
    .Y(_05920_));
 sg13g2_buf_1 _23824_ (.A(_05920_),
    .X(_05921_));
 sg13g2_buf_1 _23825_ (.A(_05921_),
    .X(_05922_));
 sg13g2_mux2_1 _23826_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net466),
    .S(net338),
    .X(_01409_));
 sg13g2_mux2_1 _23827_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(_05916_),
    .S(net338),
    .X(_01410_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net736),
    .S(net338),
    .X(_01411_));
 sg13g2_mux2_1 _23829_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(_05912_),
    .S(net338),
    .X(_01412_));
 sg13g2_mux2_1 _23830_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net842),
    .S(_05922_),
    .X(_01413_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(_05878_),
    .S(_05922_),
    .X(_01414_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net963),
    .S(net338),
    .X(_01415_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(_05880_),
    .S(net338),
    .X(_01416_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(_05881_),
    .S(net338),
    .X(_01417_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(net980),
    .S(net338),
    .X(_01418_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net587),
    .S(_05921_),
    .X(_01419_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net588),
    .S(_05921_),
    .X(_01420_));
 sg13g2_nor3_1 _23838_ (.A(_05758_),
    .B(net468),
    .C(_05907_),
    .Y(_05923_));
 sg13g2_buf_1 _23839_ (.A(_05923_),
    .X(_05924_));
 sg13g2_buf_1 _23840_ (.A(_05924_),
    .X(_05925_));
 sg13g2_mux2_1 _23841_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net466),
    .S(net337),
    .X(_01421_));
 sg13g2_mux2_1 _23842_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(_05916_),
    .S(net337),
    .X(_01422_));
 sg13g2_mux2_1 _23843_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net736),
    .S(net337),
    .X(_01423_));
 sg13g2_mux2_1 _23844_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(_05912_),
    .S(net337),
    .X(_01424_));
 sg13g2_mux2_1 _23845_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net860),
    .S(net337),
    .X(_01425_));
 sg13g2_mux2_1 _23846_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net859),
    .S(_05925_),
    .X(_01426_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(_02949_),
    .S(_05925_),
    .X(_01427_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(net985),
    .S(net337),
    .X(_01428_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net984),
    .S(net337),
    .X(_01429_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(net980),
    .S(net337),
    .X(_01430_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net587),
    .S(_05924_),
    .X(_01431_));
 sg13g2_mux2_1 _23852_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net588),
    .S(_05924_),
    .X(_01432_));
 sg13g2_nor3_1 _23853_ (.A(_05758_),
    .B(_05783_),
    .C(net468),
    .Y(_05926_));
 sg13g2_buf_1 _23854_ (.A(_05926_),
    .X(_05927_));
 sg13g2_buf_1 _23855_ (.A(_05927_),
    .X(_05928_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net466),
    .S(net336),
    .X(_01433_));
 sg13g2_mux2_1 _23857_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net660),
    .S(net336),
    .X(_01434_));
 sg13g2_mux2_1 _23858_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(net736),
    .S(net336),
    .X(_01435_));
 sg13g2_mux2_1 _23859_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net586),
    .S(net336),
    .X(_01436_));
 sg13g2_mux2_1 _23860_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(_02945_),
    .S(net336),
    .X(_01437_));
 sg13g2_mux2_1 _23861_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(net859),
    .S(_05928_),
    .X(_01438_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net986),
    .S(_05928_),
    .X(_01439_));
 sg13g2_mux2_1 _23863_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net985),
    .S(net336),
    .X(_01440_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net984),
    .S(net336),
    .X(_01441_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(_03463_),
    .S(net336),
    .X(_01442_));
 sg13g2_mux2_1 _23866_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(_05904_),
    .S(_05927_),
    .X(_01443_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(_05893_),
    .S(_05927_),
    .X(_01444_));
 sg13g2_nand2_1 _23868_ (.Y(_05929_),
    .A(net968),
    .B(_05782_));
 sg13g2_nor2_1 _23869_ (.A(_05787_),
    .B(_05929_),
    .Y(_05930_));
 sg13g2_buf_1 _23870_ (.A(_05930_),
    .X(_05931_));
 sg13g2_buf_1 _23871_ (.A(_05931_),
    .X(_05932_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net466),
    .S(net259),
    .X(_01445_));
 sg13g2_mux2_1 _23873_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net660),
    .S(net259),
    .X(_01446_));
 sg13g2_mux2_1 _23874_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net736),
    .S(net259),
    .X(_01447_));
 sg13g2_mux2_1 _23875_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net586),
    .S(net259),
    .X(_01448_));
 sg13g2_mux2_1 _23876_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net860),
    .S(net259),
    .X(_01449_));
 sg13g2_mux2_1 _23877_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net859),
    .S(net259),
    .X(_01450_));
 sg13g2_mux2_1 _23878_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net986),
    .S(_05932_),
    .X(_01451_));
 sg13g2_mux2_1 _23879_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net985),
    .S(_05932_),
    .X(_01452_));
 sg13g2_mux2_1 _23880_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net984),
    .S(net259),
    .X(_01453_));
 sg13g2_mux2_1 _23881_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net980),
    .S(net259),
    .X(_01454_));
 sg13g2_mux2_1 _23882_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net587),
    .S(_05931_),
    .X(_01455_));
 sg13g2_mux2_1 _23883_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05893_),
    .S(_05931_),
    .X(_01456_));
 sg13g2_nor2_1 _23884_ (.A(_05817_),
    .B(_05929_),
    .Y(_05933_));
 sg13g2_buf_2 _23885_ (.A(_05933_),
    .X(_05934_));
 sg13g2_nor2b_1 _23886_ (.A(net469),
    .B_N(_05934_),
    .Y(_05935_));
 sg13g2_buf_1 _23887_ (.A(_05935_),
    .X(_05936_));
 sg13g2_buf_1 _23888_ (.A(_05936_),
    .X(_05937_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net466),
    .S(net335),
    .X(_01457_));
 sg13g2_mux2_1 _23890_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(net660),
    .S(net335),
    .X(_01458_));
 sg13g2_mux2_1 _23891_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net736),
    .S(net335),
    .X(_01459_));
 sg13g2_mux2_1 _23892_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net586),
    .S(net335),
    .X(_01460_));
 sg13g2_mux2_1 _23893_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(net860),
    .S(net335),
    .X(_01461_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net859),
    .S(_05937_),
    .X(_01462_));
 sg13g2_mux2_1 _23895_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(net986),
    .S(net335),
    .X(_01463_));
 sg13g2_mux2_1 _23896_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net985),
    .S(_05937_),
    .X(_01464_));
 sg13g2_mux2_1 _23897_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net984),
    .S(net335),
    .X(_01465_));
 sg13g2_mux2_1 _23898_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net980),
    .S(net335),
    .X(_01466_));
 sg13g2_mux2_1 _23899_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net587),
    .S(_05936_),
    .X(_01467_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net610),
    .S(_05936_),
    .X(_01468_));
 sg13g2_nor2_1 _23901_ (.A(net848),
    .B(net738),
    .Y(_05938_));
 sg13g2_and2_1 _23902_ (.A(_05782_),
    .B(_05938_),
    .X(_05939_));
 sg13g2_buf_1 _23903_ (.A(_05939_),
    .X(_05940_));
 sg13g2_nor2b_1 _23904_ (.A(_05793_),
    .B_N(_05940_),
    .Y(_05941_));
 sg13g2_buf_1 _23905_ (.A(_05941_),
    .X(_05942_));
 sg13g2_buf_1 _23906_ (.A(_05942_),
    .X(_05943_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(_05905_),
    .S(net334),
    .X(_01469_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(net660),
    .S(net334),
    .X(_01470_));
 sg13g2_mux2_1 _23909_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(_05911_),
    .S(net334),
    .X(_01471_));
 sg13g2_mux2_1 _23910_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net586),
    .S(net334),
    .X(_01472_));
 sg13g2_mux2_1 _23911_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(_02945_),
    .S(net334),
    .X(_01473_));
 sg13g2_mux2_1 _23912_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(_02947_),
    .S(_05943_),
    .X(_01474_));
 sg13g2_mux2_1 _23913_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net986),
    .S(net334),
    .X(_01475_));
 sg13g2_mux2_1 _23914_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_02951_),
    .S(_05943_),
    .X(_01476_));
 sg13g2_mux2_1 _23915_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(_02953_),
    .S(net334),
    .X(_01477_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(net980),
    .S(net334),
    .X(_01478_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net587),
    .S(_05942_),
    .X(_01479_));
 sg13g2_mux2_1 _23918_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net610),
    .S(_05942_),
    .X(_01480_));
 sg13g2_and2_1 _23919_ (.A(_05759_),
    .B(_05782_),
    .X(_05944_));
 sg13g2_buf_2 _23920_ (.A(_05944_),
    .X(_05945_));
 sg13g2_nor2b_1 _23921_ (.A(_05793_),
    .B_N(_05945_),
    .Y(_05946_));
 sg13g2_buf_1 _23922_ (.A(_05946_),
    .X(_05947_));
 sg13g2_buf_1 _23923_ (.A(_05947_),
    .X(_05948_));
 sg13g2_mux2_1 _23924_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_05905_),
    .S(net333),
    .X(_01481_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(net660),
    .S(net333),
    .X(_01482_));
 sg13g2_mux2_1 _23926_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(_05911_),
    .S(net333),
    .X(_01483_));
 sg13g2_mux2_1 _23927_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net586),
    .S(net333),
    .X(_01484_));
 sg13g2_mux2_1 _23928_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net860),
    .S(net333),
    .X(_01485_));
 sg13g2_mux2_1 _23929_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(_02947_),
    .S(_05948_),
    .X(_01486_));
 sg13g2_mux2_1 _23930_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(_02949_),
    .S(net333),
    .X(_01487_));
 sg13g2_mux2_1 _23931_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(_02951_),
    .S(_05948_),
    .X(_01488_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net984),
    .S(net333),
    .X(_01489_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net980),
    .S(net333),
    .X(_01490_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(net611),
    .S(_05947_),
    .X(_01491_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net610),
    .S(_05947_),
    .X(_01492_));
 sg13g2_nor3_1 _23936_ (.A(net468),
    .B(_05798_),
    .C(_05837_),
    .Y(_05949_));
 sg13g2_buf_1 _23937_ (.A(_05949_),
    .X(_05950_));
 sg13g2_buf_1 _23938_ (.A(_05950_),
    .X(_05951_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_03478_),
    .S(net332),
    .X(_01493_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(net660),
    .S(net332),
    .X(_01494_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_09446_),
    .S(net332),
    .X(_01495_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(net613),
    .S(net332),
    .X(_01496_));
 sg13g2_mux2_1 _23943_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(net860),
    .S(net332),
    .X(_01497_));
 sg13g2_mux2_1 _23944_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(net859),
    .S(_05951_),
    .X(_01498_));
 sg13g2_mux2_1 _23945_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net986),
    .S(_05951_),
    .X(_01499_));
 sg13g2_mux2_1 _23946_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net985),
    .S(net332),
    .X(_01500_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net984),
    .S(net332),
    .X(_01501_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net980),
    .S(net332),
    .X(_01502_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net611),
    .S(_05950_),
    .X(_01503_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03467_),
    .S(_05950_),
    .X(_01504_));
 sg13g2_nor3_1 _23951_ (.A(_05760_),
    .B(_05798_),
    .C(_05819_),
    .Y(_05952_));
 sg13g2_buf_1 _23952_ (.A(_05952_),
    .X(_05953_));
 sg13g2_buf_1 _23953_ (.A(_05953_),
    .X(_05954_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(_03478_),
    .S(net258),
    .X(_01505_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(net783),
    .S(net258),
    .X(_01506_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(_09446_),
    .S(net258),
    .X(_01507_));
 sg13g2_mux2_1 _23957_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_02910_),
    .S(net258),
    .X(_01508_));
 sg13g2_mux2_1 _23958_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(net860),
    .S(net258),
    .X(_01509_));
 sg13g2_mux2_1 _23959_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(net859),
    .S(_05954_),
    .X(_01510_));
 sg13g2_mux2_1 _23960_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(net986),
    .S(_05954_),
    .X(_01511_));
 sg13g2_mux2_1 _23961_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(net985),
    .S(net258),
    .X(_01512_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(net984),
    .S(net258),
    .X(_01513_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(net980),
    .S(net258),
    .X(_01514_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_03465_),
    .S(_05953_),
    .X(_01515_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03467_),
    .S(_05953_),
    .X(_01516_));
 sg13g2_and2_1 _23966_ (.A(_05780_),
    .B(_05782_),
    .X(_05955_));
 sg13g2_buf_1 _23967_ (.A(_05955_),
    .X(_05956_));
 sg13g2_and3_1 _23968_ (.X(_05957_),
    .A(net1134),
    .B(_10505_),
    .C(_05733_));
 sg13g2_buf_1 _23969_ (.A(_05957_),
    .X(_05958_));
 sg13g2_and2_1 _23970_ (.A(_05748_),
    .B(_05958_),
    .X(_05959_));
 sg13g2_buf_1 _23971_ (.A(_05959_),
    .X(_05960_));
 sg13g2_nand2_1 _23972_ (.Y(_05961_),
    .A(_05956_),
    .B(_05960_));
 sg13g2_buf_1 _23973_ (.A(_05961_),
    .X(_05962_));
 sg13g2_buf_1 _23974_ (.A(_05961_),
    .X(_05963_));
 sg13g2_nand2_1 _23975_ (.Y(_05964_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(net330));
 sg13g2_o21ai_1 _23976_ (.B1(_05964_),
    .Y(_01517_),
    .A1(net543),
    .A2(net331));
 sg13g2_nand2_1 _23977_ (.Y(_05965_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .B(net330));
 sg13g2_o21ai_1 _23978_ (.B1(_05965_),
    .Y(_01518_),
    .A1(net545),
    .A2(net331));
 sg13g2_nand2_1 _23979_ (.Y(_05966_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .B(net330));
 sg13g2_o21ai_1 _23980_ (.B1(_05966_),
    .Y(_01519_),
    .A1(net544),
    .A2(net331));
 sg13g2_mux2_1 _23981_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .S(net331),
    .X(_01520_));
 sg13g2_nand2_1 _23982_ (.Y(_05967_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .B(_05963_));
 sg13g2_o21ai_1 _23983_ (.B1(_05967_),
    .Y(_01521_),
    .A1(net675),
    .A2(_05962_));
 sg13g2_nand2_1 _23984_ (.Y(_05968_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .B(net330));
 sg13g2_o21ai_1 _23985_ (.B1(_05968_),
    .Y(_01522_),
    .A1(net750),
    .A2(net331));
 sg13g2_nand2_1 _23986_ (.Y(_05969_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .B(net330));
 sg13g2_o21ai_1 _23987_ (.B1(_05969_),
    .Y(_01523_),
    .A1(net749),
    .A2(net331));
 sg13g2_nand2_1 _23988_ (.Y(_05970_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .B(net330));
 sg13g2_o21ai_1 _23989_ (.B1(_05970_),
    .Y(_01524_),
    .A1(net748),
    .A2(net331));
 sg13g2_nand2_1 _23990_ (.Y(_05971_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .B(net330));
 sg13g2_o21ai_1 _23991_ (.B1(_05971_),
    .Y(_01525_),
    .A1(net747),
    .A2(_05962_));
 sg13g2_buf_1 _23992_ (.A(_02955_),
    .X(_05972_));
 sg13g2_mux2_1 _23993_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net331),
    .X(_01526_));
 sg13g2_buf_1 _23994_ (.A(net611),
    .X(_05973_));
 sg13g2_mux2_1 _23995_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(net330),
    .X(_01527_));
 sg13g2_mux2_1 _23996_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_05963_),
    .X(_01528_));
 sg13g2_buf_1 _23997_ (.A(_05958_),
    .X(_05974_));
 sg13g2_nand2_1 _23998_ (.Y(_05975_),
    .A(_05799_),
    .B(net465));
 sg13g2_buf_1 _23999_ (.A(_05975_),
    .X(_05976_));
 sg13g2_buf_1 _24000_ (.A(_05975_),
    .X(_05977_));
 sg13g2_nand2_1 _24001_ (.Y(_05978_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(net384));
 sg13g2_o21ai_1 _24002_ (.B1(_05978_),
    .Y(_01529_),
    .A1(_03545_),
    .A2(_05976_));
 sg13g2_nand2_1 _24003_ (.Y(_05979_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .B(net384));
 sg13g2_o21ai_1 _24004_ (.B1(_05979_),
    .Y(_01530_),
    .A1(net545),
    .A2(net385));
 sg13g2_nand2_1 _24005_ (.Y(_05980_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .B(net384));
 sg13g2_o21ai_1 _24006_ (.B1(_05980_),
    .Y(_01531_),
    .A1(_03539_),
    .A2(net385));
 sg13g2_mux2_1 _24007_ (.A0(_02911_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .S(net385),
    .X(_01532_));
 sg13g2_nand2_1 _24008_ (.Y(_05981_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .B(net384));
 sg13g2_o21ai_1 _24009_ (.B1(_05981_),
    .Y(_01533_),
    .A1(_02920_),
    .A2(net385));
 sg13g2_nand2_1 _24010_ (.Y(_05982_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .B(net384));
 sg13g2_o21ai_1 _24011_ (.B1(_05982_),
    .Y(_01534_),
    .A1(net750),
    .A2(net385));
 sg13g2_nand2_1 _24012_ (.Y(_05983_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .B(_05977_));
 sg13g2_o21ai_1 _24013_ (.B1(_05983_),
    .Y(_01535_),
    .A1(net749),
    .A2(net385));
 sg13g2_nand2_1 _24014_ (.Y(_05984_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .B(net384));
 sg13g2_o21ai_1 _24015_ (.B1(_05984_),
    .Y(_01536_),
    .A1(_02929_),
    .A2(net385));
 sg13g2_nand2_1 _24016_ (.Y(_05985_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .B(_05977_));
 sg13g2_o21ai_1 _24017_ (.B1(_05985_),
    .Y(_01537_),
    .A1(net747),
    .A2(_05976_));
 sg13g2_mux2_1 _24018_ (.A0(_05972_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(net385),
    .X(_01538_));
 sg13g2_mux2_1 _24019_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(net384),
    .X(_01539_));
 sg13g2_mux2_1 _24020_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(net384),
    .X(_01540_));
 sg13g2_nand2_1 _24021_ (.Y(_05986_),
    .A(_05805_),
    .B(_05974_));
 sg13g2_buf_1 _24022_ (.A(_05986_),
    .X(_05987_));
 sg13g2_buf_1 _24023_ (.A(_05986_),
    .X(_05988_));
 sg13g2_nand2_1 _24024_ (.Y(_05989_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(net382));
 sg13g2_o21ai_1 _24025_ (.B1(_05989_),
    .Y(_01541_),
    .A1(_03545_),
    .A2(_05987_));
 sg13g2_nand2_1 _24026_ (.Y(_05990_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .B(_05988_));
 sg13g2_o21ai_1 _24027_ (.B1(_05990_),
    .Y(_01542_),
    .A1(net545),
    .A2(net383));
 sg13g2_nand2_1 _24028_ (.Y(_05991_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .B(net382));
 sg13g2_o21ai_1 _24029_ (.B1(_05991_),
    .Y(_01543_),
    .A1(_03539_),
    .A2(net383));
 sg13g2_mux2_1 _24030_ (.A0(_02911_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S(net383),
    .X(_01544_));
 sg13g2_nand2_1 _24031_ (.Y(_05992_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .B(net382));
 sg13g2_o21ai_1 _24032_ (.B1(_05992_),
    .Y(_01545_),
    .A1(_02920_),
    .A2(net383));
 sg13g2_nand2_1 _24033_ (.Y(_05993_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .B(net382));
 sg13g2_o21ai_1 _24034_ (.B1(_05993_),
    .Y(_01546_),
    .A1(net750),
    .A2(net383));
 sg13g2_nand2_1 _24035_ (.Y(_05994_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .B(net382));
 sg13g2_o21ai_1 _24036_ (.B1(_05994_),
    .Y(_01547_),
    .A1(_02926_),
    .A2(net383));
 sg13g2_nand2_1 _24037_ (.Y(_05995_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .B(net382));
 sg13g2_o21ai_1 _24038_ (.B1(_05995_),
    .Y(_01548_),
    .A1(_02929_),
    .A2(net383));
 sg13g2_nand2_1 _24039_ (.Y(_05996_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .B(_05988_));
 sg13g2_o21ai_1 _24040_ (.B1(_05996_),
    .Y(_01549_),
    .A1(net747),
    .A2(_05987_));
 sg13g2_mux2_1 _24041_ (.A0(_05972_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(net383),
    .X(_01550_));
 sg13g2_mux2_1 _24042_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(net382),
    .X(_01551_));
 sg13g2_mux2_1 _24043_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(net382),
    .X(_01552_));
 sg13g2_nor2_2 _24044_ (.A(_05780_),
    .B(_05798_),
    .Y(_05997_));
 sg13g2_nand2_1 _24045_ (.Y(_05998_),
    .A(_05997_),
    .B(_05960_));
 sg13g2_buf_1 _24046_ (.A(_05998_),
    .X(_05999_));
 sg13g2_buf_1 _24047_ (.A(_05998_),
    .X(_06000_));
 sg13g2_nand2_1 _24048_ (.Y(_06001_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(net328));
 sg13g2_o21ai_1 _24049_ (.B1(_06001_),
    .Y(_01553_),
    .A1(net543),
    .A2(net329));
 sg13g2_nand2_1 _24050_ (.Y(_06002_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .B(net328));
 sg13g2_o21ai_1 _24051_ (.B1(_06002_),
    .Y(_01554_),
    .A1(net545),
    .A2(net329));
 sg13g2_nand2_1 _24052_ (.Y(_06003_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .B(net328));
 sg13g2_o21ai_1 _24053_ (.B1(_06003_),
    .Y(_01555_),
    .A1(net544),
    .A2(net329));
 sg13g2_mux2_1 _24054_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .S(net329),
    .X(_01556_));
 sg13g2_nand2_1 _24055_ (.Y(_06004_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .B(net328));
 sg13g2_o21ai_1 _24056_ (.B1(_06004_),
    .Y(_01557_),
    .A1(net675),
    .A2(net329));
 sg13g2_nand2_1 _24057_ (.Y(_06005_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .B(net328));
 sg13g2_o21ai_1 _24058_ (.B1(_06005_),
    .Y(_01558_),
    .A1(net750),
    .A2(_05999_));
 sg13g2_nand2_1 _24059_ (.Y(_06006_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .B(net328));
 sg13g2_o21ai_1 _24060_ (.B1(_06006_),
    .Y(_01559_),
    .A1(net749),
    .A2(net329));
 sg13g2_nand2_1 _24061_ (.Y(_06007_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .B(net328));
 sg13g2_o21ai_1 _24062_ (.B1(_06007_),
    .Y(_01560_),
    .A1(net748),
    .A2(net329));
 sg13g2_nand2_1 _24063_ (.Y(_06008_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .B(_06000_));
 sg13g2_o21ai_1 _24064_ (.B1(_06008_),
    .Y(_01561_),
    .A1(net747),
    .A2(_05999_));
 sg13g2_mux2_1 _24065_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(net329),
    .X(_01562_));
 sg13g2_mux2_1 _24066_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_06000_),
    .X(_01563_));
 sg13g2_mux2_1 _24067_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(net328),
    .X(_01564_));
 sg13g2_nor2b_1 _24068_ (.A(_05817_),
    .B_N(_05958_),
    .Y(_06009_));
 sg13g2_buf_2 _24069_ (.A(_06009_),
    .X(_06010_));
 sg13g2_nand2_1 _24070_ (.Y(_06011_),
    .A(_05997_),
    .B(_06010_));
 sg13g2_buf_1 _24071_ (.A(_06011_),
    .X(_06012_));
 sg13g2_buf_1 _24072_ (.A(_06011_),
    .X(_06013_));
 sg13g2_nand2_1 _24073_ (.Y(_06014_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(net326));
 sg13g2_o21ai_1 _24074_ (.B1(_06014_),
    .Y(_01565_),
    .A1(net543),
    .A2(net327));
 sg13g2_nand2_1 _24075_ (.Y(_06015_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .B(net326));
 sg13g2_o21ai_1 _24076_ (.B1(_06015_),
    .Y(_01566_),
    .A1(net545),
    .A2(net327));
 sg13g2_nand2_1 _24077_ (.Y(_06016_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .B(net326));
 sg13g2_o21ai_1 _24078_ (.B1(_06016_),
    .Y(_01567_),
    .A1(net544),
    .A2(net327));
 sg13g2_mux2_1 _24079_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .S(net327),
    .X(_01568_));
 sg13g2_nand2_1 _24080_ (.Y(_06017_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .B(net326));
 sg13g2_o21ai_1 _24081_ (.B1(_06017_),
    .Y(_01569_),
    .A1(net675),
    .A2(net327));
 sg13g2_nand2_1 _24082_ (.Y(_06018_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .B(net326));
 sg13g2_o21ai_1 _24083_ (.B1(_06018_),
    .Y(_01570_),
    .A1(net750),
    .A2(_06012_));
 sg13g2_nand2_1 _24084_ (.Y(_06019_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .B(net326));
 sg13g2_o21ai_1 _24085_ (.B1(_06019_),
    .Y(_01571_),
    .A1(net749),
    .A2(net327));
 sg13g2_nand2_1 _24086_ (.Y(_06020_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .B(net326));
 sg13g2_o21ai_1 _24087_ (.B1(_06020_),
    .Y(_01572_),
    .A1(net748),
    .A2(net327));
 sg13g2_nand2_1 _24088_ (.Y(_06021_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .B(_06013_));
 sg13g2_o21ai_1 _24089_ (.B1(_06021_),
    .Y(_01573_),
    .A1(_02933_),
    .A2(_06012_));
 sg13g2_mux2_1 _24090_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(net327),
    .X(_01574_));
 sg13g2_mux2_1 _24091_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_06013_),
    .X(_01575_));
 sg13g2_mux2_1 _24092_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(net326),
    .X(_01576_));
 sg13g2_nor2b_2 _24093_ (.A(net970),
    .B_N(net969),
    .Y(_06022_));
 sg13g2_nand3_1 _24094_ (.B(_05997_),
    .C(net465),
    .A(_06022_),
    .Y(_06023_));
 sg13g2_buf_1 _24095_ (.A(_06023_),
    .X(_06024_));
 sg13g2_buf_1 _24096_ (.A(_06024_),
    .X(_06025_));
 sg13g2_buf_1 _24097_ (.A(_06024_),
    .X(_06026_));
 sg13g2_nand2_1 _24098_ (.Y(_06027_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(net324));
 sg13g2_o21ai_1 _24099_ (.B1(_06027_),
    .Y(_01577_),
    .A1(net543),
    .A2(net325));
 sg13g2_nand2_1 _24100_ (.Y(_06028_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .B(net324));
 sg13g2_o21ai_1 _24101_ (.B1(_06028_),
    .Y(_01578_),
    .A1(net545),
    .A2(net325));
 sg13g2_nand2_1 _24102_ (.Y(_06029_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .B(net324));
 sg13g2_o21ai_1 _24103_ (.B1(_06029_),
    .Y(_01579_),
    .A1(net544),
    .A2(net325));
 sg13g2_mux2_1 _24104_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .S(net325),
    .X(_01580_));
 sg13g2_nand2_1 _24105_ (.Y(_06030_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .B(net324));
 sg13g2_o21ai_1 _24106_ (.B1(_06030_),
    .Y(_01581_),
    .A1(net675),
    .A2(_06025_));
 sg13g2_nand2_1 _24107_ (.Y(_06031_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .B(_06026_));
 sg13g2_o21ai_1 _24108_ (.B1(_06031_),
    .Y(_01582_),
    .A1(net750),
    .A2(net325));
 sg13g2_nand2_1 _24109_ (.Y(_06032_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .B(net324));
 sg13g2_o21ai_1 _24110_ (.B1(_06032_),
    .Y(_01583_),
    .A1(net749),
    .A2(net325));
 sg13g2_nand2_1 _24111_ (.Y(_06033_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .B(net324));
 sg13g2_o21ai_1 _24112_ (.B1(_06033_),
    .Y(_01584_),
    .A1(net748),
    .A2(net325));
 sg13g2_nand2_1 _24113_ (.Y(_06034_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .B(net324));
 sg13g2_o21ai_1 _24114_ (.B1(_06034_),
    .Y(_01585_),
    .A1(_02933_),
    .A2(_06025_));
 sg13g2_mux2_1 _24115_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(net325),
    .X(_01586_));
 sg13g2_mux2_1 _24116_ (.A0(_05973_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_06026_),
    .X(_01587_));
 sg13g2_mux2_1 _24117_ (.A0(_03535_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(net324),
    .X(_01588_));
 sg13g2_buf_1 _24118_ (.A(_05958_),
    .X(_06035_));
 sg13g2_nand3_1 _24119_ (.B(_05997_),
    .C(net464),
    .A(_05746_),
    .Y(_06036_));
 sg13g2_buf_1 _24120_ (.A(_06036_),
    .X(_06037_));
 sg13g2_buf_1 _24121_ (.A(_06037_),
    .X(_06038_));
 sg13g2_buf_1 _24122_ (.A(_06037_),
    .X(_06039_));
 sg13g2_nand2_1 _24123_ (.Y(_06040_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(net322));
 sg13g2_o21ai_1 _24124_ (.B1(_06040_),
    .Y(_01589_),
    .A1(net543),
    .A2(net323));
 sg13g2_nand2_1 _24125_ (.Y(_06041_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .B(net322));
 sg13g2_o21ai_1 _24126_ (.B1(_06041_),
    .Y(_01590_),
    .A1(_03537_),
    .A2(net323));
 sg13g2_nand2_1 _24127_ (.Y(_06042_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .B(net322));
 sg13g2_o21ai_1 _24128_ (.B1(_06042_),
    .Y(_01591_),
    .A1(net544),
    .A2(net323));
 sg13g2_mux2_1 _24129_ (.A0(net558),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S(net323),
    .X(_01592_));
 sg13g2_buf_1 _24130_ (.A(net751),
    .X(_06043_));
 sg13g2_nand2_1 _24131_ (.Y(_06044_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .B(net322));
 sg13g2_o21ai_1 _24132_ (.B1(_06044_),
    .Y(_01593_),
    .A1(_06043_),
    .A2(_06038_));
 sg13g2_nand2_1 _24133_ (.Y(_06045_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .B(_06039_));
 sg13g2_o21ai_1 _24134_ (.B1(_06045_),
    .Y(_01594_),
    .A1(net750),
    .A2(_06038_));
 sg13g2_buf_1 _24135_ (.A(net863),
    .X(_06046_));
 sg13g2_nand2_1 _24136_ (.Y(_06047_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .B(net322));
 sg13g2_o21ai_1 _24137_ (.B1(_06047_),
    .Y(_01595_),
    .A1(_06046_),
    .A2(net323));
 sg13g2_buf_1 _24138_ (.A(net862),
    .X(_06048_));
 sg13g2_nand2_1 _24139_ (.Y(_06049_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .B(net322));
 sg13g2_o21ai_1 _24140_ (.B1(_06049_),
    .Y(_01596_),
    .A1(net734),
    .A2(net323));
 sg13g2_buf_1 _24141_ (.A(net861),
    .X(_06050_));
 sg13g2_nand2_1 _24142_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .B(net322));
 sg13g2_o21ai_1 _24143_ (.B1(_06051_),
    .Y(_01597_),
    .A1(_06050_),
    .A2(net323));
 sg13g2_mux2_1 _24144_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net323),
    .X(_01598_));
 sg13g2_mux2_1 _24145_ (.A0(_05973_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_06039_),
    .X(_01599_));
 sg13g2_mux2_1 _24146_ (.A0(_03535_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(net322),
    .X(_01600_));
 sg13g2_nor3_2 _24147_ (.A(net970),
    .B(net969),
    .C(net847),
    .Y(_06052_));
 sg13g2_nand3b_1 _24148_ (.B(_06052_),
    .C(_06035_),
    .Y(_06053_),
    .A_N(_05836_));
 sg13g2_buf_1 _24149_ (.A(_06053_),
    .X(_06054_));
 sg13g2_buf_1 _24150_ (.A(_06054_),
    .X(_06055_));
 sg13g2_buf_1 _24151_ (.A(_06054_),
    .X(_06056_));
 sg13g2_nand2_1 _24152_ (.Y(_06057_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(net320));
 sg13g2_o21ai_1 _24153_ (.B1(_06057_),
    .Y(_01601_),
    .A1(net543),
    .A2(net321));
 sg13g2_nand2_1 _24154_ (.Y(_06058_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .B(net320));
 sg13g2_o21ai_1 _24155_ (.B1(_06058_),
    .Y(_01602_),
    .A1(net545),
    .A2(net321));
 sg13g2_nand2_1 _24156_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .B(net320));
 sg13g2_o21ai_1 _24157_ (.B1(_06059_),
    .Y(_01603_),
    .A1(net544),
    .A2(net321));
 sg13g2_buf_1 _24158_ (.A(net613),
    .X(_06060_));
 sg13g2_mux2_1 _24159_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .S(net321),
    .X(_01604_));
 sg13g2_nand2_1 _24160_ (.Y(_06061_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .B(net320));
 sg13g2_o21ai_1 _24161_ (.B1(_06061_),
    .Y(_01605_),
    .A1(net659),
    .A2(net321));
 sg13g2_buf_1 _24162_ (.A(net864),
    .X(_06062_));
 sg13g2_nand2_1 _24163_ (.Y(_06063_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .B(net320));
 sg13g2_o21ai_1 _24164_ (.B1(_06063_),
    .Y(_01606_),
    .A1(net732),
    .A2(_06055_));
 sg13g2_nand2_1 _24165_ (.Y(_06064_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .B(net320));
 sg13g2_o21ai_1 _24166_ (.B1(_06064_),
    .Y(_01607_),
    .A1(net735),
    .A2(net321));
 sg13g2_nand2_1 _24167_ (.Y(_06065_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .B(net320));
 sg13g2_o21ai_1 _24168_ (.B1(_06065_),
    .Y(_01608_),
    .A1(_06048_),
    .A2(net321));
 sg13g2_nand2_1 _24169_ (.Y(_06066_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .B(_06056_));
 sg13g2_o21ai_1 _24170_ (.B1(_06066_),
    .Y(_01609_),
    .A1(net733),
    .A2(_06055_));
 sg13g2_mux2_1 _24171_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(net321),
    .X(_01610_));
 sg13g2_mux2_1 _24172_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_06056_),
    .X(_01611_));
 sg13g2_mux2_1 _24173_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(net320),
    .X(_01612_));
 sg13g2_nand3b_1 _24174_ (.B(_06010_),
    .C(net848),
    .Y(_06067_),
    .A_N(_05836_));
 sg13g2_buf_1 _24175_ (.A(_06067_),
    .X(_06068_));
 sg13g2_buf_1 _24176_ (.A(_06068_),
    .X(_06069_));
 sg13g2_buf_1 _24177_ (.A(_06068_),
    .X(_06070_));
 sg13g2_nand2_1 _24178_ (.Y(_06071_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(net256));
 sg13g2_o21ai_1 _24179_ (.B1(_06071_),
    .Y(_01613_),
    .A1(net543),
    .A2(net257));
 sg13g2_buf_1 _24180_ (.A(net600),
    .X(_06072_));
 sg13g2_nand2_1 _24181_ (.Y(_06073_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .B(net256));
 sg13g2_o21ai_1 _24182_ (.B1(_06073_),
    .Y(_01614_),
    .A1(_06072_),
    .A2(net257));
 sg13g2_nand2_1 _24183_ (.Y(_06074_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .B(net256));
 sg13g2_o21ai_1 _24184_ (.B1(_06074_),
    .Y(_01615_),
    .A1(net544),
    .A2(net257));
 sg13g2_mux2_1 _24185_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .S(net257),
    .X(_01616_));
 sg13g2_nand2_1 _24186_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .B(net256));
 sg13g2_o21ai_1 _24187_ (.B1(_06075_),
    .Y(_01617_),
    .A1(net659),
    .A2(net257));
 sg13g2_nand2_1 _24188_ (.Y(_06076_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .B(net256));
 sg13g2_o21ai_1 _24189_ (.B1(_06076_),
    .Y(_01618_),
    .A1(net732),
    .A2(_06069_));
 sg13g2_nand2_1 _24190_ (.Y(_06077_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .B(net256));
 sg13g2_o21ai_1 _24191_ (.B1(_06077_),
    .Y(_01619_),
    .A1(net735),
    .A2(net257));
 sg13g2_nand2_1 _24192_ (.Y(_06078_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .B(net256));
 sg13g2_o21ai_1 _24193_ (.B1(_06078_),
    .Y(_01620_),
    .A1(_06048_),
    .A2(net257));
 sg13g2_nand2_1 _24194_ (.Y(_06079_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .B(_06070_));
 sg13g2_o21ai_1 _24195_ (.B1(_06079_),
    .Y(_01621_),
    .A1(net733),
    .A2(_06069_));
 sg13g2_mux2_1 _24196_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(net257),
    .X(_01622_));
 sg13g2_mux2_1 _24197_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(net256),
    .X(_01623_));
 sg13g2_mux2_1 _24198_ (.A0(net546),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06070_),
    .X(_01624_));
 sg13g2_buf_1 _24199_ (.A(net599),
    .X(_06080_));
 sg13g2_nand2_1 _24200_ (.Y(_06081_),
    .A(_05848_),
    .B(net465));
 sg13g2_buf_1 _24201_ (.A(_06081_),
    .X(_06082_));
 sg13g2_buf_1 _24202_ (.A(_06081_),
    .X(_06083_));
 sg13g2_nand2_1 _24203_ (.Y(_06084_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(net380));
 sg13g2_o21ai_1 _24204_ (.B1(_06084_),
    .Y(_01625_),
    .A1(net528),
    .A2(net381));
 sg13g2_nand2_1 _24205_ (.Y(_06085_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .B(net380));
 sg13g2_o21ai_1 _24206_ (.B1(_06085_),
    .Y(_01626_),
    .A1(net529),
    .A2(net381));
 sg13g2_buf_1 _24207_ (.A(net630),
    .X(_06086_));
 sg13g2_nand2_1 _24208_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .B(net380));
 sg13g2_o21ai_1 _24209_ (.B1(_06087_),
    .Y(_01627_),
    .A1(net527),
    .A2(_06082_));
 sg13g2_mux2_1 _24210_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .S(net381),
    .X(_01628_));
 sg13g2_nand2_1 _24211_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .B(net380));
 sg13g2_o21ai_1 _24212_ (.B1(_06088_),
    .Y(_01629_),
    .A1(net659),
    .A2(_06082_));
 sg13g2_nand2_1 _24213_ (.Y(_06089_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .B(net380));
 sg13g2_o21ai_1 _24214_ (.B1(_06089_),
    .Y(_01630_),
    .A1(net732),
    .A2(net381));
 sg13g2_nand2_1 _24215_ (.Y(_06090_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .B(net380));
 sg13g2_o21ai_1 _24216_ (.B1(_06090_),
    .Y(_01631_),
    .A1(net735),
    .A2(net381));
 sg13g2_nand2_1 _24217_ (.Y(_06091_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .B(net380));
 sg13g2_o21ai_1 _24218_ (.B1(_06091_),
    .Y(_01632_),
    .A1(net734),
    .A2(net381));
 sg13g2_nand2_1 _24219_ (.Y(_06092_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .B(net380));
 sg13g2_o21ai_1 _24220_ (.B1(_06092_),
    .Y(_01633_),
    .A1(net733),
    .A2(net381));
 sg13g2_mux2_1 _24221_ (.A0(net840),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(net381),
    .X(_01634_));
 sg13g2_mux2_1 _24222_ (.A0(net531),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_06083_),
    .X(_01635_));
 sg13g2_buf_1 _24223_ (.A(net610),
    .X(_06093_));
 sg13g2_mux2_1 _24224_ (.A0(_06093_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06083_),
    .X(_01636_));
 sg13g2_nand2_1 _24225_ (.Y(_06094_),
    .A(_05855_),
    .B(net465));
 sg13g2_buf_1 _24226_ (.A(_06094_),
    .X(_06095_));
 sg13g2_buf_1 _24227_ (.A(_06094_),
    .X(_06096_));
 sg13g2_nand2_1 _24228_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(net378));
 sg13g2_o21ai_1 _24229_ (.B1(_06097_),
    .Y(_01637_),
    .A1(_06080_),
    .A2(net379));
 sg13g2_nand2_1 _24230_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .B(net378));
 sg13g2_o21ai_1 _24231_ (.B1(_06098_),
    .Y(_01638_),
    .A1(net529),
    .A2(net379));
 sg13g2_nand2_1 _24232_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .B(net378));
 sg13g2_o21ai_1 _24233_ (.B1(_06099_),
    .Y(_01639_),
    .A1(_06086_),
    .A2(_06095_));
 sg13g2_mux2_1 _24234_ (.A0(_06060_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S(net379),
    .X(_01640_));
 sg13g2_nand2_1 _24235_ (.Y(_06100_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .B(_06096_));
 sg13g2_o21ai_1 _24236_ (.B1(_06100_),
    .Y(_01641_),
    .A1(net659),
    .A2(_06095_));
 sg13g2_nand2_1 _24237_ (.Y(_06101_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .B(net378));
 sg13g2_o21ai_1 _24238_ (.B1(_06101_),
    .Y(_01642_),
    .A1(_06062_),
    .A2(net379));
 sg13g2_nand2_1 _24239_ (.Y(_06102_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .B(net378));
 sg13g2_o21ai_1 _24240_ (.B1(_06102_),
    .Y(_01643_),
    .A1(net735),
    .A2(net379));
 sg13g2_nand2_1 _24241_ (.Y(_06103_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .B(net378));
 sg13g2_o21ai_1 _24242_ (.B1(_06103_),
    .Y(_01644_),
    .A1(net734),
    .A2(net379));
 sg13g2_nand2_1 _24243_ (.Y(_06104_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .B(net378));
 sg13g2_o21ai_1 _24244_ (.B1(_06104_),
    .Y(_01645_),
    .A1(net733),
    .A2(net379));
 sg13g2_buf_1 _24245_ (.A(_02955_),
    .X(_06105_));
 sg13g2_mux2_1 _24246_ (.A0(_06105_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net379),
    .X(_01646_));
 sg13g2_buf_1 _24247_ (.A(net611),
    .X(_06106_));
 sg13g2_mux2_1 _24248_ (.A0(_06106_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(net378),
    .X(_01647_));
 sg13g2_mux2_1 _24249_ (.A0(_06093_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06096_),
    .X(_01648_));
 sg13g2_nand2_1 _24250_ (.Y(_06107_),
    .A(_05956_),
    .B(_06010_));
 sg13g2_buf_1 _24251_ (.A(_06107_),
    .X(_06108_));
 sg13g2_buf_1 _24252_ (.A(_06107_),
    .X(_06109_));
 sg13g2_nand2_1 _24253_ (.Y(_06110_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(net318));
 sg13g2_o21ai_1 _24254_ (.B1(_06110_),
    .Y(_01649_),
    .A1(_06080_),
    .A2(net319));
 sg13g2_nand2_1 _24255_ (.Y(_06111_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .B(net318));
 sg13g2_o21ai_1 _24256_ (.B1(_06111_),
    .Y(_01650_),
    .A1(_06072_),
    .A2(net319));
 sg13g2_nand2_1 _24257_ (.Y(_06112_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .B(net318));
 sg13g2_o21ai_1 _24258_ (.B1(_06112_),
    .Y(_01651_),
    .A1(_06086_),
    .A2(net319));
 sg13g2_mux2_1 _24259_ (.A0(_06060_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .S(net319),
    .X(_01652_));
 sg13g2_nand2_1 _24260_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .B(net318));
 sg13g2_o21ai_1 _24261_ (.B1(_06113_),
    .Y(_01653_),
    .A1(_06043_),
    .A2(_06108_));
 sg13g2_nand2_1 _24262_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .B(net318));
 sg13g2_o21ai_1 _24263_ (.B1(_06114_),
    .Y(_01654_),
    .A1(_06062_),
    .A2(_06108_));
 sg13g2_nand2_1 _24264_ (.Y(_06115_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .B(net318));
 sg13g2_o21ai_1 _24265_ (.B1(_06115_),
    .Y(_01655_),
    .A1(_06046_),
    .A2(net319));
 sg13g2_nand2_1 _24266_ (.Y(_06116_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .B(net318));
 sg13g2_o21ai_1 _24267_ (.B1(_06116_),
    .Y(_01656_),
    .A1(net734),
    .A2(net319));
 sg13g2_nand2_1 _24268_ (.Y(_06117_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .B(net318));
 sg13g2_o21ai_1 _24269_ (.B1(_06117_),
    .Y(_01657_),
    .A1(_06050_),
    .A2(net319));
 sg13g2_mux2_1 _24270_ (.A0(_06105_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net319),
    .X(_01658_));
 sg13g2_mux2_1 _24271_ (.A0(_06106_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_06109_),
    .X(_01659_));
 sg13g2_mux2_1 _24272_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_06109_),
    .X(_01660_));
 sg13g2_nor2_1 _24273_ (.A(_05780_),
    .B(_05836_),
    .Y(_06118_));
 sg13g2_nand2_1 _24274_ (.Y(_06119_),
    .A(_06118_),
    .B(_05960_));
 sg13g2_buf_1 _24275_ (.A(_06119_),
    .X(_06120_));
 sg13g2_buf_1 _24276_ (.A(_06119_),
    .X(_06121_));
 sg13g2_nand2_1 _24277_ (.Y(_06122_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(net316));
 sg13g2_o21ai_1 _24278_ (.B1(_06122_),
    .Y(_01661_),
    .A1(net528),
    .A2(net317));
 sg13g2_nand2_1 _24279_ (.Y(_06123_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .B(_06121_));
 sg13g2_o21ai_1 _24280_ (.B1(_06123_),
    .Y(_01662_),
    .A1(net529),
    .A2(net317));
 sg13g2_nand2_1 _24281_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .B(_06121_));
 sg13g2_o21ai_1 _24282_ (.B1(_06124_),
    .Y(_01663_),
    .A1(net527),
    .A2(net317));
 sg13g2_mux2_1 _24283_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .S(net317),
    .X(_01664_));
 sg13g2_nand2_1 _24284_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .B(net316));
 sg13g2_o21ai_1 _24285_ (.B1(_06125_),
    .Y(_01665_),
    .A1(net659),
    .A2(_06120_));
 sg13g2_nand2_1 _24286_ (.Y(_06126_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .B(net316));
 sg13g2_o21ai_1 _24287_ (.B1(_06126_),
    .Y(_01666_),
    .A1(net732),
    .A2(_06120_));
 sg13g2_nand2_1 _24288_ (.Y(_06127_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .B(net316));
 sg13g2_o21ai_1 _24289_ (.B1(_06127_),
    .Y(_01667_),
    .A1(net735),
    .A2(net317));
 sg13g2_nand2_1 _24290_ (.Y(_06128_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .B(net316));
 sg13g2_o21ai_1 _24291_ (.B1(_06128_),
    .Y(_01668_),
    .A1(net734),
    .A2(net317));
 sg13g2_nand2_1 _24292_ (.Y(_06129_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .B(net316));
 sg13g2_o21ai_1 _24293_ (.B1(_06129_),
    .Y(_01669_),
    .A1(net733),
    .A2(net317));
 sg13g2_mux2_1 _24294_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(net317),
    .X(_01670_));
 sg13g2_mux2_1 _24295_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(net316),
    .X(_01671_));
 sg13g2_mux2_1 _24296_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(net316),
    .X(_01672_));
 sg13g2_nand2_1 _24297_ (.Y(_06130_),
    .A(_06118_),
    .B(_06010_));
 sg13g2_buf_1 _24298_ (.A(_06130_),
    .X(_06131_));
 sg13g2_buf_1 _24299_ (.A(_06130_),
    .X(_06132_));
 sg13g2_nand2_1 _24300_ (.Y(_06133_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(net314));
 sg13g2_o21ai_1 _24301_ (.B1(_06133_),
    .Y(_01673_),
    .A1(net528),
    .A2(net315));
 sg13g2_nand2_1 _24302_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24303_ (.B1(_06134_),
    .Y(_01674_),
    .A1(net529),
    .A2(net315));
 sg13g2_nand2_1 _24304_ (.Y(_06135_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .B(_06132_));
 sg13g2_o21ai_1 _24305_ (.B1(_06135_),
    .Y(_01675_),
    .A1(net527),
    .A2(net315));
 sg13g2_mux2_1 _24306_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .S(net315),
    .X(_01676_));
 sg13g2_nand2_1 _24307_ (.Y(_06136_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .B(net314));
 sg13g2_o21ai_1 _24308_ (.B1(_06136_),
    .Y(_01677_),
    .A1(net659),
    .A2(_06131_));
 sg13g2_nand2_1 _24309_ (.Y(_06137_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .B(net314));
 sg13g2_o21ai_1 _24310_ (.B1(_06137_),
    .Y(_01678_),
    .A1(net732),
    .A2(_06131_));
 sg13g2_nand2_1 _24311_ (.Y(_06138_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .B(net314));
 sg13g2_o21ai_1 _24312_ (.B1(_06138_),
    .Y(_01679_),
    .A1(net735),
    .A2(net315));
 sg13g2_nand2_1 _24313_ (.Y(_06139_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .B(net314));
 sg13g2_o21ai_1 _24314_ (.B1(_06139_),
    .Y(_01680_),
    .A1(net734),
    .A2(net315));
 sg13g2_nand2_1 _24315_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .B(net314));
 sg13g2_o21ai_1 _24316_ (.B1(_06140_),
    .Y(_01681_),
    .A1(net733),
    .A2(net315));
 sg13g2_mux2_1 _24317_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(net315),
    .X(_01682_));
 sg13g2_mux2_1 _24318_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(net314),
    .X(_01683_));
 sg13g2_mux2_1 _24319_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(net314),
    .X(_01684_));
 sg13g2_nand3_1 _24320_ (.B(_06118_),
    .C(net464),
    .A(_06022_),
    .Y(_06141_));
 sg13g2_buf_1 _24321_ (.A(_06141_),
    .X(_06142_));
 sg13g2_buf_1 _24322_ (.A(_06142_),
    .X(_06143_));
 sg13g2_buf_1 _24323_ (.A(_06142_),
    .X(_06144_));
 sg13g2_nand2_1 _24324_ (.Y(_06145_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(net312));
 sg13g2_o21ai_1 _24325_ (.B1(_06145_),
    .Y(_01685_),
    .A1(net528),
    .A2(net313));
 sg13g2_nand2_1 _24326_ (.Y(_06146_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24327_ (.B1(_06146_),
    .Y(_01686_),
    .A1(net529),
    .A2(net313));
 sg13g2_nand2_1 _24328_ (.Y(_06147_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24329_ (.B1(_06147_),
    .Y(_01687_),
    .A1(net527),
    .A2(net313));
 sg13g2_mux2_1 _24330_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .S(net313),
    .X(_01688_));
 sg13g2_nand2_1 _24331_ (.Y(_06148_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .B(net312));
 sg13g2_o21ai_1 _24332_ (.B1(_06148_),
    .Y(_01689_),
    .A1(net659),
    .A2(_06143_));
 sg13g2_nand2_1 _24333_ (.Y(_06149_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .B(net312));
 sg13g2_o21ai_1 _24334_ (.B1(_06149_),
    .Y(_01690_),
    .A1(net732),
    .A2(_06143_));
 sg13g2_nand2_1 _24335_ (.Y(_06150_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .B(net312));
 sg13g2_o21ai_1 _24336_ (.B1(_06150_),
    .Y(_01691_),
    .A1(net735),
    .A2(net313));
 sg13g2_nand2_1 _24337_ (.Y(_06151_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .B(net312));
 sg13g2_o21ai_1 _24338_ (.B1(_06151_),
    .Y(_01692_),
    .A1(net734),
    .A2(net313));
 sg13g2_nand2_1 _24339_ (.Y(_06152_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .B(net312));
 sg13g2_o21ai_1 _24340_ (.B1(_06152_),
    .Y(_01693_),
    .A1(net733),
    .A2(net313));
 sg13g2_mux2_1 _24341_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(net313),
    .X(_01694_));
 sg13g2_mux2_1 _24342_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(net312),
    .X(_01695_));
 sg13g2_mux2_1 _24343_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(net312),
    .X(_01696_));
 sg13g2_nand3_1 _24344_ (.B(_06118_),
    .C(net464),
    .A(_05746_),
    .Y(_06153_));
 sg13g2_buf_1 _24345_ (.A(_06153_),
    .X(_06154_));
 sg13g2_buf_1 _24346_ (.A(_06154_),
    .X(_06155_));
 sg13g2_buf_1 _24347_ (.A(_06154_),
    .X(_06156_));
 sg13g2_nand2_1 _24348_ (.Y(_06157_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(net310));
 sg13g2_o21ai_1 _24349_ (.B1(_06157_),
    .Y(_01697_),
    .A1(net528),
    .A2(net311));
 sg13g2_nand2_1 _24350_ (.Y(_06158_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .B(_06156_));
 sg13g2_o21ai_1 _24351_ (.B1(_06158_),
    .Y(_01698_),
    .A1(net529),
    .A2(net311));
 sg13g2_nand2_1 _24352_ (.Y(_06159_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .B(_06156_));
 sg13g2_o21ai_1 _24353_ (.B1(_06159_),
    .Y(_01699_),
    .A1(net527),
    .A2(net311));
 sg13g2_mux2_1 _24354_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S(net311),
    .X(_01700_));
 sg13g2_nand2_1 _24355_ (.Y(_06160_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .B(net310));
 sg13g2_o21ai_1 _24356_ (.B1(_06160_),
    .Y(_01701_),
    .A1(net659),
    .A2(_06155_));
 sg13g2_nand2_1 _24357_ (.Y(_06161_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .B(net310));
 sg13g2_o21ai_1 _24358_ (.B1(_06161_),
    .Y(_01702_),
    .A1(net732),
    .A2(net311));
 sg13g2_nand2_1 _24359_ (.Y(_06162_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .B(net310));
 sg13g2_o21ai_1 _24360_ (.B1(_06162_),
    .Y(_01703_),
    .A1(net735),
    .A2(net311));
 sg13g2_nand2_1 _24361_ (.Y(_06163_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .B(net310));
 sg13g2_o21ai_1 _24362_ (.B1(_06163_),
    .Y(_01704_),
    .A1(net734),
    .A2(net311));
 sg13g2_nand2_1 _24363_ (.Y(_06164_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .B(net310));
 sg13g2_o21ai_1 _24364_ (.B1(_06164_),
    .Y(_01705_),
    .A1(net733),
    .A2(_06155_));
 sg13g2_mux2_1 _24365_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(net311),
    .X(_01706_));
 sg13g2_mux2_1 _24366_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(net310),
    .X(_01707_));
 sg13g2_mux2_1 _24367_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(net310),
    .X(_01708_));
 sg13g2_inv_1 _24368_ (.Y(_06165_),
    .A(_05886_));
 sg13g2_nand3_1 _24369_ (.B(_06165_),
    .C(net464),
    .A(_06052_),
    .Y(_06166_));
 sg13g2_buf_1 _24370_ (.A(_06166_),
    .X(_06167_));
 sg13g2_buf_1 _24371_ (.A(_06167_),
    .X(_06168_));
 sg13g2_buf_1 _24372_ (.A(_06167_),
    .X(_06169_));
 sg13g2_nand2_1 _24373_ (.Y(_06170_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(net308));
 sg13g2_o21ai_1 _24374_ (.B1(_06170_),
    .Y(_01709_),
    .A1(net528),
    .A2(net309));
 sg13g2_nand2_1 _24375_ (.Y(_06171_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .B(net308));
 sg13g2_o21ai_1 _24376_ (.B1(_06171_),
    .Y(_01710_),
    .A1(net529),
    .A2(net309));
 sg13g2_nand2_1 _24377_ (.Y(_06172_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .B(net308));
 sg13g2_o21ai_1 _24378_ (.B1(_06172_),
    .Y(_01711_),
    .A1(net527),
    .A2(net309));
 sg13g2_mux2_1 _24379_ (.A0(net530),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .S(net309),
    .X(_01712_));
 sg13g2_buf_1 _24380_ (.A(net751),
    .X(_06173_));
 sg13g2_nand2_1 _24381_ (.Y(_06174_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .B(net308));
 sg13g2_o21ai_1 _24382_ (.B1(_06174_),
    .Y(_01713_),
    .A1(net658),
    .A2(net309));
 sg13g2_nand2_1 _24383_ (.Y(_06175_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .B(_06169_));
 sg13g2_o21ai_1 _24384_ (.B1(_06175_),
    .Y(_01714_),
    .A1(net732),
    .A2(_06168_));
 sg13g2_buf_1 _24385_ (.A(net863),
    .X(_06176_));
 sg13g2_nand2_1 _24386_ (.Y(_06177_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .B(net308));
 sg13g2_o21ai_1 _24387_ (.B1(_06177_),
    .Y(_01715_),
    .A1(net731),
    .A2(net309));
 sg13g2_buf_1 _24388_ (.A(net862),
    .X(_06178_));
 sg13g2_nand2_1 _24389_ (.Y(_06179_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .B(net308));
 sg13g2_o21ai_1 _24390_ (.B1(_06179_),
    .Y(_01716_),
    .A1(net730),
    .A2(net309));
 sg13g2_buf_1 _24391_ (.A(net861),
    .X(_06180_));
 sg13g2_nand2_1 _24392_ (.Y(_06181_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .B(net308));
 sg13g2_o21ai_1 _24393_ (.B1(_06181_),
    .Y(_01717_),
    .A1(net729),
    .A2(_06168_));
 sg13g2_mux2_1 _24394_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net309),
    .X(_01718_));
 sg13g2_mux2_1 _24395_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_06169_),
    .X(_01719_));
 sg13g2_mux2_1 _24396_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(net308),
    .X(_01720_));
 sg13g2_nand3_1 _24397_ (.B(_06165_),
    .C(_06010_),
    .A(net848),
    .Y(_06182_));
 sg13g2_buf_1 _24398_ (.A(_06182_),
    .X(_06183_));
 sg13g2_buf_1 _24399_ (.A(_06183_),
    .X(_06184_));
 sg13g2_buf_1 _24400_ (.A(_06183_),
    .X(_06185_));
 sg13g2_nand2_1 _24401_ (.Y(_06186_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(net254));
 sg13g2_o21ai_1 _24402_ (.B1(_06186_),
    .Y(_01721_),
    .A1(net528),
    .A2(net255));
 sg13g2_nand2_1 _24403_ (.Y(_06187_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .B(net254));
 sg13g2_o21ai_1 _24404_ (.B1(_06187_),
    .Y(_01722_),
    .A1(net529),
    .A2(net255));
 sg13g2_nand2_1 _24405_ (.Y(_06188_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .B(net254));
 sg13g2_o21ai_1 _24406_ (.B1(_06188_),
    .Y(_01723_),
    .A1(net527),
    .A2(net255));
 sg13g2_buf_1 _24407_ (.A(net613),
    .X(_06189_));
 sg13g2_mux2_1 _24408_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .S(net255),
    .X(_01724_));
 sg13g2_nand2_1 _24409_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .B(net254));
 sg13g2_o21ai_1 _24410_ (.B1(_06190_),
    .Y(_01725_),
    .A1(net658),
    .A2(net255));
 sg13g2_buf_1 _24411_ (.A(net864),
    .X(_06191_));
 sg13g2_nand2_1 _24412_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24413_ (.B1(_06192_),
    .Y(_01726_),
    .A1(net728),
    .A2(_06184_));
 sg13g2_nand2_1 _24414_ (.Y(_06193_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .B(net254));
 sg13g2_o21ai_1 _24415_ (.B1(_06193_),
    .Y(_01727_),
    .A1(net731),
    .A2(net255));
 sg13g2_nand2_1 _24416_ (.Y(_06194_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .B(net254));
 sg13g2_o21ai_1 _24417_ (.B1(_06194_),
    .Y(_01728_),
    .A1(net730),
    .A2(net255));
 sg13g2_nand2_1 _24418_ (.Y(_06195_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .B(net254));
 sg13g2_o21ai_1 _24419_ (.B1(_06195_),
    .Y(_01729_),
    .A1(net729),
    .A2(_06184_));
 sg13g2_mux2_1 _24420_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net255),
    .X(_01730_));
 sg13g2_mux2_1 _24421_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(_06185_),
    .X(_01731_));
 sg13g2_mux2_1 _24422_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(net254),
    .X(_01732_));
 sg13g2_nand2_1 _24423_ (.Y(_06196_),
    .A(_05895_),
    .B(net465));
 sg13g2_buf_1 _24424_ (.A(_06196_),
    .X(_06197_));
 sg13g2_buf_1 _24425_ (.A(_06196_),
    .X(_06198_));
 sg13g2_nand2_1 _24426_ (.Y(_06199_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(net376));
 sg13g2_o21ai_1 _24427_ (.B1(_06199_),
    .Y(_01733_),
    .A1(net528),
    .A2(net377));
 sg13g2_buf_1 _24428_ (.A(net600),
    .X(_06200_));
 sg13g2_nand2_1 _24429_ (.Y(_06201_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .B(_06198_));
 sg13g2_o21ai_1 _24430_ (.B1(_06201_),
    .Y(_01734_),
    .A1(net523),
    .A2(net377));
 sg13g2_nand2_1 _24431_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .B(net376));
 sg13g2_o21ai_1 _24432_ (.B1(_06202_),
    .Y(_01735_),
    .A1(net527),
    .A2(net377));
 sg13g2_mux2_1 _24433_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .S(net377),
    .X(_01736_));
 sg13g2_nand2_1 _24434_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .B(net376));
 sg13g2_o21ai_1 _24435_ (.B1(_06203_),
    .Y(_01737_),
    .A1(net658),
    .A2(net377));
 sg13g2_nand2_1 _24436_ (.Y(_06204_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .B(net376));
 sg13g2_o21ai_1 _24437_ (.B1(_06204_),
    .Y(_01738_),
    .A1(net728),
    .A2(_06197_));
 sg13g2_nand2_1 _24438_ (.Y(_06205_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .B(net376));
 sg13g2_o21ai_1 _24439_ (.B1(_06205_),
    .Y(_01739_),
    .A1(net731),
    .A2(net377));
 sg13g2_nand2_1 _24440_ (.Y(_06206_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .B(net376));
 sg13g2_o21ai_1 _24441_ (.B1(_06206_),
    .Y(_01740_),
    .A1(net730),
    .A2(net377));
 sg13g2_nand2_1 _24442_ (.Y(_06207_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .B(net376));
 sg13g2_o21ai_1 _24443_ (.B1(_06207_),
    .Y(_01741_),
    .A1(net729),
    .A2(_06197_));
 sg13g2_mux2_1 _24444_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net377),
    .X(_01742_));
 sg13g2_mux2_1 _24445_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_06198_),
    .X(_01743_));
 sg13g2_mux2_1 _24446_ (.A0(net526),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(net376),
    .X(_01744_));
 sg13g2_buf_1 _24447_ (.A(net599),
    .X(_06208_));
 sg13g2_nand2_1 _24448_ (.Y(_06209_),
    .A(_05900_),
    .B(net465));
 sg13g2_buf_1 _24449_ (.A(_06209_),
    .X(_06210_));
 sg13g2_buf_1 _24450_ (.A(_06209_),
    .X(_06211_));
 sg13g2_nand2_1 _24451_ (.Y(_06212_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(net374));
 sg13g2_o21ai_1 _24452_ (.B1(_06212_),
    .Y(_01745_),
    .A1(net522),
    .A2(net375));
 sg13g2_nand2_1 _24453_ (.Y(_06213_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .B(net374));
 sg13g2_o21ai_1 _24454_ (.B1(_06213_),
    .Y(_01746_),
    .A1(net523),
    .A2(net375));
 sg13g2_buf_1 _24455_ (.A(net630),
    .X(_06214_));
 sg13g2_nand2_1 _24456_ (.Y(_06215_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .B(net374));
 sg13g2_o21ai_1 _24457_ (.B1(_06215_),
    .Y(_01747_),
    .A1(net521),
    .A2(net375));
 sg13g2_mux2_1 _24458_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S(net375),
    .X(_01748_));
 sg13g2_nand2_1 _24459_ (.Y(_06216_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .B(net374));
 sg13g2_o21ai_1 _24460_ (.B1(_06216_),
    .Y(_01749_),
    .A1(net658),
    .A2(_06210_));
 sg13g2_nand2_1 _24461_ (.Y(_06217_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .B(_06211_));
 sg13g2_o21ai_1 _24462_ (.B1(_06217_),
    .Y(_01750_),
    .A1(net728),
    .A2(net375));
 sg13g2_nand2_1 _24463_ (.Y(_06218_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .B(net374));
 sg13g2_o21ai_1 _24464_ (.B1(_06218_),
    .Y(_01751_),
    .A1(net731),
    .A2(net375));
 sg13g2_nand2_1 _24465_ (.Y(_06219_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .B(net374));
 sg13g2_o21ai_1 _24466_ (.B1(_06219_),
    .Y(_01752_),
    .A1(net730),
    .A2(net375));
 sg13g2_nand2_1 _24467_ (.Y(_06220_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .B(net374));
 sg13g2_o21ai_1 _24468_ (.B1(_06220_),
    .Y(_01753_),
    .A1(net729),
    .A2(_06210_));
 sg13g2_mux2_1 _24469_ (.A0(net839),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net375),
    .X(_01754_));
 sg13g2_mux2_1 _24470_ (.A0(net525),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(_06211_),
    .X(_01755_));
 sg13g2_buf_1 _24471_ (.A(net610),
    .X(_06221_));
 sg13g2_mux2_1 _24472_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(net374),
    .X(_01756_));
 sg13g2_nor2_2 _24473_ (.A(_05780_),
    .B(_05886_),
    .Y(_06222_));
 sg13g2_nand2_1 _24474_ (.Y(_06223_),
    .A(_06222_),
    .B(_05960_));
 sg13g2_buf_1 _24475_ (.A(_06223_),
    .X(_06224_));
 sg13g2_buf_1 _24476_ (.A(_06223_),
    .X(_06225_));
 sg13g2_nand2_1 _24477_ (.Y(_06226_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(net306));
 sg13g2_o21ai_1 _24478_ (.B1(_06226_),
    .Y(_01757_),
    .A1(net522),
    .A2(net307));
 sg13g2_nand2_1 _24479_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .B(_06225_));
 sg13g2_o21ai_1 _24480_ (.B1(_06227_),
    .Y(_01758_),
    .A1(net523),
    .A2(net307));
 sg13g2_nand2_1 _24481_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .B(net306));
 sg13g2_o21ai_1 _24482_ (.B1(_06228_),
    .Y(_01759_),
    .A1(net521),
    .A2(_06224_));
 sg13g2_mux2_1 _24483_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .S(net307),
    .X(_01760_));
 sg13g2_nand2_1 _24484_ (.Y(_06229_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .B(net306));
 sg13g2_o21ai_1 _24485_ (.B1(_06229_),
    .Y(_01761_),
    .A1(net658),
    .A2(net307));
 sg13g2_nand2_1 _24486_ (.Y(_06230_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .B(net306));
 sg13g2_o21ai_1 _24487_ (.B1(_06230_),
    .Y(_01762_),
    .A1(net728),
    .A2(_06224_));
 sg13g2_nand2_1 _24488_ (.Y(_06231_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .B(net306));
 sg13g2_o21ai_1 _24489_ (.B1(_06231_),
    .Y(_01763_),
    .A1(net731),
    .A2(net307));
 sg13g2_nand2_1 _24490_ (.Y(_06232_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .B(net306));
 sg13g2_o21ai_1 _24491_ (.B1(_06232_),
    .Y(_01764_),
    .A1(net730),
    .A2(net307));
 sg13g2_nand2_1 _24492_ (.Y(_06233_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .B(net306));
 sg13g2_o21ai_1 _24493_ (.B1(_06233_),
    .Y(_01765_),
    .A1(net729),
    .A2(net307));
 sg13g2_buf_1 _24494_ (.A(_02955_),
    .X(_06234_));
 sg13g2_mux2_1 _24495_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(net307),
    .X(_01766_));
 sg13g2_buf_1 _24496_ (.A(net611),
    .X(_06235_));
 sg13g2_mux2_1 _24497_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06225_),
    .X(_01767_));
 sg13g2_mux2_1 _24498_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(net306),
    .X(_01768_));
 sg13g2_nand2_1 _24499_ (.Y(_06236_),
    .A(_06222_),
    .B(_06010_));
 sg13g2_buf_1 _24500_ (.A(_06236_),
    .X(_06237_));
 sg13g2_buf_1 _24501_ (.A(_06236_),
    .X(_06238_));
 sg13g2_nand2_1 _24502_ (.Y(_06239_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(net304));
 sg13g2_o21ai_1 _24503_ (.B1(_06239_),
    .Y(_01769_),
    .A1(net522),
    .A2(net305));
 sg13g2_nand2_1 _24504_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24505_ (.B1(_06240_),
    .Y(_01770_),
    .A1(net523),
    .A2(net305));
 sg13g2_nand2_1 _24506_ (.Y(_06241_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .B(net304));
 sg13g2_o21ai_1 _24507_ (.B1(_06241_),
    .Y(_01771_),
    .A1(net521),
    .A2(_06237_));
 sg13g2_mux2_1 _24508_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .S(net305),
    .X(_01772_));
 sg13g2_nand2_1 _24509_ (.Y(_06242_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .B(net304));
 sg13g2_o21ai_1 _24510_ (.B1(_06242_),
    .Y(_01773_),
    .A1(net658),
    .A2(net305));
 sg13g2_nand2_1 _24511_ (.Y(_06243_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .B(net304));
 sg13g2_o21ai_1 _24512_ (.B1(_06243_),
    .Y(_01774_),
    .A1(net728),
    .A2(_06237_));
 sg13g2_nand2_1 _24513_ (.Y(_06244_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .B(net304));
 sg13g2_o21ai_1 _24514_ (.B1(_06244_),
    .Y(_01775_),
    .A1(net731),
    .A2(net305));
 sg13g2_nand2_1 _24515_ (.Y(_06245_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .B(net304));
 sg13g2_o21ai_1 _24516_ (.B1(_06245_),
    .Y(_01776_),
    .A1(net730),
    .A2(net305));
 sg13g2_nand2_1 _24517_ (.Y(_06246_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .B(net304));
 sg13g2_o21ai_1 _24518_ (.B1(_06246_),
    .Y(_01777_),
    .A1(net729),
    .A2(net305));
 sg13g2_mux2_1 _24519_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(net305),
    .X(_01778_));
 sg13g2_mux2_1 _24520_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06238_),
    .X(_01779_));
 sg13g2_mux2_1 _24521_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(net304),
    .X(_01780_));
 sg13g2_nand3_1 _24522_ (.B(_05956_),
    .C(net464),
    .A(_06022_),
    .Y(_06247_));
 sg13g2_buf_1 _24523_ (.A(_06247_),
    .X(_06248_));
 sg13g2_buf_1 _24524_ (.A(_06248_),
    .X(_06249_));
 sg13g2_buf_1 _24525_ (.A(_06248_),
    .X(_06250_));
 sg13g2_nand2_1 _24526_ (.Y(_06251_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(net302));
 sg13g2_o21ai_1 _24527_ (.B1(_06251_),
    .Y(_01781_),
    .A1(net522),
    .A2(net303));
 sg13g2_nand2_1 _24528_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .B(_06250_));
 sg13g2_o21ai_1 _24529_ (.B1(_06252_),
    .Y(_01782_),
    .A1(net523),
    .A2(net303));
 sg13g2_nand2_1 _24530_ (.Y(_06253_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .B(net302));
 sg13g2_o21ai_1 _24531_ (.B1(_06253_),
    .Y(_01783_),
    .A1(net521),
    .A2(_06249_));
 sg13g2_mux2_1 _24532_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .S(net303),
    .X(_01784_));
 sg13g2_nand2_1 _24533_ (.Y(_06254_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .B(_06250_));
 sg13g2_o21ai_1 _24534_ (.B1(_06254_),
    .Y(_01785_),
    .A1(_06173_),
    .A2(net303));
 sg13g2_nand2_1 _24535_ (.Y(_06255_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .B(net302));
 sg13g2_o21ai_1 _24536_ (.B1(_06255_),
    .Y(_01786_),
    .A1(_06191_),
    .A2(_06249_));
 sg13g2_nand2_1 _24537_ (.Y(_06256_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .B(net302));
 sg13g2_o21ai_1 _24538_ (.B1(_06256_),
    .Y(_01787_),
    .A1(_06176_),
    .A2(net303));
 sg13g2_nand2_1 _24539_ (.Y(_06257_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .B(net302));
 sg13g2_o21ai_1 _24540_ (.B1(_06257_),
    .Y(_01788_),
    .A1(_06178_),
    .A2(net303));
 sg13g2_nand2_1 _24541_ (.Y(_06258_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .B(net302));
 sg13g2_o21ai_1 _24542_ (.B1(_06258_),
    .Y(_01789_),
    .A1(_06180_),
    .A2(net303));
 sg13g2_mux2_1 _24543_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net303),
    .X(_01790_));
 sg13g2_mux2_1 _24544_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(net302),
    .X(_01791_));
 sg13g2_mux2_1 _24545_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(net302),
    .X(_01792_));
 sg13g2_nand3_1 _24546_ (.B(_06222_),
    .C(net464),
    .A(_06022_),
    .Y(_06259_));
 sg13g2_buf_1 _24547_ (.A(_06259_),
    .X(_06260_));
 sg13g2_buf_1 _24548_ (.A(_06260_),
    .X(_06261_));
 sg13g2_buf_1 _24549_ (.A(_06260_),
    .X(_06262_));
 sg13g2_nand2_1 _24550_ (.Y(_06263_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(net300));
 sg13g2_o21ai_1 _24551_ (.B1(_06263_),
    .Y(_01793_),
    .A1(net522),
    .A2(net301));
 sg13g2_nand2_1 _24552_ (.Y(_06264_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24553_ (.B1(_06264_),
    .Y(_01794_),
    .A1(net523),
    .A2(net301));
 sg13g2_nand2_1 _24554_ (.Y(_06265_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .B(net300));
 sg13g2_o21ai_1 _24555_ (.B1(_06265_),
    .Y(_01795_),
    .A1(net521),
    .A2(_06261_));
 sg13g2_mux2_1 _24556_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .S(net301),
    .X(_01796_));
 sg13g2_nand2_1 _24557_ (.Y(_06266_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .B(net300));
 sg13g2_o21ai_1 _24558_ (.B1(_06266_),
    .Y(_01797_),
    .A1(net658),
    .A2(net301));
 sg13g2_nand2_1 _24559_ (.Y(_06267_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .B(net300));
 sg13g2_o21ai_1 _24560_ (.B1(_06267_),
    .Y(_01798_),
    .A1(net728),
    .A2(_06261_));
 sg13g2_nand2_1 _24561_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .B(net300));
 sg13g2_o21ai_1 _24562_ (.B1(_06268_),
    .Y(_01799_),
    .A1(net731),
    .A2(net301));
 sg13g2_nand2_1 _24563_ (.Y(_06269_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .B(net300));
 sg13g2_o21ai_1 _24564_ (.B1(_06269_),
    .Y(_01800_),
    .A1(net730),
    .A2(net301));
 sg13g2_nand2_1 _24565_ (.Y(_06270_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .B(net300));
 sg13g2_o21ai_1 _24566_ (.B1(_06270_),
    .Y(_01801_),
    .A1(net729),
    .A2(net301));
 sg13g2_mux2_1 _24567_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(net301),
    .X(_01802_));
 sg13g2_mux2_1 _24568_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06262_),
    .X(_01803_));
 sg13g2_mux2_1 _24569_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(net300),
    .X(_01804_));
 sg13g2_nand3_1 _24570_ (.B(_06222_),
    .C(net464),
    .A(_05746_),
    .Y(_06271_));
 sg13g2_buf_1 _24571_ (.A(_06271_),
    .X(_06272_));
 sg13g2_buf_1 _24572_ (.A(_06272_),
    .X(_06273_));
 sg13g2_buf_1 _24573_ (.A(_06272_),
    .X(_06274_));
 sg13g2_nand2_1 _24574_ (.Y(_06275_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(net298));
 sg13g2_o21ai_1 _24575_ (.B1(_06275_),
    .Y(_01805_),
    .A1(net522),
    .A2(net299));
 sg13g2_nand2_1 _24576_ (.Y(_06276_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .B(_06274_));
 sg13g2_o21ai_1 _24577_ (.B1(_06276_),
    .Y(_01806_),
    .A1(net523),
    .A2(net299));
 sg13g2_nand2_1 _24578_ (.Y(_06277_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .B(net298));
 sg13g2_o21ai_1 _24579_ (.B1(_06277_),
    .Y(_01807_),
    .A1(net521),
    .A2(net299));
 sg13g2_mux2_1 _24580_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S(net299),
    .X(_01808_));
 sg13g2_nand2_1 _24581_ (.Y(_06278_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .B(net298));
 sg13g2_o21ai_1 _24582_ (.B1(_06278_),
    .Y(_01809_),
    .A1(net658),
    .A2(net299));
 sg13g2_nand2_1 _24583_ (.Y(_06279_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .B(net298));
 sg13g2_o21ai_1 _24584_ (.B1(_06279_),
    .Y(_01810_),
    .A1(net728),
    .A2(_06273_));
 sg13g2_nand2_1 _24585_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .B(net298));
 sg13g2_o21ai_1 _24586_ (.B1(_06280_),
    .Y(_01811_),
    .A1(net731),
    .A2(net299));
 sg13g2_nand2_1 _24587_ (.Y(_06281_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .B(net298));
 sg13g2_o21ai_1 _24588_ (.B1(_06281_),
    .Y(_01812_),
    .A1(net730),
    .A2(net299));
 sg13g2_nand2_1 _24589_ (.Y(_06282_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .B(net298));
 sg13g2_o21ai_1 _24590_ (.B1(_06282_),
    .Y(_01813_),
    .A1(net729),
    .A2(_06273_));
 sg13g2_mux2_1 _24591_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(net299),
    .X(_01814_));
 sg13g2_mux2_1 _24592_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06274_),
    .X(_01815_));
 sg13g2_mux2_1 _24593_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(net298),
    .X(_01816_));
 sg13g2_nand3_1 _24594_ (.B(_05956_),
    .C(net464),
    .A(_05746_),
    .Y(_06283_));
 sg13g2_buf_1 _24595_ (.A(_06283_),
    .X(_06284_));
 sg13g2_buf_1 _24596_ (.A(_06284_),
    .X(_06285_));
 sg13g2_buf_1 _24597_ (.A(_06284_),
    .X(_06286_));
 sg13g2_nand2_1 _24598_ (.Y(_06287_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(net296));
 sg13g2_o21ai_1 _24599_ (.B1(_06287_),
    .Y(_01817_),
    .A1(net522),
    .A2(net297));
 sg13g2_nand2_1 _24600_ (.Y(_06288_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24601_ (.B1(_06288_),
    .Y(_01818_),
    .A1(net523),
    .A2(net297));
 sg13g2_nand2_1 _24602_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .B(net296));
 sg13g2_o21ai_1 _24603_ (.B1(_06289_),
    .Y(_01819_),
    .A1(net521),
    .A2(net297));
 sg13g2_mux2_1 _24604_ (.A0(_06189_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S(net297),
    .X(_01820_));
 sg13g2_nand2_1 _24605_ (.Y(_06290_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .B(net296));
 sg13g2_o21ai_1 _24606_ (.B1(_06290_),
    .Y(_01821_),
    .A1(_06173_),
    .A2(net297));
 sg13g2_nand2_1 _24607_ (.Y(_06291_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .B(net296));
 sg13g2_o21ai_1 _24608_ (.B1(_06291_),
    .Y(_01822_),
    .A1(net728),
    .A2(_06285_));
 sg13g2_nand2_1 _24609_ (.Y(_06292_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .B(net296));
 sg13g2_o21ai_1 _24610_ (.B1(_06292_),
    .Y(_01823_),
    .A1(_06176_),
    .A2(net297));
 sg13g2_nand2_1 _24611_ (.Y(_06293_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .B(net296));
 sg13g2_o21ai_1 _24612_ (.B1(_06293_),
    .Y(_01824_),
    .A1(_06178_),
    .A2(net297));
 sg13g2_nand2_1 _24613_ (.Y(_06294_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .B(net296));
 sg13g2_o21ai_1 _24614_ (.B1(_06294_),
    .Y(_01825_),
    .A1(_06180_),
    .A2(_06285_));
 sg13g2_mux2_1 _24615_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net297),
    .X(_01826_));
 sg13g2_mux2_1 _24616_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(net296),
    .X(_01827_));
 sg13g2_mux2_1 _24617_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06286_),
    .X(_01828_));
 sg13g2_nand2b_1 _24618_ (.Y(_06295_),
    .B(_05960_),
    .A_N(_05929_));
 sg13g2_buf_1 _24619_ (.A(_06295_),
    .X(_06296_));
 sg13g2_buf_1 _24620_ (.A(_06296_),
    .X(_06297_));
 sg13g2_buf_1 _24621_ (.A(_06296_),
    .X(_06298_));
 sg13g2_nand2_1 _24622_ (.Y(_06299_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(net252));
 sg13g2_o21ai_1 _24623_ (.B1(_06299_),
    .Y(_01829_),
    .A1(net522),
    .A2(_06297_));
 sg13g2_nand2_1 _24624_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .B(net252));
 sg13g2_o21ai_1 _24625_ (.B1(_06300_),
    .Y(_01830_),
    .A1(_06200_),
    .A2(net253));
 sg13g2_nand2_1 _24626_ (.Y(_06301_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24627_ (.B1(_06301_),
    .Y(_01831_),
    .A1(net521),
    .A2(net253));
 sg13g2_mux2_1 _24628_ (.A0(_06189_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .S(net253),
    .X(_01832_));
 sg13g2_nand2_1 _24629_ (.Y(_06302_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .B(net252));
 sg13g2_o21ai_1 _24630_ (.B1(_06302_),
    .Y(_01833_),
    .A1(net751),
    .A2(net253));
 sg13g2_nand2_1 _24631_ (.Y(_06303_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .B(_06298_));
 sg13g2_o21ai_1 _24632_ (.B1(_06303_),
    .Y(_01834_),
    .A1(_06191_),
    .A2(net253));
 sg13g2_nand2_1 _24633_ (.Y(_06304_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .B(net252));
 sg13g2_o21ai_1 _24634_ (.B1(_06304_),
    .Y(_01835_),
    .A1(net863),
    .A2(net253));
 sg13g2_nand2_1 _24635_ (.Y(_06305_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .B(net252));
 sg13g2_o21ai_1 _24636_ (.B1(_06305_),
    .Y(_01836_),
    .A1(net862),
    .A2(_06297_));
 sg13g2_nand2_1 _24637_ (.Y(_06306_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .B(net252));
 sg13g2_o21ai_1 _24638_ (.B1(_06306_),
    .Y(_01837_),
    .A1(net861),
    .A2(net253));
 sg13g2_mux2_1 _24639_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(net253),
    .X(_01838_));
 sg13g2_mux2_1 _24640_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(net252),
    .X(_01839_));
 sg13g2_mux2_1 _24641_ (.A0(net520),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(net252),
    .X(_01840_));
 sg13g2_nand2_1 _24642_ (.Y(_06307_),
    .A(_05934_),
    .B(net465));
 sg13g2_buf_1 _24643_ (.A(_06307_),
    .X(_06308_));
 sg13g2_buf_1 _24644_ (.A(_06307_),
    .X(_06309_));
 sg13g2_nand2_1 _24645_ (.Y(_06310_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(net372));
 sg13g2_o21ai_1 _24646_ (.B1(_06310_),
    .Y(_01841_),
    .A1(_06208_),
    .A2(net373));
 sg13g2_nand2_1 _24647_ (.Y(_06311_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .B(net372));
 sg13g2_o21ai_1 _24648_ (.B1(_06311_),
    .Y(_01842_),
    .A1(_06200_),
    .A2(net373));
 sg13g2_nand2_1 _24649_ (.Y(_06312_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .B(_06309_));
 sg13g2_o21ai_1 _24650_ (.B1(_06312_),
    .Y(_01843_),
    .A1(_06214_),
    .A2(net373));
 sg13g2_mux2_1 _24651_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .S(net373),
    .X(_01844_));
 sg13g2_nand2_1 _24652_ (.Y(_06313_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .B(net372));
 sg13g2_o21ai_1 _24653_ (.B1(_06313_),
    .Y(_01845_),
    .A1(net751),
    .A2(_06308_));
 sg13g2_nand2_1 _24654_ (.Y(_06314_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .B(_06309_));
 sg13g2_o21ai_1 _24655_ (.B1(_06314_),
    .Y(_01846_),
    .A1(net864),
    .A2(net373));
 sg13g2_nand2_1 _24656_ (.Y(_06315_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .B(net372));
 sg13g2_o21ai_1 _24657_ (.B1(_06315_),
    .Y(_01847_),
    .A1(net863),
    .A2(net373));
 sg13g2_nand2_1 _24658_ (.Y(_06316_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .B(net372));
 sg13g2_o21ai_1 _24659_ (.B1(_06316_),
    .Y(_01848_),
    .A1(net862),
    .A2(_06308_));
 sg13g2_nand2_1 _24660_ (.Y(_06317_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .B(net372));
 sg13g2_o21ai_1 _24661_ (.B1(_06317_),
    .Y(_01849_),
    .A1(net861),
    .A2(net373));
 sg13g2_mux2_1 _24662_ (.A0(net838),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(net373),
    .X(_01850_));
 sg13g2_mux2_1 _24663_ (.A0(net519),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(net372),
    .X(_01851_));
 sg13g2_mux2_1 _24664_ (.A0(_06221_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(net372),
    .X(_01852_));
 sg13g2_nand2_1 _24665_ (.Y(_06318_),
    .A(_05940_),
    .B(_05974_));
 sg13g2_buf_1 _24666_ (.A(_06318_),
    .X(_06319_));
 sg13g2_buf_1 _24667_ (.A(_06318_),
    .X(_06320_));
 sg13g2_nand2_1 _24668_ (.Y(_06321_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(net370));
 sg13g2_o21ai_1 _24669_ (.B1(_06321_),
    .Y(_01853_),
    .A1(_06208_),
    .A2(net371));
 sg13g2_nand2_1 _24670_ (.Y(_06322_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .B(net370));
 sg13g2_o21ai_1 _24671_ (.B1(_06322_),
    .Y(_01854_),
    .A1(net600),
    .A2(net371));
 sg13g2_nand2_1 _24672_ (.Y(_06323_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .B(_06320_));
 sg13g2_o21ai_1 _24673_ (.B1(_06323_),
    .Y(_01855_),
    .A1(_06214_),
    .A2(net371));
 sg13g2_mux2_1 _24674_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .S(net371),
    .X(_01856_));
 sg13g2_nand2_1 _24675_ (.Y(_06324_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .B(net370));
 sg13g2_o21ai_1 _24676_ (.B1(_06324_),
    .Y(_01857_),
    .A1(net751),
    .A2(_06319_));
 sg13g2_nand2_1 _24677_ (.Y(_06325_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .B(_06320_));
 sg13g2_o21ai_1 _24678_ (.B1(_06325_),
    .Y(_01858_),
    .A1(net864),
    .A2(net371));
 sg13g2_nand2_1 _24679_ (.Y(_06326_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .B(net370));
 sg13g2_o21ai_1 _24680_ (.B1(_06326_),
    .Y(_01859_),
    .A1(net863),
    .A2(net371));
 sg13g2_nand2_1 _24681_ (.Y(_06327_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .B(net370));
 sg13g2_o21ai_1 _24682_ (.B1(_06327_),
    .Y(_01860_),
    .A1(net862),
    .A2(_06319_));
 sg13g2_nand2_1 _24683_ (.Y(_06328_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .B(net370));
 sg13g2_o21ai_1 _24684_ (.B1(_06328_),
    .Y(_01861_),
    .A1(net861),
    .A2(net371));
 sg13g2_mux2_1 _24685_ (.A0(_06234_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(net371),
    .X(_01862_));
 sg13g2_mux2_1 _24686_ (.A0(_06235_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(net370),
    .X(_01863_));
 sg13g2_mux2_1 _24687_ (.A0(_06221_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(net370),
    .X(_01864_));
 sg13g2_nand2_1 _24688_ (.Y(_06329_),
    .A(_05945_),
    .B(net465));
 sg13g2_buf_1 _24689_ (.A(_06329_),
    .X(_06330_));
 sg13g2_buf_1 _24690_ (.A(_06329_),
    .X(_06331_));
 sg13g2_nand2_1 _24691_ (.Y(_06332_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(net368));
 sg13g2_o21ai_1 _24692_ (.B1(_06332_),
    .Y(_01865_),
    .A1(net599),
    .A2(_06330_));
 sg13g2_nand2_1 _24693_ (.Y(_06333_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .B(net368));
 sg13g2_o21ai_1 _24694_ (.B1(_06333_),
    .Y(_01866_),
    .A1(net600),
    .A2(net369));
 sg13g2_nand2_1 _24695_ (.Y(_06334_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .B(_06331_));
 sg13g2_o21ai_1 _24696_ (.B1(_06334_),
    .Y(_01867_),
    .A1(net630),
    .A2(net369));
 sg13g2_mux2_1 _24697_ (.A0(net557),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S(net369),
    .X(_01868_));
 sg13g2_nand2_1 _24698_ (.Y(_06335_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .B(net368));
 sg13g2_o21ai_1 _24699_ (.B1(_06335_),
    .Y(_01869_),
    .A1(net751),
    .A2(net369));
 sg13g2_nand2_1 _24700_ (.Y(_06336_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .B(net368));
 sg13g2_o21ai_1 _24701_ (.B1(_06336_),
    .Y(_01870_),
    .A1(net864),
    .A2(net369));
 sg13g2_nand2_1 _24702_ (.Y(_06337_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .B(net368));
 sg13g2_o21ai_1 _24703_ (.B1(_06337_),
    .Y(_01871_),
    .A1(net863),
    .A2(net369));
 sg13g2_nand2_1 _24704_ (.Y(_06338_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .B(net368));
 sg13g2_o21ai_1 _24705_ (.B1(_06338_),
    .Y(_01872_),
    .A1(net862),
    .A2(_06330_));
 sg13g2_nand2_1 _24706_ (.Y(_06339_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .B(net368));
 sg13g2_o21ai_1 _24707_ (.B1(_06339_),
    .Y(_01873_),
    .A1(net861),
    .A2(net369));
 sg13g2_mux2_1 _24708_ (.A0(_06234_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(net369),
    .X(_01874_));
 sg13g2_mux2_1 _24709_ (.A0(_06235_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(net368),
    .X(_01875_));
 sg13g2_mux2_1 _24710_ (.A0(_03468_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06331_),
    .X(_01876_));
 sg13g2_nand3_1 _24711_ (.B(_06052_),
    .C(_06035_),
    .A(_05809_),
    .Y(_06340_));
 sg13g2_buf_1 _24712_ (.A(_06340_),
    .X(_06341_));
 sg13g2_buf_1 _24713_ (.A(_06341_),
    .X(_06342_));
 sg13g2_buf_1 _24714_ (.A(_06341_),
    .X(_06343_));
 sg13g2_nand2_1 _24715_ (.Y(_06344_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(net294));
 sg13g2_o21ai_1 _24716_ (.B1(_06344_),
    .Y(_01877_),
    .A1(net599),
    .A2(net295));
 sg13g2_nand2_1 _24717_ (.Y(_06345_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .B(_06343_));
 sg13g2_o21ai_1 _24718_ (.B1(_06345_),
    .Y(_01878_),
    .A1(net600),
    .A2(net295));
 sg13g2_nand2_1 _24719_ (.Y(_06346_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .B(net294));
 sg13g2_o21ai_1 _24720_ (.B1(_06346_),
    .Y(_01879_),
    .A1(net630),
    .A2(_06342_));
 sg13g2_mux2_1 _24721_ (.A0(_02938_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .S(net295),
    .X(_01880_));
 sg13g2_nand2_1 _24722_ (.Y(_06347_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .B(net294));
 sg13g2_o21ai_1 _24723_ (.B1(_06347_),
    .Y(_01881_),
    .A1(net751),
    .A2(net295));
 sg13g2_nand2_1 _24724_ (.Y(_06348_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .B(net294));
 sg13g2_o21ai_1 _24725_ (.B1(_06348_),
    .Y(_01882_),
    .A1(_02922_),
    .A2(net295));
 sg13g2_nand2_1 _24726_ (.Y(_06349_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .B(net294));
 sg13g2_o21ai_1 _24727_ (.B1(_06349_),
    .Y(_01883_),
    .A1(net863),
    .A2(net295));
 sg13g2_nand2_1 _24728_ (.Y(_06350_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .B(net294));
 sg13g2_o21ai_1 _24729_ (.B1(_06350_),
    .Y(_01884_),
    .A1(net862),
    .A2(net295));
 sg13g2_nand2_1 _24730_ (.Y(_06351_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .B(_06343_));
 sg13g2_o21ai_1 _24731_ (.B1(_06351_),
    .Y(_01885_),
    .A1(net861),
    .A2(_06342_));
 sg13g2_mux2_1 _24732_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(net295),
    .X(_01886_));
 sg13g2_mux2_1 _24733_ (.A0(_03466_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(net294),
    .X(_01887_));
 sg13g2_mux2_1 _24734_ (.A0(_03468_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(net294),
    .X(_01888_));
 sg13g2_nand3_1 _24735_ (.B(_05809_),
    .C(_06010_),
    .A(net848),
    .Y(_06352_));
 sg13g2_buf_1 _24736_ (.A(_06352_),
    .X(_06353_));
 sg13g2_buf_1 _24737_ (.A(_06353_),
    .X(_06354_));
 sg13g2_buf_1 _24738_ (.A(_06353_),
    .X(_06355_));
 sg13g2_nand2_1 _24739_ (.Y(_06356_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(net250));
 sg13g2_o21ai_1 _24740_ (.B1(_06356_),
    .Y(_01889_),
    .A1(_03544_),
    .A2(_06354_));
 sg13g2_nand2_1 _24741_ (.Y(_06357_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .B(_06355_));
 sg13g2_o21ai_1 _24742_ (.B1(_06357_),
    .Y(_01890_),
    .A1(net600),
    .A2(net251));
 sg13g2_nand2_1 _24743_ (.Y(_06358_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .B(net250));
 sg13g2_o21ai_1 _24744_ (.B1(_06358_),
    .Y(_01891_),
    .A1(net630),
    .A2(net251));
 sg13g2_mux2_1 _24745_ (.A0(_02938_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .S(net251),
    .X(_01892_));
 sg13g2_nand2_1 _24746_ (.Y(_06359_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .B(net250));
 sg13g2_o21ai_1 _24747_ (.B1(_06359_),
    .Y(_01893_),
    .A1(net751),
    .A2(net251));
 sg13g2_nand2_1 _24748_ (.Y(_06360_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .B(net250));
 sg13g2_o21ai_1 _24749_ (.B1(_06360_),
    .Y(_01894_),
    .A1(_02922_),
    .A2(net251));
 sg13g2_nand2_1 _24750_ (.Y(_06361_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .B(net250));
 sg13g2_o21ai_1 _24751_ (.B1(_06361_),
    .Y(_01895_),
    .A1(net863),
    .A2(net251));
 sg13g2_nand2_1 _24752_ (.Y(_06362_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .B(net250));
 sg13g2_o21ai_1 _24753_ (.B1(_06362_),
    .Y(_01896_),
    .A1(net862),
    .A2(net251));
 sg13g2_nand2_1 _24754_ (.Y(_06363_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .B(_06355_));
 sg13g2_o21ai_1 _24755_ (.B1(_06363_),
    .Y(_01897_),
    .A1(net861),
    .A2(_06354_));
 sg13g2_mux2_1 _24756_ (.A0(net855),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(net251),
    .X(_01898_));
 sg13g2_mux2_1 _24757_ (.A0(_03466_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(net250),
    .X(_01899_));
 sg13g2_mux2_1 _24758_ (.A0(net553),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(net250),
    .X(_01900_));
 sg13g2_mux2_1 _24759_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(_03483_),
    .S(_05789_),
    .X(_01901_));
 sg13g2_buf_1 _24760_ (.A(net506),
    .X(_06364_));
 sg13g2_mux2_1 _24761_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net426),
    .S(_05801_),
    .X(_01902_));
 sg13g2_mux2_1 _24762_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net426),
    .S(_05807_),
    .X(_01903_));
 sg13g2_mux2_1 _24763_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net426),
    .S(_05813_),
    .X(_01904_));
 sg13g2_mux2_1 _24764_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(_06364_),
    .S(_05821_),
    .X(_01905_));
 sg13g2_mux2_1 _24765_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06364_),
    .S(_05830_),
    .X(_01906_));
 sg13g2_mux2_1 _24766_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(net426),
    .S(_05833_),
    .X(_01907_));
 sg13g2_mux2_1 _24767_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net426),
    .S(_05839_),
    .X(_01908_));
 sg13g2_mux2_1 _24768_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net426),
    .S(_05843_),
    .X(_01909_));
 sg13g2_mux2_1 _24769_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net426),
    .S(_05850_),
    .X(_01910_));
 sg13g2_mux2_1 _24770_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net426),
    .S(_05857_),
    .X(_01911_));
 sg13g2_buf_1 _24771_ (.A(net506),
    .X(_06365_));
 sg13g2_mux2_1 _24772_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(_06365_),
    .S(_05862_),
    .X(_01912_));
 sg13g2_mux2_1 _24773_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net425),
    .S(_05868_),
    .X(_01913_));
 sg13g2_mux2_1 _24774_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net425),
    .S(_05871_),
    .X(_01914_));
 sg13g2_mux2_1 _24775_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net425),
    .S(_05875_),
    .X(_01915_));
 sg13g2_mux2_1 _24776_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net425),
    .S(_05883_),
    .X(_01916_));
 sg13g2_mux2_1 _24777_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net425),
    .S(_05888_),
    .X(_01917_));
 sg13g2_mux2_1 _24778_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net425),
    .S(_05891_),
    .X(_01918_));
 sg13g2_mux2_1 _24779_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net425),
    .S(_05897_),
    .X(_01919_));
 sg13g2_mux2_1 _24780_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(net425),
    .S(_05902_),
    .X(_01920_));
 sg13g2_mux2_1 _24781_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(_06365_),
    .S(_05909_),
    .X(_01921_));
 sg13g2_buf_1 _24782_ (.A(net506),
    .X(_06366_));
 sg13g2_mux2_1 _24783_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net424),
    .S(_05914_),
    .X(_01922_));
 sg13g2_mux2_1 _24784_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(_06366_),
    .S(_05918_),
    .X(_01923_));
 sg13g2_mux2_1 _24785_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net424),
    .S(_05921_),
    .X(_01924_));
 sg13g2_mux2_1 _24786_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net424),
    .S(_05924_),
    .X(_01925_));
 sg13g2_mux2_1 _24787_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net424),
    .S(_05927_),
    .X(_01926_));
 sg13g2_mux2_1 _24788_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net424),
    .S(_05931_),
    .X(_01927_));
 sg13g2_mux2_1 _24789_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net424),
    .S(_05936_),
    .X(_01928_));
 sg13g2_mux2_1 _24790_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net424),
    .S(_05942_),
    .X(_01929_));
 sg13g2_mux2_1 _24791_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(_06366_),
    .S(_05947_),
    .X(_01930_));
 sg13g2_mux2_1 _24792_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(net424),
    .S(_05950_),
    .X(_01931_));
 sg13g2_mux2_1 _24793_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_09243_),
    .S(_05953_),
    .X(_01932_));
 sg13g2_nor2_2 _24794_ (.A(net1058),
    .B(_09168_),
    .Y(_06367_));
 sg13g2_nand3_1 _24795_ (.B(_00215_),
    .C(_06367_),
    .A(net1057),
    .Y(_06368_));
 sg13g2_buf_1 _24796_ (.A(_06368_),
    .X(_06369_));
 sg13g2_nor2_1 _24797_ (.A(net1053),
    .B(net129),
    .Y(_06370_));
 sg13g2_buf_2 _24798_ (.A(_06370_),
    .X(_06371_));
 sg13g2_nand3_1 _24799_ (.B(net387),
    .C(_06371_),
    .A(net971),
    .Y(_06372_));
 sg13g2_buf_2 _24800_ (.A(_06372_),
    .X(_06373_));
 sg13g2_mux2_1 _24801_ (.A0(net994),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .S(_06373_),
    .X(_01949_));
 sg13g2_mux2_1 _24802_ (.A0(net993),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .S(_06373_),
    .X(_01950_));
 sg13g2_nand2_1 _24803_ (.Y(_06374_),
    .A(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .B(_06373_));
 sg13g2_o21ai_1 _24804_ (.B1(_06374_),
    .Y(_01951_),
    .A1(net753),
    .A2(_06373_));
 sg13g2_nand2_1 _24805_ (.Y(_06375_),
    .A(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .B(_06373_));
 sg13g2_o21ai_1 _24806_ (.B1(_06375_),
    .Y(_01952_),
    .A1(net752),
    .A2(_06373_));
 sg13g2_nand3_1 _24807_ (.B(_10045_),
    .C(_06371_),
    .A(net971),
    .Y(_06376_));
 sg13g2_buf_2 _24808_ (.A(_06376_),
    .X(_06377_));
 sg13g2_nand2_1 _24809_ (.Y(_06378_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(_06377_));
 sg13g2_o21ai_1 _24810_ (.B1(_06378_),
    .Y(_01953_),
    .A1(net866),
    .A2(_06377_));
 sg13g2_mux2_1 _24811_ (.A0(net994),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06377_),
    .X(_01954_));
 sg13g2_mux2_1 _24812_ (.A0(net993),
    .A1(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .S(_06377_),
    .X(_01955_));
 sg13g2_nand2_1 _24813_ (.Y(_06379_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_06377_));
 sg13g2_o21ai_1 _24814_ (.B1(_06379_),
    .Y(_01956_),
    .A1(net753),
    .A2(_06377_));
 sg13g2_nand2_1 _24815_ (.Y(_06380_),
    .A(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .B(_06377_));
 sg13g2_o21ai_1 _24816_ (.B1(_06380_),
    .Y(_01957_),
    .A1(net752),
    .A2(_06377_));
 sg13g2_buf_1 _24817_ (.A(net1047),
    .X(_06381_));
 sg13g2_nand2_1 _24818_ (.Y(_06382_),
    .A(_04828_),
    .B(_06371_));
 sg13g2_buf_1 _24819_ (.A(_06382_),
    .X(_06383_));
 sg13g2_mux2_1 _24820_ (.A0(net837),
    .A1(_04826_),
    .S(net68),
    .X(_01958_));
 sg13g2_buf_1 _24821_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06384_));
 sg13g2_mux2_1 _24822_ (.A0(net900),
    .A1(_06384_),
    .S(_06383_),
    .X(_01959_));
 sg13g2_buf_1 _24823_ (.A(net1045),
    .X(_06385_));
 sg13g2_mux2_1 _24824_ (.A0(net836),
    .A1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .S(net68),
    .X(_01960_));
 sg13g2_buf_1 _24825_ (.A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .X(_06386_));
 sg13g2_nand2_1 _24826_ (.Y(_06387_),
    .A(_06386_),
    .B(net68));
 sg13g2_o21ai_1 _24827_ (.B1(_06387_),
    .Y(_01961_),
    .A1(_12631_),
    .A2(net68));
 sg13g2_mux2_1 _24828_ (.A0(net994),
    .A1(_05511_),
    .S(net68),
    .X(_01962_));
 sg13g2_mux2_1 _24829_ (.A0(net993),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .S(_06383_),
    .X(_01963_));
 sg13g2_nand2_1 _24830_ (.Y(_06388_),
    .A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B(net68));
 sg13g2_o21ai_1 _24831_ (.B1(_06388_),
    .Y(_01964_),
    .A1(_12645_),
    .A2(net68));
 sg13g2_buf_1 _24832_ (.A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .X(_06389_));
 sg13g2_nand2_1 _24833_ (.Y(_06390_),
    .A(_06389_),
    .B(_06382_));
 sg13g2_o21ai_1 _24834_ (.B1(_06390_),
    .Y(_01965_),
    .A1(_12024_),
    .A2(net68));
 sg13g2_nand2_1 _24835_ (.Y(_06391_),
    .A(_05353_),
    .B(_06371_));
 sg13g2_buf_1 _24836_ (.A(_06391_),
    .X(_06392_));
 sg13g2_mux2_1 _24837_ (.A0(net837),
    .A1(_04812_),
    .S(net67),
    .X(_01966_));
 sg13g2_mux2_1 _24838_ (.A0(net900),
    .A1(_05269_),
    .S(net67),
    .X(_01967_));
 sg13g2_mux2_1 _24839_ (.A0(net836),
    .A1(_05351_),
    .S(net67),
    .X(_01968_));
 sg13g2_nand2_1 _24840_ (.Y(_06393_),
    .A(_05389_),
    .B(net67));
 sg13g2_o21ai_1 _24841_ (.B1(_06393_),
    .Y(_01969_),
    .A1(net866),
    .A2(net67));
 sg13g2_mux2_1 _24842_ (.A0(net994),
    .A1(_05504_),
    .S(_06392_),
    .X(_01970_));
 sg13g2_mux2_1 _24843_ (.A0(net993),
    .A1(_05538_),
    .S(_06392_),
    .X(_01971_));
 sg13g2_nand2_1 _24844_ (.Y(_06394_),
    .A(_05630_),
    .B(net67));
 sg13g2_o21ai_1 _24845_ (.B1(_06394_),
    .Y(_01972_),
    .A1(_12018_),
    .A2(net67));
 sg13g2_nand2_1 _24846_ (.Y(_06395_),
    .A(_05018_),
    .B(_06391_));
 sg13g2_o21ai_1 _24847_ (.B1(_06395_),
    .Y(_01973_),
    .A1(_12024_),
    .A2(net67));
 sg13g2_nor3_1 _24848_ (.A(net916),
    .B(_05350_),
    .C(net129),
    .Y(_06396_));
 sg13g2_buf_4 _24849_ (.X(_06397_),
    .A(_06396_));
 sg13g2_mux2_1 _24850_ (.A0(_04813_),
    .A1(net837),
    .S(_06397_),
    .X(_01974_));
 sg13g2_buf_1 _24851_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06398_));
 sg13g2_mux2_1 _24852_ (.A0(_06398_),
    .A1(net900),
    .S(_06397_),
    .X(_01975_));
 sg13g2_mux2_1 _24853_ (.A0(\cpu.gpio.r_src_io[6][2] ),
    .A1(net836),
    .S(_06397_),
    .X(_01976_));
 sg13g2_mux2_1 _24854_ (.A0(\cpu.gpio.r_src_io[6][3] ),
    .A1(net1039),
    .S(_06397_),
    .X(_01977_));
 sg13g2_mux2_1 _24855_ (.A0(_05505_),
    .A1(net1006),
    .S(_06397_),
    .X(_01978_));
 sg13g2_buf_1 _24856_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06399_));
 sg13g2_mux2_1 _24857_ (.A0(_06399_),
    .A1(net1005),
    .S(_06397_),
    .X(_01979_));
 sg13g2_mux2_1 _24858_ (.A0(\cpu.gpio.r_src_io[7][2] ),
    .A1(net1038),
    .S(_06397_),
    .X(_01980_));
 sg13g2_mux2_1 _24859_ (.A0(\cpu.gpio.r_src_io[7][3] ),
    .A1(_10034_),
    .S(_06397_),
    .X(_01981_));
 sg13g2_nand2b_1 _24860_ (.Y(_06400_),
    .B(_06371_),
    .A_N(_05022_));
 sg13g2_buf_2 _24861_ (.A(_06400_),
    .X(_06401_));
 sg13g2_mux2_1 _24862_ (.A0(net994),
    .A1(_05498_),
    .S(_06401_),
    .X(_01982_));
 sg13g2_buf_1 _24863_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06402_));
 sg13g2_mux2_1 _24864_ (.A0(net993),
    .A1(_06402_),
    .S(_06401_),
    .X(_01983_));
 sg13g2_nand2_1 _24865_ (.Y(_06403_),
    .A(\cpu.gpio.r_src_o[3][2] ),
    .B(_06401_));
 sg13g2_o21ai_1 _24866_ (.B1(_06403_),
    .Y(_01984_),
    .A1(_12018_),
    .A2(_06401_));
 sg13g2_nand2_1 _24867_ (.Y(_06404_),
    .A(\cpu.gpio.r_src_o[3][3] ),
    .B(_06401_));
 sg13g2_o21ai_1 _24868_ (.B1(_06404_),
    .Y(_01985_),
    .A1(_12024_),
    .A2(_06401_));
 sg13g2_nand2_1 _24869_ (.Y(_06405_),
    .A(_04818_),
    .B(_06371_));
 sg13g2_buf_1 _24870_ (.A(_06405_),
    .X(_06406_));
 sg13g2_mux2_1 _24871_ (.A0(_06381_),
    .A1(_04816_),
    .S(net66),
    .X(_01986_));
 sg13g2_buf_1 _24872_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06407_));
 sg13g2_mux2_1 _24873_ (.A0(net900),
    .A1(_06407_),
    .S(net66),
    .X(_01987_));
 sg13g2_mux2_1 _24874_ (.A0(_06385_),
    .A1(\cpu.gpio.r_src_o[4][2] ),
    .S(_06406_),
    .X(_01988_));
 sg13g2_nand2_1 _24875_ (.Y(_06408_),
    .A(\cpu.gpio.r_src_o[4][3] ),
    .B(net66));
 sg13g2_o21ai_1 _24876_ (.B1(_06408_),
    .Y(_01989_),
    .A1(_11996_),
    .A2(net66));
 sg13g2_mux2_1 _24877_ (.A0(_12409_),
    .A1(_05503_),
    .S(net66),
    .X(_01990_));
 sg13g2_buf_1 _24878_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06409_));
 sg13g2_mux2_1 _24879_ (.A0(_12411_),
    .A1(_06409_),
    .S(net66),
    .X(_01991_));
 sg13g2_nand2_1 _24880_ (.Y(_06410_),
    .A(\cpu.gpio.r_src_o[5][2] ),
    .B(net66));
 sg13g2_o21ai_1 _24881_ (.B1(_06410_),
    .Y(_01992_),
    .A1(_12018_),
    .A2(_06406_));
 sg13g2_nand2_1 _24882_ (.Y(_06411_),
    .A(\cpu.gpio.r_src_o[5][3] ),
    .B(_06405_));
 sg13g2_o21ai_1 _24883_ (.B1(_06411_),
    .Y(_01993_),
    .A1(_12024_),
    .A2(net66));
 sg13g2_nand2_1 _24884_ (.Y(_06412_),
    .A(_04823_),
    .B(_06371_));
 sg13g2_buf_2 _24885_ (.A(_06412_),
    .X(_06413_));
 sg13g2_mux2_1 _24886_ (.A0(_12409_),
    .A1(_05500_),
    .S(_06413_),
    .X(_01998_));
 sg13g2_buf_1 _24887_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06414_));
 sg13g2_mux2_1 _24888_ (.A0(_12411_),
    .A1(_06414_),
    .S(_06413_),
    .X(_01999_));
 sg13g2_nand2_1 _24889_ (.Y(_06415_),
    .A(\cpu.gpio.r_src_o[7][2] ),
    .B(_06413_));
 sg13g2_o21ai_1 _24890_ (.B1(_06415_),
    .Y(_02000_),
    .A1(_12018_),
    .A2(_06413_));
 sg13g2_nand2_1 _24891_ (.Y(_06416_),
    .A(\cpu.gpio.r_src_o[7][3] ),
    .B(_06413_));
 sg13g2_o21ai_1 _24892_ (.B1(_06416_),
    .Y(_02001_),
    .A1(_12024_),
    .A2(_06413_));
 sg13g2_buf_1 _24893_ (.A(_02842_),
    .X(_06417_));
 sg13g2_and2_1 _24894_ (.A(net721),
    .B(_08822_),
    .X(_06418_));
 sg13g2_buf_4 _24895_ (.X(_06419_),
    .A(_06418_));
 sg13g2_nor2_1 _24896_ (.A(\cpu.icache.r_offset[2] ),
    .B(_00233_),
    .Y(_06420_));
 sg13g2_buf_1 _24897_ (.A(_06420_),
    .X(_06421_));
 sg13g2_buf_1 _24898_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06422_));
 sg13g2_buf_1 _24899_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06423_));
 sg13g2_nor2b_1 _24900_ (.A(_06422_),
    .B_N(_06423_),
    .Y(_06424_));
 sg13g2_buf_1 _24901_ (.A(_06424_),
    .X(_06425_));
 sg13g2_and2_1 _24902_ (.A(_06421_),
    .B(_06425_),
    .X(_06426_));
 sg13g2_buf_1 _24903_ (.A(_06426_),
    .X(_06427_));
 sg13g2_nand2_2 _24904_ (.Y(_06428_),
    .A(_06419_),
    .B(_06427_));
 sg13g2_mux2_1 _24905_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06428_),
    .X(_02005_));
 sg13g2_buf_1 _24906_ (.A(_12043_),
    .X(_06429_));
 sg13g2_inv_1 _24907_ (.Y(_06430_),
    .A(_00233_));
 sg13g2_buf_1 _24908_ (.A(_00234_),
    .X(_06431_));
 sg13g2_nand4_1 _24909_ (.B(_06423_),
    .C(_06430_),
    .A(_06422_),
    .Y(_06432_),
    .D(_06431_));
 sg13g2_buf_2 _24910_ (.A(_06432_),
    .X(_06433_));
 sg13g2_inv_1 _24911_ (.Y(_06434_),
    .A(_06433_));
 sg13g2_nand2_2 _24912_ (.Y(_06435_),
    .A(_06419_),
    .B(_06434_));
 sg13g2_mux2_1 _24913_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06435_),
    .X(_02006_));
 sg13g2_buf_1 _24914_ (.A(net988),
    .X(_06436_));
 sg13g2_mux2_1 _24915_ (.A0(_06436_),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06435_),
    .X(_02007_));
 sg13g2_nor2b_1 _24916_ (.A(_06423_),
    .B_N(_06422_),
    .Y(_06437_));
 sg13g2_buf_1 _24917_ (.A(_06437_),
    .X(_06438_));
 sg13g2_and2_1 _24918_ (.A(_06421_),
    .B(_06438_),
    .X(_06439_));
 sg13g2_buf_1 _24919_ (.A(_06439_),
    .X(_06440_));
 sg13g2_nand2_2 _24920_ (.Y(_06441_),
    .A(_06419_),
    .B(_06440_));
 sg13g2_mux2_1 _24921_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06441_),
    .X(_02008_));
 sg13g2_buf_1 _24922_ (.A(_02848_),
    .X(_06442_));
 sg13g2_mux2_1 _24923_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06441_),
    .X(_02009_));
 sg13g2_mux2_1 _24924_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06441_),
    .X(_02010_));
 sg13g2_mux2_1 _24925_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06441_),
    .X(_02011_));
 sg13g2_nor2_1 _24926_ (.A(_00233_),
    .B(_06431_),
    .Y(_06443_));
 sg13g2_buf_1 _24927_ (.A(_06443_),
    .X(_06444_));
 sg13g2_and2_1 _24928_ (.A(_06425_),
    .B(_06444_),
    .X(_06445_));
 sg13g2_buf_1 _24929_ (.A(_06445_),
    .X(_06446_));
 sg13g2_nand2_2 _24930_ (.Y(_06447_),
    .A(_06419_),
    .B(_06446_));
 sg13g2_mux2_1 _24931_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06447_),
    .X(_02012_));
 sg13g2_mux2_1 _24932_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06447_),
    .X(_02013_));
 sg13g2_mux2_1 _24933_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06447_),
    .X(_02014_));
 sg13g2_mux2_1 _24934_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06447_),
    .X(_02015_));
 sg13g2_mux2_1 _24935_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06428_),
    .X(_02016_));
 sg13g2_nor2_1 _24936_ (.A(_06422_),
    .B(_06423_),
    .Y(_06448_));
 sg13g2_and2_1 _24937_ (.A(_06444_),
    .B(_06448_),
    .X(_06449_));
 sg13g2_buf_1 _24938_ (.A(_06449_),
    .X(_06450_));
 sg13g2_nand2_2 _24939_ (.Y(_06451_),
    .A(_06419_),
    .B(_06450_));
 sg13g2_mux2_1 _24940_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06451_),
    .X(_02017_));
 sg13g2_mux2_1 _24941_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06451_),
    .X(_02018_));
 sg13g2_mux2_1 _24942_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06451_),
    .X(_02019_));
 sg13g2_mux2_1 _24943_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06451_),
    .X(_02020_));
 sg13g2_inv_1 _24944_ (.Y(_06452_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nand2_1 _24945_ (.Y(_06453_),
    .A(_06422_),
    .B(_06423_));
 sg13g2_nor3_1 _24946_ (.A(_06431_),
    .B(_06452_),
    .C(_06453_),
    .Y(_06454_));
 sg13g2_nand2_1 _24947_ (.Y(_06455_),
    .A(_06419_),
    .B(_06454_));
 sg13g2_buf_1 _24948_ (.A(_06455_),
    .X(_06456_));
 sg13g2_buf_1 _24949_ (.A(net423),
    .X(_06457_));
 sg13g2_mux2_1 _24950_ (.A0(_06417_),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net367),
    .X(_02021_));
 sg13g2_mux2_1 _24951_ (.A0(_06442_),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net367),
    .X(_02022_));
 sg13g2_mux2_1 _24952_ (.A0(_06429_),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(net367),
    .X(_02023_));
 sg13g2_mux2_1 _24953_ (.A0(_06436_),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(net367),
    .X(_02024_));
 sg13g2_and2_1 _24954_ (.A(_06438_),
    .B(_06444_),
    .X(_06458_));
 sg13g2_buf_1 _24955_ (.A(_06458_),
    .X(_06459_));
 sg13g2_nand2_2 _24956_ (.Y(_06460_),
    .A(_06419_),
    .B(_06459_));
 sg13g2_mux2_1 _24957_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06460_),
    .X(_02025_));
 sg13g2_mux2_1 _24958_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06460_),
    .X(_02026_));
 sg13g2_mux2_1 _24959_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06428_),
    .X(_02027_));
 sg13g2_mux2_1 _24960_ (.A0(_06429_),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06460_),
    .X(_02028_));
 sg13g2_mux2_1 _24961_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06460_),
    .X(_02029_));
 sg13g2_mux2_1 _24962_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06428_),
    .X(_02030_));
 sg13g2_and2_1 _24963_ (.A(_06421_),
    .B(_06448_),
    .X(_06461_));
 sg13g2_buf_1 _24964_ (.A(_06461_),
    .X(_06462_));
 sg13g2_nand2_2 _24965_ (.Y(_06463_),
    .A(_06419_),
    .B(_06462_));
 sg13g2_mux2_1 _24966_ (.A0(net960),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06463_),
    .X(_02031_));
 sg13g2_mux2_1 _24967_ (.A0(net958),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06463_),
    .X(_02032_));
 sg13g2_mux2_1 _24968_ (.A0(net959),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06463_),
    .X(_02033_));
 sg13g2_mux2_1 _24969_ (.A0(net835),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06463_),
    .X(_02034_));
 sg13g2_mux2_1 _24970_ (.A0(_06417_),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06435_),
    .X(_02035_));
 sg13g2_mux2_1 _24971_ (.A0(_06442_),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06435_),
    .X(_02036_));
 sg13g2_buf_1 _24972_ (.A(_02842_),
    .X(_06464_));
 sg13g2_nand2_1 _24973_ (.Y(_06465_),
    .A(_08444_),
    .B(_08658_));
 sg13g2_buf_4 _24974_ (.X(_06466_),
    .A(_06465_));
 sg13g2_nand2_1 _24975_ (.Y(_06467_),
    .A(_06421_),
    .B(_06425_));
 sg13g2_buf_2 _24976_ (.A(_06467_),
    .X(_06468_));
 sg13g2_nor2_2 _24977_ (.A(_06466_),
    .B(_06468_),
    .Y(_06469_));
 sg13g2_mux2_1 _24978_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(net957),
    .S(_06469_),
    .X(_02037_));
 sg13g2_buf_1 _24979_ (.A(_12043_),
    .X(_06470_));
 sg13g2_nor2_2 _24980_ (.A(_06466_),
    .B(_06433_),
    .Y(_06471_));
 sg13g2_mux2_1 _24981_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(_06470_),
    .S(_06471_),
    .X(_02038_));
 sg13g2_buf_1 _24982_ (.A(net988),
    .X(_06472_));
 sg13g2_mux2_1 _24983_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(_06472_),
    .S(_06471_),
    .X(_02039_));
 sg13g2_nand2_1 _24984_ (.Y(_06473_),
    .A(_06421_),
    .B(_06438_));
 sg13g2_buf_2 _24985_ (.A(_06473_),
    .X(_06474_));
 sg13g2_nor2_2 _24986_ (.A(_06466_),
    .B(_06474_),
    .Y(_06475_));
 sg13g2_mux2_1 _24987_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net957),
    .S(_06475_),
    .X(_02040_));
 sg13g2_buf_1 _24988_ (.A(_02848_),
    .X(_06476_));
 sg13g2_mux2_1 _24989_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net955),
    .S(_06475_),
    .X(_02041_));
 sg13g2_mux2_1 _24990_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net956),
    .S(_06475_),
    .X(_02042_));
 sg13g2_mux2_1 _24991_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net834),
    .S(_06475_),
    .X(_02043_));
 sg13g2_nand2_1 _24992_ (.Y(_06477_),
    .A(_06425_),
    .B(_06444_));
 sg13g2_buf_2 _24993_ (.A(_06477_),
    .X(_06478_));
 sg13g2_nor2_2 _24994_ (.A(_06466_),
    .B(_06478_),
    .Y(_06479_));
 sg13g2_mux2_1 _24995_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net957),
    .S(_06479_),
    .X(_02044_));
 sg13g2_mux2_1 _24996_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net955),
    .S(_06479_),
    .X(_02045_));
 sg13g2_mux2_1 _24997_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net956),
    .S(_06479_),
    .X(_02046_));
 sg13g2_mux2_1 _24998_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net834),
    .S(_06479_),
    .X(_02047_));
 sg13g2_mux2_1 _24999_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net955),
    .S(_06469_),
    .X(_02048_));
 sg13g2_nand2_1 _25000_ (.Y(_06480_),
    .A(_06444_),
    .B(_06448_));
 sg13g2_buf_2 _25001_ (.A(_06480_),
    .X(_06481_));
 sg13g2_nor2_2 _25002_ (.A(_06466_),
    .B(_06481_),
    .Y(_06482_));
 sg13g2_mux2_1 _25003_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net957),
    .S(_06482_),
    .X(_02049_));
 sg13g2_mux2_1 _25004_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(_06476_),
    .S(_06482_),
    .X(_02050_));
 sg13g2_mux2_1 _25005_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net956),
    .S(_06482_),
    .X(_02051_));
 sg13g2_mux2_1 _25006_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net834),
    .S(_06482_),
    .X(_02052_));
 sg13g2_or3_1 _25007_ (.A(_06431_),
    .B(_06452_),
    .C(_06453_),
    .X(_06483_));
 sg13g2_buf_1 _25008_ (.A(_06483_),
    .X(_06484_));
 sg13g2_nor2_1 _25009_ (.A(_06466_),
    .B(_06484_),
    .Y(_06485_));
 sg13g2_buf_2 _25010_ (.A(_06485_),
    .X(_06486_));
 sg13g2_mux2_1 _25011_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net957),
    .S(_06486_),
    .X(_02053_));
 sg13g2_mux2_1 _25012_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net955),
    .S(_06486_),
    .X(_02054_));
 sg13g2_mux2_1 _25013_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(_06470_),
    .S(_06486_),
    .X(_02055_));
 sg13g2_mux2_1 _25014_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net834),
    .S(_06486_),
    .X(_02056_));
 sg13g2_nand2_1 _25015_ (.Y(_06487_),
    .A(_06438_),
    .B(_06444_));
 sg13g2_buf_2 _25016_ (.A(_06487_),
    .X(_06488_));
 sg13g2_nor2_2 _25017_ (.A(_06466_),
    .B(_06488_),
    .Y(_06489_));
 sg13g2_mux2_1 _25018_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net957),
    .S(_06489_),
    .X(_02057_));
 sg13g2_mux2_1 _25019_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net955),
    .S(_06489_),
    .X(_02058_));
 sg13g2_mux2_1 _25020_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(net956),
    .S(_06469_),
    .X(_02059_));
 sg13g2_mux2_1 _25021_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(net956),
    .S(_06489_),
    .X(_02060_));
 sg13g2_mux2_1 _25022_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(_06472_),
    .S(_06489_),
    .X(_02061_));
 sg13g2_mux2_1 _25023_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(net834),
    .S(_06469_),
    .X(_02062_));
 sg13g2_nand2_1 _25024_ (.Y(_06490_),
    .A(_06421_),
    .B(_06448_));
 sg13g2_buf_2 _25025_ (.A(_06490_),
    .X(_06491_));
 sg13g2_nor2_2 _25026_ (.A(_06466_),
    .B(_06491_),
    .Y(_06492_));
 sg13g2_mux2_1 _25027_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(_06464_),
    .S(_06492_),
    .X(_02063_));
 sg13g2_mux2_1 _25028_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net955),
    .S(_06492_),
    .X(_02064_));
 sg13g2_mux2_1 _25029_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net956),
    .S(_06492_),
    .X(_02065_));
 sg13g2_mux2_1 _25030_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(net834),
    .S(_06492_),
    .X(_02066_));
 sg13g2_mux2_1 _25031_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net957),
    .S(_06471_),
    .X(_02067_));
 sg13g2_mux2_1 _25032_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(_06476_),
    .S(_06471_),
    .X(_02068_));
 sg13g2_nand2_1 _25033_ (.Y(_06493_),
    .A(_08444_),
    .B(_08517_));
 sg13g2_buf_4 _25034_ (.X(_06494_),
    .A(_06493_));
 sg13g2_nor2_2 _25035_ (.A(_06494_),
    .B(_06468_),
    .Y(_06495_));
 sg13g2_mux2_1 _25036_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(net957),
    .S(_06495_),
    .X(_02069_));
 sg13g2_nor2_2 _25037_ (.A(_06494_),
    .B(_06433_),
    .Y(_06496_));
 sg13g2_mux2_1 _25038_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net956),
    .S(_06496_),
    .X(_02070_));
 sg13g2_mux2_1 _25039_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(net834),
    .S(_06496_),
    .X(_02071_));
 sg13g2_buf_1 _25040_ (.A(_02842_),
    .X(_06497_));
 sg13g2_nor2_2 _25041_ (.A(_06494_),
    .B(_06474_),
    .Y(_06498_));
 sg13g2_mux2_1 _25042_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(net954),
    .S(_06498_),
    .X(_02072_));
 sg13g2_mux2_1 _25043_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(net955),
    .S(_06498_),
    .X(_02073_));
 sg13g2_buf_1 _25044_ (.A(_12043_),
    .X(_06499_));
 sg13g2_mux2_1 _25045_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net953),
    .S(_06498_),
    .X(_02074_));
 sg13g2_buf_1 _25046_ (.A(net988),
    .X(_06500_));
 sg13g2_mux2_1 _25047_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net833),
    .S(_06498_),
    .X(_02075_));
 sg13g2_nor2_2 _25048_ (.A(_06494_),
    .B(_06478_),
    .Y(_06501_));
 sg13g2_mux2_1 _25049_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net954),
    .S(_06501_),
    .X(_02076_));
 sg13g2_buf_1 _25050_ (.A(_02848_),
    .X(_06502_));
 sg13g2_mux2_1 _25051_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(net952),
    .S(_06501_),
    .X(_02077_));
 sg13g2_mux2_1 _25052_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net953),
    .S(_06501_),
    .X(_02078_));
 sg13g2_mux2_1 _25053_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net833),
    .S(_06501_),
    .X(_02079_));
 sg13g2_mux2_1 _25054_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net952),
    .S(_06495_),
    .X(_02080_));
 sg13g2_nor2_2 _25055_ (.A(_06494_),
    .B(_06481_),
    .Y(_06503_));
 sg13g2_mux2_1 _25056_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net954),
    .S(_06503_),
    .X(_02081_));
 sg13g2_mux2_1 _25057_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(_06502_),
    .S(_06503_),
    .X(_02082_));
 sg13g2_mux2_1 _25058_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net953),
    .S(_06503_),
    .X(_02083_));
 sg13g2_mux2_1 _25059_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net833),
    .S(_06503_),
    .X(_02084_));
 sg13g2_nor2_1 _25060_ (.A(_06494_),
    .B(_06484_),
    .Y(_06504_));
 sg13g2_buf_2 _25061_ (.A(_06504_),
    .X(_06505_));
 sg13g2_mux2_1 _25062_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net954),
    .S(_06505_),
    .X(_02085_));
 sg13g2_mux2_1 _25063_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net952),
    .S(_06505_),
    .X(_02086_));
 sg13g2_mux2_1 _25064_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net953),
    .S(_06505_),
    .X(_02087_));
 sg13g2_mux2_1 _25065_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net833),
    .S(_06505_),
    .X(_02088_));
 sg13g2_nor2_2 _25066_ (.A(_06494_),
    .B(_06488_),
    .Y(_06506_));
 sg13g2_mux2_1 _25067_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(net954),
    .S(_06506_),
    .X(_02089_));
 sg13g2_mux2_1 _25068_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net952),
    .S(_06506_),
    .X(_02090_));
 sg13g2_mux2_1 _25069_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(net953),
    .S(_06495_),
    .X(_02091_));
 sg13g2_mux2_1 _25070_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(net953),
    .S(_06506_),
    .X(_02092_));
 sg13g2_mux2_1 _25071_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(net833),
    .S(_06506_),
    .X(_02093_));
 sg13g2_mux2_1 _25072_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(net833),
    .S(_06495_),
    .X(_02094_));
 sg13g2_nor2_2 _25073_ (.A(_06494_),
    .B(_06491_),
    .Y(_06507_));
 sg13g2_mux2_1 _25074_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net954),
    .S(_06507_),
    .X(_02095_));
 sg13g2_mux2_1 _25075_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(_06502_),
    .S(_06507_),
    .X(_02096_));
 sg13g2_mux2_1 _25076_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net953),
    .S(_06507_),
    .X(_02097_));
 sg13g2_mux2_1 _25077_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net833),
    .S(_06507_),
    .X(_02098_));
 sg13g2_mux2_1 _25078_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net954),
    .S(_06496_),
    .X(_02099_));
 sg13g2_mux2_1 _25079_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net952),
    .S(_06496_),
    .X(_02100_));
 sg13g2_nand2_2 _25080_ (.Y(_06508_),
    .A(net451),
    .B(_06427_));
 sg13g2_mux2_1 _25081_ (.A0(net960),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06508_),
    .X(_02101_));
 sg13g2_and2_1 _25082_ (.A(_08996_),
    .B(_06434_),
    .X(_06509_));
 sg13g2_buf_1 _25083_ (.A(_06509_),
    .X(_06510_));
 sg13g2_mux2_1 _25084_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net953),
    .S(_06510_),
    .X(_02102_));
 sg13g2_mux2_1 _25085_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(_06500_),
    .S(_06510_),
    .X(_02103_));
 sg13g2_nand2_2 _25086_ (.Y(_06511_),
    .A(net451),
    .B(_06440_));
 sg13g2_mux2_1 _25087_ (.A0(net960),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06511_),
    .X(_02104_));
 sg13g2_mux2_1 _25088_ (.A0(net958),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06511_),
    .X(_02105_));
 sg13g2_mux2_1 _25089_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06511_),
    .X(_02106_));
 sg13g2_mux2_1 _25090_ (.A0(net835),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06511_),
    .X(_02107_));
 sg13g2_buf_1 _25091_ (.A(_02842_),
    .X(_06512_));
 sg13g2_nand2_2 _25092_ (.Y(_06513_),
    .A(net451),
    .B(_06446_));
 sg13g2_mux2_1 _25093_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06513_),
    .X(_02108_));
 sg13g2_mux2_1 _25094_ (.A0(net958),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06513_),
    .X(_02109_));
 sg13g2_mux2_1 _25095_ (.A0(net959),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06513_),
    .X(_02110_));
 sg13g2_mux2_1 _25096_ (.A0(net835),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06513_),
    .X(_02111_));
 sg13g2_buf_1 _25097_ (.A(_02848_),
    .X(_06514_));
 sg13g2_mux2_1 _25098_ (.A0(net950),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06508_),
    .X(_02112_));
 sg13g2_nand2_2 _25099_ (.Y(_06515_),
    .A(net451),
    .B(_06450_));
 sg13g2_mux2_1 _25100_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06515_),
    .X(_02113_));
 sg13g2_mux2_1 _25101_ (.A0(net950),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06515_),
    .X(_02114_));
 sg13g2_buf_1 _25102_ (.A(_12043_),
    .X(_06516_));
 sg13g2_mux2_1 _25103_ (.A0(_06516_),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06515_),
    .X(_02115_));
 sg13g2_buf_1 _25104_ (.A(net988),
    .X(_06517_));
 sg13g2_mux2_1 _25105_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06515_),
    .X(_02116_));
 sg13g2_nand2_1 _25106_ (.Y(_06518_),
    .A(net451),
    .B(_06454_));
 sg13g2_buf_1 _25107_ (.A(_06518_),
    .X(_06519_));
 sg13g2_buf_1 _25108_ (.A(net293),
    .X(_06520_));
 sg13g2_mux2_1 _25109_ (.A0(_06512_),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net249),
    .X(_02117_));
 sg13g2_mux2_1 _25110_ (.A0(net950),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net249),
    .X(_02118_));
 sg13g2_mux2_1 _25111_ (.A0(_06516_),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(net249),
    .X(_02119_));
 sg13g2_mux2_1 _25112_ (.A0(_06517_),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(net249),
    .X(_02120_));
 sg13g2_nand2_2 _25113_ (.Y(_06521_),
    .A(net451),
    .B(_06459_));
 sg13g2_mux2_1 _25114_ (.A0(_06512_),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06521_),
    .X(_02121_));
 sg13g2_mux2_1 _25115_ (.A0(net950),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06521_),
    .X(_02122_));
 sg13g2_mux2_1 _25116_ (.A0(net949),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06508_),
    .X(_02123_));
 sg13g2_mux2_1 _25117_ (.A0(net949),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06521_),
    .X(_02124_));
 sg13g2_mux2_1 _25118_ (.A0(_06517_),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06521_),
    .X(_02125_));
 sg13g2_mux2_1 _25119_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06508_),
    .X(_02126_));
 sg13g2_nand2_2 _25120_ (.Y(_06522_),
    .A(net451),
    .B(_06462_));
 sg13g2_mux2_1 _25121_ (.A0(net951),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06522_),
    .X(_02127_));
 sg13g2_mux2_1 _25122_ (.A0(_06514_),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06522_),
    .X(_02128_));
 sg13g2_mux2_1 _25123_ (.A0(net949),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06522_),
    .X(_02129_));
 sg13g2_mux2_1 _25124_ (.A0(net832),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06522_),
    .X(_02130_));
 sg13g2_mux2_1 _25125_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net954),
    .S(_06510_),
    .X(_02131_));
 sg13g2_mux2_1 _25126_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net952),
    .S(_06510_),
    .X(_02132_));
 sg13g2_nand2_2 _25127_ (.Y(_06523_),
    .A(net638),
    .B(_06427_));
 sg13g2_mux2_1 _25128_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06523_),
    .X(_02133_));
 sg13g2_and2_1 _25129_ (.A(net638),
    .B(_06434_),
    .X(_06524_));
 sg13g2_buf_1 _25130_ (.A(_06524_),
    .X(_06525_));
 sg13g2_mux2_1 _25131_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(_06499_),
    .S(_06525_),
    .X(_02134_));
 sg13g2_mux2_1 _25132_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net833),
    .S(_06525_),
    .X(_02135_));
 sg13g2_nand2_2 _25133_ (.Y(_06526_),
    .A(net638),
    .B(_06440_));
 sg13g2_mux2_1 _25134_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06526_),
    .X(_02136_));
 sg13g2_mux2_1 _25135_ (.A0(net950),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06526_),
    .X(_02137_));
 sg13g2_mux2_1 _25136_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06526_),
    .X(_02138_));
 sg13g2_mux2_1 _25137_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06526_),
    .X(_02139_));
 sg13g2_nand2_2 _25138_ (.Y(_06527_),
    .A(net638),
    .B(_06446_));
 sg13g2_mux2_1 _25139_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06527_),
    .X(_02140_));
 sg13g2_mux2_1 _25140_ (.A0(net950),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06527_),
    .X(_02141_));
 sg13g2_mux2_1 _25141_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06527_),
    .X(_02142_));
 sg13g2_mux2_1 _25142_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06527_),
    .X(_02143_));
 sg13g2_mux2_1 _25143_ (.A0(net950),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06523_),
    .X(_02144_));
 sg13g2_nand2_2 _25144_ (.Y(_06528_),
    .A(net638),
    .B(_06450_));
 sg13g2_mux2_1 _25145_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06528_),
    .X(_02145_));
 sg13g2_mux2_1 _25146_ (.A0(_06514_),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06528_),
    .X(_02146_));
 sg13g2_mux2_1 _25147_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06528_),
    .X(_02147_));
 sg13g2_mux2_1 _25148_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06528_),
    .X(_02148_));
 sg13g2_and2_1 _25149_ (.A(_08511_),
    .B(_06454_),
    .X(_06529_));
 sg13g2_buf_2 _25150_ (.A(_06529_),
    .X(_06530_));
 sg13g2_mux2_1 _25151_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(_06497_),
    .S(_06530_),
    .X(_02149_));
 sg13g2_mux2_1 _25152_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net952),
    .S(_06530_),
    .X(_02150_));
 sg13g2_mux2_1 _25153_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(_06499_),
    .S(_06530_),
    .X(_02151_));
 sg13g2_mux2_1 _25154_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(_06500_),
    .S(_06530_),
    .X(_02152_));
 sg13g2_nand2_2 _25155_ (.Y(_06531_),
    .A(net638),
    .B(_06459_));
 sg13g2_mux2_1 _25156_ (.A0(net951),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06531_),
    .X(_02153_));
 sg13g2_mux2_1 _25157_ (.A0(net950),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06531_),
    .X(_02154_));
 sg13g2_mux2_1 _25158_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06523_),
    .X(_02155_));
 sg13g2_mux2_1 _25159_ (.A0(net949),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06531_),
    .X(_02156_));
 sg13g2_mux2_1 _25160_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06531_),
    .X(_02157_));
 sg13g2_mux2_1 _25161_ (.A0(net832),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06523_),
    .X(_02158_));
 sg13g2_nand2_2 _25162_ (.Y(_06532_),
    .A(net638),
    .B(_06462_));
 sg13g2_mux2_1 _25163_ (.A0(_06464_),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06532_),
    .X(_02159_));
 sg13g2_mux2_1 _25164_ (.A0(net955),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06532_),
    .X(_02160_));
 sg13g2_mux2_1 _25165_ (.A0(net956),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06532_),
    .X(_02161_));
 sg13g2_mux2_1 _25166_ (.A0(net834),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06532_),
    .X(_02162_));
 sg13g2_mux2_1 _25167_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(_06497_),
    .S(_06525_),
    .X(_02163_));
 sg13g2_mux2_1 _25168_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(net952),
    .S(_06525_),
    .X(_02164_));
 sg13g2_buf_1 _25169_ (.A(_02842_),
    .X(_06533_));
 sg13g2_nand2_1 _25170_ (.Y(_06534_),
    .A(net817),
    .B(_08658_));
 sg13g2_buf_4 _25171_ (.X(_06535_),
    .A(_06534_));
 sg13g2_nor2_2 _25172_ (.A(_06535_),
    .B(_06468_),
    .Y(_06536_));
 sg13g2_mux2_1 _25173_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(net948),
    .S(_06536_),
    .X(_02165_));
 sg13g2_buf_1 _25174_ (.A(_12043_),
    .X(_06537_));
 sg13g2_nor2_2 _25175_ (.A(_06535_),
    .B(_06433_),
    .Y(_06538_));
 sg13g2_mux2_1 _25176_ (.A0(\cpu.icache.r_data[5][10] ),
    .A1(_06537_),
    .S(_06538_),
    .X(_02166_));
 sg13g2_buf_1 _25177_ (.A(_02779_),
    .X(_06539_));
 sg13g2_mux2_1 _25178_ (.A0(\cpu.icache.r_data[5][11] ),
    .A1(_06539_),
    .S(_06538_),
    .X(_02167_));
 sg13g2_nor2_2 _25179_ (.A(_06535_),
    .B(_06474_),
    .Y(_06540_));
 sg13g2_mux2_1 _25180_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(net948),
    .S(_06540_),
    .X(_02168_));
 sg13g2_buf_1 _25181_ (.A(_02848_),
    .X(_06541_));
 sg13g2_mux2_1 _25182_ (.A0(\cpu.icache.r_data[5][13] ),
    .A1(net946),
    .S(_06540_),
    .X(_02169_));
 sg13g2_mux2_1 _25183_ (.A0(\cpu.icache.r_data[5][14] ),
    .A1(net947),
    .S(_06540_),
    .X(_02170_));
 sg13g2_mux2_1 _25184_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(net831),
    .S(_06540_),
    .X(_02171_));
 sg13g2_nor2_2 _25185_ (.A(_06535_),
    .B(_06478_),
    .Y(_06542_));
 sg13g2_mux2_1 _25186_ (.A0(\cpu.icache.r_data[5][16] ),
    .A1(net948),
    .S(_06542_),
    .X(_02172_));
 sg13g2_mux2_1 _25187_ (.A0(\cpu.icache.r_data[5][17] ),
    .A1(net946),
    .S(_06542_),
    .X(_02173_));
 sg13g2_mux2_1 _25188_ (.A0(\cpu.icache.r_data[5][18] ),
    .A1(net947),
    .S(_06542_),
    .X(_02174_));
 sg13g2_mux2_1 _25189_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(net831),
    .S(_06542_),
    .X(_02175_));
 sg13g2_mux2_1 _25190_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(net946),
    .S(_06536_),
    .X(_02176_));
 sg13g2_nor2_2 _25191_ (.A(_06535_),
    .B(_06481_),
    .Y(_06543_));
 sg13g2_mux2_1 _25192_ (.A0(\cpu.icache.r_data[5][20] ),
    .A1(net948),
    .S(_06543_),
    .X(_02177_));
 sg13g2_mux2_1 _25193_ (.A0(\cpu.icache.r_data[5][21] ),
    .A1(net946),
    .S(_06543_),
    .X(_02178_));
 sg13g2_mux2_1 _25194_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(net947),
    .S(_06543_),
    .X(_02179_));
 sg13g2_mux2_1 _25195_ (.A0(\cpu.icache.r_data[5][23] ),
    .A1(net831),
    .S(_06543_),
    .X(_02180_));
 sg13g2_nor2_1 _25196_ (.A(_06535_),
    .B(_06484_),
    .Y(_06544_));
 sg13g2_buf_2 _25197_ (.A(_06544_),
    .X(_06545_));
 sg13g2_mux2_1 _25198_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(_06533_),
    .S(_06545_),
    .X(_02181_));
 sg13g2_mux2_1 _25199_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(_06541_),
    .S(_06545_),
    .X(_02182_));
 sg13g2_mux2_1 _25200_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(net947),
    .S(_06545_),
    .X(_02183_));
 sg13g2_mux2_1 _25201_ (.A0(\cpu.icache.r_data[5][27] ),
    .A1(net831),
    .S(_06545_),
    .X(_02184_));
 sg13g2_nor2_2 _25202_ (.A(_06535_),
    .B(_06488_),
    .Y(_06546_));
 sg13g2_mux2_1 _25203_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(net948),
    .S(_06546_),
    .X(_02185_));
 sg13g2_mux2_1 _25204_ (.A0(\cpu.icache.r_data[5][29] ),
    .A1(net946),
    .S(_06546_),
    .X(_02186_));
 sg13g2_mux2_1 _25205_ (.A0(\cpu.icache.r_data[5][2] ),
    .A1(net947),
    .S(_06536_),
    .X(_02187_));
 sg13g2_mux2_1 _25206_ (.A0(\cpu.icache.r_data[5][30] ),
    .A1(net947),
    .S(_06546_),
    .X(_02188_));
 sg13g2_mux2_1 _25207_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(net831),
    .S(_06546_),
    .X(_02189_));
 sg13g2_mux2_1 _25208_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(net831),
    .S(_06536_),
    .X(_02190_));
 sg13g2_nor2_2 _25209_ (.A(_06535_),
    .B(_06491_),
    .Y(_06547_));
 sg13g2_mux2_1 _25210_ (.A0(\cpu.icache.r_data[5][4] ),
    .A1(net948),
    .S(_06547_),
    .X(_02191_));
 sg13g2_mux2_1 _25211_ (.A0(\cpu.icache.r_data[5][5] ),
    .A1(net946),
    .S(_06547_),
    .X(_02192_));
 sg13g2_mux2_1 _25212_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(net947),
    .S(_06547_),
    .X(_02193_));
 sg13g2_mux2_1 _25213_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(net831),
    .S(_06547_),
    .X(_02194_));
 sg13g2_mux2_1 _25214_ (.A0(\cpu.icache.r_data[5][8] ),
    .A1(_06533_),
    .S(_06538_),
    .X(_02195_));
 sg13g2_mux2_1 _25215_ (.A0(\cpu.icache.r_data[5][9] ),
    .A1(_06541_),
    .S(_06538_),
    .X(_02196_));
 sg13g2_nand2_1 _25216_ (.Y(_06548_),
    .A(net817),
    .B(_08517_));
 sg13g2_buf_4 _25217_ (.X(_06549_),
    .A(_06548_));
 sg13g2_nor2_2 _25218_ (.A(_06549_),
    .B(_06468_),
    .Y(_06550_));
 sg13g2_mux2_1 _25219_ (.A0(\cpu.icache.r_data[6][0] ),
    .A1(net948),
    .S(_06550_),
    .X(_02197_));
 sg13g2_nor2_2 _25220_ (.A(_06549_),
    .B(_06433_),
    .Y(_06551_));
 sg13g2_mux2_1 _25221_ (.A0(\cpu.icache.r_data[6][10] ),
    .A1(_06537_),
    .S(_06551_),
    .X(_02198_));
 sg13g2_mux2_1 _25222_ (.A0(\cpu.icache.r_data[6][11] ),
    .A1(_06539_),
    .S(_06551_),
    .X(_02199_));
 sg13g2_nor2_2 _25223_ (.A(_06549_),
    .B(_06474_),
    .Y(_06552_));
 sg13g2_mux2_1 _25224_ (.A0(\cpu.icache.r_data[6][12] ),
    .A1(net948),
    .S(_06552_),
    .X(_02200_));
 sg13g2_mux2_1 _25225_ (.A0(\cpu.icache.r_data[6][13] ),
    .A1(net946),
    .S(_06552_),
    .X(_02201_));
 sg13g2_mux2_1 _25226_ (.A0(\cpu.icache.r_data[6][14] ),
    .A1(net947),
    .S(_06552_),
    .X(_02202_));
 sg13g2_mux2_1 _25227_ (.A0(\cpu.icache.r_data[6][15] ),
    .A1(net831),
    .S(_06552_),
    .X(_02203_));
 sg13g2_buf_1 _25228_ (.A(_02842_),
    .X(_06553_));
 sg13g2_nor2_2 _25229_ (.A(_06549_),
    .B(_06478_),
    .Y(_06554_));
 sg13g2_mux2_1 _25230_ (.A0(\cpu.icache.r_data[6][16] ),
    .A1(net945),
    .S(_06554_),
    .X(_02204_));
 sg13g2_mux2_1 _25231_ (.A0(\cpu.icache.r_data[6][17] ),
    .A1(net946),
    .S(_06554_),
    .X(_02205_));
 sg13g2_buf_1 _25232_ (.A(_12043_),
    .X(_06555_));
 sg13g2_mux2_1 _25233_ (.A0(\cpu.icache.r_data[6][18] ),
    .A1(net944),
    .S(_06554_),
    .X(_02206_));
 sg13g2_buf_2 _25234_ (.A(_11998_),
    .X(_06556_));
 sg13g2_mux2_1 _25235_ (.A0(\cpu.icache.r_data[6][19] ),
    .A1(net943),
    .S(_06554_),
    .X(_02207_));
 sg13g2_buf_1 _25236_ (.A(_02848_),
    .X(_06557_));
 sg13g2_mux2_1 _25237_ (.A0(\cpu.icache.r_data[6][1] ),
    .A1(net942),
    .S(_06550_),
    .X(_02208_));
 sg13g2_nor2_2 _25238_ (.A(_06549_),
    .B(_06481_),
    .Y(_06558_));
 sg13g2_mux2_1 _25239_ (.A0(\cpu.icache.r_data[6][20] ),
    .A1(net945),
    .S(_06558_),
    .X(_02209_));
 sg13g2_mux2_1 _25240_ (.A0(\cpu.icache.r_data[6][21] ),
    .A1(net942),
    .S(_06558_),
    .X(_02210_));
 sg13g2_mux2_1 _25241_ (.A0(\cpu.icache.r_data[6][22] ),
    .A1(net944),
    .S(_06558_),
    .X(_02211_));
 sg13g2_mux2_1 _25242_ (.A0(\cpu.icache.r_data[6][23] ),
    .A1(net943),
    .S(_06558_),
    .X(_02212_));
 sg13g2_nor2_1 _25243_ (.A(_06549_),
    .B(_06484_),
    .Y(_06559_));
 sg13g2_buf_2 _25244_ (.A(_06559_),
    .X(_06560_));
 sg13g2_mux2_1 _25245_ (.A0(\cpu.icache.r_data[6][24] ),
    .A1(_06553_),
    .S(_06560_),
    .X(_02213_));
 sg13g2_mux2_1 _25246_ (.A0(\cpu.icache.r_data[6][25] ),
    .A1(net942),
    .S(_06560_),
    .X(_02214_));
 sg13g2_mux2_1 _25247_ (.A0(\cpu.icache.r_data[6][26] ),
    .A1(_06555_),
    .S(_06560_),
    .X(_02215_));
 sg13g2_mux2_1 _25248_ (.A0(\cpu.icache.r_data[6][27] ),
    .A1(_06556_),
    .S(_06560_),
    .X(_02216_));
 sg13g2_nor2_2 _25249_ (.A(_06549_),
    .B(_06488_),
    .Y(_06561_));
 sg13g2_mux2_1 _25250_ (.A0(\cpu.icache.r_data[6][28] ),
    .A1(_06553_),
    .S(_06561_),
    .X(_02217_));
 sg13g2_mux2_1 _25251_ (.A0(\cpu.icache.r_data[6][29] ),
    .A1(net942),
    .S(_06561_),
    .X(_02218_));
 sg13g2_mux2_1 _25252_ (.A0(\cpu.icache.r_data[6][2] ),
    .A1(net944),
    .S(_06550_),
    .X(_02219_));
 sg13g2_mux2_1 _25253_ (.A0(\cpu.icache.r_data[6][30] ),
    .A1(net944),
    .S(_06561_),
    .X(_02220_));
 sg13g2_mux2_1 _25254_ (.A0(\cpu.icache.r_data[6][31] ),
    .A1(_06556_),
    .S(_06561_),
    .X(_02221_));
 sg13g2_mux2_1 _25255_ (.A0(\cpu.icache.r_data[6][3] ),
    .A1(net943),
    .S(_06550_),
    .X(_02222_));
 sg13g2_nor2_2 _25256_ (.A(_06549_),
    .B(_06491_),
    .Y(_06562_));
 sg13g2_mux2_1 _25257_ (.A0(\cpu.icache.r_data[6][4] ),
    .A1(net945),
    .S(_06562_),
    .X(_02223_));
 sg13g2_mux2_1 _25258_ (.A0(\cpu.icache.r_data[6][5] ),
    .A1(_06557_),
    .S(_06562_),
    .X(_02224_));
 sg13g2_mux2_1 _25259_ (.A0(\cpu.icache.r_data[6][6] ),
    .A1(net944),
    .S(_06562_),
    .X(_02225_));
 sg13g2_mux2_1 _25260_ (.A0(\cpu.icache.r_data[6][7] ),
    .A1(net943),
    .S(_06562_),
    .X(_02226_));
 sg13g2_mux2_1 _25261_ (.A0(\cpu.icache.r_data[6][8] ),
    .A1(net945),
    .S(_06551_),
    .X(_02227_));
 sg13g2_mux2_1 _25262_ (.A0(\cpu.icache.r_data[6][9] ),
    .A1(net942),
    .S(_06551_),
    .X(_02228_));
 sg13g2_nand2_1 _25263_ (.Y(_06563_),
    .A(net817),
    .B(_08778_));
 sg13g2_buf_4 _25264_ (.X(_06564_),
    .A(_06563_));
 sg13g2_nor2_2 _25265_ (.A(_06564_),
    .B(_06468_),
    .Y(_06565_));
 sg13g2_mux2_1 _25266_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(net945),
    .S(_06565_),
    .X(_02229_));
 sg13g2_nor2_2 _25267_ (.A(_06564_),
    .B(_06433_),
    .Y(_06566_));
 sg13g2_mux2_1 _25268_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(_06555_),
    .S(_06566_),
    .X(_02230_));
 sg13g2_mux2_1 _25269_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net943),
    .S(_06566_),
    .X(_02231_));
 sg13g2_nor2_2 _25270_ (.A(_06564_),
    .B(_06474_),
    .Y(_06567_));
 sg13g2_mux2_1 _25271_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(net945),
    .S(_06567_),
    .X(_02232_));
 sg13g2_mux2_1 _25272_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(net942),
    .S(_06567_),
    .X(_02233_));
 sg13g2_mux2_1 _25273_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net944),
    .S(_06567_),
    .X(_02234_));
 sg13g2_mux2_1 _25274_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(net943),
    .S(_06567_),
    .X(_02235_));
 sg13g2_nor2_2 _25275_ (.A(_06564_),
    .B(_06478_),
    .Y(_06568_));
 sg13g2_mux2_1 _25276_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(net945),
    .S(_06568_),
    .X(_02236_));
 sg13g2_mux2_1 _25277_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net942),
    .S(_06568_),
    .X(_02237_));
 sg13g2_mux2_1 _25278_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(net944),
    .S(_06568_),
    .X(_02238_));
 sg13g2_mux2_1 _25279_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(net943),
    .S(_06568_),
    .X(_02239_));
 sg13g2_mux2_1 _25280_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net942),
    .S(_06565_),
    .X(_02240_));
 sg13g2_nor2_2 _25281_ (.A(_06564_),
    .B(_06481_),
    .Y(_06569_));
 sg13g2_mux2_1 _25282_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net945),
    .S(_06569_),
    .X(_02241_));
 sg13g2_mux2_1 _25283_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(_06557_),
    .S(_06569_),
    .X(_02242_));
 sg13g2_mux2_1 _25284_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net944),
    .S(_06569_),
    .X(_02243_));
 sg13g2_mux2_1 _25285_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net943),
    .S(_06569_),
    .X(_02244_));
 sg13g2_nor2_1 _25286_ (.A(_06564_),
    .B(_06484_),
    .Y(_06570_));
 sg13g2_buf_2 _25287_ (.A(_06570_),
    .X(_06571_));
 sg13g2_mux2_1 _25288_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1015),
    .S(_06571_),
    .X(_02245_));
 sg13g2_mux2_1 _25289_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net1008),
    .S(_06571_),
    .X(_02246_));
 sg13g2_mux2_1 _25290_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net1011),
    .S(_06571_),
    .X(_02247_));
 sg13g2_mux2_1 _25291_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net1010),
    .S(_06571_),
    .X(_02248_));
 sg13g2_nor2_2 _25292_ (.A(_06564_),
    .B(_06488_),
    .Y(_06572_));
 sg13g2_mux2_1 _25293_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1015),
    .S(_06572_),
    .X(_02249_));
 sg13g2_mux2_1 _25294_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net1008),
    .S(_06572_),
    .X(_02250_));
 sg13g2_mux2_1 _25295_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net1011),
    .S(_06565_),
    .X(_02251_));
 sg13g2_mux2_1 _25296_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_11926_),
    .S(_06572_),
    .X(_02252_));
 sg13g2_mux2_1 _25297_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net1010),
    .S(_06572_),
    .X(_02253_));
 sg13g2_mux2_1 _25298_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_11941_),
    .S(_06565_),
    .X(_02254_));
 sg13g2_nor2_2 _25299_ (.A(_06564_),
    .B(_06491_),
    .Y(_06573_));
 sg13g2_mux2_1 _25300_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_11905_),
    .S(_06573_),
    .X(_02255_));
 sg13g2_mux2_1 _25301_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_11960_),
    .S(_06573_),
    .X(_02256_));
 sg13g2_mux2_1 _25302_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_11926_),
    .S(_06573_),
    .X(_02257_));
 sg13g2_mux2_1 _25303_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_11941_),
    .S(_06573_),
    .X(_02258_));
 sg13g2_mux2_1 _25304_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_11905_),
    .S(_06566_),
    .X(_02259_));
 sg13g2_mux2_1 _25305_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_11960_),
    .S(_06566_),
    .X(_02260_));
 sg13g2_mux2_1 _25306_ (.A0(net977),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(_06457_),
    .X(_02264_));
 sg13g2_buf_1 _25307_ (.A(_06456_),
    .X(_06574_));
 sg13g2_buf_1 _25308_ (.A(_06455_),
    .X(_06575_));
 sg13g2_nand2_1 _25309_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net422));
 sg13g2_o21ai_1 _25310_ (.B1(_06576_),
    .Y(_02265_),
    .A1(net453),
    .A2(net366));
 sg13g2_nand2_1 _25311_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(net422));
 sg13g2_o21ai_1 _25312_ (.B1(_06577_),
    .Y(_02266_),
    .A1(net454),
    .A2(net366));
 sg13g2_nand2_1 _25313_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net422));
 sg13g2_o21ai_1 _25314_ (.B1(_06578_),
    .Y(_02267_),
    .A1(net413),
    .A2(net366));
 sg13g2_nand2_1 _25315_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net422));
 sg13g2_o21ai_1 _25316_ (.B1(_06579_),
    .Y(_02268_),
    .A1(net415),
    .A2(net366));
 sg13g2_nand2_1 _25317_ (.Y(_06580_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(_06575_));
 sg13g2_o21ai_1 _25318_ (.B1(_06580_),
    .Y(_02269_),
    .A1(net455),
    .A2(_06574_));
 sg13g2_nand2_1 _25319_ (.Y(_06581_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net422));
 sg13g2_o21ai_1 _25320_ (.B1(_06581_),
    .Y(_02270_),
    .A1(net411),
    .A2(net366));
 sg13g2_nand2_1 _25321_ (.Y(_06582_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net423));
 sg13g2_o21ai_1 _25322_ (.B1(_06582_),
    .Y(_02271_),
    .A1(net414),
    .A2(_06574_));
 sg13g2_nand2_1 _25323_ (.Y(_06583_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net423));
 sg13g2_o21ai_1 _25324_ (.B1(_06583_),
    .Y(_02272_),
    .A1(net412),
    .A2(net366));
 sg13g2_nand2_1 _25325_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net423));
 sg13g2_o21ai_1 _25326_ (.B1(_06584_),
    .Y(_02273_),
    .A1(net510),
    .A2(net366));
 sg13g2_mux2_1 _25327_ (.A0(net976),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net422),
    .X(_02274_));
 sg13g2_mux2_1 _25328_ (.A0(net975),
    .A1(\cpu.icache.r_tag[0][7] ),
    .S(_06575_),
    .X(_02275_));
 sg13g2_nand2_1 _25329_ (.Y(_06585_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(_06456_));
 sg13g2_o21ai_1 _25330_ (.B1(_06585_),
    .Y(_02276_),
    .A1(net1064),
    .A2(net367));
 sg13g2_mux2_1 _25331_ (.A0(net974),
    .A1(\cpu.icache.r_tag[0][9] ),
    .S(net422),
    .X(_02277_));
 sg13g2_mux2_1 _25332_ (.A0(net973),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net422),
    .X(_02278_));
 sg13g2_nand2_1 _25333_ (.Y(_06586_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net423));
 sg13g2_o21ai_1 _25334_ (.B1(_06586_),
    .Y(_02279_),
    .A1(net1063),
    .A2(_06457_));
 sg13g2_nand2_1 _25335_ (.Y(_06587_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(net423));
 sg13g2_o21ai_1 _25336_ (.B1(_06587_),
    .Y(_02280_),
    .A1(net362),
    .A2(net367));
 sg13g2_nand2_1 _25337_ (.Y(_06588_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(net423));
 sg13g2_o21ai_1 _25338_ (.B1(_06588_),
    .Y(_02281_),
    .A1(net361),
    .A2(net367));
 sg13g2_nand2_1 _25339_ (.Y(_06589_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net423));
 sg13g2_o21ai_1 _25340_ (.B1(_06589_),
    .Y(_02282_),
    .A1(net452),
    .A2(net367));
 sg13g2_nor2b_1 _25341_ (.A(_06453_),
    .B_N(_06444_),
    .Y(_06590_));
 sg13g2_buf_1 _25342_ (.A(_06590_),
    .X(_06591_));
 sg13g2_nand2_1 _25343_ (.Y(_06592_),
    .A(_08474_),
    .B(_06591_));
 sg13g2_buf_1 _25344_ (.A(_06592_),
    .X(_06593_));
 sg13g2_buf_1 _25345_ (.A(_06593_),
    .X(_06594_));
 sg13g2_mux2_1 _25346_ (.A0(net977),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net248),
    .X(_02283_));
 sg13g2_buf_1 _25347_ (.A(_06593_),
    .X(_06595_));
 sg13g2_nand2_1 _25348_ (.Y(_06596_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net248));
 sg13g2_o21ai_1 _25349_ (.B1(_06596_),
    .Y(_02284_),
    .A1(net453),
    .A2(net247));
 sg13g2_buf_1 _25350_ (.A(_06593_),
    .X(_06597_));
 sg13g2_nand2_1 _25351_ (.Y(_06598_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net246));
 sg13g2_o21ai_1 _25352_ (.B1(_06598_),
    .Y(_02285_),
    .A1(net454),
    .A2(net247));
 sg13g2_nand2_1 _25353_ (.Y(_06599_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(net246));
 sg13g2_o21ai_1 _25354_ (.B1(_06599_),
    .Y(_02286_),
    .A1(net413),
    .A2(net247));
 sg13g2_nand2_1 _25355_ (.Y(_06600_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net246));
 sg13g2_o21ai_1 _25356_ (.B1(_06600_),
    .Y(_02287_),
    .A1(net415),
    .A2(_06595_));
 sg13g2_nand2_1 _25357_ (.Y(_06601_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net246));
 sg13g2_o21ai_1 _25358_ (.B1(_06601_),
    .Y(_02288_),
    .A1(net455),
    .A2(net247));
 sg13g2_nand2_1 _25359_ (.Y(_06602_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net246));
 sg13g2_o21ai_1 _25360_ (.B1(_06602_),
    .Y(_02289_),
    .A1(_08841_),
    .A2(net247));
 sg13g2_nand2_1 _25361_ (.Y(_06603_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(net246));
 sg13g2_o21ai_1 _25362_ (.B1(_06603_),
    .Y(_02290_),
    .A1(_08581_),
    .A2(net247));
 sg13g2_nand2_1 _25363_ (.Y(_06604_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net246));
 sg13g2_o21ai_1 _25364_ (.B1(_06604_),
    .Y(_02291_),
    .A1(net412),
    .A2(net247));
 sg13g2_nand2_1 _25365_ (.Y(_06605_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net246));
 sg13g2_o21ai_1 _25366_ (.B1(_06605_),
    .Y(_02292_),
    .A1(net510),
    .A2(net247));
 sg13g2_mux2_1 _25367_ (.A0(net976),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net248),
    .X(_02293_));
 sg13g2_mux2_1 _25368_ (.A0(net975),
    .A1(\cpu.icache.r_tag[1][7] ),
    .S(_06594_),
    .X(_02294_));
 sg13g2_nand2_1 _25369_ (.Y(_06606_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(_06597_));
 sg13g2_o21ai_1 _25370_ (.B1(_06606_),
    .Y(_02295_),
    .A1(net1064),
    .A2(_06595_));
 sg13g2_mux2_1 _25371_ (.A0(net974),
    .A1(\cpu.icache.r_tag[1][9] ),
    .S(_06594_),
    .X(_02296_));
 sg13g2_mux2_1 _25372_ (.A0(net973),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net248),
    .X(_02297_));
 sg13g2_nand2_1 _25373_ (.Y(_06607_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(_06597_));
 sg13g2_o21ai_1 _25374_ (.B1(_06607_),
    .Y(_02298_),
    .A1(net1063),
    .A2(net248));
 sg13g2_nand2_1 _25375_ (.Y(_06608_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06593_));
 sg13g2_o21ai_1 _25376_ (.B1(_06608_),
    .Y(_02299_),
    .A1(net362),
    .A2(net248));
 sg13g2_nand2_1 _25377_ (.Y(_06609_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06593_));
 sg13g2_o21ai_1 _25378_ (.B1(_06609_),
    .Y(_02300_),
    .A1(net361),
    .A2(net248));
 sg13g2_nand2_1 _25379_ (.Y(_06610_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06593_));
 sg13g2_o21ai_1 _25380_ (.B1(_06610_),
    .Y(_02301_),
    .A1(net452),
    .A2(net248));
 sg13g2_nand2_1 _25381_ (.Y(_06611_),
    .A(_08488_),
    .B(_06591_));
 sg13g2_buf_1 _25382_ (.A(_06611_),
    .X(_06612_));
 sg13g2_buf_1 _25383_ (.A(_06612_),
    .X(_06613_));
 sg13g2_mux2_1 _25384_ (.A0(net977),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net292),
    .X(_02302_));
 sg13g2_buf_1 _25385_ (.A(_06612_),
    .X(_06614_));
 sg13g2_nand2_1 _25386_ (.Y(_06615_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(net292));
 sg13g2_o21ai_1 _25387_ (.B1(_06615_),
    .Y(_02303_),
    .A1(net453),
    .A2(net291));
 sg13g2_buf_1 _25388_ (.A(_06612_),
    .X(_06616_));
 sg13g2_nand2_1 _25389_ (.Y(_06617_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net290));
 sg13g2_o21ai_1 _25390_ (.B1(_06617_),
    .Y(_02304_),
    .A1(net454),
    .A2(net291));
 sg13g2_nand2_1 _25391_ (.Y(_06618_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net290));
 sg13g2_o21ai_1 _25392_ (.B1(_06618_),
    .Y(_02305_),
    .A1(net413),
    .A2(net291));
 sg13g2_nand2_1 _25393_ (.Y(_06619_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(_06616_));
 sg13g2_o21ai_1 _25394_ (.B1(_06619_),
    .Y(_02306_),
    .A1(net415),
    .A2(_06614_));
 sg13g2_nand2_1 _25395_ (.Y(_06620_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net290));
 sg13g2_o21ai_1 _25396_ (.B1(_06620_),
    .Y(_02307_),
    .A1(net455),
    .A2(net291));
 sg13g2_nand2_1 _25397_ (.Y(_06621_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net290));
 sg13g2_o21ai_1 _25398_ (.B1(_06621_),
    .Y(_02308_),
    .A1(net411),
    .A2(net291));
 sg13g2_nand2_1 _25399_ (.Y(_06622_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net290));
 sg13g2_o21ai_1 _25400_ (.B1(_06622_),
    .Y(_02309_),
    .A1(net414),
    .A2(_06614_));
 sg13g2_nand2_1 _25401_ (.Y(_06623_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net290));
 sg13g2_o21ai_1 _25402_ (.B1(_06623_),
    .Y(_02310_),
    .A1(net412),
    .A2(net291));
 sg13g2_nand2_1 _25403_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(_06616_));
 sg13g2_o21ai_1 _25404_ (.B1(_06624_),
    .Y(_02311_),
    .A1(net510),
    .A2(net291));
 sg13g2_mux2_1 _25405_ (.A0(net976),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net292),
    .X(_02312_));
 sg13g2_mux2_1 _25406_ (.A0(net975),
    .A1(\cpu.icache.r_tag[2][7] ),
    .S(net292),
    .X(_02313_));
 sg13g2_nand2_1 _25407_ (.Y(_06625_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(net290));
 sg13g2_o21ai_1 _25408_ (.B1(_06625_),
    .Y(_02314_),
    .A1(net1064),
    .A2(net291));
 sg13g2_mux2_1 _25409_ (.A0(net974),
    .A1(\cpu.icache.r_tag[2][9] ),
    .S(_06613_),
    .X(_02315_));
 sg13g2_mux2_1 _25410_ (.A0(net973),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net292),
    .X(_02316_));
 sg13g2_nand2_1 _25411_ (.Y(_06626_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(net290));
 sg13g2_o21ai_1 _25412_ (.B1(_06626_),
    .Y(_02317_),
    .A1(net1063),
    .A2(_06613_));
 sg13g2_nand2_1 _25413_ (.Y(_06627_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06612_));
 sg13g2_o21ai_1 _25414_ (.B1(_06627_),
    .Y(_02318_),
    .A1(net362),
    .A2(net292));
 sg13g2_nand2_1 _25415_ (.Y(_06628_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06612_));
 sg13g2_o21ai_1 _25416_ (.B1(_06628_),
    .Y(_02319_),
    .A1(net361),
    .A2(net292));
 sg13g2_nand2_1 _25417_ (.Y(_06629_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06612_));
 sg13g2_o21ai_1 _25418_ (.B1(_06629_),
    .Y(_02320_),
    .A1(net452),
    .A2(net292));
 sg13g2_mux2_1 _25419_ (.A0(net977),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net249),
    .X(_02321_));
 sg13g2_buf_1 _25420_ (.A(net293),
    .X(_06630_));
 sg13g2_buf_1 _25421_ (.A(_06518_),
    .X(_06631_));
 sg13g2_nand2_1 _25422_ (.Y(_06632_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net289));
 sg13g2_o21ai_1 _25423_ (.B1(_06632_),
    .Y(_02322_),
    .A1(net453),
    .A2(net245));
 sg13g2_nand2_1 _25424_ (.Y(_06633_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net289));
 sg13g2_o21ai_1 _25425_ (.B1(_06633_),
    .Y(_02323_),
    .A1(net454),
    .A2(net245));
 sg13g2_nand2_1 _25426_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net289));
 sg13g2_o21ai_1 _25427_ (.B1(_06634_),
    .Y(_02324_),
    .A1(net413),
    .A2(net245));
 sg13g2_nand2_1 _25428_ (.Y(_06635_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net289));
 sg13g2_o21ai_1 _25429_ (.B1(_06635_),
    .Y(_02325_),
    .A1(net415),
    .A2(net245));
 sg13g2_nand2_1 _25430_ (.Y(_06636_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net289));
 sg13g2_o21ai_1 _25431_ (.B1(_06636_),
    .Y(_02326_),
    .A1(net455),
    .A2(net245));
 sg13g2_nand2_1 _25432_ (.Y(_06637_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net289));
 sg13g2_o21ai_1 _25433_ (.B1(_06637_),
    .Y(_02327_),
    .A1(net411),
    .A2(_06630_));
 sg13g2_nand2_1 _25434_ (.Y(_06638_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net293));
 sg13g2_o21ai_1 _25435_ (.B1(_06638_),
    .Y(_02328_),
    .A1(net414),
    .A2(_06630_));
 sg13g2_nand2_1 _25436_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net293));
 sg13g2_o21ai_1 _25437_ (.B1(_06639_),
    .Y(_02329_),
    .A1(net412),
    .A2(net245));
 sg13g2_nand2_1 _25438_ (.Y(_06640_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net293));
 sg13g2_o21ai_1 _25439_ (.B1(_06640_),
    .Y(_02330_),
    .A1(net510),
    .A2(net245));
 sg13g2_mux2_1 _25440_ (.A0(net976),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net289),
    .X(_02331_));
 sg13g2_mux2_1 _25441_ (.A0(net975),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net289),
    .X(_02332_));
 sg13g2_nand2_1 _25442_ (.Y(_06641_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(_06519_));
 sg13g2_o21ai_1 _25443_ (.B1(_06641_),
    .Y(_02333_),
    .A1(net1064),
    .A2(_06520_));
 sg13g2_mux2_1 _25444_ (.A0(net974),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(_06631_),
    .X(_02334_));
 sg13g2_mux2_1 _25445_ (.A0(net973),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(_06631_),
    .X(_02335_));
 sg13g2_nand2_1 _25446_ (.Y(_06642_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(_06519_));
 sg13g2_o21ai_1 _25447_ (.B1(_06642_),
    .Y(_02336_),
    .A1(net1063),
    .A2(_06520_));
 sg13g2_nand2_1 _25448_ (.Y(_06643_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net293));
 sg13g2_o21ai_1 _25449_ (.B1(_06643_),
    .Y(_02337_),
    .A1(net362),
    .A2(net249));
 sg13g2_nand2_1 _25450_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net293));
 sg13g2_o21ai_1 _25451_ (.B1(_06644_),
    .Y(_02338_),
    .A1(net361),
    .A2(net249));
 sg13g2_nand2_1 _25452_ (.Y(_06645_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(net293));
 sg13g2_o21ai_1 _25453_ (.B1(_06645_),
    .Y(_02339_),
    .A1(net452),
    .A2(net249));
 sg13g2_nand2_1 _25454_ (.Y(_06646_),
    .A(_08511_),
    .B(_06591_));
 sg13g2_buf_1 _25455_ (.A(_06646_),
    .X(_06647_));
 sg13g2_buf_1 _25456_ (.A(_06647_),
    .X(_06648_));
 sg13g2_mux2_1 _25457_ (.A0(net977),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net421),
    .X(_02340_));
 sg13g2_buf_1 _25458_ (.A(_06647_),
    .X(_06649_));
 sg13g2_nand2_1 _25459_ (.Y(_06650_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(net421));
 sg13g2_o21ai_1 _25460_ (.B1(_06650_),
    .Y(_02341_),
    .A1(net453),
    .A2(_06649_));
 sg13g2_buf_1 _25461_ (.A(_06647_),
    .X(_06651_));
 sg13g2_nand2_1 _25462_ (.Y(_06652_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net419));
 sg13g2_o21ai_1 _25463_ (.B1(_06652_),
    .Y(_02342_),
    .A1(net454),
    .A2(net420));
 sg13g2_nand2_1 _25464_ (.Y(_06653_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net419));
 sg13g2_o21ai_1 _25465_ (.B1(_06653_),
    .Y(_02343_),
    .A1(net413),
    .A2(net420));
 sg13g2_nand2_1 _25466_ (.Y(_06654_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(net419));
 sg13g2_o21ai_1 _25467_ (.B1(_06654_),
    .Y(_02344_),
    .A1(net415),
    .A2(net420));
 sg13g2_nand2_1 _25468_ (.Y(_06655_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net419));
 sg13g2_o21ai_1 _25469_ (.B1(_06655_),
    .Y(_02345_),
    .A1(net455),
    .A2(net420));
 sg13g2_nand2_1 _25470_ (.Y(_06656_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net419));
 sg13g2_o21ai_1 _25471_ (.B1(_06656_),
    .Y(_02346_),
    .A1(net411),
    .A2(net420));
 sg13g2_nand2_1 _25472_ (.Y(_06657_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(_06651_));
 sg13g2_o21ai_1 _25473_ (.B1(_06657_),
    .Y(_02347_),
    .A1(net414),
    .A2(_06649_));
 sg13g2_nand2_1 _25474_ (.Y(_06658_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net419));
 sg13g2_o21ai_1 _25475_ (.B1(_06658_),
    .Y(_02348_),
    .A1(net412),
    .A2(net420));
 sg13g2_nand2_1 _25476_ (.Y(_06659_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net419));
 sg13g2_o21ai_1 _25477_ (.B1(_06659_),
    .Y(_02349_),
    .A1(net510),
    .A2(net420));
 sg13g2_mux2_1 _25478_ (.A0(net976),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net421),
    .X(_02350_));
 sg13g2_mux2_1 _25479_ (.A0(net975),
    .A1(\cpu.icache.r_tag[4][7] ),
    .S(net421),
    .X(_02351_));
 sg13g2_nand2_1 _25480_ (.Y(_06660_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(_06651_));
 sg13g2_o21ai_1 _25481_ (.B1(_06660_),
    .Y(_02352_),
    .A1(net1064),
    .A2(net420));
 sg13g2_mux2_1 _25482_ (.A0(net974),
    .A1(\cpu.icache.r_tag[4][9] ),
    .S(_06648_),
    .X(_02353_));
 sg13g2_mux2_1 _25483_ (.A0(net973),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net421),
    .X(_02354_));
 sg13g2_nand2_1 _25484_ (.Y(_06661_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(net419));
 sg13g2_o21ai_1 _25485_ (.B1(_06661_),
    .Y(_02355_),
    .A1(net1063),
    .A2(_06648_));
 sg13g2_nand2_1 _25486_ (.Y(_06662_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25487_ (.B1(_06662_),
    .Y(_02356_),
    .A1(net362),
    .A2(net421));
 sg13g2_nand2_1 _25488_ (.Y(_06663_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25489_ (.B1(_06663_),
    .Y(_02357_),
    .A1(net361),
    .A2(net421));
 sg13g2_nand2_1 _25490_ (.Y(_06664_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06647_));
 sg13g2_o21ai_1 _25491_ (.B1(_06664_),
    .Y(_02358_),
    .A1(net452),
    .A2(net421));
 sg13g2_nand2_1 _25492_ (.Y(_06665_),
    .A(_08564_),
    .B(_06591_));
 sg13g2_buf_1 _25493_ (.A(_06665_),
    .X(_06666_));
 sg13g2_buf_1 _25494_ (.A(_06666_),
    .X(_06667_));
 sg13g2_mux2_1 _25495_ (.A0(net977),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(_06667_),
    .X(_02359_));
 sg13g2_buf_1 _25496_ (.A(_06666_),
    .X(_06668_));
 sg13g2_nand2_1 _25497_ (.Y(_06669_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net365));
 sg13g2_o21ai_1 _25498_ (.B1(_06669_),
    .Y(_02360_),
    .A1(net453),
    .A2(_06668_));
 sg13g2_buf_1 _25499_ (.A(_06666_),
    .X(_06670_));
 sg13g2_nand2_1 _25500_ (.Y(_06671_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net363));
 sg13g2_o21ai_1 _25501_ (.B1(_06671_),
    .Y(_02361_),
    .A1(net454),
    .A2(net364));
 sg13g2_nand2_1 _25502_ (.Y(_06672_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(net363));
 sg13g2_o21ai_1 _25503_ (.B1(_06672_),
    .Y(_02362_),
    .A1(net413),
    .A2(net364));
 sg13g2_nand2_1 _25504_ (.Y(_06673_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(_06670_));
 sg13g2_o21ai_1 _25505_ (.B1(_06673_),
    .Y(_02363_),
    .A1(net415),
    .A2(_06668_));
 sg13g2_nand2_1 _25506_ (.Y(_06674_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net363));
 sg13g2_o21ai_1 _25507_ (.B1(_06674_),
    .Y(_02364_),
    .A1(net455),
    .A2(net364));
 sg13g2_nand2_1 _25508_ (.Y(_06675_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net363));
 sg13g2_o21ai_1 _25509_ (.B1(_06675_),
    .Y(_02365_),
    .A1(net411),
    .A2(net364));
 sg13g2_nand2_1 _25510_ (.Y(_06676_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(net363));
 sg13g2_o21ai_1 _25511_ (.B1(_06676_),
    .Y(_02366_),
    .A1(net414),
    .A2(net364));
 sg13g2_nand2_1 _25512_ (.Y(_06677_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(net363));
 sg13g2_o21ai_1 _25513_ (.B1(_06677_),
    .Y(_02367_),
    .A1(net412),
    .A2(net364));
 sg13g2_nand2_1 _25514_ (.Y(_06678_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net363));
 sg13g2_o21ai_1 _25515_ (.B1(_06678_),
    .Y(_02368_),
    .A1(net510),
    .A2(net364));
 sg13g2_mux2_1 _25516_ (.A0(net976),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(_06667_),
    .X(_02369_));
 sg13g2_mux2_1 _25517_ (.A0(net975),
    .A1(\cpu.icache.r_tag[5][7] ),
    .S(net365),
    .X(_02370_));
 sg13g2_nand2_1 _25518_ (.Y(_06679_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(_06670_));
 sg13g2_o21ai_1 _25519_ (.B1(_06679_),
    .Y(_02371_),
    .A1(net1064),
    .A2(net364));
 sg13g2_mux2_1 _25520_ (.A0(net974),
    .A1(\cpu.icache.r_tag[5][9] ),
    .S(net365),
    .X(_02372_));
 sg13g2_mux2_1 _25521_ (.A0(net973),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net365),
    .X(_02373_));
 sg13g2_nand2_1 _25522_ (.Y(_06680_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(net363));
 sg13g2_o21ai_1 _25523_ (.B1(_06680_),
    .Y(_02374_),
    .A1(net1063),
    .A2(net365));
 sg13g2_nand2_1 _25524_ (.Y(_06681_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06666_));
 sg13g2_o21ai_1 _25525_ (.B1(_06681_),
    .Y(_02375_),
    .A1(net362),
    .A2(net365));
 sg13g2_nand2_1 _25526_ (.Y(_06682_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06666_));
 sg13g2_o21ai_1 _25527_ (.B1(_06682_),
    .Y(_02376_),
    .A1(net361),
    .A2(net365));
 sg13g2_nand2_1 _25528_ (.Y(_06683_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06666_));
 sg13g2_o21ai_1 _25529_ (.B1(_06683_),
    .Y(_02377_),
    .A1(net452),
    .A2(net365));
 sg13g2_nand2_1 _25530_ (.Y(_06684_),
    .A(_08559_),
    .B(_06591_));
 sg13g2_buf_1 _25531_ (.A(_06684_),
    .X(_06685_));
 sg13g2_buf_1 _25532_ (.A(_06685_),
    .X(_06686_));
 sg13g2_mux2_1 _25533_ (.A0(_04534_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net418),
    .X(_02378_));
 sg13g2_buf_1 _25534_ (.A(_06685_),
    .X(_06687_));
 sg13g2_nand2_1 _25535_ (.Y(_06688_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(net418));
 sg13g2_o21ai_1 _25536_ (.B1(_06688_),
    .Y(_02379_),
    .A1(net453),
    .A2(net417));
 sg13g2_buf_1 _25537_ (.A(_06685_),
    .X(_06689_));
 sg13g2_nand2_1 _25538_ (.Y(_06690_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net416));
 sg13g2_o21ai_1 _25539_ (.B1(_06690_),
    .Y(_02380_),
    .A1(net454),
    .A2(net417));
 sg13g2_nand2_1 _25540_ (.Y(_06691_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net416));
 sg13g2_o21ai_1 _25541_ (.B1(_06691_),
    .Y(_02381_),
    .A1(net413),
    .A2(net417));
 sg13g2_nand2_1 _25542_ (.Y(_06692_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net416));
 sg13g2_o21ai_1 _25543_ (.B1(_06692_),
    .Y(_02382_),
    .A1(net415),
    .A2(net417));
 sg13g2_nand2_1 _25544_ (.Y(_06693_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net416));
 sg13g2_o21ai_1 _25545_ (.B1(_06693_),
    .Y(_02383_),
    .A1(net455),
    .A2(_06687_));
 sg13g2_nand2_1 _25546_ (.Y(_06694_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net416));
 sg13g2_o21ai_1 _25547_ (.B1(_06694_),
    .Y(_02384_),
    .A1(net411),
    .A2(net417));
 sg13g2_nand2_1 _25548_ (.Y(_06695_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net416));
 sg13g2_o21ai_1 _25549_ (.B1(_06695_),
    .Y(_02385_),
    .A1(net414),
    .A2(net417));
 sg13g2_nand2_1 _25550_ (.Y(_06696_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net416));
 sg13g2_o21ai_1 _25551_ (.B1(_06696_),
    .Y(_02386_),
    .A1(_08819_),
    .A2(net417));
 sg13g2_nand2_1 _25552_ (.Y(_06697_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net416));
 sg13g2_o21ai_1 _25553_ (.B1(_06697_),
    .Y(_02387_),
    .A1(net510),
    .A2(net417));
 sg13g2_mux2_1 _25554_ (.A0(_04562_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net418),
    .X(_02388_));
 sg13g2_mux2_1 _25555_ (.A0(_04589_),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(_06686_),
    .X(_02389_));
 sg13g2_nand2_1 _25556_ (.Y(_06698_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(_06689_));
 sg13g2_o21ai_1 _25557_ (.B1(_06698_),
    .Y(_02390_),
    .A1(net1064),
    .A2(_06687_));
 sg13g2_mux2_1 _25558_ (.A0(_04648_),
    .A1(\cpu.icache.r_tag[6][9] ),
    .S(_06686_),
    .X(_02391_));
 sg13g2_mux2_1 _25559_ (.A0(_04688_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net418),
    .X(_02392_));
 sg13g2_nand2_1 _25560_ (.Y(_06699_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06689_));
 sg13g2_o21ai_1 _25561_ (.B1(_06699_),
    .Y(_02393_),
    .A1(net1063),
    .A2(net418));
 sg13g2_nand2_1 _25562_ (.Y(_06700_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06685_));
 sg13g2_o21ai_1 _25563_ (.B1(_06700_),
    .Y(_02394_),
    .A1(net362),
    .A2(net418));
 sg13g2_nand2_1 _25564_ (.Y(_06701_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06685_));
 sg13g2_o21ai_1 _25565_ (.B1(_06701_),
    .Y(_02395_),
    .A1(net361),
    .A2(net418));
 sg13g2_nand2_1 _25566_ (.Y(_06702_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06685_));
 sg13g2_o21ai_1 _25567_ (.B1(_06702_),
    .Y(_02396_),
    .A1(net452),
    .A2(net418));
 sg13g2_nand2_1 _25568_ (.Y(_06703_),
    .A(_08553_),
    .B(_06591_));
 sg13g2_buf_1 _25569_ (.A(_06703_),
    .X(_06704_));
 sg13g2_buf_1 _25570_ (.A(_06704_),
    .X(_06705_));
 sg13g2_mux2_1 _25571_ (.A0(_04534_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net463),
    .X(_02397_));
 sg13g2_buf_1 _25572_ (.A(_06704_),
    .X(_06706_));
 sg13g2_nand2_1 _25573_ (.Y(_06707_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(net463));
 sg13g2_o21ai_1 _25574_ (.B1(_06707_),
    .Y(_02398_),
    .A1(_08752_),
    .A2(net462));
 sg13g2_buf_1 _25575_ (.A(_06704_),
    .X(_06708_));
 sg13g2_nand2_1 _25576_ (.Y(_06709_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net461));
 sg13g2_o21ai_1 _25577_ (.B1(_06709_),
    .Y(_02399_),
    .A1(net454),
    .A2(net462));
 sg13g2_nand2_1 _25578_ (.Y(_06710_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net461));
 sg13g2_o21ai_1 _25579_ (.B1(_06710_),
    .Y(_02400_),
    .A1(_08798_),
    .A2(net462));
 sg13g2_nand2_1 _25580_ (.Y(_06711_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(net461));
 sg13g2_o21ai_1 _25581_ (.B1(_06711_),
    .Y(_02401_),
    .A1(_08547_),
    .A2(_06706_));
 sg13g2_nand2_1 _25582_ (.Y(_06712_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(_06708_));
 sg13g2_o21ai_1 _25583_ (.B1(_06712_),
    .Y(_02402_),
    .A1(_08706_),
    .A2(_06706_));
 sg13g2_nand2_1 _25584_ (.Y(_06713_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net461));
 sg13g2_o21ai_1 _25585_ (.B1(_06713_),
    .Y(_02403_),
    .A1(net411),
    .A2(net462));
 sg13g2_nand2_1 _25586_ (.Y(_06714_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net461));
 sg13g2_o21ai_1 _25587_ (.B1(_06714_),
    .Y(_02404_),
    .A1(net414),
    .A2(net462));
 sg13g2_nand2_1 _25588_ (.Y(_06715_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net461));
 sg13g2_o21ai_1 _25589_ (.B1(_06715_),
    .Y(_02405_),
    .A1(net412),
    .A2(net462));
 sg13g2_nand2_1 _25590_ (.Y(_06716_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net461));
 sg13g2_o21ai_1 _25591_ (.B1(_06716_),
    .Y(_02406_),
    .A1(net510),
    .A2(net462));
 sg13g2_mux2_1 _25592_ (.A0(_04562_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net463),
    .X(_02407_));
 sg13g2_mux2_1 _25593_ (.A0(_04589_),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(_06705_),
    .X(_02408_));
 sg13g2_nand2_1 _25594_ (.Y(_06717_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(net461));
 sg13g2_o21ai_1 _25595_ (.B1(_06717_),
    .Y(_02409_),
    .A1(_08615_),
    .A2(net462));
 sg13g2_mux2_1 _25596_ (.A0(_04648_),
    .A1(\cpu.icache.r_tag[7][9] ),
    .S(_06705_),
    .X(_02410_));
 sg13g2_mux2_1 _25597_ (.A0(_04688_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net463),
    .X(_02411_));
 sg13g2_nand2_1 _25598_ (.Y(_06718_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(_06708_));
 sg13g2_o21ai_1 _25599_ (.B1(_06718_),
    .Y(_02412_),
    .A1(net1063),
    .A2(net463));
 sg13g2_nand2_1 _25600_ (.Y(_06719_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06704_));
 sg13g2_o21ai_1 _25601_ (.B1(_06719_),
    .Y(_02413_),
    .A1(_08439_),
    .A2(net463));
 sg13g2_nand2_1 _25602_ (.Y(_06720_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06704_));
 sg13g2_o21ai_1 _25603_ (.B1(_06720_),
    .Y(_02414_),
    .A1(_08507_),
    .A2(net463));
 sg13g2_nand2_1 _25604_ (.Y(_06721_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06704_));
 sg13g2_o21ai_1 _25605_ (.B1(_06721_),
    .Y(_02415_),
    .A1(net452),
    .A2(net463));
 sg13g2_buf_1 _25606_ (.A(_10038_),
    .X(_06722_));
 sg13g2_and2_1 _25607_ (.A(net128),
    .B(net594),
    .X(_06723_));
 sg13g2_buf_2 _25608_ (.A(_06723_),
    .X(_06724_));
 sg13g2_buf_1 _25609_ (.A(_06724_),
    .X(_06725_));
 sg13g2_mux2_1 _25610_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(_06381_),
    .S(net81),
    .X(_02425_));
 sg13g2_mux2_1 _25611_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(_10099_),
    .S(net81),
    .X(_02426_));
 sg13g2_mux2_1 _25612_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(_10105_),
    .S(net81),
    .X(_02427_));
 sg13g2_mux2_1 _25613_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(_10113_),
    .S(net81),
    .X(_02428_));
 sg13g2_mux2_1 _25614_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(_10119_),
    .S(net81),
    .X(_02429_));
 sg13g2_mux2_1 _25615_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(_10125_),
    .S(net81),
    .X(_02430_));
 sg13g2_mux2_1 _25616_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(_10130_),
    .S(_06725_),
    .X(_02431_));
 sg13g2_nor3_1 _25617_ (.A(_09168_),
    .B(net692),
    .C(_04827_),
    .Y(_06726_));
 sg13g2_buf_2 _25618_ (.A(_06726_),
    .X(_06727_));
 sg13g2_buf_1 _25619_ (.A(_06727_),
    .X(_06728_));
 sg13g2_mux2_1 _25620_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(net837),
    .S(net127),
    .X(_02432_));
 sg13g2_mux2_1 _25621_ (.A0(\cpu.intr.r_clock_cmp[17] ),
    .A1(net900),
    .S(net127),
    .X(_02433_));
 sg13g2_mux2_1 _25622_ (.A0(\cpu.intr.r_clock_cmp[18] ),
    .A1(net836),
    .S(net127),
    .X(_02434_));
 sg13g2_mux2_1 _25623_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(net1039),
    .S(net127),
    .X(_02435_));
 sg13g2_mux2_1 _25624_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(_09997_),
    .S(net81),
    .X(_02436_));
 sg13g2_mux2_1 _25625_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(_12011_),
    .S(_06728_),
    .X(_02437_));
 sg13g2_mux2_1 _25626_ (.A0(\cpu.intr.r_clock_cmp[21] ),
    .A1(_12015_),
    .S(_06728_),
    .X(_02438_));
 sg13g2_mux2_1 _25627_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(net1038),
    .S(net127),
    .X(_02439_));
 sg13g2_mux2_1 _25628_ (.A0(\cpu.intr.r_clock_cmp[23] ),
    .A1(net1041),
    .S(net127),
    .X(_02440_));
 sg13g2_mux2_1 _25629_ (.A0(\cpu.intr.r_clock_cmp[24] ),
    .A1(_10087_),
    .S(net127),
    .X(_02441_));
 sg13g2_mux2_1 _25630_ (.A0(\cpu.intr.r_clock_cmp[25] ),
    .A1(_10094_),
    .S(net127),
    .X(_02442_));
 sg13g2_mux2_1 _25631_ (.A0(\cpu.intr.r_clock_cmp[26] ),
    .A1(_10099_),
    .S(_06727_),
    .X(_02443_));
 sg13g2_mux2_1 _25632_ (.A0(\cpu.intr.r_clock_cmp[27] ),
    .A1(_10105_),
    .S(_06727_),
    .X(_02444_));
 sg13g2_mux2_1 _25633_ (.A0(\cpu.intr.r_clock_cmp[28] ),
    .A1(_10113_),
    .S(_06727_),
    .X(_02445_));
 sg13g2_mux2_1 _25634_ (.A0(\cpu.intr.r_clock_cmp[29] ),
    .A1(_10119_),
    .S(_06727_),
    .X(_02446_));
 sg13g2_mux2_1 _25635_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(_06385_),
    .S(net81),
    .X(_02447_));
 sg13g2_mux2_1 _25636_ (.A0(\cpu.intr.r_clock_cmp[30] ),
    .A1(_10125_),
    .S(_06727_),
    .X(_02448_));
 sg13g2_mux2_1 _25637_ (.A0(\cpu.intr.r_clock_cmp[31] ),
    .A1(_10130_),
    .S(_06727_),
    .X(_02449_));
 sg13g2_mux2_1 _25638_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(net1039),
    .S(_06725_),
    .X(_02450_));
 sg13g2_mux2_1 _25639_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(_12011_),
    .S(_06724_),
    .X(_02451_));
 sg13g2_mux2_1 _25640_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(_12015_),
    .S(_06724_),
    .X(_02452_));
 sg13g2_mux2_1 _25641_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(net1038),
    .S(_06724_),
    .X(_02453_));
 sg13g2_mux2_1 _25642_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(_10034_),
    .S(_06724_),
    .X(_02454_));
 sg13g2_mux2_1 _25643_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(_10087_),
    .S(_06724_),
    .X(_02455_));
 sg13g2_mux2_1 _25644_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(_10094_),
    .S(_06724_),
    .X(_02456_));
 sg13g2_and2_1 _25645_ (.A(net128),
    .B(_04974_),
    .X(_06729_));
 sg13g2_buf_2 _25646_ (.A(_06729_),
    .X(_06730_));
 sg13g2_buf_1 _25647_ (.A(_06730_),
    .X(_06731_));
 sg13g2_mux2_1 _25648_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net837),
    .S(_06731_),
    .X(_02480_));
 sg13g2_mux2_1 _25649_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10099_),
    .S(net80),
    .X(_02481_));
 sg13g2_mux2_1 _25650_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10105_),
    .S(net80),
    .X(_02482_));
 sg13g2_mux2_1 _25651_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10113_),
    .S(net80),
    .X(_02483_));
 sg13g2_mux2_1 _25652_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10119_),
    .S(net80),
    .X(_02484_));
 sg13g2_mux2_1 _25653_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10125_),
    .S(net80),
    .X(_02485_));
 sg13g2_mux2_1 _25654_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10130_),
    .S(net80),
    .X(_02486_));
 sg13g2_o21ai_1 _25655_ (.B1(_09990_),
    .Y(_02487_),
    .A1(_09983_),
    .A2(net144));
 sg13g2_nand2_1 _25656_ (.Y(_06732_),
    .A(net1040),
    .B(net143));
 sg13g2_o21ai_1 _25657_ (.B1(_06732_),
    .Y(_02488_),
    .A1(_09991_),
    .A2(net144));
 sg13g2_o21ai_1 _25658_ (.B1(_10003_),
    .Y(_02489_),
    .A1(_05363_),
    .A2(net144));
 sg13g2_inv_1 _25659_ (.Y(_06733_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25660_ (.B1(_10009_),
    .Y(_02490_),
    .A1(_06733_),
    .A2(net144));
 sg13g2_mux2_1 _25661_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(_09997_),
    .S(net80),
    .X(_02491_));
 sg13g2_o21ai_1 _25662_ (.B1(_10015_),
    .Y(_02492_),
    .A1(_05478_),
    .A2(_09980_));
 sg13g2_inv_1 _25663_ (.Y(_06734_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25664_ (.B1(_10021_),
    .Y(_02493_),
    .A1(_06734_),
    .A2(net144));
 sg13g2_inv_1 _25665_ (.Y(_06735_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25666_ (.B1(_10028_),
    .Y(_02494_),
    .A1(_06735_),
    .A2(net144));
 sg13g2_mux2_1 _25667_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net1041),
    .S(net143),
    .X(_02495_));
 sg13g2_mux2_1 _25668_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(net836),
    .S(net80),
    .X(_02496_));
 sg13g2_mux2_1 _25669_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(_10062_),
    .S(_06731_),
    .X(_02497_));
 sg13g2_mux2_1 _25670_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(net1006),
    .S(_06730_),
    .X(_02498_));
 sg13g2_mux2_1 _25671_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(net1005),
    .S(_06730_),
    .X(_02499_));
 sg13g2_mux2_1 _25672_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net1038),
    .S(_06730_),
    .X(_02500_));
 sg13g2_mux2_1 _25673_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(net1041),
    .S(_06730_),
    .X(_02501_));
 sg13g2_mux2_1 _25674_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10087_),
    .S(_06730_),
    .X(_02502_));
 sg13g2_mux2_1 _25675_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10094_),
    .S(_06730_),
    .X(_02503_));
 sg13g2_o21ai_1 _25676_ (.B1(\cpu.qspi.r_state[17] ),
    .Y(_06736_),
    .A1(_09776_),
    .A2(_11783_));
 sg13g2_nor2_1 _25677_ (.A(_09788_),
    .B(_09778_),
    .Y(_06737_));
 sg13g2_nor4_1 _25678_ (.A(_11800_),
    .B(_09798_),
    .C(_11780_),
    .D(_11775_),
    .Y(_06738_));
 sg13g2_nor2b_1 _25679_ (.A(_11798_),
    .B_N(_06738_),
    .Y(_06739_));
 sg13g2_nor2_1 _25680_ (.A(_11778_),
    .B(\cpu.qspi.r_state[11] ),
    .Y(_06740_));
 sg13g2_and4_1 _25681_ (.A(_06736_),
    .B(_06737_),
    .C(_06739_),
    .D(_06740_),
    .X(_06741_));
 sg13g2_buf_1 _25682_ (.A(_06741_),
    .X(_06742_));
 sg13g2_mux2_1 _25683_ (.A0(\cpu.qspi.r_read_delay[0][0] ),
    .A1(\cpu.qspi.r_read_delay[1][0] ),
    .S(_09814_),
    .X(_06743_));
 sg13g2_mux2_1 _25684_ (.A0(_06743_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .S(_09808_),
    .X(_06744_));
 sg13g2_or4_1 _25685_ (.A(_09787_),
    .B(_09797_),
    .C(net1122),
    .D(_09790_),
    .X(_06745_));
 sg13g2_buf_1 _25686_ (.A(_06745_),
    .X(_06746_));
 sg13g2_inv_1 _25687_ (.Y(_06747_),
    .A(_09780_));
 sg13g2_a21o_1 _25688_ (.A2(_06747_),
    .A1(_09827_),
    .B1(_09795_),
    .X(_06748_));
 sg13g2_a221oi_1 _25689_ (.B2(_00168_),
    .C1(_06748_),
    .B1(_06746_),
    .A1(_09842_),
    .Y(_06749_),
    .A2(_06744_));
 sg13g2_nor2_1 _25690_ (.A(_09780_),
    .B(net29),
    .Y(_06750_));
 sg13g2_a21oi_1 _25691_ (.A1(net29),
    .A2(_06749_),
    .Y(_02504_),
    .B1(_06750_));
 sg13g2_mux2_1 _25692_ (.A0(\cpu.qspi.r_read_delay[0][1] ),
    .A1(\cpu.qspi.r_read_delay[1][1] ),
    .S(_09814_),
    .X(_06751_));
 sg13g2_mux2_1 _25693_ (.A0(_06751_),
    .A1(\cpu.qspi.r_read_delay[2][1] ),
    .S(_09808_),
    .X(_06752_));
 sg13g2_nor2_1 _25694_ (.A(_09827_),
    .B(_06746_),
    .Y(_06753_));
 sg13g2_nand2_1 _25695_ (.Y(_06754_),
    .A(_09842_),
    .B(_06753_));
 sg13g2_nand2_1 _25696_ (.Y(_06755_),
    .A(_06747_),
    .B(_09781_));
 sg13g2_nand2b_1 _25697_ (.Y(_06756_),
    .B(_09780_),
    .A_N(_09781_));
 sg13g2_a21o_1 _25698_ (.A2(_06756_),
    .A1(_06755_),
    .B1(_06753_),
    .X(_06757_));
 sg13g2_a221oi_1 _25699_ (.B2(_06757_),
    .C1(_09795_),
    .B1(_06754_),
    .A1(_09842_),
    .Y(_06758_),
    .A2(_06752_));
 sg13g2_nor2_1 _25700_ (.A(_09781_),
    .B(net29),
    .Y(_06759_));
 sg13g2_a21oi_1 _25701_ (.A1(net29),
    .A2(_06758_),
    .Y(_02505_),
    .B1(_06759_));
 sg13g2_mux2_1 _25702_ (.A0(\cpu.qspi.r_read_delay[0][2] ),
    .A1(\cpu.qspi.r_read_delay[1][2] ),
    .S(_09814_),
    .X(_06760_));
 sg13g2_mux2_1 _25703_ (.A0(_06760_),
    .A1(\cpu.qspi.r_read_delay[2][2] ),
    .S(_09808_),
    .X(_06761_));
 sg13g2_nor2_1 _25704_ (.A(_09780_),
    .B(_09781_),
    .Y(_06762_));
 sg13g2_xor2_1 _25705_ (.B(_06762_),
    .A(_00167_),
    .X(_06763_));
 sg13g2_mux2_1 _25706_ (.A0(_06746_),
    .A1(_09792_),
    .S(_09827_),
    .X(_06764_));
 sg13g2_nand2_1 _25707_ (.Y(_06765_),
    .A(_06763_),
    .B(_06764_));
 sg13g2_a221oi_1 _25708_ (.B2(_06754_),
    .C1(_09795_),
    .B1(_06765_),
    .A1(_09842_),
    .Y(_06766_),
    .A2(_06761_));
 sg13g2_nor2_1 _25709_ (.A(\cpu.qspi.r_count[2] ),
    .B(net29),
    .Y(_06767_));
 sg13g2_a21oi_1 _25710_ (.A1(_06742_),
    .A2(_06766_),
    .Y(_02506_),
    .B1(_06767_));
 sg13g2_a21oi_1 _25711_ (.A1(_09827_),
    .A2(_09791_),
    .Y(_06768_),
    .B1(_06746_));
 sg13g2_o21ai_1 _25712_ (.B1(net29),
    .Y(_06769_),
    .A1(_09782_),
    .A2(_06768_));
 sg13g2_inv_1 _25713_ (.Y(_06770_),
    .A(_06768_));
 sg13g2_mux2_1 _25714_ (.A0(\cpu.qspi.r_read_delay[0][3] ),
    .A1(\cpu.qspi.r_read_delay[1][3] ),
    .S(_09814_),
    .X(_06771_));
 sg13g2_mux2_1 _25715_ (.A0(_06771_),
    .A1(\cpu.qspi.r_read_delay[2][3] ),
    .S(_09808_),
    .X(_06772_));
 sg13g2_a22oi_1 _25716_ (.Y(_06773_),
    .B1(_06772_),
    .B2(_09842_),
    .A2(_06770_),
    .A1(_09784_));
 sg13g2_inv_1 _25717_ (.Y(_06774_),
    .A(_06773_));
 sg13g2_a22oi_1 _25718_ (.Y(_06775_),
    .B1(_06774_),
    .B2(net29),
    .A2(_06769_),
    .A1(\cpu.qspi.r_count[3] ));
 sg13g2_inv_1 _25719_ (.Y(_02507_),
    .A(_06775_));
 sg13g2_or2_1 _25720_ (.X(_06776_),
    .B(_09784_),
    .A(_00232_));
 sg13g2_a21oi_1 _25721_ (.A1(_09792_),
    .A2(_06776_),
    .Y(_06777_),
    .B1(_06768_));
 sg13g2_mux2_1 _25722_ (.A0(\cpu.qspi.r_count[4] ),
    .A1(_06777_),
    .S(net29),
    .X(_02508_));
 sg13g2_nand2_1 _25723_ (.Y(_06778_),
    .A(_09908_),
    .B(_06367_));
 sg13g2_buf_2 _25724_ (.A(_06778_),
    .X(_06779_));
 sg13g2_nor3_1 _25725_ (.A(net506),
    .B(net609),
    .C(_06779_),
    .Y(_06780_));
 sg13g2_buf_1 _25726_ (.A(_06780_),
    .X(_06781_));
 sg13g2_nand2_1 _25727_ (.Y(_06782_),
    .A(net865),
    .B(_06781_));
 sg13g2_nand3_1 _25728_ (.B(_09908_),
    .C(_06367_),
    .A(_09144_),
    .Y(_06783_));
 sg13g2_buf_1 _25729_ (.A(_06783_),
    .X(_06784_));
 sg13g2_nand2_1 _25730_ (.Y(_06785_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06784_));
 sg13g2_a21oi_1 _25731_ (.A1(_06782_),
    .A2(_06785_),
    .Y(_02519_),
    .B1(net712));
 sg13g2_nand2_1 _25732_ (.Y(_06786_),
    .A(net1040),
    .B(_06781_));
 sg13g2_nand2_1 _25733_ (.Y(_06787_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06784_));
 sg13g2_a21oi_1 _25734_ (.A1(_06786_),
    .A2(_06787_),
    .Y(_02520_),
    .B1(net712));
 sg13g2_nand2_1 _25735_ (.Y(_06788_),
    .A(net898),
    .B(_06781_));
 sg13g2_nand2_1 _25736_ (.Y(_06789_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06784_));
 sg13g2_nand3_1 _25737_ (.B(_06788_),
    .C(_06789_),
    .A(net694),
    .Y(_02521_));
 sg13g2_nand2_1 _25738_ (.Y(_06790_),
    .A(net1039),
    .B(_06781_));
 sg13g2_nand2_1 _25739_ (.Y(_06791_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06784_));
 sg13g2_a21oi_1 _25740_ (.A1(_06790_),
    .A2(_06791_),
    .Y(_02522_),
    .B1(net712));
 sg13g2_nor2_1 _25741_ (.A(net595),
    .B(_06779_),
    .Y(_06792_));
 sg13g2_nand2_1 _25742_ (.Y(_06793_),
    .A(net865),
    .B(_06792_));
 sg13g2_nand3_1 _25743_ (.B(_04854_),
    .C(_06367_),
    .A(_09908_),
    .Y(_06794_));
 sg13g2_buf_1 _25744_ (.A(_06794_),
    .X(_06795_));
 sg13g2_nand2_1 _25745_ (.Y(_06796_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06795_));
 sg13g2_a21oi_1 _25746_ (.A1(_06793_),
    .A2(_06796_),
    .Y(_02523_),
    .B1(_09233_));
 sg13g2_nand2_1 _25747_ (.Y(_06797_),
    .A(net1040),
    .B(_06792_));
 sg13g2_nand2_1 _25748_ (.Y(_06798_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06795_));
 sg13g2_buf_2 _25749_ (.A(net916),
    .X(_06799_));
 sg13g2_buf_1 _25750_ (.A(_06799_),
    .X(_06800_));
 sg13g2_a21oi_1 _25751_ (.A1(_06797_),
    .A2(_06798_),
    .Y(_02524_),
    .B1(net657));
 sg13g2_nand2_1 _25752_ (.Y(_06801_),
    .A(_10057_),
    .B(_06792_));
 sg13g2_nand2_1 _25753_ (.Y(_06802_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06795_));
 sg13g2_nand3_1 _25754_ (.B(_06801_),
    .C(_06802_),
    .A(net694),
    .Y(_02525_));
 sg13g2_nand2_1 _25755_ (.Y(_06803_),
    .A(net1044),
    .B(_06792_));
 sg13g2_nand2_1 _25756_ (.Y(_06804_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06795_));
 sg13g2_a21oi_1 _25757_ (.A1(_06803_),
    .A2(_06804_),
    .Y(_02526_),
    .B1(net657));
 sg13g2_nor2_1 _25758_ (.A(net534),
    .B(_06779_),
    .Y(_06805_));
 sg13g2_buf_1 _25759_ (.A(_06805_),
    .X(_06806_));
 sg13g2_nand2_1 _25760_ (.Y(_06807_),
    .A(_02804_),
    .B(_06806_));
 sg13g2_or2_1 _25761_ (.X(_06808_),
    .B(_06779_),
    .A(net534));
 sg13g2_buf_1 _25762_ (.A(_06808_),
    .X(_06809_));
 sg13g2_nand2_1 _25763_ (.Y(_06810_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06809_));
 sg13g2_a21oi_1 _25764_ (.A1(_06807_),
    .A2(_06810_),
    .Y(_02527_),
    .B1(net657));
 sg13g2_nand2_1 _25765_ (.Y(_06811_),
    .A(_10051_),
    .B(_06806_));
 sg13g2_nand2_1 _25766_ (.Y(_06812_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06809_));
 sg13g2_a21oi_1 _25767_ (.A1(_06811_),
    .A2(_06812_),
    .Y(_02528_),
    .B1(net657));
 sg13g2_nand2_1 _25768_ (.Y(_06813_),
    .A(net898),
    .B(_06806_));
 sg13g2_nand2_1 _25769_ (.Y(_06814_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06809_));
 sg13g2_nand3_1 _25770_ (.B(_06813_),
    .C(_06814_),
    .A(net715),
    .Y(_02529_));
 sg13g2_nand2_1 _25771_ (.Y(_06815_),
    .A(net1044),
    .B(_06806_));
 sg13g2_nand2_1 _25772_ (.Y(_06816_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06809_));
 sg13g2_a21oi_1 _25773_ (.A1(_06815_),
    .A2(_06816_),
    .Y(_02530_),
    .B1(net657));
 sg13g2_buf_1 _25774_ (.A(net1137),
    .X(_06817_));
 sg13g2_buf_1 _25775_ (.A(_06817_),
    .X(_06818_));
 sg13g2_nand2b_1 _25776_ (.Y(_06819_),
    .B(_09765_),
    .A_N(_09768_));
 sg13g2_buf_1 _25777_ (.A(_06819_),
    .X(_06820_));
 sg13g2_buf_1 _25778_ (.A(_06820_),
    .X(_06821_));
 sg13g2_mux2_1 _25779_ (.A0(_00215_),
    .A1(_09709_),
    .S(net92),
    .X(_06822_));
 sg13g2_nand2b_1 _25780_ (.Y(_06823_),
    .B(net941),
    .A_N(_10427_));
 sg13g2_o21ai_1 _25781_ (.B1(_06823_),
    .Y(_06824_),
    .A1(net830),
    .A2(_06822_));
 sg13g2_buf_1 _25782_ (.A(_08284_),
    .X(_06825_));
 sg13g2_mux2_1 _25783_ (.A0(_09661_),
    .A1(_09667_),
    .S(net92),
    .X(_06826_));
 sg13g2_nand2_1 _25784_ (.Y(_06827_),
    .A(net829),
    .B(_06826_));
 sg13g2_o21ai_1 _25785_ (.B1(_06827_),
    .Y(_06828_),
    .A1(net829),
    .A2(_08728_));
 sg13g2_a22oi_1 _25786_ (.Y(_06829_),
    .B1(_06828_),
    .B2(_11800_),
    .A2(_06824_),
    .A1(_11798_));
 sg13g2_nand3_1 _25787_ (.B(_09780_),
    .C(_09779_),
    .A(net1122),
    .Y(_06830_));
 sg13g2_o21ai_1 _25788_ (.B1(_06830_),
    .Y(_06831_),
    .A1(_09779_),
    .A2(_06755_));
 sg13g2_nand2b_1 _25789_ (.Y(_06832_),
    .B(_09794_),
    .A_N(_09781_));
 sg13g2_a21oi_1 _25790_ (.A1(_06755_),
    .A2(_06832_),
    .Y(_06833_),
    .B1(net1122));
 sg13g2_inv_1 _25791_ (.Y(_06834_),
    .A(\cpu.qspi.r_count[2] ));
 sg13g2_o21ai_1 _25792_ (.B1(_06834_),
    .Y(_06835_),
    .A1(_06831_),
    .A2(_06833_));
 sg13g2_nand2_1 _25793_ (.Y(_06836_),
    .A(net1122),
    .B(_09779_));
 sg13g2_a21oi_1 _25794_ (.A1(_00168_),
    .A2(_06836_),
    .Y(_06837_),
    .B1(_09781_));
 sg13g2_nor2_1 _25795_ (.A(_06834_),
    .B(_06837_),
    .Y(_06838_));
 sg13g2_mux2_1 _25796_ (.A0(_06755_),
    .A1(_09781_),
    .S(_09794_),
    .X(_06839_));
 sg13g2_nand2_1 _25797_ (.Y(_06840_),
    .A(net1122),
    .B(_06838_));
 sg13g2_o21ai_1 _25798_ (.B1(_06840_),
    .Y(_06841_),
    .A1(_09797_),
    .A2(_09801_));
 sg13g2_a21oi_1 _25799_ (.A1(_06838_),
    .A2(_06839_),
    .Y(_06842_),
    .B1(_06841_));
 sg13g2_buf_1 _25800_ (.A(_08284_),
    .X(_06843_));
 sg13g2_buf_1 _25801_ (.A(_06820_),
    .X(_06844_));
 sg13g2_mux2_1 _25802_ (.A0(_09590_),
    .A1(_09574_),
    .S(net91),
    .X(_06845_));
 sg13g2_nand2_1 _25803_ (.Y(_06846_),
    .A(net828),
    .B(_06845_));
 sg13g2_o21ai_1 _25804_ (.B1(_06846_),
    .Y(_06847_),
    .A1(net829),
    .A2(_08439_));
 sg13g2_inv_1 _25805_ (.Y(_06848_),
    .A(_09794_));
 sg13g2_nor4_1 _25806_ (.A(_09797_),
    .B(_09795_),
    .C(net1122),
    .D(_09790_),
    .Y(_06849_));
 sg13g2_and3_1 _25807_ (.X(_06850_),
    .A(_06739_),
    .B(_06740_),
    .C(_06849_));
 sg13g2_and2_1 _25808_ (.A(_09800_),
    .B(_06850_),
    .X(_06851_));
 sg13g2_buf_1 _25809_ (.A(_06851_),
    .X(_06852_));
 sg13g2_or2_1 _25810_ (.X(_06853_),
    .B(_06852_),
    .A(_11778_));
 sg13g2_buf_1 _25811_ (.A(_06853_),
    .X(_06854_));
 sg13g2_a21oi_1 _25812_ (.A1(_09798_),
    .A2(_06848_),
    .Y(_06855_),
    .B1(_06854_));
 sg13g2_inv_1 _25813_ (.Y(_06856_),
    .A(_09779_));
 sg13g2_nand2_1 _25814_ (.Y(_06857_),
    .A(_08442_),
    .B(net1137));
 sg13g2_o21ai_1 _25815_ (.B1(_06857_),
    .Y(_06858_),
    .A1(net1137),
    .A2(_11839_));
 sg13g2_a22oi_1 _25816_ (.Y(_06859_),
    .B1(_06858_),
    .B2(_11775_),
    .A2(\cpu.qspi.r_state[0] ),
    .A1(_06856_));
 sg13g2_inv_1 _25817_ (.Y(_06860_),
    .A(_04786_));
 sg13g2_a22oi_1 _25818_ (.Y(_06861_),
    .B1(_06860_),
    .B2(net1100),
    .A2(_04793_),
    .A1(net1014));
 sg13g2_a221oi_1 _25819_ (.B2(net1014),
    .C1(net1009),
    .B1(_05147_),
    .A1(net1100),
    .Y(_06862_),
    .A2(_05141_));
 sg13g2_a21oi_1 _25820_ (.A1(net1009),
    .A2(_06861_),
    .Y(_06863_),
    .B1(_06862_));
 sg13g2_inv_1 _25821_ (.Y(_06864_),
    .A(_11908_));
 sg13g2_nor2_1 _25822_ (.A(_11885_),
    .B(_06864_),
    .Y(_06865_));
 sg13g2_buf_1 _25823_ (.A(_06865_),
    .X(_06866_));
 sg13g2_inv_1 _25824_ (.Y(_06867_),
    .A(net1100));
 sg13g2_nor2_1 _25825_ (.A(_11884_),
    .B(_06867_),
    .Y(_06868_));
 sg13g2_a22oi_1 _25826_ (.Y(_06869_),
    .B1(_06868_),
    .B2(_05465_),
    .A2(_06866_),
    .A1(_04763_));
 sg13g2_nor2_1 _25827_ (.A(_06864_),
    .B(_12004_),
    .Y(_06870_));
 sg13g2_nor2_1 _25828_ (.A(net1100),
    .B(_06870_),
    .Y(_06871_));
 sg13g2_and2_1 _25829_ (.A(net1100),
    .B(_11911_),
    .X(_06872_));
 sg13g2_a22oi_1 _25830_ (.Y(_06873_),
    .B1(_06872_),
    .B2(_04772_),
    .A2(_06871_),
    .A1(_05458_));
 sg13g2_o21ai_1 _25831_ (.B1(_06873_),
    .Y(_06874_),
    .A1(net1013),
    .A2(_06869_));
 sg13g2_a21oi_1 _25832_ (.A1(net1013),
    .A2(_06863_),
    .Y(_06875_),
    .B1(_06874_));
 sg13g2_nand2b_1 _25833_ (.Y(_06876_),
    .B(_09790_),
    .A_N(_06875_));
 sg13g2_nand3_1 _25834_ (.B(_06859_),
    .C(_06876_),
    .A(_06855_),
    .Y(_06877_));
 sg13g2_a221oi_1 _25835_ (.B2(_11780_),
    .C1(_06877_),
    .B1(_06847_),
    .A1(_06835_),
    .Y(_06878_),
    .A2(_06842_));
 sg13g2_xnor2_1 _25836_ (.Y(_06879_),
    .A(_06848_),
    .B(_11783_));
 sg13g2_a22oi_1 _25837_ (.Y(_06880_),
    .B1(_06879_),
    .B2(_06852_),
    .A2(_06878_),
    .A1(_06829_));
 sg13g2_inv_1 _25838_ (.Y(_06881_),
    .A(\cpu.qspi.r_mask[0] ));
 sg13g2_a22oi_1 _25839_ (.Y(_06882_),
    .B1(_09814_),
    .B2(\cpu.qspi.r_mask[1] ),
    .A2(_09808_),
    .A1(\cpu.qspi.r_mask[2] ));
 sg13g2_o21ai_1 _25840_ (.B1(_06882_),
    .Y(_06883_),
    .A1(_06881_),
    .A2(_09818_));
 sg13g2_or2_1 _25841_ (.X(_06884_),
    .B(_06883_),
    .A(_11779_));
 sg13g2_nor3_2 _25842_ (.A(_09787_),
    .B(_09788_),
    .C(_09778_),
    .Y(_06885_));
 sg13g2_nor2_1 _25843_ (.A(_09842_),
    .B(_09827_),
    .Y(_06886_));
 sg13g2_and4_1 _25844_ (.A(_09777_),
    .B(_06884_),
    .C(_06885_),
    .D(_06886_),
    .X(_06887_));
 sg13g2_buf_1 _25845_ (.A(_06887_),
    .X(_06888_));
 sg13g2_mux2_1 _25846_ (.A0(net12),
    .A1(_06880_),
    .S(_06888_),
    .X(_02535_));
 sg13g2_nand2_1 _25847_ (.Y(_06889_),
    .A(_09676_),
    .B(_09679_));
 sg13g2_nor2_1 _25848_ (.A(_00217_),
    .B(_06821_),
    .Y(_06890_));
 sg13g2_a21oi_1 _25849_ (.A1(_06889_),
    .A2(_06821_),
    .Y(_06891_),
    .B1(_06890_));
 sg13g2_nand2_1 _25850_ (.Y(_06892_),
    .A(net830),
    .B(_11011_));
 sg13g2_o21ai_1 _25851_ (.B1(_06892_),
    .Y(_06893_),
    .A1(net830),
    .A2(_06891_));
 sg13g2_nand2_1 _25852_ (.Y(_06894_),
    .A(_06867_),
    .B(net1014));
 sg13g2_mux2_1 _25853_ (.A0(_05242_),
    .A1(_05574_),
    .S(_11885_),
    .X(_06895_));
 sg13g2_nand2_1 _25854_ (.Y(_06896_),
    .A(_11883_),
    .B(_06895_));
 sg13g2_nand2b_1 _25855_ (.Y(_06897_),
    .B(_11887_),
    .A_N(_05250_));
 sg13g2_nand3_1 _25856_ (.B(_06896_),
    .C(_06897_),
    .A(net1100),
    .Y(_06898_));
 sg13g2_a22oi_1 _25857_ (.Y(_06899_),
    .B1(_05172_),
    .B2(_11909_),
    .A2(_05166_),
    .A1(net1007));
 sg13g2_nand2b_1 _25858_ (.Y(_06900_),
    .B(_06866_),
    .A_N(_05257_));
 sg13g2_o21ai_1 _25859_ (.B1(_06900_),
    .Y(_06901_),
    .A1(net1009),
    .A2(_06899_));
 sg13g2_a22oi_1 _25860_ (.Y(_06902_),
    .B1(_06898_),
    .B2(_11885_),
    .A2(_06866_),
    .A1(_05234_));
 sg13g2_nor2_1 _25861_ (.A(net1013),
    .B(_06902_),
    .Y(_06903_));
 sg13g2_a221oi_1 _25862_ (.B2(net1013),
    .C1(_06903_),
    .B1(_06901_),
    .A1(_06894_),
    .Y(_06904_),
    .A2(_06898_));
 sg13g2_inv_1 _25863_ (.Y(_06905_),
    .A(_06871_));
 sg13g2_o21ai_1 _25864_ (.B1(_09790_),
    .Y(_06906_),
    .A1(_05568_),
    .A2(_06905_));
 sg13g2_o21ai_1 _25865_ (.B1(_06855_),
    .Y(_06907_),
    .A1(_06904_),
    .A2(_06906_));
 sg13g2_a21oi_1 _25866_ (.A1(_11798_),
    .A2(_06893_),
    .Y(_06908_),
    .B1(_06907_));
 sg13g2_mux2_1 _25867_ (.A0(_09566_),
    .A1(_09550_),
    .S(net91),
    .X(_06909_));
 sg13g2_nand2_1 _25868_ (.Y(_06910_),
    .A(net828),
    .B(_06909_));
 sg13g2_o21ai_1 _25869_ (.B1(_06910_),
    .Y(_06911_),
    .A1(net829),
    .A2(_08507_));
 sg13g2_nor2_1 _25870_ (.A(_09359_),
    .B(_09383_),
    .Y(_06912_));
 sg13g2_mux2_1 _25871_ (.A0(net449),
    .A1(_06912_),
    .S(net91),
    .X(_06913_));
 sg13g2_nand2_1 _25872_ (.Y(_06914_),
    .A(net828),
    .B(_06913_));
 sg13g2_o21ai_1 _25873_ (.B1(_06914_),
    .Y(_06915_),
    .A1(net829),
    .A2(_08798_));
 sg13g2_nand2_1 _25874_ (.Y(_06916_),
    .A(_09751_),
    .B(_06844_));
 sg13g2_o21ai_1 _25875_ (.B1(_06916_),
    .Y(_06917_),
    .A1(_09741_),
    .A2(net92));
 sg13g2_nand2b_1 _25876_ (.Y(_06918_),
    .B(net1137),
    .A_N(_10629_));
 sg13g2_o21ai_1 _25877_ (.B1(_06918_),
    .Y(_06919_),
    .A1(net941),
    .A2(_06917_));
 sg13g2_and2_1 _25878_ (.A(_11775_),
    .B(_06919_),
    .X(_06920_));
 sg13g2_a221oi_1 _25879_ (.B2(_11800_),
    .C1(_06920_),
    .B1(_06915_),
    .A1(_11780_),
    .Y(_06921_),
    .A2(_06911_));
 sg13g2_a22oi_1 _25880_ (.Y(_06922_),
    .B1(_06908_),
    .B2(_06921_),
    .A2(_06852_),
    .A1(_09821_));
 sg13g2_mux2_1 _25881_ (.A0(net13),
    .A1(_06922_),
    .S(_06888_),
    .X(_02536_));
 sg13g2_nand2_1 _25882_ (.Y(_06923_),
    .A(net724),
    .B(net830));
 sg13g2_nand2_1 _25883_ (.Y(_06924_),
    .A(net829),
    .B(net506));
 sg13g2_a21oi_1 _25884_ (.A1(_06923_),
    .A2(_06924_),
    .Y(_06925_),
    .B1(_00169_));
 sg13g2_a22oi_1 _25885_ (.Y(_06926_),
    .B1(_05199_),
    .B2(net1014),
    .A2(_05192_),
    .A1(net1007));
 sg13g2_nand2_1 _25886_ (.Y(_06927_),
    .A(_04999_),
    .B(_06866_));
 sg13g2_o21ai_1 _25887_ (.B1(_06927_),
    .Y(_06928_),
    .A1(net1009),
    .A2(_06926_));
 sg13g2_nand2b_1 _25888_ (.Y(_06929_),
    .B(net1007),
    .A_N(_05329_));
 sg13g2_a221oi_1 _25889_ (.B2(net1009),
    .C1(net1013),
    .B1(_06929_),
    .A1(_05598_),
    .Y(_06930_),
    .A2(_06868_));
 sg13g2_a21oi_1 _25890_ (.A1(_11910_),
    .A2(_06928_),
    .Y(_06931_),
    .B1(_06930_));
 sg13g2_nand2_1 _25891_ (.Y(_06932_),
    .A(_11883_),
    .B(_11909_));
 sg13g2_nand3_1 _25892_ (.B(net1007),
    .C(_04991_),
    .A(_11910_),
    .Y(_06933_));
 sg13g2_o21ai_1 _25893_ (.B1(_06933_),
    .Y(_06934_),
    .A1(_05321_),
    .A2(_06932_));
 sg13g2_a22oi_1 _25894_ (.Y(_06935_),
    .B1(_06934_),
    .B2(_11947_),
    .A2(_06864_),
    .A1(_06867_));
 sg13g2_a221oi_1 _25895_ (.B2(_06935_),
    .C1(_11781_),
    .B1(_06931_),
    .A1(_05605_),
    .Y(_06936_),
    .A2(_06871_));
 sg13g2_mux2_1 _25896_ (.A0(_00219_),
    .A1(_09691_),
    .S(net91),
    .X(_06937_));
 sg13g2_nand2b_1 _25897_ (.Y(_06938_),
    .B(net941),
    .A_N(_10365_));
 sg13g2_o21ai_1 _25898_ (.B1(_06938_),
    .Y(_06939_),
    .A1(net941),
    .A2(_06937_));
 sg13g2_mux2_1 _25899_ (.A0(_09532_),
    .A1(_09540_),
    .S(net91),
    .X(_06940_));
 sg13g2_nand2_1 _25900_ (.Y(_06941_),
    .A(net828),
    .B(_06940_));
 sg13g2_o21ai_1 _25901_ (.B1(_06941_),
    .Y(_06942_),
    .A1(net828),
    .A2(_08547_));
 sg13g2_a22oi_1 _25902_ (.Y(_06943_),
    .B1(_06942_),
    .B2(_11800_),
    .A2(_06939_),
    .A1(_11798_));
 sg13g2_mux2_1 _25903_ (.A0(net355),
    .A1(_09516_),
    .S(_06820_),
    .X(_06944_));
 sg13g2_nand2_1 _25904_ (.Y(_06945_),
    .A(net828),
    .B(_06944_));
 sg13g2_o21ai_1 _25905_ (.B1(_06945_),
    .Y(_06946_),
    .A1(_06843_),
    .A2(_08776_));
 sg13g2_nand3b_1 _25906_ (.B(_09720_),
    .C(net91),
    .Y(_06947_),
    .A_N(_09713_));
 sg13g2_o21ai_1 _25907_ (.B1(_06947_),
    .Y(_06948_),
    .A1(_09723_),
    .A2(net92));
 sg13g2_nand2b_1 _25908_ (.Y(_06949_),
    .B(net941),
    .A_N(_10330_));
 sg13g2_o21ai_1 _25909_ (.B1(_06949_),
    .Y(_06950_),
    .A1(net941),
    .A2(_06948_));
 sg13g2_a22oi_1 _25910_ (.Y(_06951_),
    .B1(_06950_),
    .B2(_11775_),
    .A2(_06946_),
    .A1(_11780_));
 sg13g2_nand2_1 _25911_ (.Y(_06952_),
    .A(_06943_),
    .B(_06951_));
 sg13g2_nor4_1 _25912_ (.A(_06854_),
    .B(_06925_),
    .C(_06936_),
    .D(_06952_),
    .Y(_06953_));
 sg13g2_o21ai_1 _25913_ (.B1(_06852_),
    .Y(_06954_),
    .A1(_09794_),
    .A2(_09821_));
 sg13g2_nand2_1 _25914_ (.Y(_06955_),
    .A(_06888_),
    .B(_06954_));
 sg13g2_nand2b_1 _25915_ (.Y(_06956_),
    .B(net14),
    .A_N(_06888_));
 sg13g2_o21ai_1 _25916_ (.B1(_06956_),
    .Y(_02537_),
    .A1(_06953_),
    .A2(_06955_));
 sg13g2_nand3b_1 _25917_ (.B(_09735_),
    .C(_06844_),
    .Y(_06957_),
    .A_N(_09727_));
 sg13g2_o21ai_1 _25918_ (.B1(_06957_),
    .Y(_06958_),
    .A1(_09738_),
    .A2(net92));
 sg13g2_nand2_1 _25919_ (.Y(_06959_),
    .A(net941),
    .B(_11031_));
 sg13g2_o21ai_1 _25920_ (.B1(_06959_),
    .Y(_06960_),
    .A1(net830),
    .A2(_06958_));
 sg13g2_mux2_1 _25921_ (.A0(net356),
    .A1(_09458_),
    .S(net91),
    .X(_06961_));
 sg13g2_nand2_1 _25922_ (.Y(_06962_),
    .A(_06843_),
    .B(_06961_));
 sg13g2_o21ai_1 _25923_ (.B1(_06962_),
    .Y(_06963_),
    .A1(net829),
    .A2(_08752_));
 sg13g2_a22oi_1 _25924_ (.Y(_06964_),
    .B1(_06963_),
    .B2(_11780_),
    .A2(_06960_),
    .A1(_11798_));
 sg13g2_mux2_1 _25925_ (.A0(_00213_),
    .A1(_09700_),
    .S(net92),
    .X(_06965_));
 sg13g2_nand2b_1 _25926_ (.Y(_06966_),
    .B(net941),
    .A_N(_10457_));
 sg13g2_o21ai_1 _25927_ (.B1(_06966_),
    .Y(_06967_),
    .A1(net830),
    .A2(_06965_));
 sg13g2_mux2_1 _25928_ (.A0(_09804_),
    .A1(_09489_),
    .S(net91),
    .X(_06968_));
 sg13g2_a21oi_1 _25929_ (.A1(net828),
    .A2(_06968_),
    .Y(_06969_),
    .B1(_09805_));
 sg13g2_nor4_1 _25930_ (.A(_09810_),
    .B(_09803_),
    .C(_11777_),
    .D(_06969_),
    .Y(_06970_));
 sg13g2_a21oi_1 _25931_ (.A1(_11775_),
    .A2(_06967_),
    .Y(_06971_),
    .B1(_06970_));
 sg13g2_nand2_1 _25932_ (.Y(_06972_),
    .A(net642),
    .B(_06817_));
 sg13g2_nand2_1 _25933_ (.Y(_06973_),
    .A(net828),
    .B(_09166_));
 sg13g2_a21oi_1 _25934_ (.A1(_06972_),
    .A2(_06973_),
    .Y(_06974_),
    .B1(_00169_));
 sg13g2_mux2_1 _25935_ (.A0(_05055_),
    .A1(_05429_),
    .S(net1009),
    .X(_06975_));
 sg13g2_a21oi_1 _25936_ (.A1(_11887_),
    .A2(_05115_),
    .Y(_06976_),
    .B1(_06867_));
 sg13g2_o21ai_1 _25937_ (.B1(_06976_),
    .Y(_06977_),
    .A1(net1013),
    .A2(_06975_));
 sg13g2_nand2_1 _25938_ (.Y(_06978_),
    .A(_06894_),
    .B(_06977_));
 sg13g2_a22oi_1 _25939_ (.Y(_06979_),
    .B1(_05063_),
    .B2(_11881_),
    .A2(_05082_),
    .A1(_11908_));
 sg13g2_nor2_1 _25940_ (.A(_11947_),
    .B(_06979_),
    .Y(_06980_));
 sg13g2_a21oi_1 _25941_ (.A1(_05123_),
    .A2(_06866_),
    .Y(_06981_),
    .B1(_06980_));
 sg13g2_a21oi_1 _25942_ (.A1(net1007),
    .A2(_05055_),
    .Y(_06982_),
    .B1(net1009));
 sg13g2_a21oi_1 _25943_ (.A1(_05436_),
    .A2(_06866_),
    .Y(_06983_),
    .B1(_06982_));
 sg13g2_mux2_1 _25944_ (.A0(_06981_),
    .A1(_06983_),
    .S(_11883_),
    .X(_06984_));
 sg13g2_a221oi_1 _25945_ (.B2(_06984_),
    .C1(_11781_),
    .B1(_06978_),
    .A1(_05075_),
    .Y(_06985_),
    .A2(_06871_));
 sg13g2_nor4_1 _25946_ (.A(_09798_),
    .B(_06854_),
    .C(_06974_),
    .D(_06985_),
    .Y(_06986_));
 sg13g2_nor2_1 _25947_ (.A(net829),
    .B(_08706_),
    .Y(_06987_));
 sg13g2_nand2_1 _25948_ (.Y(_06988_),
    .A(_09339_),
    .B(net92));
 sg13g2_o21ai_1 _25949_ (.B1(_06988_),
    .Y(_06989_),
    .A1(net409),
    .A2(net92));
 sg13g2_nor2_1 _25950_ (.A(net830),
    .B(_06989_),
    .Y(_06990_));
 sg13g2_o21ai_1 _25951_ (.B1(_11800_),
    .Y(_06991_),
    .A1(_06987_),
    .A2(_06990_));
 sg13g2_and4_1 _25952_ (.A(_06964_),
    .B(_06971_),
    .C(_06986_),
    .D(_06991_),
    .X(_06992_));
 sg13g2_nand2b_1 _25953_ (.Y(_06993_),
    .B(net15),
    .A_N(_06888_));
 sg13g2_o21ai_1 _25954_ (.B1(_06993_),
    .Y(_02538_),
    .A1(_06955_),
    .A2(_06992_));
 sg13g2_nand2_1 _25955_ (.Y(_06994_),
    .A(net680),
    .B(_09086_));
 sg13g2_nor3_1 _25956_ (.A(_09170_),
    .B(net595),
    .C(_06994_),
    .Y(_06995_));
 sg13g2_nor2b_1 _25957_ (.A(net757),
    .B_N(_06995_),
    .Y(_06996_));
 sg13g2_buf_4 _25958_ (.X(_06997_),
    .A(_06996_));
 sg13g2_mux2_1 _25959_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(net837),
    .S(_06997_),
    .X(_02543_));
 sg13g2_mux2_1 _25960_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(net872),
    .S(_06997_),
    .X(_02544_));
 sg13g2_mux2_1 _25961_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(net836),
    .S(_06997_),
    .X(_02545_));
 sg13g2_mux2_1 _25962_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(net1039),
    .S(_06997_),
    .X(_02546_));
 sg13g2_mux2_1 _25963_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(net1006),
    .S(_06997_),
    .X(_02547_));
 sg13g2_mux2_1 _25964_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(net1005),
    .S(_06997_),
    .X(_02548_));
 sg13g2_mux2_1 _25965_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(net1038),
    .S(_06997_),
    .X(_02549_));
 sg13g2_mux2_1 _25966_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(net1041),
    .S(_06997_),
    .X(_02550_));
 sg13g2_nand3b_1 _25967_ (.B(net681),
    .C(_09086_),
    .Y(_06998_),
    .A_N(net874));
 sg13g2_nor3_1 _25968_ (.A(_09170_),
    .B(net595),
    .C(_06998_),
    .Y(_06999_));
 sg13g2_buf_4 _25969_ (.X(_07000_),
    .A(_06999_));
 sg13g2_mux2_1 _25970_ (.A0(\cpu.spi.r_clk_count[1][0] ),
    .A1(net899),
    .S(_07000_),
    .X(_02551_));
 sg13g2_mux2_1 _25971_ (.A0(\cpu.spi.r_clk_count[1][1] ),
    .A1(net872),
    .S(_07000_),
    .X(_02552_));
 sg13g2_mux2_1 _25972_ (.A0(\cpu.spi.r_clk_count[1][2] ),
    .A1(net871),
    .S(_07000_),
    .X(_02553_));
 sg13g2_mux2_1 _25973_ (.A0(\cpu.spi.r_clk_count[1][3] ),
    .A1(net1039),
    .S(_07000_),
    .X(_02554_));
 sg13g2_mux2_1 _25974_ (.A0(\cpu.spi.r_clk_count[1][4] ),
    .A1(net1006),
    .S(_07000_),
    .X(_02555_));
 sg13g2_mux2_1 _25975_ (.A0(\cpu.spi.r_clk_count[1][5] ),
    .A1(net1005),
    .S(_07000_),
    .X(_02556_));
 sg13g2_mux2_1 _25976_ (.A0(\cpu.spi.r_clk_count[1][6] ),
    .A1(net1038),
    .S(_07000_),
    .X(_02557_));
 sg13g2_mux2_1 _25977_ (.A0(\cpu.spi.r_clk_count[1][7] ),
    .A1(net1041),
    .S(_07000_),
    .X(_02558_));
 sg13g2_nand2_1 _25978_ (.Y(_07001_),
    .A(net676),
    .B(_06995_));
 sg13g2_buf_1 _25979_ (.A(_07001_),
    .X(_07002_));
 sg13g2_mux2_1 _25980_ (.A0(net837),
    .A1(_04853_),
    .S(net90),
    .X(_02559_));
 sg13g2_mux2_1 _25981_ (.A0(net900),
    .A1(_05281_),
    .S(_07002_),
    .X(_02560_));
 sg13g2_mux2_1 _25982_ (.A0(net836),
    .A1(_05338_),
    .S(_07002_),
    .X(_02561_));
 sg13g2_nand2_1 _25983_ (.Y(_07003_),
    .A(_05401_),
    .B(net90));
 sg13g2_o21ai_1 _25984_ (.B1(_07003_),
    .Y(_02562_),
    .A1(_11996_),
    .A2(net90));
 sg13g2_mux2_1 _25985_ (.A0(net994),
    .A1(_05490_),
    .S(net90),
    .X(_02563_));
 sg13g2_mux2_1 _25986_ (.A0(net993),
    .A1(_05553_),
    .S(net90),
    .X(_02564_));
 sg13g2_nand2_1 _25987_ (.Y(_07004_),
    .A(_05641_),
    .B(net90));
 sg13g2_o21ai_1 _25988_ (.B1(_07004_),
    .Y(_02565_),
    .A1(_12018_),
    .A2(net90));
 sg13g2_nand2_1 _25989_ (.Y(_07005_),
    .A(_05034_),
    .B(_07001_));
 sg13g2_o21ai_1 _25990_ (.B1(_07005_),
    .Y(_02566_),
    .A1(_12024_),
    .A2(net90));
 sg13g2_buf_1 _25991_ (.A(_00206_),
    .X(_07006_));
 sg13g2_nor2_1 _25992_ (.A(_07006_),
    .B(net410),
    .Y(_07007_));
 sg13g2_nor4_1 _25993_ (.A(\cpu.spi.r_state[5] ),
    .B(net1125),
    .C(_09236_),
    .D(_11802_),
    .Y(_07008_));
 sg13g2_buf_1 _25994_ (.A(_07008_),
    .X(_07009_));
 sg13g2_nand2_1 _25995_ (.Y(_07010_),
    .A(_07006_),
    .B(net656));
 sg13g2_buf_2 _25996_ (.A(_07010_),
    .X(_07011_));
 sg13g2_nor2_1 _25997_ (.A(_09239_),
    .B(_07011_),
    .Y(_07012_));
 sg13g2_a21oi_1 _25998_ (.A1(_09219_),
    .A2(_07007_),
    .Y(_07013_),
    .B1(_07012_));
 sg13g2_o21ai_1 _25999_ (.B1(_09235_),
    .Y(_07014_),
    .A1(_09158_),
    .A2(net410));
 sg13g2_nand3_1 _26000_ (.B(_07013_),
    .C(_07014_),
    .A(_09280_),
    .Y(_07015_));
 sg13g2_buf_2 _26001_ (.A(_07015_),
    .X(_07016_));
 sg13g2_buf_1 _26002_ (.A(_07016_),
    .X(_07017_));
 sg13g2_buf_1 _26003_ (.A(_07011_),
    .X(_07018_));
 sg13g2_buf_1 _26004_ (.A(_11835_),
    .X(_07019_));
 sg13g2_nand2b_1 _26005_ (.Y(_07020_),
    .B(_07019_),
    .A_N(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_o21ai_1 _26006_ (.B1(_07020_),
    .Y(_07021_),
    .A1(net551),
    .A2(_04853_));
 sg13g2_mux2_1 _26007_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(_03477_),
    .X(_07022_));
 sg13g2_nor2_1 _26008_ (.A(net676),
    .B(_07022_),
    .Y(_07023_));
 sg13g2_a21oi_1 _26009_ (.A1(net668),
    .A2(_07021_),
    .Y(_07024_),
    .B1(_07023_));
 sg13g2_nor2_1 _26010_ (.A(net875),
    .B(_04853_),
    .Y(_07025_));
 sg13g2_a21oi_1 _26011_ (.A1(net875),
    .A2(_00298_),
    .Y(_07026_),
    .B1(_07025_));
 sg13g2_mux2_1 _26012_ (.A0(_00298_),
    .A1(_00297_),
    .S(net1019),
    .X(_07027_));
 sg13g2_nor2_1 _26013_ (.A(net876),
    .B(_07027_),
    .Y(_07028_));
 sg13g2_a21oi_1 _26014_ (.A1(net876),
    .A2(_07026_),
    .Y(_07029_),
    .B1(_07028_));
 sg13g2_nand2_1 _26015_ (.Y(_07030_),
    .A(net360),
    .B(_07029_));
 sg13g2_nor2_1 _26016_ (.A(_09201_),
    .B(net656),
    .Y(_07031_));
 sg13g2_nor2b_1 _26017_ (.A(net106),
    .B_N(_09201_),
    .Y(_07032_));
 sg13g2_a21oi_1 _26018_ (.A1(net88),
    .A2(_07029_),
    .Y(_07033_),
    .B1(_07032_));
 sg13g2_a22oi_1 _26019_ (.Y(_07034_),
    .B1(_07033_),
    .B2(net1051),
    .A2(_07031_),
    .A1(_07030_));
 sg13g2_nand2_1 _26020_ (.Y(_07035_),
    .A(net460),
    .B(_07034_));
 sg13g2_o21ai_1 _26021_ (.B1(_07035_),
    .Y(_07036_),
    .A1(_07018_),
    .A2(_07024_));
 sg13g2_nand2_1 _26022_ (.Y(_07037_),
    .A(_09201_),
    .B(net31));
 sg13g2_o21ai_1 _26023_ (.B1(_07037_),
    .Y(_02567_),
    .A1(_07017_),
    .A2(_07036_));
 sg13g2_nand2b_1 _26024_ (.Y(_07038_),
    .B(net585),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _26025_ (.B1(_07038_),
    .Y(_07039_),
    .A1(net551),
    .A2(_05281_));
 sg13g2_mux2_1 _26026_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net608),
    .X(_07040_));
 sg13g2_nor2_1 _26027_ (.A(net676),
    .B(_07040_),
    .Y(_07041_));
 sg13g2_a21oi_1 _26028_ (.A1(net668),
    .A2(_07039_),
    .Y(_07042_),
    .B1(_07041_));
 sg13g2_nor2_1 _26029_ (.A(net1019),
    .B(_05281_),
    .Y(_07043_));
 sg13g2_a21oi_1 _26030_ (.A1(net875),
    .A2(_00303_),
    .Y(_07044_),
    .B1(_07043_));
 sg13g2_nand2_1 _26031_ (.Y(_07045_),
    .A(net1017),
    .B(_00302_));
 sg13g2_o21ai_1 _26032_ (.B1(_07045_),
    .Y(_07046_),
    .A1(net1018),
    .A2(_05282_));
 sg13g2_nor2_1 _26033_ (.A(net1020),
    .B(_07046_),
    .Y(_07047_));
 sg13g2_a21oi_1 _26034_ (.A1(net876),
    .A2(_07044_),
    .Y(_07048_),
    .B1(_07047_));
 sg13g2_nand2_1 _26035_ (.Y(_07049_),
    .A(net360),
    .B(_07048_));
 sg13g2_xor2_1 _26036_ (.B(\cpu.spi.r_count[1] ),
    .A(_09201_),
    .X(_07050_));
 sg13g2_nor2_1 _26037_ (.A(net656),
    .B(_07050_),
    .Y(_07051_));
 sg13g2_nand2b_1 _26038_ (.Y(_07052_),
    .B(net106),
    .A_N(_07048_));
 sg13g2_o21ai_1 _26039_ (.B1(_07052_),
    .Y(_07053_),
    .A1(net88),
    .A2(_07050_));
 sg13g2_a22oi_1 _26040_ (.Y(_07054_),
    .B1(_07053_),
    .B2(net1051),
    .A2(_07051_),
    .A1(_07049_));
 sg13g2_nand2_1 _26041_ (.Y(_07055_),
    .A(_07018_),
    .B(_07054_));
 sg13g2_o21ai_1 _26042_ (.B1(_07055_),
    .Y(_07056_),
    .A1(net460),
    .A2(_07042_));
 sg13g2_nand2_1 _26043_ (.Y(_07057_),
    .A(\cpu.spi.r_count[1] ),
    .B(net31));
 sg13g2_o21ai_1 _26044_ (.B1(_07057_),
    .Y(_02568_),
    .A1(net31),
    .A2(_07056_));
 sg13g2_nand2b_1 _26045_ (.Y(_07058_),
    .B(net585),
    .A_N(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_o21ai_1 _26046_ (.B1(_07058_),
    .Y(_07059_),
    .A1(net585),
    .A2(_05338_));
 sg13g2_mux2_1 _26047_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net608),
    .X(_07060_));
 sg13g2_nor2_1 _26048_ (.A(net676),
    .B(_07060_),
    .Y(_07061_));
 sg13g2_a21oi_1 _26049_ (.A1(net668),
    .A2(_07059_),
    .Y(_07062_),
    .B1(_07061_));
 sg13g2_nor2_1 _26050_ (.A(_11814_),
    .B(_05338_),
    .Y(_07063_));
 sg13g2_a21oi_1 _26051_ (.A1(net875),
    .A2(_00093_),
    .Y(_07064_),
    .B1(_07063_));
 sg13g2_nand2_1 _26052_ (.Y(_07065_),
    .A(_11817_),
    .B(_00092_));
 sg13g2_o21ai_1 _26053_ (.B1(_07065_),
    .Y(_07066_),
    .A1(net1018),
    .A2(_05339_));
 sg13g2_nor2_1 _26054_ (.A(net1020),
    .B(_07066_),
    .Y(_07067_));
 sg13g2_a21oi_1 _26055_ (.A1(net876),
    .A2(_07064_),
    .Y(_07068_),
    .B1(_07067_));
 sg13g2_nand2_1 _26056_ (.Y(_07069_),
    .A(net360),
    .B(_07068_));
 sg13g2_xnor2_1 _26057_ (.Y(_07070_),
    .A(\cpu.spi.r_count[2] ),
    .B(_09202_));
 sg13g2_nor2_1 _26058_ (.A(net656),
    .B(_07070_),
    .Y(_07071_));
 sg13g2_nand2b_1 _26059_ (.Y(_07072_),
    .B(net106),
    .A_N(_07068_));
 sg13g2_o21ai_1 _26060_ (.B1(_07072_),
    .Y(_07073_),
    .A1(net88),
    .A2(_07070_));
 sg13g2_a22oi_1 _26061_ (.Y(_07074_),
    .B1(_07073_),
    .B2(net1051),
    .A2(_07071_),
    .A1(_07069_));
 sg13g2_nand2_1 _26062_ (.Y(_07075_),
    .A(net460),
    .B(_07074_));
 sg13g2_o21ai_1 _26063_ (.B1(_07075_),
    .Y(_07076_),
    .A1(net460),
    .A2(_07062_));
 sg13g2_nand2_1 _26064_ (.Y(_07077_),
    .A(\cpu.spi.r_count[2] ),
    .B(_07016_));
 sg13g2_o21ai_1 _26065_ (.B1(_07077_),
    .Y(_02569_),
    .A1(net31),
    .A2(_07076_));
 sg13g2_nand2b_1 _26066_ (.Y(_07078_),
    .B(net585),
    .A_N(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_o21ai_1 _26067_ (.B1(_07078_),
    .Y(_07079_),
    .A1(net585),
    .A2(_05401_));
 sg13g2_mux2_1 _26068_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net608),
    .X(_07080_));
 sg13g2_nor2_1 _26069_ (.A(net757),
    .B(_07080_),
    .Y(_07081_));
 sg13g2_a21oi_1 _26070_ (.A1(net668),
    .A2(_07079_),
    .Y(_07082_),
    .B1(_07081_));
 sg13g2_xor2_1 _26071_ (.B(_09203_),
    .A(_09200_),
    .X(_07083_));
 sg13g2_nor2_1 _26072_ (.A(net656),
    .B(_07083_),
    .Y(_07084_));
 sg13g2_nor2_1 _26073_ (.A(net1019),
    .B(_05401_),
    .Y(_07085_));
 sg13g2_a21oi_1 _26074_ (.A1(net1019),
    .A2(_00103_),
    .Y(_07086_),
    .B1(_07085_));
 sg13g2_nand2_1 _26075_ (.Y(_07087_),
    .A(net1017),
    .B(_00102_));
 sg13g2_o21ai_1 _26076_ (.B1(_07087_),
    .Y(_07088_),
    .A1(net1018),
    .A2(_05402_));
 sg13g2_nor2_1 _26077_ (.A(net1020),
    .B(_07088_),
    .Y(_07089_));
 sg13g2_a21oi_1 _26078_ (.A1(net876),
    .A2(_07086_),
    .Y(_07090_),
    .B1(_07089_));
 sg13g2_nand2_1 _26079_ (.Y(_07091_),
    .A(net410),
    .B(_07090_));
 sg13g2_nand2b_1 _26080_ (.Y(_07092_),
    .B(net106),
    .A_N(_07090_));
 sg13g2_o21ai_1 _26081_ (.B1(_07092_),
    .Y(_07093_),
    .A1(net88),
    .A2(_07083_));
 sg13g2_a22oi_1 _26082_ (.Y(_07094_),
    .B1(_07093_),
    .B2(net1051),
    .A2(_07091_),
    .A1(_07084_));
 sg13g2_nand2_1 _26083_ (.Y(_07095_),
    .A(_07011_),
    .B(_07094_));
 sg13g2_o21ai_1 _26084_ (.B1(_07095_),
    .Y(_07096_),
    .A1(net460),
    .A2(_07082_));
 sg13g2_nand2_1 _26085_ (.Y(_07097_),
    .A(_09200_),
    .B(_07016_));
 sg13g2_o21ai_1 _26086_ (.B1(_07097_),
    .Y(_02570_),
    .A1(net31),
    .A2(_07096_));
 sg13g2_nand2b_1 _26087_ (.Y(_07098_),
    .B(net585),
    .A_N(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_o21ai_1 _26088_ (.B1(_07098_),
    .Y(_07099_),
    .A1(_07019_),
    .A2(_05490_));
 sg13g2_mux2_1 _26089_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(_03477_),
    .X(_07100_));
 sg13g2_nor2_1 _26090_ (.A(net757),
    .B(_07100_),
    .Y(_07101_));
 sg13g2_a21oi_1 _26091_ (.A1(net668),
    .A2(_07099_),
    .Y(_07102_),
    .B1(_07101_));
 sg13g2_nor2_1 _26092_ (.A(_09200_),
    .B(_09203_),
    .Y(_07103_));
 sg13g2_xnor2_1 _26093_ (.Y(_07104_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07103_));
 sg13g2_nor2_1 _26094_ (.A(net656),
    .B(_07104_),
    .Y(_07105_));
 sg13g2_nor2_1 _26095_ (.A(_11816_),
    .B(_05490_),
    .Y(_07106_));
 sg13g2_a21oi_1 _26096_ (.A1(_11814_),
    .A2(_00113_),
    .Y(_07107_),
    .B1(_07106_));
 sg13g2_nand2_1 _26097_ (.Y(_07108_),
    .A(_11817_),
    .B(_00112_));
 sg13g2_o21ai_1 _26098_ (.B1(_07108_),
    .Y(_07109_),
    .A1(_11816_),
    .A2(_05491_));
 sg13g2_nor2_1 _26099_ (.A(_11809_),
    .B(_07109_),
    .Y(_07110_));
 sg13g2_a21oi_1 _26100_ (.A1(net876),
    .A2(_07107_),
    .Y(_07111_),
    .B1(_07110_));
 sg13g2_nand2_1 _26101_ (.Y(_07112_),
    .A(net410),
    .B(_07111_));
 sg13g2_nand2b_1 _26102_ (.Y(_07113_),
    .B(net106),
    .A_N(_07111_));
 sg13g2_o21ai_1 _26103_ (.B1(_07113_),
    .Y(_07114_),
    .A1(net88),
    .A2(_07104_));
 sg13g2_a22oi_1 _26104_ (.Y(_07115_),
    .B1(_07114_),
    .B2(net1051),
    .A2(_07112_),
    .A1(_07105_));
 sg13g2_nand2_1 _26105_ (.Y(_07116_),
    .A(_07011_),
    .B(_07115_));
 sg13g2_o21ai_1 _26106_ (.B1(_07116_),
    .Y(_07117_),
    .A1(net460),
    .A2(_07102_));
 sg13g2_nand2_1 _26107_ (.Y(_07118_),
    .A(\cpu.spi.r_count[4] ),
    .B(_07016_));
 sg13g2_o21ai_1 _26108_ (.B1(_07118_),
    .Y(_02571_),
    .A1(net31),
    .A2(_07117_));
 sg13g2_nand2b_1 _26109_ (.Y(_07119_),
    .B(net608),
    .A_N(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_o21ai_1 _26110_ (.B1(_07119_),
    .Y(_07120_),
    .A1(net585),
    .A2(_05553_));
 sg13g2_mux2_1 _26111_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net608),
    .X(_07121_));
 sg13g2_nor2_1 _26112_ (.A(net757),
    .B(_07121_),
    .Y(_07122_));
 sg13g2_a21oi_1 _26113_ (.A1(net676),
    .A2(_07120_),
    .Y(_07123_),
    .B1(_07122_));
 sg13g2_nor2_1 _26114_ (.A(net1018),
    .B(_05553_),
    .Y(_07124_));
 sg13g2_a21oi_1 _26115_ (.A1(net1019),
    .A2(_00119_),
    .Y(_07125_),
    .B1(_07124_));
 sg13g2_nand2_1 _26116_ (.Y(_07126_),
    .A(net1017),
    .B(_00118_));
 sg13g2_o21ai_1 _26117_ (.B1(_07126_),
    .Y(_07127_),
    .A1(net1018),
    .A2(_05554_));
 sg13g2_nor2_1 _26118_ (.A(net1020),
    .B(_07127_),
    .Y(_07128_));
 sg13g2_a21oi_1 _26119_ (.A1(net876),
    .A2(_07125_),
    .Y(_07129_),
    .B1(_07128_));
 sg13g2_nand2_1 _26120_ (.Y(_07130_),
    .A(net360),
    .B(_07129_));
 sg13g2_xnor2_1 _26121_ (.Y(_07131_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09204_));
 sg13g2_nor2_1 _26122_ (.A(net656),
    .B(_07131_),
    .Y(_07132_));
 sg13g2_nand2b_1 _26123_ (.Y(_07133_),
    .B(net106),
    .A_N(_07129_));
 sg13g2_o21ai_1 _26124_ (.B1(_07133_),
    .Y(_07134_),
    .A1(net88),
    .A2(_07131_));
 sg13g2_a22oi_1 _26125_ (.Y(_07135_),
    .B1(_07134_),
    .B2(net1051),
    .A2(_07132_),
    .A1(_07130_));
 sg13g2_nand2_1 _26126_ (.Y(_07136_),
    .A(_07011_),
    .B(_07135_));
 sg13g2_o21ai_1 _26127_ (.B1(_07136_),
    .Y(_07137_),
    .A1(net460),
    .A2(_07123_));
 sg13g2_nand2_1 _26128_ (.Y(_07138_),
    .A(\cpu.spi.r_count[5] ),
    .B(_07016_));
 sg13g2_o21ai_1 _26129_ (.B1(_07138_),
    .Y(_02572_),
    .A1(net31),
    .A2(_07137_));
 sg13g2_nand2b_1 _26130_ (.Y(_07139_),
    .B(net608),
    .A_N(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_o21ai_1 _26131_ (.B1(_07139_),
    .Y(_07140_),
    .A1(net585),
    .A2(_05641_));
 sg13g2_mux2_1 _26132_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net608),
    .X(_07141_));
 sg13g2_nor2_1 _26133_ (.A(net757),
    .B(_07141_),
    .Y(_07142_));
 sg13g2_a21oi_1 _26134_ (.A1(net676),
    .A2(_07140_),
    .Y(_07143_),
    .B1(_07142_));
 sg13g2_nor2_1 _26135_ (.A(net1018),
    .B(_05641_),
    .Y(_07144_));
 sg13g2_a21oi_1 _26136_ (.A1(net1019),
    .A2(_00130_),
    .Y(_07145_),
    .B1(_07144_));
 sg13g2_nand2_1 _26137_ (.Y(_07146_),
    .A(net1017),
    .B(_00129_));
 sg13g2_o21ai_1 _26138_ (.B1(_07146_),
    .Y(_07147_),
    .A1(net1018),
    .A2(_05642_));
 sg13g2_nor2_1 _26139_ (.A(net1020),
    .B(_07147_),
    .Y(_07148_));
 sg13g2_a21oi_1 _26140_ (.A1(net876),
    .A2(_07145_),
    .Y(_07149_),
    .B1(_07148_));
 sg13g2_nand2_1 _26141_ (.Y(_07150_),
    .A(net360),
    .B(_07149_));
 sg13g2_xnor2_1 _26142_ (.Y(_07151_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09205_));
 sg13g2_nor2_1 _26143_ (.A(_07009_),
    .B(_07151_),
    .Y(_07152_));
 sg13g2_nand2b_1 _26144_ (.Y(_07153_),
    .B(net106),
    .A_N(_07149_));
 sg13g2_o21ai_1 _26145_ (.B1(_07153_),
    .Y(_07154_),
    .A1(_09221_),
    .A2(_07151_));
 sg13g2_a22oi_1 _26146_ (.Y(_07155_),
    .B1(_07154_),
    .B2(_09250_),
    .A2(_07152_),
    .A1(_07150_));
 sg13g2_nand2_1 _26147_ (.Y(_07156_),
    .A(_07011_),
    .B(_07155_));
 sg13g2_o21ai_1 _26148_ (.B1(_07156_),
    .Y(_07157_),
    .A1(net460),
    .A2(_07143_));
 sg13g2_nand2_1 _26149_ (.Y(_07158_),
    .A(\cpu.spi.r_count[6] ),
    .B(_07016_));
 sg13g2_o21ai_1 _26150_ (.B1(_07158_),
    .Y(_02573_),
    .A1(_07017_),
    .A2(_07157_));
 sg13g2_nand2b_1 _26151_ (.Y(_07159_),
    .B(net681),
    .A_N(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_o21ai_1 _26152_ (.B1(_07159_),
    .Y(_07160_),
    .A1(net681),
    .A2(_05034_));
 sg13g2_mux2_1 _26153_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(net681),
    .X(_07161_));
 sg13g2_nor2_1 _26154_ (.A(net874),
    .B(_07161_),
    .Y(_07162_));
 sg13g2_a21oi_1 _26155_ (.A1(net874),
    .A2(_07160_),
    .Y(_07163_),
    .B1(_07162_));
 sg13g2_nor2_1 _26156_ (.A(_07011_),
    .B(_07163_),
    .Y(_07164_));
 sg13g2_nor2_1 _26157_ (.A(net1017),
    .B(_05034_),
    .Y(_07165_));
 sg13g2_a21oi_1 _26158_ (.A1(net1019),
    .A2(_00141_),
    .Y(_07166_),
    .B1(_07165_));
 sg13g2_nand2_1 _26159_ (.Y(_07167_),
    .A(_11813_),
    .B(_00140_));
 sg13g2_o21ai_1 _26160_ (.B1(_07167_),
    .Y(_07168_),
    .A1(net1017),
    .A2(_05036_));
 sg13g2_nor2_1 _26161_ (.A(_11808_),
    .B(_07168_),
    .Y(_07169_));
 sg13g2_a21oi_1 _26162_ (.A1(net1020),
    .A2(_07166_),
    .Y(_07170_),
    .B1(_07169_));
 sg13g2_nor2_1 _26163_ (.A(_09220_),
    .B(_09210_),
    .Y(_07171_));
 sg13g2_a21oi_1 _26164_ (.A1(net88),
    .A2(_07170_),
    .Y(_07172_),
    .B1(_07171_));
 sg13g2_nor2_1 _26165_ (.A(_09199_),
    .B(_07170_),
    .Y(_07173_));
 sg13g2_nor2b_1 _26166_ (.A(_09207_),
    .B_N(_09199_),
    .Y(_07174_));
 sg13g2_a21oi_1 _26167_ (.A1(_09207_),
    .A2(_07173_),
    .Y(_07175_),
    .B1(_07174_));
 sg13g2_o21ai_1 _26168_ (.B1(_07011_),
    .Y(_07176_),
    .A1(net656),
    .A2(_07175_));
 sg13g2_a21oi_1 _26169_ (.A1(net1054),
    .A2(_07172_),
    .Y(_07177_),
    .B1(_07176_));
 sg13g2_or2_1 _26170_ (.X(_07178_),
    .B(_07177_),
    .A(_07164_));
 sg13g2_nor3_1 _26171_ (.A(_09172_),
    .B(_09207_),
    .C(_07164_),
    .Y(_07179_));
 sg13g2_o21ai_1 _26172_ (.B1(_09199_),
    .Y(_07180_),
    .A1(_07016_),
    .A2(_07179_));
 sg13g2_o21ai_1 _26173_ (.B1(_07180_),
    .Y(_02574_),
    .A1(net31),
    .A2(_07178_));
 sg13g2_inv_1 _26174_ (.Y(_07181_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_mux4_1 _26175_ (.S0(_05511_),
    .A0(_09107_),
    .A1(_09094_),
    .A2(_09091_),
    .A3(_09114_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07182_));
 sg13g2_nand2_1 _26176_ (.Y(_07183_),
    .A(net3),
    .B(_05511_));
 sg13g2_nand2b_1 _26177_ (.Y(_07184_),
    .B(_09104_),
    .A_N(_05511_));
 sg13g2_nand3_1 _26178_ (.B(_07183_),
    .C(_07184_),
    .A(_06389_),
    .Y(_07185_));
 sg13g2_o21ai_1 _26179_ (.B1(_07185_),
    .Y(_07186_),
    .A1(_06389_),
    .A2(_07182_));
 sg13g2_nand2b_1 _26180_ (.Y(_07187_),
    .B(_05511_),
    .A_N(_09096_));
 sg13g2_o21ai_1 _26181_ (.B1(_07187_),
    .Y(_07188_),
    .A1(_09101_),
    .A2(_05511_));
 sg13g2_a21o_1 _26182_ (.A2(_07188_),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B1(_00135_),
    .X(_07189_));
 sg13g2_mux4_1 _26183_ (.S0(_05511_),
    .A0(_09089_),
    .A1(_09112_),
    .A2(_09100_),
    .A3(_09109_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07190_));
 sg13g2_nor3_1 _26184_ (.A(_07181_),
    .B(_06389_),
    .C(_07190_),
    .Y(_07191_));
 sg13g2_a221oi_1 _26185_ (.B2(_06389_),
    .C1(_07191_),
    .B1(_07189_),
    .A1(_07181_),
    .Y(_07192_),
    .A2(_07186_));
 sg13g2_mux4_1 _26186_ (.S0(_04826_),
    .A0(_09089_),
    .A1(_09112_),
    .A2(_09100_),
    .A3(_09109_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07193_));
 sg13g2_nand2_1 _26187_ (.Y(_07194_),
    .A(_09096_),
    .B(_04826_));
 sg13g2_nand2b_1 _26188_ (.Y(_07195_),
    .B(_09101_),
    .A_N(_04826_));
 sg13g2_nand3_1 _26189_ (.B(_07194_),
    .C(_07195_),
    .A(_06386_),
    .Y(_07196_));
 sg13g2_o21ai_1 _26190_ (.B1(_07196_),
    .Y(_07197_),
    .A1(_06386_),
    .A2(_07193_));
 sg13g2_nor2_1 _26191_ (.A(_09104_),
    .B(_04826_),
    .Y(_07198_));
 sg13g2_a21oi_1 _26192_ (.A1(_05542_),
    .A2(_04826_),
    .Y(_07199_),
    .B1(_07198_));
 sg13g2_o21ai_1 _26193_ (.B1(_05357_),
    .Y(_07200_),
    .A1(_06384_),
    .A2(_07199_));
 sg13g2_mux4_1 _26194_ (.S0(_04826_),
    .A0(_09107_),
    .A1(_09094_),
    .A2(_09091_),
    .A3(_09114_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07201_));
 sg13g2_nor3_1 _26195_ (.A(_06384_),
    .B(_06386_),
    .C(_07201_),
    .Y(_07202_));
 sg13g2_a221oi_1 _26196_ (.B2(_06386_),
    .C1(_07202_),
    .B1(_07200_),
    .A1(_06384_),
    .Y(_07203_),
    .A2(_07197_));
 sg13g2_mux2_1 _26197_ (.A0(_07192_),
    .A1(_07203_),
    .S(_11821_),
    .X(_07204_));
 sg13g2_nor2_1 _26198_ (.A(net1126),
    .B(_11866_),
    .Y(_07205_));
 sg13g2_nor2b_1 _26199_ (.A(_09174_),
    .B_N(net1126),
    .Y(_07206_));
 sg13g2_a22oi_1 _26200_ (.Y(_07207_),
    .B1(_07206_),
    .B2(_11866_),
    .A2(_07205_),
    .A1(_09174_));
 sg13g2_nand3b_1 _26201_ (.B(_09211_),
    .C(net919),
    .Y(_07208_),
    .A_N(_07207_));
 sg13g2_buf_4 _26202_ (.X(_07209_),
    .A(_07208_));
 sg13g2_mux2_1 _26203_ (.A0(_07204_),
    .A1(_09189_),
    .S(_07209_),
    .X(_02578_));
 sg13g2_mux2_1 _26204_ (.A0(_09189_),
    .A1(_09188_),
    .S(_07209_),
    .X(_02579_));
 sg13g2_mux2_1 _26205_ (.A0(_09188_),
    .A1(_09192_),
    .S(_07209_),
    .X(_02580_));
 sg13g2_mux2_1 _26206_ (.A0(_09192_),
    .A1(_09186_),
    .S(_07209_),
    .X(_02581_));
 sg13g2_mux2_1 _26207_ (.A0(_09186_),
    .A1(_09194_),
    .S(_07209_),
    .X(_02582_));
 sg13g2_mux2_1 _26208_ (.A0(_09194_),
    .A1(_09193_),
    .S(_07209_),
    .X(_02583_));
 sg13g2_mux2_1 _26209_ (.A0(_09193_),
    .A1(_09187_),
    .S(_07209_),
    .X(_02584_));
 sg13g2_mux2_1 _26210_ (.A0(_09187_),
    .A1(\cpu.spi.r_in[7] ),
    .S(_07209_),
    .X(_02585_));
 sg13g2_inv_1 _26211_ (.Y(_07210_),
    .A(_09247_));
 sg13g2_nor3_2 _26212_ (.A(net668),
    .B(_07210_),
    .C(_06994_),
    .Y(_07211_));
 sg13g2_mux2_1 _26213_ (.A0(\cpu.spi.r_mode[0][0] ),
    .A1(net899),
    .S(_07211_),
    .X(_02587_));
 sg13g2_mux2_1 _26214_ (.A0(_11825_),
    .A1(net872),
    .S(_07211_),
    .X(_02588_));
 sg13g2_nor2_2 _26215_ (.A(_07210_),
    .B(_06998_),
    .Y(_07212_));
 sg13g2_mux2_1 _26216_ (.A0(\cpu.spi.r_mode[1][0] ),
    .A1(net899),
    .S(_07212_),
    .X(_02589_));
 sg13g2_mux2_1 _26217_ (.A0(_11826_),
    .A1(net872),
    .S(_07212_),
    .X(_02590_));
 sg13g2_nand4_1 _26218_ (.B(net680),
    .C(_09086_),
    .A(net676),
    .Y(_07213_),
    .D(_09247_));
 sg13g2_buf_1 _26219_ (.A(_07213_),
    .X(_07214_));
 sg13g2_mux2_1 _26220_ (.A0(net837),
    .A1(\cpu.spi.r_mode[2][0] ),
    .S(_07214_),
    .X(_02591_));
 sg13g2_mux2_1 _26221_ (.A0(net900),
    .A1(_11830_),
    .S(_07214_),
    .X(_02592_));
 sg13g2_nand2_1 _26222_ (.Y(_07215_),
    .A(_09239_),
    .B(_09248_));
 sg13g2_nor2_1 _26223_ (.A(net1127),
    .B(_09239_),
    .Y(_07216_));
 sg13g2_a22oi_1 _26224_ (.Y(_07217_),
    .B1(_07216_),
    .B2(_11807_),
    .A2(_11867_),
    .A1(net1125));
 sg13g2_nand4_1 _26225_ (.B(_11862_),
    .C(_11871_),
    .A(_07215_),
    .Y(_07218_),
    .D(_07217_));
 sg13g2_buf_1 _26226_ (.A(_07218_),
    .X(_07219_));
 sg13g2_buf_1 _26227_ (.A(_11866_),
    .X(_07220_));
 sg13g2_nor2b_1 _26228_ (.A(_07220_),
    .B_N(_00204_),
    .Y(_07221_));
 sg13g2_o21ai_1 _26229_ (.B1(_09250_),
    .Y(_07222_),
    .A1(_07006_),
    .A2(_07221_));
 sg13g2_o21ai_1 _26230_ (.B1(_07222_),
    .Y(_07223_),
    .A1(_09217_),
    .A2(_09987_));
 sg13g2_a21oi_1 _26231_ (.A1(_11807_),
    .A2(_07223_),
    .Y(_07224_),
    .B1(net33));
 sg13g2_a21o_1 _26232_ (.A2(_07219_),
    .A1(\cpu.spi.r_out[0] ),
    .B1(_07224_),
    .X(_02593_));
 sg13g2_buf_1 _26233_ (.A(_09234_),
    .X(_07225_));
 sg13g2_mux2_1 _26234_ (.A0(_00162_),
    .A1(_00204_),
    .S(_07220_),
    .X(_07226_));
 sg13g2_nor2_1 _26235_ (.A(_09171_),
    .B(_11855_),
    .Y(_07227_));
 sg13g2_buf_2 _26236_ (.A(_07227_),
    .X(_07228_));
 sg13g2_a22oi_1 _26237_ (.Y(_07229_),
    .B1(_07228_),
    .B2(_09995_),
    .A2(net873),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26238_ (.B1(_07229_),
    .Y(_07230_),
    .A1(net827),
    .A2(_07226_));
 sg13g2_mux2_1 _26239_ (.A0(_07230_),
    .A1(\cpu.spi.r_out[1] ),
    .S(net33),
    .X(_02594_));
 sg13g2_mux2_1 _26240_ (.A0(_00163_),
    .A1(_00162_),
    .S(net584),
    .X(_07231_));
 sg13g2_a22oi_1 _26241_ (.Y(_07232_),
    .B1(_07228_),
    .B2(_10002_),
    .A2(net873),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26242_ (.B1(_07232_),
    .Y(_07233_),
    .A1(net827),
    .A2(_07231_));
 sg13g2_mux2_1 _26243_ (.A0(_07233_),
    .A1(\cpu.spi.r_out[2] ),
    .S(net33),
    .X(_02595_));
 sg13g2_mux2_1 _26244_ (.A0(_00268_),
    .A1(_00163_),
    .S(net584),
    .X(_07234_));
 sg13g2_a22oi_1 _26245_ (.Y(_07235_),
    .B1(_07228_),
    .B2(_10007_),
    .A2(net873),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26246_ (.B1(_07235_),
    .Y(_07236_),
    .A1(net827),
    .A2(_07234_));
 sg13g2_mux2_1 _26247_ (.A0(_07236_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net33),
    .X(_02596_));
 sg13g2_mux2_1 _26248_ (.A0(_00164_),
    .A1(_00268_),
    .S(net584),
    .X(_07237_));
 sg13g2_a22oi_1 _26249_ (.Y(_07238_),
    .B1(_07228_),
    .B2(_10013_),
    .A2(net873),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26250_ (.B1(_07238_),
    .Y(_07239_),
    .A1(net827),
    .A2(_07237_));
 sg13g2_mux2_1 _26251_ (.A0(_07239_),
    .A1(\cpu.spi.r_out[4] ),
    .S(net33),
    .X(_02597_));
 sg13g2_mux2_1 _26252_ (.A0(_00165_),
    .A1(_00164_),
    .S(net584),
    .X(_07240_));
 sg13g2_a22oi_1 _26253_ (.Y(_07241_),
    .B1(_07228_),
    .B2(_10019_),
    .A2(net873),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26254_ (.B1(_07241_),
    .Y(_07242_),
    .A1(net827),
    .A2(_07240_));
 sg13g2_mux2_1 _26255_ (.A0(_07242_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net33),
    .X(_02598_));
 sg13g2_inv_1 _26256_ (.Y(_07243_),
    .A(_00166_));
 sg13g2_nand2_1 _26257_ (.Y(_07244_),
    .A(_00165_),
    .B(net584));
 sg13g2_o21ai_1 _26258_ (.B1(_07244_),
    .Y(_07245_),
    .A1(_07243_),
    .A2(net584));
 sg13g2_a22oi_1 _26259_ (.Y(_07246_),
    .B1(_07228_),
    .B2(net1119),
    .A2(net873),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26260_ (.B1(_07246_),
    .Y(_07247_),
    .A1(_07225_),
    .A2(_07245_));
 sg13g2_mux2_1 _26261_ (.A0(_07247_),
    .A1(\cpu.spi.r_out[6] ),
    .S(net33),
    .X(_02599_));
 sg13g2_buf_1 _26262_ (.A(_00262_),
    .X(_07248_));
 sg13g2_nor2_1 _26263_ (.A(_07248_),
    .B(net584),
    .Y(_07249_));
 sg13g2_a21oi_1 _26264_ (.A1(_07243_),
    .A2(net584),
    .Y(_07250_),
    .B1(_07249_));
 sg13g2_a22oi_1 _26265_ (.Y(_07251_),
    .B1(_07228_),
    .B2(net1118),
    .A2(net873),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26266_ (.B1(_07251_),
    .Y(_07252_),
    .A1(_07225_),
    .A2(_07250_));
 sg13g2_mux2_1 _26267_ (.A0(_07252_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net33),
    .X(_02600_));
 sg13g2_mux2_1 _26268_ (.A0(_11827_),
    .A1(net551),
    .S(_09249_),
    .X(_02603_));
 sg13g2_nand2_1 _26269_ (.Y(_07253_),
    .A(net613),
    .B(_09249_));
 sg13g2_o21ai_1 _26270_ (.B1(_07253_),
    .Y(_02604_),
    .A1(_11824_),
    .A2(_09249_));
 sg13g2_mux2_1 _26271_ (.A0(\cpu.spi.r_src[0] ),
    .A1(net871),
    .S(_07211_),
    .X(_02605_));
 sg13g2_mux2_1 _26272_ (.A0(\cpu.spi.r_src[1] ),
    .A1(net871),
    .S(_07212_),
    .X(_02606_));
 sg13g2_mux2_1 _26273_ (.A0(net836),
    .A1(_11811_),
    .S(_07214_),
    .X(_02607_));
 sg13g2_nor2b_1 _26274_ (.A(_09170_),
    .B_N(_05038_),
    .Y(_07254_));
 sg13g2_buf_4 _26275_ (.X(_07255_),
    .A(_07254_));
 sg13g2_mux2_1 _26276_ (.A0(\cpu.spi.r_timeout[0] ),
    .A1(net899),
    .S(_07255_),
    .X(_02608_));
 sg13g2_mux2_1 _26277_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(net872),
    .S(_07255_),
    .X(_02609_));
 sg13g2_mux2_1 _26278_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(net871),
    .S(_07255_),
    .X(_02610_));
 sg13g2_mux2_1 _26279_ (.A0(\cpu.spi.r_timeout[3] ),
    .A1(net1039),
    .S(_07255_),
    .X(_02611_));
 sg13g2_mux2_1 _26280_ (.A0(\cpu.spi.r_timeout[4] ),
    .A1(net1006),
    .S(_07255_),
    .X(_02612_));
 sg13g2_mux2_1 _26281_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(net1005),
    .S(_07255_),
    .X(_02613_));
 sg13g2_mux2_1 _26282_ (.A0(\cpu.spi.r_timeout[6] ),
    .A1(net1038),
    .S(_07255_),
    .X(_02614_));
 sg13g2_mux2_1 _26283_ (.A0(\cpu.spi.r_timeout[7] ),
    .A1(net1041),
    .S(_07255_),
    .X(_02615_));
 sg13g2_inv_1 _26284_ (.Y(_07256_),
    .A(\cpu.spi.r_timeout_count[0] ));
 sg13g2_nand3_1 _26285_ (.B(_09197_),
    .C(_09209_),
    .A(_09185_),
    .Y(_07257_));
 sg13g2_nor3_1 _26286_ (.A(_00207_),
    .B(_09177_),
    .C(_07257_),
    .Y(_07258_));
 sg13g2_nand2_1 _26287_ (.Y(_07259_),
    .A(_09173_),
    .B(_07257_));
 sg13g2_o21ai_1 _26288_ (.B1(_07259_),
    .Y(_07260_),
    .A1(_09173_),
    .A2(net1127));
 sg13g2_nor4_1 _26289_ (.A(net1053),
    .B(_09235_),
    .C(_07258_),
    .D(_07260_),
    .Y(_07261_));
 sg13g2_buf_2 _26290_ (.A(_07261_),
    .X(_07262_));
 sg13g2_buf_1 _26291_ (.A(_07262_),
    .X(_07263_));
 sg13g2_mux2_1 _26292_ (.A0(_00265_),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(net1054),
    .X(_07264_));
 sg13g2_nand2_1 _26293_ (.Y(_07265_),
    .A(net32),
    .B(_07264_));
 sg13g2_o21ai_1 _26294_ (.B1(_07265_),
    .Y(_02616_),
    .A1(_07256_),
    .A2(net32));
 sg13g2_o21ai_1 _26295_ (.B1(net32),
    .Y(_07266_),
    .A1(_07256_),
    .A2(net914));
 sg13g2_nor2_1 _26296_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .Y(_07267_));
 sg13g2_mux2_1 _26297_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(_07267_),
    .S(net827),
    .X(_07268_));
 sg13g2_a22oi_1 _26298_ (.Y(_07269_),
    .B1(_07268_),
    .B2(net32),
    .A2(_07266_),
    .A1(\cpu.spi.r_timeout_count[1] ));
 sg13g2_inv_1 _26299_ (.Y(_02617_),
    .A(_07269_));
 sg13g2_o21ai_1 _26300_ (.B1(_07262_),
    .Y(_07270_),
    .A1(net914),
    .A2(_07267_));
 sg13g2_mux2_1 _26301_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(_09178_),
    .S(net827),
    .X(_07271_));
 sg13g2_a22oi_1 _26302_ (.Y(_07272_),
    .B1(_07271_),
    .B2(net32),
    .A2(_07270_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_inv_1 _26303_ (.Y(_02618_),
    .A(_07272_));
 sg13g2_o21ai_1 _26304_ (.B1(_07262_),
    .Y(_07273_),
    .A1(net914),
    .A2(_09178_));
 sg13g2_nand2b_1 _26305_ (.Y(_07274_),
    .B(_09178_),
    .A_N(\cpu.spi.r_timeout_count[3] ));
 sg13g2_nand2_1 _26306_ (.Y(_07275_),
    .A(net1054),
    .B(\cpu.spi.r_timeout[3] ));
 sg13g2_o21ai_1 _26307_ (.B1(_07275_),
    .Y(_07276_),
    .A1(net914),
    .A2(_07274_));
 sg13g2_a22oi_1 _26308_ (.Y(_07277_),
    .B1(_07276_),
    .B2(net32),
    .A2(_07273_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_inv_1 _26309_ (.Y(_02619_),
    .A(_07277_));
 sg13g2_o21ai_1 _26310_ (.B1(_07262_),
    .Y(_07278_),
    .A1(net914),
    .A2(_09179_));
 sg13g2_nand2_1 _26311_ (.Y(_07279_),
    .A(net1054),
    .B(\cpu.spi.r_timeout[4] ));
 sg13g2_o21ai_1 _26312_ (.B1(_07279_),
    .Y(_07280_),
    .A1(net914),
    .A2(_09180_));
 sg13g2_a22oi_1 _26313_ (.Y(_07281_),
    .B1(_07280_),
    .B2(net32),
    .A2(_07278_),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_inv_1 _26314_ (.Y(_02620_),
    .A(_07281_));
 sg13g2_nor2_1 _26315_ (.A(\cpu.spi.r_timeout_count[4] ),
    .B(_07274_),
    .Y(_07282_));
 sg13g2_o21ai_1 _26316_ (.B1(_07262_),
    .Y(_07283_),
    .A1(net914),
    .A2(_07282_));
 sg13g2_mux2_1 _26317_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(_09181_),
    .S(net827),
    .X(_07284_));
 sg13g2_a22oi_1 _26318_ (.Y(_07285_),
    .B1(_07284_),
    .B2(net32),
    .A2(_07283_),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_inv_1 _26319_ (.Y(_02621_),
    .A(_07285_));
 sg13g2_o21ai_1 _26320_ (.B1(_07262_),
    .Y(_07286_),
    .A1(net1054),
    .A2(_09181_));
 sg13g2_nand2_1 _26321_ (.Y(_07287_),
    .A(net1054),
    .B(\cpu.spi.r_timeout[6] ));
 sg13g2_o21ai_1 _26322_ (.B1(_07287_),
    .Y(_07288_),
    .A1(_09251_),
    .A2(_09183_));
 sg13g2_a22oi_1 _26323_ (.Y(_07289_),
    .B1(_07288_),
    .B2(_07263_),
    .A2(_07286_),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_inv_1 _26324_ (.Y(_02622_),
    .A(_07289_));
 sg13g2_inv_1 _26325_ (.Y(_07290_),
    .A(_09183_));
 sg13g2_o21ai_1 _26326_ (.B1(_07262_),
    .Y(_07291_),
    .A1(net1054),
    .A2(_07290_));
 sg13g2_nor3_1 _26327_ (.A(\cpu.spi.r_timeout_count[7] ),
    .B(net1051),
    .C(_09183_),
    .Y(_07292_));
 sg13g2_a21o_1 _26328_ (.A2(\cpu.spi.r_timeout[7] ),
    .A1(_09251_),
    .B1(_07292_),
    .X(_07293_));
 sg13g2_a22oi_1 _26329_ (.Y(_07294_),
    .B1(_07293_),
    .B2(_07263_),
    .A2(_07291_),
    .A1(\cpu.spi.r_timeout_count[7] ));
 sg13g2_inv_1 _26330_ (.Y(_02623_),
    .A(_07294_));
 sg13g2_buf_1 _26331_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07295_));
 sg13g2_nor2_1 _26332_ (.A(_07295_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07296_));
 sg13g2_nand2_1 _26333_ (.Y(_07297_),
    .A(_09869_),
    .B(_07296_));
 sg13g2_nor2_1 _26334_ (.A(net1053),
    .B(_07297_),
    .Y(_07298_));
 sg13g2_buf_1 _26335_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07299_));
 sg13g2_buf_1 _26336_ (.A(net1085),
    .X(_07300_));
 sg13g2_buf_1 _26337_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07301_));
 sg13g2_buf_1 _26338_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07302_));
 sg13g2_buf_1 _26339_ (.A(_07302_),
    .X(_07303_));
 sg13g2_nor2_2 _26340_ (.A(_07301_),
    .B(_07303_),
    .Y(_07304_));
 sg13g2_buf_2 _26341_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07305_));
 sg13g2_inv_1 _26342_ (.Y(_07306_),
    .A(_07305_));
 sg13g2_nand3_1 _26343_ (.B(net940),
    .C(_07304_),
    .A(_07306_),
    .Y(_07307_));
 sg13g2_o21ai_1 _26344_ (.B1(_07307_),
    .Y(_07308_),
    .A1(net940),
    .A2(_07304_));
 sg13g2_and2_1 _26345_ (.A(_07298_),
    .B(_07308_),
    .X(_07309_));
 sg13g2_buf_2 _26346_ (.A(_07309_),
    .X(_07310_));
 sg13g2_mux2_1 _26347_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07310_),
    .X(_02636_));
 sg13g2_mux2_1 _26348_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07310_),
    .X(_02637_));
 sg13g2_mux2_1 _26349_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07310_),
    .X(_02638_));
 sg13g2_mux2_1 _26350_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07310_),
    .X(_02639_));
 sg13g2_mux2_1 _26351_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07310_),
    .X(_02640_));
 sg13g2_mux2_1 _26352_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07310_),
    .X(_02641_));
 sg13g2_xor2_1 _26353_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07311_));
 sg13g2_mux2_1 _26354_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07311_),
    .S(_07310_),
    .X(_02642_));
 sg13g2_and4_1 _26355_ (.A(_07305_),
    .B(net940),
    .C(_07298_),
    .D(_07304_),
    .X(_07312_));
 sg13g2_buf_1 _26356_ (.A(_07312_),
    .X(_07313_));
 sg13g2_mux2_1 _26357_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net173),
    .X(_02643_));
 sg13g2_mux2_1 _26358_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net173),
    .X(_02644_));
 sg13g2_mux2_1 _26359_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net173),
    .X(_02645_));
 sg13g2_mux2_1 _26360_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net173),
    .X(_02646_));
 sg13g2_mux2_1 _26361_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net173),
    .X(_02647_));
 sg13g2_mux2_1 _26362_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net173),
    .X(_02648_));
 sg13g2_mux2_1 _26363_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07313_),
    .X(_02649_));
 sg13g2_mux2_1 _26364_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07311_),
    .S(net173),
    .X(_02650_));
 sg13g2_buf_1 _26365_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07314_));
 sg13g2_buf_1 _26366_ (.A(_07314_),
    .X(_07315_));
 sg13g2_buf_1 _26367_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07316_));
 sg13g2_buf_1 _26368_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07317_));
 sg13g2_and2_1 _26369_ (.A(net1083),
    .B(_07317_),
    .X(_07318_));
 sg13g2_buf_1 _26370_ (.A(_07318_),
    .X(_07319_));
 sg13g2_nor2_1 _26371_ (.A(_09152_),
    .B(net1057),
    .Y(_07320_));
 sg13g2_and3_1 _26372_ (.X(_07321_),
    .A(_11833_),
    .B(_07320_),
    .C(_06367_));
 sg13g2_buf_2 _26373_ (.A(_07321_),
    .X(_07322_));
 sg13g2_nand2_2 _26374_ (.Y(_07323_),
    .A(net430),
    .B(_07322_));
 sg13g2_nand3_1 _26375_ (.B(_07319_),
    .C(_07323_),
    .A(net938),
    .Y(_07324_));
 sg13g2_buf_1 _26376_ (.A(_07317_),
    .X(_07325_));
 sg13g2_nor2_1 _26377_ (.A(net1083),
    .B(net938),
    .Y(_07326_));
 sg13g2_o21ai_1 _26378_ (.B1(_07326_),
    .Y(_07327_),
    .A1(net937),
    .A2(_07323_));
 sg13g2_buf_1 _26379_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07328_));
 sg13g2_buf_1 _26380_ (.A(_07328_),
    .X(_07329_));
 sg13g2_a21oi_1 _26381_ (.A1(_07324_),
    .A2(_07327_),
    .Y(_07330_),
    .B1(net936));
 sg13g2_buf_1 _26382_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07331_));
 sg13g2_nor2_1 _26383_ (.A(_07331_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07332_));
 sg13g2_nand2_1 _26384_ (.Y(_07333_),
    .A(_09869_),
    .B(_07332_));
 sg13g2_buf_1 _26385_ (.A(_07333_),
    .X(_07334_));
 sg13g2_nor2_1 _26386_ (.A(net938),
    .B(_07334_),
    .Y(_07335_));
 sg13g2_nand2_1 _26387_ (.Y(_07336_),
    .A(_07314_),
    .B(_07319_));
 sg13g2_inv_1 _26388_ (.Y(_07337_),
    .A(_07316_));
 sg13g2_nand2_1 _26389_ (.Y(_07338_),
    .A(net938),
    .B(_07334_));
 sg13g2_nand2_1 _26390_ (.Y(_07339_),
    .A(_07337_),
    .B(_07338_));
 sg13g2_a21oi_1 _26391_ (.A1(_07336_),
    .A2(_07339_),
    .Y(_07340_),
    .B1(net936));
 sg13g2_o21ai_1 _26392_ (.B1(net919),
    .Y(_07341_),
    .A1(_07335_),
    .A2(_07340_));
 sg13g2_nor2_1 _26393_ (.A(_07330_),
    .B(_07341_),
    .Y(_07342_));
 sg13g2_buf_2 _26394_ (.A(_07342_),
    .X(_07343_));
 sg13g2_buf_1 _26395_ (.A(_07343_),
    .X(_07344_));
 sg13g2_nor2_1 _26396_ (.A(net1083),
    .B(net936),
    .Y(_07345_));
 sg13g2_xnor2_1 _26397_ (.Y(_07346_),
    .A(net938),
    .B(_07345_));
 sg13g2_buf_1 _26398_ (.A(_07346_),
    .X(_07347_));
 sg13g2_buf_1 _26399_ (.A(_07347_),
    .X(_07348_));
 sg13g2_nor2b_1 _26400_ (.A(_07347_),
    .B_N(_09988_),
    .Y(_07349_));
 sg13g2_a21oi_1 _26401_ (.A1(\cpu.uart.r_out[1] ),
    .A2(_07348_),
    .Y(_07350_),
    .B1(_07349_));
 sg13g2_nor2_1 _26402_ (.A(\cpu.uart.r_out[0] ),
    .B(_07344_),
    .Y(_07351_));
 sg13g2_a21oi_1 _26403_ (.A1(_07344_),
    .A2(_07350_),
    .Y(_02651_),
    .B1(_07351_));
 sg13g2_nor2b_1 _26404_ (.A(_07347_),
    .B_N(_09995_),
    .Y(_07352_));
 sg13g2_a21oi_1 _26405_ (.A1(\cpu.uart.r_out[2] ),
    .A2(net583),
    .Y(_07353_),
    .B1(_07352_));
 sg13g2_nor2_1 _26406_ (.A(\cpu.uart.r_out[1] ),
    .B(net30),
    .Y(_07354_));
 sg13g2_a21oi_1 _26407_ (.A1(net30),
    .A2(_07353_),
    .Y(_02652_),
    .B1(_07354_));
 sg13g2_nor2b_1 _26408_ (.A(_07347_),
    .B_N(net1045),
    .Y(_07355_));
 sg13g2_a21oi_1 _26409_ (.A1(\cpu.uart.r_out[3] ),
    .A2(_07348_),
    .Y(_07356_),
    .B1(_07355_));
 sg13g2_nor2_1 _26410_ (.A(\cpu.uart.r_out[2] ),
    .B(_07343_),
    .Y(_07357_));
 sg13g2_a21oi_1 _26411_ (.A1(net30),
    .A2(_07356_),
    .Y(_02653_),
    .B1(_07357_));
 sg13g2_nor2_1 _26412_ (.A(_11996_),
    .B(net583),
    .Y(_07358_));
 sg13g2_a21oi_1 _26413_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net583),
    .Y(_07359_),
    .B1(_07358_));
 sg13g2_nor2_1 _26414_ (.A(\cpu.uart.r_out[3] ),
    .B(_07343_),
    .Y(_07360_));
 sg13g2_a21oi_1 _26415_ (.A1(net30),
    .A2(_07359_),
    .Y(_02654_),
    .B1(_07360_));
 sg13g2_nor2b_1 _26416_ (.A(_07347_),
    .B_N(_10013_),
    .Y(_07361_));
 sg13g2_a21oi_1 _26417_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net583),
    .Y(_07362_),
    .B1(_07361_));
 sg13g2_nor2_1 _26418_ (.A(\cpu.uart.r_out[4] ),
    .B(_07343_),
    .Y(_07363_));
 sg13g2_a21oi_1 _26419_ (.A1(net30),
    .A2(_07362_),
    .Y(_02655_),
    .B1(_07363_));
 sg13g2_nor2b_1 _26420_ (.A(_07347_),
    .B_N(_10019_),
    .Y(_07364_));
 sg13g2_a21oi_1 _26421_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net583),
    .Y(_07365_),
    .B1(_07364_));
 sg13g2_nor2_1 _26422_ (.A(\cpu.uart.r_out[5] ),
    .B(_07343_),
    .Y(_07366_));
 sg13g2_a21oi_1 _26423_ (.A1(net30),
    .A2(_07365_),
    .Y(_02656_),
    .B1(_07366_));
 sg13g2_nor2_1 _26424_ (.A(_12018_),
    .B(net583),
    .Y(_07367_));
 sg13g2_a21oi_1 _26425_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net583),
    .Y(_07368_),
    .B1(_07367_));
 sg13g2_nor2_1 _26426_ (.A(\cpu.uart.r_out[6] ),
    .B(_07343_),
    .Y(_07369_));
 sg13g2_a21oi_1 _26427_ (.A1(net30),
    .A2(_07368_),
    .Y(_02657_),
    .B1(_07369_));
 sg13g2_nor2_1 _26428_ (.A(_07248_),
    .B(net583),
    .Y(_07370_));
 sg13g2_mux2_1 _26429_ (.A0(\cpu.uart.r_out[7] ),
    .A1(_07370_),
    .S(net30),
    .X(_02658_));
 sg13g2_nand2b_1 _26430_ (.Y(_07371_),
    .B(_09897_),
    .A_N(_09858_));
 sg13g2_nor3_1 _26431_ (.A(net1084),
    .B(_07302_),
    .C(net1085),
    .Y(_07372_));
 sg13g2_a22oi_1 _26432_ (.Y(_07373_),
    .B1(_07371_),
    .B2(_07372_),
    .A2(net1085),
    .A1(net1084));
 sg13g2_nor4_1 _26433_ (.A(_07305_),
    .B(\cpu.uart.r_rstate[1] ),
    .C(_07302_),
    .D(net1085),
    .Y(_07374_));
 sg13g2_a21o_1 _26434_ (.A2(_07371_),
    .A1(net1084),
    .B1(_07302_),
    .X(_07375_));
 sg13g2_a22oi_1 _26435_ (.Y(_07376_),
    .B1(_07375_),
    .B2(net1085),
    .A2(_07374_),
    .A1(_07311_));
 sg13g2_o21ai_1 _26436_ (.B1(_07376_),
    .Y(_07377_),
    .A1(_07306_),
    .A2(_07373_));
 sg13g2_nor2_1 _26437_ (.A(_07306_),
    .B(net1084),
    .Y(_07378_));
 sg13g2_nor2b_1 _26438_ (.A(net1085),
    .B_N(_07311_),
    .Y(_07379_));
 sg13g2_nand2_1 _26439_ (.Y(_07380_),
    .A(net1084),
    .B(net1085));
 sg13g2_nor2_1 _26440_ (.A(_07305_),
    .B(_07380_),
    .Y(_07381_));
 sg13g2_a21oi_1 _26441_ (.A1(_07378_),
    .A2(_07379_),
    .Y(_07382_),
    .B1(_07381_));
 sg13g2_nor3_1 _26442_ (.A(net939),
    .B(_07297_),
    .C(_07382_),
    .Y(_07383_));
 sg13g2_xor2_1 _26443_ (.B(_07304_),
    .A(_07300_),
    .X(_07384_));
 sg13g2_o21ai_1 _26444_ (.B1(net919),
    .Y(_07385_),
    .A1(_09869_),
    .A2(_07384_));
 sg13g2_nor3_1 _26445_ (.A(_07377_),
    .B(_07383_),
    .C(_07385_),
    .Y(_07386_));
 sg13g2_and2_1 _26446_ (.A(_07305_),
    .B(_07301_),
    .X(_07387_));
 sg13g2_buf_1 _26447_ (.A(_07387_),
    .X(_07388_));
 sg13g2_o21ai_1 _26448_ (.B1(net940),
    .Y(_07389_),
    .A1(net939),
    .A2(_07388_));
 sg13g2_nor2b_1 _26449_ (.A(_07374_),
    .B_N(_07389_),
    .Y(_07390_));
 sg13g2_and2_1 _26450_ (.A(_07386_),
    .B(_07390_),
    .X(_07391_));
 sg13g2_nor2_1 _26451_ (.A(_07295_),
    .B(_07386_),
    .Y(_07392_));
 sg13g2_a21oi_1 _26452_ (.A1(_07295_),
    .A2(_07391_),
    .Y(_02661_),
    .B1(_07392_));
 sg13g2_nand2_1 _26453_ (.Y(_07393_),
    .A(_07295_),
    .B(_07390_));
 sg13g2_inv_1 _26454_ (.Y(_07394_),
    .A(\cpu.uart.r_rcnt[1] ));
 sg13g2_a21oi_1 _26455_ (.A1(_07386_),
    .A2(_07393_),
    .Y(_07395_),
    .B1(_07394_));
 sg13g2_a21o_1 _26456_ (.A2(_07391_),
    .A1(_07296_),
    .B1(_07395_),
    .X(_02662_));
 sg13g2_nand2_1 _26457_ (.Y(_07396_),
    .A(\cpu.uart.r_out[0] ),
    .B(_07347_));
 sg13g2_xnor2_1 _26458_ (.Y(_07397_),
    .A(\cpu.uart.r_x_invert ),
    .B(_07396_));
 sg13g2_nor2b_1 _26459_ (.A(_07328_),
    .B_N(_07314_),
    .Y(_07398_));
 sg13g2_nand2_1 _26460_ (.Y(_07399_),
    .A(net1083),
    .B(_07398_));
 sg13g2_or2_1 _26461_ (.X(_07400_),
    .B(_07328_),
    .A(_07314_));
 sg13g2_nand2_1 _26462_ (.Y(_07401_),
    .A(_07314_),
    .B(_07328_));
 sg13g2_a21oi_1 _26463_ (.A1(_07400_),
    .A2(_07401_),
    .Y(_07402_),
    .B1(_07317_));
 sg13g2_nand2_1 _26464_ (.Y(_07403_),
    .A(_07337_),
    .B(_07402_));
 sg13g2_nand3_1 _26465_ (.B(_07399_),
    .C(_07403_),
    .A(net919),
    .Y(_07404_));
 sg13g2_mux2_1 _26466_ (.A0(_07397_),
    .A1(_00261_),
    .S(_07404_),
    .X(_07405_));
 sg13g2_buf_1 _26467_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07406_));
 sg13g2_inv_1 _26468_ (.Y(_07407_),
    .A(_07323_));
 sg13g2_nand4_1 _26469_ (.B(net937),
    .C(_07407_),
    .A(net1083),
    .Y(_07408_),
    .D(_07398_));
 sg13g2_buf_1 _26470_ (.A(_07408_),
    .X(_07409_));
 sg13g2_nor2_1 _26471_ (.A(_07371_),
    .B(_07400_),
    .Y(_07410_));
 sg13g2_o21ai_1 _26472_ (.B1(_07337_),
    .Y(_07411_),
    .A1(_07402_),
    .A2(_07410_));
 sg13g2_a21oi_1 _26473_ (.A1(_07334_),
    .A2(_07336_),
    .Y(_07412_),
    .B1(_07328_));
 sg13g2_nor2_1 _26474_ (.A(_07335_),
    .B(_07412_),
    .Y(_07413_));
 sg13g2_nand2_1 _26475_ (.Y(_07414_),
    .A(_07411_),
    .B(_07413_));
 sg13g2_a21oi_1 _26476_ (.A1(_07409_),
    .A2(_07414_),
    .Y(_07415_),
    .B1(net798));
 sg13g2_mux2_1 _26477_ (.A0(_07405_),
    .A1(_07406_),
    .S(_07415_),
    .X(_02667_));
 sg13g2_a21oi_1 _26478_ (.A1(net937),
    .A2(_07332_),
    .Y(_07416_),
    .B1(_07328_));
 sg13g2_o21ai_1 _26479_ (.B1(net936),
    .Y(_07417_),
    .A1(net937),
    .A2(_07332_));
 sg13g2_o21ai_1 _26480_ (.B1(_07417_),
    .Y(_07418_),
    .A1(_07337_),
    .A2(_07416_));
 sg13g2_nand2_1 _26481_ (.Y(_07419_),
    .A(net938),
    .B(_07418_));
 sg13g2_nor4_2 _26482_ (.A(net1083),
    .B(net937),
    .C(net938),
    .Y(_07420_),
    .D(net936));
 sg13g2_nor2_1 _26483_ (.A(net1053),
    .B(_07420_),
    .Y(_07421_));
 sg13g2_and4_1 _26484_ (.A(_09869_),
    .B(_07409_),
    .C(_07419_),
    .D(_07421_),
    .X(_07422_));
 sg13g2_buf_1 _26485_ (.A(_07422_),
    .X(_07423_));
 sg13g2_inv_1 _26486_ (.Y(_07424_),
    .A(_07328_));
 sg13g2_nor2_1 _26487_ (.A(net1083),
    .B(net937),
    .Y(_07425_));
 sg13g2_nor2_1 _26488_ (.A(_07401_),
    .B(_07425_),
    .Y(_07426_));
 sg13g2_a21oi_1 _26489_ (.A1(_07424_),
    .A2(_07326_),
    .Y(_07427_),
    .B1(_07426_));
 sg13g2_nand2_1 _26490_ (.Y(_07428_),
    .A(_07423_),
    .B(_07427_));
 sg13g2_nor2b_1 _26491_ (.A(_07331_),
    .B_N(_07423_),
    .Y(_07429_));
 sg13g2_a21oi_1 _26492_ (.A1(_07331_),
    .A2(_07428_),
    .Y(_07430_),
    .B1(_07429_));
 sg13g2_inv_1 _26493_ (.Y(_02670_),
    .A(_07430_));
 sg13g2_nand2_1 _26494_ (.Y(_07431_),
    .A(_07331_),
    .B(_07427_));
 sg13g2_nand2_1 _26495_ (.Y(_07432_),
    .A(_07423_),
    .B(_07431_));
 sg13g2_o21ai_1 _26496_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07433_),
    .A1(_07331_),
    .A2(_07428_));
 sg13g2_o21ai_1 _26497_ (.B1(_07433_),
    .Y(_02671_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07432_));
 sg13g2_nor3_1 _26498_ (.A(_09168_),
    .B(_10042_),
    .C(net692),
    .Y(_07434_));
 sg13g2_buf_1 _26499_ (.A(_07434_),
    .X(_07435_));
 sg13g2_buf_1 _26500_ (.A(net153),
    .X(_07436_));
 sg13g2_nand2_1 _26501_ (.Y(_07437_),
    .A(_10114_),
    .B(_10116_));
 sg13g2_nand3_1 _26502_ (.B(_10126_),
    .C(_10131_),
    .A(_10120_),
    .Y(_07438_));
 sg13g2_buf_1 _26503_ (.A(_07438_),
    .X(_07439_));
 sg13g2_nor2_1 _26504_ (.A(_07437_),
    .B(_07439_),
    .Y(_07440_));
 sg13g2_nand2_1 _26505_ (.Y(_07441_),
    .A(_10038_),
    .B(_10045_));
 sg13g2_buf_1 _26506_ (.A(_07441_),
    .X(_07442_));
 sg13g2_o21ai_1 _26507_ (.B1(net110),
    .Y(_07443_),
    .A1(net126),
    .A2(_07440_));
 sg13g2_nand2_1 _26508_ (.Y(_07444_),
    .A(_04897_),
    .B(_07443_));
 sg13g2_and2_1 _26509_ (.A(_10038_),
    .B(net387),
    .X(_07445_));
 sg13g2_buf_1 _26510_ (.A(_07445_),
    .X(_07446_));
 sg13g2_buf_1 _26511_ (.A(_07446_),
    .X(_07447_));
 sg13g2_nor3_1 _26512_ (.A(_04897_),
    .B(_07437_),
    .C(_07439_),
    .Y(_07448_));
 sg13g2_a22oi_1 _26513_ (.Y(_07449_),
    .B1(_07448_),
    .B2(net98),
    .A2(net89),
    .A1(net1047));
 sg13g2_nand2_1 _26514_ (.Y(_02457_),
    .A(_07444_),
    .B(_07449_));
 sg13g2_and2_1 _26515_ (.A(_04897_),
    .B(_07440_),
    .X(_07450_));
 sg13g2_buf_1 _26516_ (.A(_07450_),
    .X(_07451_));
 sg13g2_o21ai_1 _26517_ (.B1(net110),
    .Y(_07452_),
    .A1(net126),
    .A2(_07451_));
 sg13g2_nand2_1 _26518_ (.Y(_07453_),
    .A(_05295_),
    .B(_07452_));
 sg13g2_nor2b_1 _26519_ (.A(_05295_),
    .B_N(_07451_),
    .Y(_07454_));
 sg13g2_a22oi_1 _26520_ (.Y(_07455_),
    .B1(_07454_),
    .B2(net98),
    .A2(_07447_),
    .A1(net1046));
 sg13g2_nand2_1 _26521_ (.Y(_02458_),
    .A(_07453_),
    .B(_07455_));
 sg13g2_and2_1 _26522_ (.A(_05295_),
    .B(_07451_),
    .X(_07456_));
 sg13g2_buf_1 _26523_ (.A(_07456_),
    .X(_07457_));
 sg13g2_o21ai_1 _26524_ (.B1(_07442_),
    .Y(_07458_),
    .A1(_07436_),
    .A2(_07457_));
 sg13g2_nand2_1 _26525_ (.Y(_07459_),
    .A(_05366_),
    .B(_07458_));
 sg13g2_nor2b_1 _26526_ (.A(_05366_),
    .B_N(_07457_),
    .Y(_07460_));
 sg13g2_a22oi_1 _26527_ (.Y(_07461_),
    .B1(_07460_),
    .B2(_10111_),
    .A2(net89),
    .A1(net1045));
 sg13g2_nand2_1 _26528_ (.Y(_02459_),
    .A(_07459_),
    .B(_07461_));
 sg13g2_nand3_1 _26529_ (.B(_05295_),
    .C(_05366_),
    .A(_04897_),
    .Y(_07462_));
 sg13g2_or3_1 _26530_ (.A(_10122_),
    .B(_07439_),
    .C(_07462_),
    .X(_07463_));
 sg13g2_buf_1 _26531_ (.A(_07463_),
    .X(_07464_));
 sg13g2_a21oi_1 _26532_ (.A1(_10040_),
    .A2(_07464_),
    .Y(_07465_),
    .B1(net99));
 sg13g2_nand2b_1 _26533_ (.Y(_07466_),
    .B(_07465_),
    .A_N(_05411_));
 sg13g2_o21ai_1 _26534_ (.B1(_05411_),
    .Y(_07467_),
    .A1(net126),
    .A2(_07464_));
 sg13g2_a22oi_1 _26535_ (.Y(_02460_),
    .B1(_07466_),
    .B2(_07467_),
    .A2(net89),
    .A1(net866));
 sg13g2_and3_1 _26536_ (.X(_07468_),
    .A(_05366_),
    .B(_05411_),
    .C(_07457_));
 sg13g2_buf_1 _26537_ (.A(_07468_),
    .X(_07469_));
 sg13g2_o21ai_1 _26538_ (.B1(net110),
    .Y(_07470_),
    .A1(net153),
    .A2(_07469_));
 sg13g2_nand2_1 _26539_ (.Y(_07471_),
    .A(net119),
    .B(_07469_));
 sg13g2_nor2_1 _26540_ (.A(_05477_),
    .B(_07471_),
    .Y(_07472_));
 sg13g2_a221oi_1 _26541_ (.B2(_05477_),
    .C1(_07472_),
    .B1(_07470_),
    .A1(net1043),
    .Y(_07473_),
    .A2(_07446_));
 sg13g2_inv_1 _26542_ (.Y(_02461_),
    .A(_07473_));
 sg13g2_nand2_1 _26543_ (.Y(_07474_),
    .A(_05411_),
    .B(_05477_));
 sg13g2_nor2_1 _26544_ (.A(_07464_),
    .B(_07474_),
    .Y(_07475_));
 sg13g2_nor2_1 _26545_ (.A(_07436_),
    .B(_07475_),
    .Y(_07476_));
 sg13g2_o21ai_1 _26546_ (.B1(_05526_),
    .Y(_07477_),
    .A1(_10100_),
    .A2(_07476_));
 sg13g2_nor3_1 _26547_ (.A(_05526_),
    .B(_07464_),
    .C(_07474_),
    .Y(_07478_));
 sg13g2_a22oi_1 _26548_ (.Y(_07479_),
    .B1(_07478_),
    .B2(_10111_),
    .A2(_07447_),
    .A1(net1042));
 sg13g2_nand2_1 _26549_ (.Y(_02462_),
    .A(_07477_),
    .B(_07479_));
 sg13g2_nand3_1 _26550_ (.B(_05526_),
    .C(_07469_),
    .A(_05477_),
    .Y(_07480_));
 sg13g2_buf_1 _26551_ (.A(_07480_),
    .X(_07481_));
 sg13g2_a21oi_1 _26552_ (.A1(_10040_),
    .A2(_07481_),
    .Y(_07482_),
    .B1(_10047_));
 sg13g2_nand2b_1 _26553_ (.Y(_07483_),
    .B(_07482_),
    .A_N(_05615_));
 sg13g2_o21ai_1 _26554_ (.B1(_05615_),
    .Y(_07484_),
    .A1(net126),
    .A2(_07481_));
 sg13g2_a22oi_1 _26555_ (.Y(_02463_),
    .B1(_07483_),
    .B2(_07484_),
    .A2(net89),
    .A1(_12645_));
 sg13g2_nand3_1 _26556_ (.B(_05615_),
    .C(_07475_),
    .A(_05526_),
    .Y(_07485_));
 sg13g2_buf_1 _26557_ (.A(_07485_),
    .X(_07486_));
 sg13g2_a21oi_1 _26558_ (.A1(net119),
    .A2(_07486_),
    .Y(_07487_),
    .B1(_10047_));
 sg13g2_nand2b_1 _26559_ (.Y(_07488_),
    .B(_07487_),
    .A_N(_05008_));
 sg13g2_o21ai_1 _26560_ (.B1(_05008_),
    .Y(_07489_),
    .A1(net126),
    .A2(_07486_));
 sg13g2_a22oi_1 _26561_ (.Y(_02464_),
    .B1(_07488_),
    .B2(_07489_),
    .A2(net89),
    .A1(net752));
 sg13g2_nand2_1 _26562_ (.Y(_07490_),
    .A(_05615_),
    .B(_05008_));
 sg13g2_nor2_1 _26563_ (.A(_07481_),
    .B(_07490_),
    .Y(_07491_));
 sg13g2_o21ai_1 _26564_ (.B1(net110),
    .Y(_07492_),
    .A1(net153),
    .A2(_07491_));
 sg13g2_inv_1 _26565_ (.Y(_07493_),
    .A(_07491_));
 sg13g2_nor3_1 _26566_ (.A(_05665_),
    .B(net153),
    .C(_07493_),
    .Y(_07494_));
 sg13g2_a221oi_1 _26567_ (.B2(_05665_),
    .C1(_07494_),
    .B1(_07492_),
    .A1(_10087_),
    .Y(_07495_),
    .A2(_07446_));
 sg13g2_inv_1 _26568_ (.Y(_02465_),
    .A(_07495_));
 sg13g2_and2_1 _26569_ (.A(_05665_),
    .B(_07491_),
    .X(_07496_));
 sg13g2_buf_1 _26570_ (.A(_07496_),
    .X(_07497_));
 sg13g2_o21ai_1 _26571_ (.B1(net110),
    .Y(_07498_),
    .A1(net126),
    .A2(_07497_));
 sg13g2_nand2_1 _26572_ (.Y(_07499_),
    .A(_05676_),
    .B(_07498_));
 sg13g2_nor2b_1 _26573_ (.A(_05676_),
    .B_N(_07497_),
    .Y(_07500_));
 sg13g2_a22oi_1 _26574_ (.Y(_07501_),
    .B1(_07500_),
    .B2(net98),
    .A2(net89),
    .A1(_10094_));
 sg13g2_nand2_1 _26575_ (.Y(_02466_),
    .A(_07499_),
    .B(_07501_));
 sg13g2_inv_1 _26576_ (.Y(_07502_),
    .A(_04983_));
 sg13g2_nand2_1 _26577_ (.Y(_07503_),
    .A(_05676_),
    .B(_07497_));
 sg13g2_a21oi_1 _26578_ (.A1(net119),
    .A2(_07503_),
    .Y(_07504_),
    .B1(net99));
 sg13g2_nor3_1 _26579_ (.A(_04983_),
    .B(net153),
    .C(_07503_),
    .Y(_07505_));
 sg13g2_a21oi_1 _26580_ (.A1(_10099_),
    .A2(_07446_),
    .Y(_07506_),
    .B1(_07505_));
 sg13g2_o21ai_1 _26581_ (.B1(_07506_),
    .Y(_02467_),
    .A1(_07502_),
    .A2(_07504_));
 sg13g2_nand4_1 _26582_ (.B(_05665_),
    .C(_05676_),
    .A(_05008_),
    .Y(_07507_),
    .D(_04983_));
 sg13g2_nor2_1 _26583_ (.A(_07486_),
    .B(_07507_),
    .Y(_07508_));
 sg13g2_o21ai_1 _26584_ (.B1(net110),
    .Y(_07509_),
    .A1(net153),
    .A2(_07508_));
 sg13g2_nor4_1 _26585_ (.A(_05105_),
    .B(net153),
    .C(_07486_),
    .D(_07507_),
    .Y(_07510_));
 sg13g2_a221oi_1 _26586_ (.B2(_05105_),
    .C1(_07510_),
    .B1(_07509_),
    .A1(_10105_),
    .Y(_07511_),
    .A2(_07446_));
 sg13g2_inv_1 _26587_ (.Y(_02468_),
    .A(_07511_));
 sg13g2_nand4_1 _26588_ (.B(_05676_),
    .C(_04983_),
    .A(_05665_),
    .Y(_07512_),
    .D(_05105_));
 sg13g2_nor2_1 _26589_ (.A(_07493_),
    .B(_07512_),
    .Y(_07513_));
 sg13g2_o21ai_1 _26590_ (.B1(net110),
    .Y(_07514_),
    .A1(net126),
    .A2(_07513_));
 sg13g2_nand2_1 _26591_ (.Y(_07515_),
    .A(_05133_),
    .B(_07514_));
 sg13g2_nor3_1 _26592_ (.A(_05133_),
    .B(_07493_),
    .C(_07512_),
    .Y(_07516_));
 sg13g2_a22oi_1 _26593_ (.Y(_07517_),
    .B1(_07516_),
    .B2(net119),
    .A2(net89),
    .A1(_10113_));
 sg13g2_nand2_1 _26594_ (.Y(_02469_),
    .A(_07515_),
    .B(_07517_));
 sg13g2_and3_1 _26595_ (.X(_07518_),
    .A(_05105_),
    .B(_05133_),
    .C(_07508_));
 sg13g2_buf_1 _26596_ (.A(_07518_),
    .X(_07519_));
 sg13g2_o21ai_1 _26597_ (.B1(net110),
    .Y(_07520_),
    .A1(net153),
    .A2(_07519_));
 sg13g2_nand2_1 _26598_ (.Y(_07521_),
    .A(_10039_),
    .B(_07519_));
 sg13g2_nor2_1 _26599_ (.A(_05158_),
    .B(_07521_),
    .Y(_07522_));
 sg13g2_a221oi_1 _26600_ (.B2(_05158_),
    .C1(_07522_),
    .B1(_07520_),
    .A1(_10119_),
    .Y(_07523_),
    .A2(_07446_));
 sg13g2_inv_1 _26601_ (.Y(_02470_),
    .A(_07523_));
 sg13g2_inv_1 _26602_ (.Y(_07524_),
    .A(_05184_));
 sg13g2_nand3_1 _26603_ (.B(_05158_),
    .C(_07513_),
    .A(_05133_),
    .Y(_07525_));
 sg13g2_a21oi_1 _26604_ (.A1(net119),
    .A2(_07525_),
    .Y(_07526_),
    .B1(_10100_));
 sg13g2_nor2_1 _26605_ (.A(net126),
    .B(_07525_),
    .Y(_07527_));
 sg13g2_a22oi_1 _26606_ (.Y(_07528_),
    .B1(_07527_),
    .B2(_07524_),
    .A2(_07446_),
    .A1(_10125_));
 sg13g2_o21ai_1 _26607_ (.B1(_07528_),
    .Y(_02471_),
    .A1(_07524_),
    .A2(_07526_));
 sg13g2_nand3_1 _26608_ (.B(_05184_),
    .C(_07519_),
    .A(_05158_),
    .Y(_07529_));
 sg13g2_inv_1 _26609_ (.Y(_07530_),
    .A(\cpu.intr.r_clock_count[31] ));
 sg13g2_a221oi_1 _26610_ (.B2(_10039_),
    .C1(_07530_),
    .B1(_07529_),
    .A1(net128),
    .Y(_07531_),
    .A2(net447));
 sg13g2_o21ai_1 _26611_ (.B1(_07530_),
    .Y(_07532_),
    .A1(_07435_),
    .A2(_07529_));
 sg13g2_nor2b_1 _26612_ (.A(_07531_),
    .B_N(_07532_),
    .Y(_07533_));
 sg13g2_a21o_1 _26613_ (.A2(net89),
    .A1(_10130_),
    .B1(_07533_),
    .X(_02472_));
 sg13g2_buf_1 _26614_ (.A(net798),
    .X(_07534_));
 sg13g2_nor2_1 _26615_ (.A(\cpu.r_clk_invert ),
    .B(net796),
    .Y(_07535_));
 sg13g2_a21oi_1 _26616_ (.A1(_09109_),
    .A2(_07534_),
    .Y(_02539_),
    .B1(_07535_));
 sg13g2_nand2b_1 _26617_ (.Y(_07536_),
    .B(net919),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26618_ (.A(_07536_),
    .X(_07537_));
 sg13g2_nor2b_1 _26619_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net400),
    .Y(_07538_));
 sg13g2_nand4_1 _26620_ (.B(_02878_),
    .C(_11980_),
    .A(_09281_),
    .Y(_07539_),
    .D(_11887_));
 sg13g2_buf_2 _26621_ (.A(_07539_),
    .X(_07540_));
 sg13g2_nor2_1 _26622_ (.A(net567),
    .B(_07540_),
    .Y(_07541_));
 sg13g2_nor3_1 _26623_ (.A(_07537_),
    .B(_07538_),
    .C(_07541_),
    .Y(_00737_));
 sg13g2_nor2_1 _26624_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net399),
    .Y(_07542_));
 sg13g2_nor2_1 _26625_ (.A(net490),
    .B(_07540_),
    .Y(_07543_));
 sg13g2_nor3_1 _26626_ (.A(_07537_),
    .B(_07542_),
    .C(_07543_),
    .Y(_00738_));
 sg13g2_nor2_1 _26627_ (.A(\cpu.dcache.r_valid[2] ),
    .B(_12300_),
    .Y(_07544_));
 sg13g2_nor2_1 _26628_ (.A(net678),
    .B(_07540_),
    .Y(_07545_));
 sg13g2_nor3_1 _26629_ (.A(_07537_),
    .B(_07544_),
    .C(_07545_),
    .Y(_00739_));
 sg13g2_nor2_1 _26630_ (.A(\cpu.dcache.r_valid[3] ),
    .B(_02961_),
    .Y(_07546_));
 sg13g2_nor2_1 _26631_ (.A(net566),
    .B(_07540_),
    .Y(_07547_));
 sg13g2_nor3_1 _26632_ (.A(_07537_),
    .B(_07546_),
    .C(_07547_),
    .Y(_00740_));
 sg13g2_inv_1 _26633_ (.Y(_07548_),
    .A(\cpu.dcache.r_valid[4] ));
 sg13g2_inv_1 _26634_ (.Y(_07549_),
    .A(_07540_));
 sg13g2_a221oi_1 _26635_ (.B2(_10036_),
    .C1(_07537_),
    .B1(_07549_),
    .A1(_07548_),
    .Y(_00741_),
    .A2(net396));
 sg13g2_nor2_1 _26636_ (.A(\cpu.dcache.r_valid[5] ),
    .B(_12655_),
    .Y(_07550_));
 sg13g2_nor2_1 _26637_ (.A(net754),
    .B(_07540_),
    .Y(_07551_));
 sg13g2_nor3_1 _26638_ (.A(_07537_),
    .B(_07550_),
    .C(_07551_),
    .Y(_00742_));
 sg13g2_nor2_1 _26639_ (.A(\cpu.dcache.r_valid[6] ),
    .B(_02712_),
    .Y(_07552_));
 sg13g2_nor2_1 _26640_ (.A(net677),
    .B(_07540_),
    .Y(_07553_));
 sg13g2_nor3_1 _26641_ (.A(_07537_),
    .B(_07552_),
    .C(_07553_),
    .Y(_00743_));
 sg13g2_nor2_1 _26642_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net393),
    .Y(_07554_));
 sg13g2_nor2_1 _26643_ (.A(net485),
    .B(_07540_),
    .Y(_07555_));
 sg13g2_nor3_1 _26644_ (.A(_07537_),
    .B(_07554_),
    .C(_07555_),
    .Y(_00744_));
 sg13g2_nand3_1 _26645_ (.B(_10162_),
    .C(_04700_),
    .A(_11375_),
    .Y(_07556_));
 sg13g2_buf_1 _26646_ (.A(_07556_),
    .X(_07557_));
 sg13g2_nand2_1 _26647_ (.Y(_07558_),
    .A(_08285_),
    .B(net518));
 sg13g2_o21ai_1 _26648_ (.B1(_07558_),
    .Y(_07559_),
    .A1(net599),
    .A2(net518));
 sg13g2_and3_1 _26649_ (.X(_00791_),
    .A(_04401_),
    .B(_11776_),
    .C(_07559_));
 sg13g2_and4_1 _26650_ (.A(_03424_),
    .B(_10550_),
    .C(\cpu.dec.do_flush_all ),
    .D(_09265_),
    .X(_00923_));
 sg13g2_and4_1 _26651_ (.A(_03424_),
    .B(_10597_),
    .C(\cpu.dec.do_flush_all ),
    .D(net710),
    .X(_00941_));
 sg13g2_nor2_1 _26652_ (.A(_11395_),
    .B(_11160_),
    .Y(_07560_));
 sg13g2_nand2_1 _26653_ (.Y(_07561_),
    .A(_06825_),
    .B(_11395_));
 sg13g2_o21ai_1 _26654_ (.B1(_07561_),
    .Y(_07562_),
    .A1(net288),
    .A2(_07560_));
 sg13g2_nand4_1 _26655_ (.B(_03830_),
    .C(net710),
    .A(net982),
    .Y(_07563_),
    .D(net621));
 sg13g2_mux2_1 _26656_ (.A0(_10586_),
    .A1(_09133_),
    .S(_07563_),
    .X(_07564_));
 sg13g2_nand2_1 _26657_ (.Y(_07565_),
    .A(net518),
    .B(_07564_));
 sg13g2_o21ai_1 _26658_ (.B1(_07565_),
    .Y(_07566_),
    .A1(_03552_),
    .A2(net518));
 sg13g2_and3_1 _26659_ (.X(_00942_),
    .A(_11776_),
    .B(_07562_),
    .C(_07566_));
 sg13g2_nand2_1 _26660_ (.Y(_07567_),
    .A(_08339_),
    .B(net710));
 sg13g2_or2_1 _26661_ (.X(_07568_),
    .B(_07567_),
    .A(_00294_));
 sg13g2_a21o_1 _26662_ (.A2(_04957_),
    .A1(net854),
    .B1(_07568_),
    .X(_07569_));
 sg13g2_nand3b_1 _26663_ (.B(_09769_),
    .C(net919),
    .Y(_07570_),
    .A_N(_11889_));
 sg13g2_a21oi_1 _26664_ (.A1(_09773_),
    .A2(_07570_),
    .Y(_07571_),
    .B1(_08339_));
 sg13g2_nand2b_1 _26665_ (.Y(_07572_),
    .B(net802),
    .A_N(_07571_));
 sg13g2_a21oi_1 _26666_ (.A1(_08326_),
    .A2(_07569_),
    .Y(_01060_),
    .B1(_07572_));
 sg13g2_nor2_1 _26667_ (.A(_00294_),
    .B(_07567_),
    .Y(_07573_));
 sg13g2_o21ai_1 _26668_ (.B1(_07573_),
    .Y(_07574_),
    .A1(_11784_),
    .A2(_04957_));
 sg13g2_a21oi_1 _26669_ (.A1(_08324_),
    .A2(_07574_),
    .Y(_01061_),
    .B1(_07572_));
 sg13g2_inv_1 _26670_ (.Y(_07575_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26671_ (.Y(_07576_),
    .B(_09082_),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26672_ (.A(_07576_),
    .X(_07577_));
 sg13g2_a21oi_1 _26673_ (.A1(_07575_),
    .A2(net366),
    .Y(_02416_),
    .B1(_07577_));
 sg13g2_nor2_1 _26674_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06486_),
    .Y(_07578_));
 sg13g2_nor2_1 _26675_ (.A(_07577_),
    .B(_07578_),
    .Y(_02417_));
 sg13g2_nor2_1 _26676_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06505_),
    .Y(_07579_));
 sg13g2_nor2_1 _26677_ (.A(_07577_),
    .B(_07579_),
    .Y(_02418_));
 sg13g2_inv_1 _26678_ (.Y(_07580_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26679_ (.A1(_07580_),
    .A2(net245),
    .Y(_02419_),
    .B1(_07577_));
 sg13g2_nor2_1 _26680_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06530_),
    .Y(_07581_));
 sg13g2_nor2_1 _26681_ (.A(_07577_),
    .B(_07581_),
    .Y(_02420_));
 sg13g2_nor2_1 _26682_ (.A(\cpu.icache.r_valid[5] ),
    .B(_06545_),
    .Y(_07582_));
 sg13g2_nor2_1 _26683_ (.A(_07577_),
    .B(_07582_),
    .Y(_02421_));
 sg13g2_nor2_1 _26684_ (.A(\cpu.icache.r_valid[6] ),
    .B(_06560_),
    .Y(_07583_));
 sg13g2_nor2_1 _26685_ (.A(_07577_),
    .B(_07583_),
    .Y(_02422_));
 sg13g2_nor2_1 _26686_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06571_),
    .Y(_07584_));
 sg13g2_nor2_1 _26687_ (.A(_07577_),
    .B(_07584_),
    .Y(_02423_));
 sg13g2_nand3_1 _26688_ (.B(net128),
    .C(_04918_),
    .A(net1044),
    .Y(_07585_));
 sg13g2_nand2_1 _26689_ (.Y(_07586_),
    .A(_09120_),
    .B(_07585_));
 sg13g2_nand3_1 _26690_ (.B(net128),
    .C(_05285_),
    .A(_10008_),
    .Y(_07587_));
 sg13g2_a21oi_1 _26691_ (.A1(_07586_),
    .A2(_07587_),
    .Y(_00313_),
    .B1(net657));
 sg13g2_nor2_1 _26692_ (.A(_02878_),
    .B(_11907_),
    .Y(_07588_));
 sg13g2_nor2b_1 _26693_ (.A(_07588_),
    .B_N(_00311_),
    .Y(_00582_));
 sg13g2_nor2_1 _26694_ (.A(_11911_),
    .B(_11948_),
    .Y(_07589_));
 sg13g2_nor2_1 _26695_ (.A(_07588_),
    .B(_07589_),
    .Y(_00583_));
 sg13g2_xnor2_1 _26696_ (.Y(_07590_),
    .A(_06864_),
    .B(_11887_));
 sg13g2_nor2_1 _26697_ (.A(_07588_),
    .B(_07590_),
    .Y(_00584_));
 sg13g2_nor2_1 _26698_ (.A(_11879_),
    .B(net518),
    .Y(_07591_));
 sg13g2_a21oi_1 _26699_ (.A1(net1070),
    .A2(net518),
    .Y(_07592_),
    .B1(_07591_));
 sg13g2_nor2_1 _26700_ (.A(net711),
    .B(_07592_),
    .Y(_00792_));
 sg13g2_a22oi_1 _26701_ (.Y(_07593_),
    .B1(net352),
    .B2(_11396_),
    .A2(net288),
    .A1(_06818_));
 sg13g2_buf_1 _26702_ (.A(_07593_),
    .X(_07594_));
 sg13g2_or2_1 _26703_ (.X(_07595_),
    .B(_07594_),
    .A(net819));
 sg13g2_nand4_1 _26704_ (.B(_03830_),
    .C(_11393_),
    .A(_11164_),
    .Y(_07596_),
    .D(net621));
 sg13g2_a21oi_1 _26705_ (.A1(net982),
    .A2(_07596_),
    .Y(_07597_),
    .B1(_09230_));
 sg13g2_nor2_1 _26706_ (.A(_03522_),
    .B(_07597_),
    .Y(_07598_));
 sg13g2_nor2_1 _26707_ (.A(_10561_),
    .B(_07598_),
    .Y(_07599_));
 sg13g2_a21oi_1 _26708_ (.A1(_03552_),
    .A2(_07598_),
    .Y(_07600_),
    .B1(_07599_));
 sg13g2_nand2_1 _26709_ (.Y(_07601_),
    .A(_07594_),
    .B(_07600_));
 sg13g2_nand3_1 _26710_ (.B(_07595_),
    .C(_07601_),
    .A(_09084_),
    .Y(_00793_));
 sg13g2_nand2_1 _26711_ (.Y(_07602_),
    .A(_10458_),
    .B(net518));
 sg13g2_o21ai_1 _26712_ (.B1(_07602_),
    .Y(_07603_),
    .A1(net864),
    .A2(net518));
 sg13g2_and2_1 _26713_ (.A(net682),
    .B(_07603_),
    .X(_00794_));
 sg13g2_nor4_1 _26714_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11385_),
    .C(_03416_),
    .D(_07567_),
    .Y(_07604_));
 sg13g2_nor3_1 _26715_ (.A(_11381_),
    .B(_07571_),
    .C(_07604_),
    .Y(_07605_));
 sg13g2_nor4_1 _26716_ (.A(_09146_),
    .B(\cpu.ex.c_div_running ),
    .C(\cpu.ex.c_mult_running ),
    .D(_07605_),
    .Y(_07606_));
 sg13g2_nor3_1 _26717_ (.A(_06818_),
    .B(_04750_),
    .C(_07606_),
    .Y(_07607_));
 sg13g2_nor2_1 _26718_ (.A(_06825_),
    .B(_09837_),
    .Y(_07608_));
 sg13g2_o21ai_1 _26719_ (.B1(_09830_),
    .Y(_00939_),
    .A1(_07607_),
    .A2(_07608_));
 sg13g2_nand2_1 _26720_ (.Y(_07609_),
    .A(_09281_),
    .B(_09263_));
 sg13g2_nand3_1 _26721_ (.B(\cpu.dec.do_flush_write ),
    .C(_11393_),
    .A(net982),
    .Y(_07610_));
 sg13g2_a21oi_1 _26722_ (.A1(_07609_),
    .A2(_07610_),
    .Y(_00940_),
    .B1(net657));
 sg13g2_nand2_1 _26723_ (.Y(_07611_),
    .A(\cpu.dec.io ),
    .B(_11393_));
 sg13g2_nand2_1 _26724_ (.Y(_07612_),
    .A(_02877_),
    .B(_09263_));
 sg13g2_a21oi_1 _26725_ (.A1(_07611_),
    .A2(_07612_),
    .Y(_00943_),
    .B1(net657));
 sg13g2_nor2_1 _26726_ (.A(net601),
    .B(_07557_),
    .Y(_07613_));
 sg13g2_a21oi_1 _26727_ (.A1(_10586_),
    .A2(_07557_),
    .Y(_07614_),
    .B1(_07613_));
 sg13g2_nand2_1 _26728_ (.Y(_07615_),
    .A(_07594_),
    .B(_07614_));
 sg13g2_o21ai_1 _26729_ (.B1(_07615_),
    .Y(_07616_),
    .A1(_09133_),
    .A2(_07594_));
 sg13g2_nor2_1 _26730_ (.A(_09254_),
    .B(_07616_),
    .Y(_00990_));
 sg13g2_a22oi_1 _26731_ (.Y(_07617_),
    .B1(_11410_),
    .B2(net1132),
    .A2(_11393_),
    .A1(_11385_));
 sg13g2_nor2_1 _26732_ (.A(_09254_),
    .B(_07617_),
    .Y(_00991_));
 sg13g2_nor2_2 _26733_ (.A(net981),
    .B(_05741_),
    .Y(_07618_));
 sg13g2_mux2_1 _26734_ (.A0(_10505_),
    .A1(net507),
    .S(_07618_),
    .X(_07619_));
 sg13g2_nand2_1 _26735_ (.Y(_07620_),
    .A(_04401_),
    .B(_07619_));
 sg13g2_a21oi_1 _26736_ (.A1(_11386_),
    .A2(_07620_),
    .Y(_01066_),
    .B1(_06800_));
 sg13g2_buf_1 _26737_ (.A(_09253_),
    .X(_07621_));
 sg13g2_nand2_1 _26738_ (.Y(_07622_),
    .A(_09243_),
    .B(_07618_));
 sg13g2_o21ai_1 _26739_ (.B1(_07622_),
    .Y(_07623_),
    .A1(_05796_),
    .A2(_07618_));
 sg13g2_nor2_1 _26740_ (.A(net707),
    .B(net391),
    .Y(_07624_));
 sg13g2_a21oi_1 _26741_ (.A1(net391),
    .A2(_07623_),
    .Y(_07625_),
    .B1(_07624_));
 sg13g2_nor2_1 _26742_ (.A(_07621_),
    .B(_07625_),
    .Y(_01067_));
 sg13g2_mux2_1 _26743_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_03472_),
    .S(_07618_),
    .X(_07626_));
 sg13g2_nand2b_1 _26744_ (.Y(_07627_),
    .B(_07626_),
    .A_N(_08330_));
 sg13g2_a21oi_1 _26745_ (.A1(net459),
    .A2(_07627_),
    .Y(_01068_),
    .B1(_06800_));
 sg13g2_nor2_1 _26746_ (.A(net1113),
    .B(_10676_),
    .Y(_07628_));
 sg13g2_nor2_1 _26747_ (.A(_10401_),
    .B(net968),
    .Y(_07629_));
 sg13g2_nand2_1 _26748_ (.Y(_07630_),
    .A(net1086),
    .B(_07629_));
 sg13g2_nor2_1 _26749_ (.A(_10192_),
    .B(_07630_),
    .Y(_07631_));
 sg13g2_and2_1 _26750_ (.A(_07628_),
    .B(_07631_),
    .X(_07632_));
 sg13g2_buf_1 _26751_ (.A(_07632_),
    .X(_07633_));
 sg13g2_nor2_1 _26752_ (.A(_03552_),
    .B(_00235_),
    .Y(_07634_));
 sg13g2_or3_1 _26753_ (.A(_00237_),
    .B(_05741_),
    .C(_07634_),
    .X(_07635_));
 sg13g2_buf_1 _26754_ (.A(_07635_),
    .X(_07636_));
 sg13g2_or2_1 _26755_ (.X(_07637_),
    .B(_07636_),
    .A(net288));
 sg13g2_buf_1 _26756_ (.A(_07637_),
    .X(_07638_));
 sg13g2_buf_1 _26757_ (.A(_07638_),
    .X(_07639_));
 sg13g2_nand2_1 _26758_ (.Y(_07640_),
    .A(_03312_),
    .B(_10550_));
 sg13g2_a21oi_1 _26759_ (.A1(_07636_),
    .A2(_07640_),
    .Y(_07641_),
    .B1(net288));
 sg13g2_buf_2 _26760_ (.A(_07641_),
    .X(_07642_));
 sg13g2_o21ai_1 _26761_ (.B1(_07642_),
    .Y(_07643_),
    .A1(_07633_),
    .A2(_07639_));
 sg13g2_nor2_1 _26762_ (.A(_03527_),
    .B(_07638_),
    .Y(_07644_));
 sg13g2_buf_2 _26763_ (.A(_07644_),
    .X(_07645_));
 sg13g2_buf_1 _26764_ (.A(_07645_),
    .X(_07646_));
 sg13g2_a22oi_1 _26765_ (.Y(_07647_),
    .B1(net125),
    .B2(_07633_),
    .A2(_07643_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26766_ (.A(net654),
    .B(_07647_),
    .Y(_01069_));
 sg13g2_nor3_1 _26767_ (.A(net847),
    .B(_04778_),
    .C(net738),
    .Y(_07648_));
 sg13g2_buf_2 _26768_ (.A(_07648_),
    .X(_07649_));
 sg13g2_and2_1 _26769_ (.A(net967),
    .B(_07630_),
    .X(_07650_));
 sg13g2_a21oi_1 _26770_ (.A1(net970),
    .A2(_07631_),
    .Y(_07651_),
    .B1(_07650_));
 sg13g2_nand2_1 _26771_ (.Y(_07652_),
    .A(_05845_),
    .B(_07631_));
 sg13g2_o21ai_1 _26772_ (.B1(_07652_),
    .Y(_07653_),
    .A1(_10516_),
    .A2(_07651_));
 sg13g2_buf_1 _26773_ (.A(_07653_),
    .X(_07654_));
 sg13g2_nor2b_2 _26774_ (.A(net172),
    .B_N(_07654_),
    .Y(_07655_));
 sg13g2_buf_1 _26775_ (.A(net172),
    .X(_07656_));
 sg13g2_buf_1 _26776_ (.A(_07642_),
    .X(_07657_));
 sg13g2_o21ai_1 _26777_ (.B1(net171),
    .Y(_07658_),
    .A1(_05799_),
    .A2(net152));
 sg13g2_a22oi_1 _26778_ (.Y(_07659_),
    .B1(_07658_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07655_),
    .A1(_07649_));
 sg13g2_nor2_1 _26779_ (.A(net654),
    .B(_07659_),
    .Y(_01070_));
 sg13g2_o21ai_1 _26780_ (.B1(net171),
    .Y(_07660_),
    .A1(_05805_),
    .A2(_07656_));
 sg13g2_a22oi_1 _26781_ (.Y(_07661_),
    .B1(_07660_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07645_),
    .A1(_05805_));
 sg13g2_nor2_1 _26782_ (.A(_07621_),
    .B(_07661_),
    .Y(_01071_));
 sg13g2_nand2_1 _26783_ (.Y(_07662_),
    .A(net847),
    .B(net1012));
 sg13g2_nor3_1 _26784_ (.A(_05740_),
    .B(net969),
    .C(_07662_),
    .Y(_07663_));
 sg13g2_buf_2 _26785_ (.A(_07663_),
    .X(_07664_));
 sg13g2_buf_1 _26786_ (.A(net172),
    .X(_07665_));
 sg13g2_nand2b_1 _26787_ (.Y(_07666_),
    .B(_05755_),
    .A_N(net969));
 sg13g2_nand2_1 _26788_ (.Y(_07667_),
    .A(net848),
    .B(_05746_));
 sg13g2_o21ai_1 _26789_ (.B1(_07667_),
    .Y(_07668_),
    .A1(net970),
    .A2(_07666_));
 sg13g2_and2_1 _26790_ (.A(_05734_),
    .B(_07668_),
    .X(_07669_));
 sg13g2_buf_1 _26791_ (.A(_07669_),
    .X(_07670_));
 sg13g2_and2_1 _26792_ (.A(_07654_),
    .B(_07670_),
    .X(_07671_));
 sg13g2_o21ai_1 _26793_ (.B1(net171),
    .Y(_07672_),
    .A1(net151),
    .A2(_07671_));
 sg13g2_a22oi_1 _26794_ (.Y(_07673_),
    .B1(_07672_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07664_),
    .A1(_07655_));
 sg13g2_nor2_1 _26795_ (.A(net654),
    .B(_07673_),
    .Y(_01072_));
 sg13g2_nor2_1 _26796_ (.A(_05756_),
    .B(_05817_),
    .Y(_07674_));
 sg13g2_and2_1 _26797_ (.A(_07654_),
    .B(_07674_),
    .X(_07675_));
 sg13g2_buf_1 _26798_ (.A(_07675_),
    .X(_07676_));
 sg13g2_o21ai_1 _26799_ (.B1(net171),
    .Y(_07677_),
    .A1(net151),
    .A2(_07676_));
 sg13g2_a22oi_1 _26800_ (.Y(_07678_),
    .B1(_07677_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07676_),
    .A1(net125));
 sg13g2_nor2_1 _26801_ (.A(net654),
    .B(_07678_),
    .Y(_01073_));
 sg13g2_nor2_1 _26802_ (.A(net738),
    .B(_07662_),
    .Y(_07679_));
 sg13g2_buf_2 _26803_ (.A(_07679_),
    .X(_07680_));
 sg13g2_and2_1 _26804_ (.A(_05938_),
    .B(_07654_),
    .X(_07681_));
 sg13g2_o21ai_1 _26805_ (.B1(net171),
    .Y(_07682_),
    .A1(net151),
    .A2(_07681_));
 sg13g2_a22oi_1 _26806_ (.Y(_07683_),
    .B1(_07682_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07680_),
    .A1(_07655_));
 sg13g2_nor2_1 _26807_ (.A(net654),
    .B(_07683_),
    .Y(_01074_));
 sg13g2_and2_1 _26808_ (.A(_05759_),
    .B(_07654_),
    .X(_07684_));
 sg13g2_buf_1 _26809_ (.A(_07684_),
    .X(_07685_));
 sg13g2_o21ai_1 _26810_ (.B1(net171),
    .Y(_07686_),
    .A1(_07665_),
    .A2(_07685_));
 sg13g2_a22oi_1 _26811_ (.Y(_07687_),
    .B1(_07686_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07685_),
    .A1(_07646_));
 sg13g2_nor2_1 _26812_ (.A(net654),
    .B(_07687_),
    .Y(_01075_));
 sg13g2_a21oi_1 _26813_ (.A1(net1086),
    .A2(_05782_),
    .Y(_07688_),
    .B1(_04778_));
 sg13g2_and2_1 _26814_ (.A(_06052_),
    .B(_07688_),
    .X(_07689_));
 sg13g2_buf_2 _26815_ (.A(_07689_),
    .X(_07690_));
 sg13g2_nand2_1 _26816_ (.Y(_07691_),
    .A(net968),
    .B(_05746_));
 sg13g2_o21ai_1 _26817_ (.B1(_07691_),
    .Y(_07692_),
    .A1(_05782_),
    .A2(_05837_));
 sg13g2_nand2_1 _26818_ (.Y(_07693_),
    .A(net1086),
    .B(_07692_));
 sg13g2_nor2b_1 _26819_ (.A(_07693_),
    .B_N(_07654_),
    .Y(_07694_));
 sg13g2_nand2_1 _26820_ (.Y(_07695_),
    .A(_03312_),
    .B(_10542_));
 sg13g2_a21oi_1 _26821_ (.A1(_07636_),
    .A2(_07695_),
    .Y(_07696_),
    .B1(net288));
 sg13g2_buf_2 _26822_ (.A(_07696_),
    .X(_07697_));
 sg13g2_buf_1 _26823_ (.A(_07697_),
    .X(_07698_));
 sg13g2_o21ai_1 _26824_ (.B1(net170),
    .Y(_07699_),
    .A1(net151),
    .A2(_07694_));
 sg13g2_a22oi_1 _26825_ (.Y(_07700_),
    .B1(_07699_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07690_),
    .A1(_07655_));
 sg13g2_nor2_1 _26826_ (.A(net654),
    .B(_07700_),
    .Y(_01076_));
 sg13g2_nor2_1 _26827_ (.A(net847),
    .B(_05817_),
    .Y(_07701_));
 sg13g2_nand2b_1 _26828_ (.Y(_07702_),
    .B(_10676_),
    .A_N(net1086));
 sg13g2_a21oi_1 _26829_ (.A1(_07629_),
    .A2(_07702_),
    .Y(_07703_),
    .B1(net967));
 sg13g2_nor2_1 _26830_ (.A(net967),
    .B(net1086),
    .Y(_07704_));
 sg13g2_a22oi_1 _26831_ (.Y(_07705_),
    .B1(_07704_),
    .B2(_07628_),
    .A2(_06165_),
    .A1(net1086));
 sg13g2_nor2b_1 _26832_ (.A(_07705_),
    .B_N(_07629_),
    .Y(_07706_));
 sg13g2_a21o_1 _26833_ (.A2(_07703_),
    .A1(_10516_),
    .B1(_07706_),
    .X(_07707_));
 sg13g2_buf_1 _26834_ (.A(_07707_),
    .X(_07708_));
 sg13g2_and2_1 _26835_ (.A(_07701_),
    .B(_07708_),
    .X(_07709_));
 sg13g2_buf_1 _26836_ (.A(_07709_),
    .X(_07710_));
 sg13g2_o21ai_1 _26837_ (.B1(net170),
    .Y(_07711_),
    .A1(net151),
    .A2(_07710_));
 sg13g2_a22oi_1 _26838_ (.Y(_07712_),
    .B1(_07711_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07710_),
    .A1(_07646_));
 sg13g2_nor2_1 _26839_ (.A(net654),
    .B(_07712_),
    .Y(_01077_));
 sg13g2_buf_1 _26840_ (.A(_09253_),
    .X(_07713_));
 sg13g2_nor2b_1 _26841_ (.A(net172),
    .B_N(_07708_),
    .Y(_07714_));
 sg13g2_o21ai_1 _26842_ (.B1(net170),
    .Y(_07715_),
    .A1(_05848_),
    .A2(net152));
 sg13g2_a22oi_1 _26843_ (.Y(_07716_),
    .B1(_07715_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07714_),
    .A1(_07649_));
 sg13g2_nor2_1 _26844_ (.A(net653),
    .B(_07716_),
    .Y(_01078_));
 sg13g2_o21ai_1 _26845_ (.B1(net170),
    .Y(_07717_),
    .A1(_05855_),
    .A2(net152));
 sg13g2_a22oi_1 _26846_ (.Y(_07718_),
    .B1(_07717_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07645_),
    .A1(_05855_));
 sg13g2_nor2_1 _26847_ (.A(net653),
    .B(_07718_),
    .Y(_01079_));
 sg13g2_a22oi_1 _26848_ (.Y(_07719_),
    .B1(_05845_),
    .B2(_07704_),
    .A2(_05809_),
    .A1(net1086));
 sg13g2_nor2b_1 _26849_ (.A(_07719_),
    .B_N(_07629_),
    .Y(_07720_));
 sg13g2_a21oi_1 _26850_ (.A1(_05796_),
    .A2(_07703_),
    .Y(_07721_),
    .B1(_07720_));
 sg13g2_buf_2 _26851_ (.A(_07721_),
    .X(_07722_));
 sg13g2_nor2b_1 _26852_ (.A(_07722_),
    .B_N(_07701_),
    .Y(_07723_));
 sg13g2_o21ai_1 _26853_ (.B1(net171),
    .Y(_07724_),
    .A1(_07665_),
    .A2(_07723_));
 sg13g2_a22oi_1 _26854_ (.Y(_07725_),
    .B1(_07724_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07723_),
    .A1(net125));
 sg13g2_nor2_1 _26855_ (.A(_07713_),
    .B(_07725_),
    .Y(_01080_));
 sg13g2_and2_1 _26856_ (.A(_07670_),
    .B(_07708_),
    .X(_07726_));
 sg13g2_o21ai_1 _26857_ (.B1(net170),
    .Y(_07727_),
    .A1(net151),
    .A2(_07726_));
 sg13g2_a22oi_1 _26858_ (.Y(_07728_),
    .B1(_07727_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07714_),
    .A1(_07664_));
 sg13g2_nor2_1 _26859_ (.A(net653),
    .B(_07728_),
    .Y(_01081_));
 sg13g2_and2_1 _26860_ (.A(_07674_),
    .B(_07708_),
    .X(_07729_));
 sg13g2_buf_1 _26861_ (.A(_07729_),
    .X(_07730_));
 sg13g2_o21ai_1 _26862_ (.B1(_07698_),
    .Y(_07731_),
    .A1(net151),
    .A2(_07730_));
 sg13g2_a22oi_1 _26863_ (.Y(_07732_),
    .B1(_07731_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07730_),
    .A1(net125));
 sg13g2_nor2_1 _26864_ (.A(net653),
    .B(_07732_),
    .Y(_01082_));
 sg13g2_and2_1 _26865_ (.A(_05938_),
    .B(_07708_),
    .X(_07733_));
 sg13g2_o21ai_1 _26866_ (.B1(net170),
    .Y(_07734_),
    .A1(net151),
    .A2(_07733_));
 sg13g2_a22oi_1 _26867_ (.Y(_07735_),
    .B1(_07734_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07714_),
    .A1(_07680_));
 sg13g2_nor2_1 _26868_ (.A(net653),
    .B(_07735_),
    .Y(_01083_));
 sg13g2_nor2_2 _26869_ (.A(_07691_),
    .B(_05836_),
    .Y(_07736_));
 sg13g2_buf_1 _26870_ (.A(net172),
    .X(_07737_));
 sg13g2_o21ai_1 _26871_ (.B1(_07698_),
    .Y(_07738_),
    .A1(net150),
    .A2(_07736_));
 sg13g2_a22oi_1 _26872_ (.Y(_07739_),
    .B1(_07738_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07736_),
    .A1(net125));
 sg13g2_nor2_1 _26873_ (.A(_07713_),
    .B(_07739_),
    .Y(_01084_));
 sg13g2_nor2b_1 _26874_ (.A(_07693_),
    .B_N(_07708_),
    .Y(_07740_));
 sg13g2_o21ai_1 _26875_ (.B1(net170),
    .Y(_07741_),
    .A1(net150),
    .A2(_07740_));
 sg13g2_a22oi_1 _26876_ (.Y(_07742_),
    .B1(_07741_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07714_),
    .A1(_07690_));
 sg13g2_nor2_1 _26877_ (.A(net653),
    .B(_07742_),
    .Y(_01085_));
 sg13g2_nor2_1 _26878_ (.A(_05796_),
    .B(_07651_),
    .Y(_07743_));
 sg13g2_or2_1 _26879_ (.X(_07744_),
    .B(_07743_),
    .A(_07633_));
 sg13g2_buf_1 _26880_ (.A(_07744_),
    .X(_07745_));
 sg13g2_and2_1 _26881_ (.A(_07701_),
    .B(_07745_),
    .X(_07746_));
 sg13g2_buf_1 _26882_ (.A(_07746_),
    .X(_07747_));
 sg13g2_o21ai_1 _26883_ (.B1(net170),
    .Y(_07748_),
    .A1(net150),
    .A2(_07747_));
 sg13g2_a22oi_1 _26884_ (.Y(_07749_),
    .B1(_07748_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07747_),
    .A1(net125));
 sg13g2_nor2_1 _26885_ (.A(net653),
    .B(_07749_),
    .Y(_01086_));
 sg13g2_nor2b_1 _26886_ (.A(net172),
    .B_N(_07745_),
    .Y(_07750_));
 sg13g2_o21ai_1 _26887_ (.B1(_07697_),
    .Y(_07751_),
    .A1(_05895_),
    .A2(net152));
 sg13g2_a22oi_1 _26888_ (.Y(_07752_),
    .B1(_07751_),
    .B2(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A2(_07750_),
    .A1(_07649_));
 sg13g2_nor2_1 _26889_ (.A(net653),
    .B(_07752_),
    .Y(_01087_));
 sg13g2_buf_1 _26890_ (.A(_06799_),
    .X(_07753_));
 sg13g2_o21ai_1 _26891_ (.B1(_07697_),
    .Y(_07754_),
    .A1(_05900_),
    .A2(net152));
 sg13g2_a22oi_1 _26892_ (.Y(_07755_),
    .B1(_07754_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07645_),
    .A1(_05900_));
 sg13g2_nor2_1 _26893_ (.A(net652),
    .B(_07755_),
    .Y(_01088_));
 sg13g2_and2_1 _26894_ (.A(_07670_),
    .B(_07745_),
    .X(_07756_));
 sg13g2_o21ai_1 _26895_ (.B1(_07697_),
    .Y(_07757_),
    .A1(net150),
    .A2(_07756_));
 sg13g2_a22oi_1 _26896_ (.Y(_07758_),
    .B1(_07757_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07750_),
    .A1(_07664_));
 sg13g2_nor2_1 _26897_ (.A(net652),
    .B(_07758_),
    .Y(_01089_));
 sg13g2_and2_1 _26898_ (.A(_07674_),
    .B(_07745_),
    .X(_07759_));
 sg13g2_buf_1 _26899_ (.A(_07759_),
    .X(_07760_));
 sg13g2_o21ai_1 _26900_ (.B1(_07697_),
    .Y(_07761_),
    .A1(net150),
    .A2(_07760_));
 sg13g2_a22oi_1 _26901_ (.Y(_07762_),
    .B1(_07761_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07760_),
    .A1(net125));
 sg13g2_nor2_1 _26902_ (.A(net652),
    .B(_07762_),
    .Y(_01090_));
 sg13g2_nor3_1 _26903_ (.A(net847),
    .B(net738),
    .C(_07722_),
    .Y(_07763_));
 sg13g2_o21ai_1 _26904_ (.B1(_07642_),
    .Y(_07764_),
    .A1(_07639_),
    .A2(_07763_));
 sg13g2_and2_1 _26905_ (.A(_11919_),
    .B(_07763_),
    .X(_07765_));
 sg13g2_inv_1 _26906_ (.Y(_07766_),
    .A(net152));
 sg13g2_a22oi_1 _26907_ (.Y(_07767_),
    .B1(_07765_),
    .B2(_07766_),
    .A2(_07764_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26908_ (.A(net652),
    .B(_07767_),
    .Y(_01091_));
 sg13g2_and2_1 _26909_ (.A(_05938_),
    .B(_07745_),
    .X(_07768_));
 sg13g2_o21ai_1 _26910_ (.B1(_07697_),
    .Y(_07769_),
    .A1(net150),
    .A2(_07768_));
 sg13g2_a22oi_1 _26911_ (.Y(_07770_),
    .B1(_07769_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07750_),
    .A1(_07680_));
 sg13g2_nor2_1 _26912_ (.A(net652),
    .B(_07770_),
    .Y(_01092_));
 sg13g2_and2_1 _26913_ (.A(_05759_),
    .B(_07745_),
    .X(_07771_));
 sg13g2_buf_1 _26914_ (.A(_07771_),
    .X(_07772_));
 sg13g2_o21ai_1 _26915_ (.B1(_07697_),
    .Y(_07773_),
    .A1(net150),
    .A2(_07772_));
 sg13g2_a22oi_1 _26916_ (.Y(_07774_),
    .B1(_07773_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07772_),
    .A1(net125));
 sg13g2_nor2_1 _26917_ (.A(net652),
    .B(_07774_),
    .Y(_01093_));
 sg13g2_nor2_2 _26918_ (.A(_07667_),
    .B(_07722_),
    .Y(_07775_));
 sg13g2_o21ai_1 _26919_ (.B1(net171),
    .Y(_07776_),
    .A1(_07737_),
    .A2(_07775_));
 sg13g2_a22oi_1 _26920_ (.Y(_07777_),
    .B1(_07776_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07775_),
    .A1(_07645_));
 sg13g2_nor2_1 _26921_ (.A(net652),
    .B(_07777_),
    .Y(_01094_));
 sg13g2_nor2_1 _26922_ (.A(net172),
    .B(_07722_),
    .Y(_07778_));
 sg13g2_nor2b_1 _26923_ (.A(_07722_),
    .B_N(_07670_),
    .Y(_07779_));
 sg13g2_o21ai_1 _26924_ (.B1(_07657_),
    .Y(_07780_),
    .A1(_07737_),
    .A2(_07779_));
 sg13g2_a22oi_1 _26925_ (.Y(_07781_),
    .B1(_07780_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07778_),
    .A1(_07664_));
 sg13g2_nor2_1 _26926_ (.A(net652),
    .B(_07781_),
    .Y(_01095_));
 sg13g2_o21ai_1 _26927_ (.B1(_07657_),
    .Y(_07782_),
    .A1(_05934_),
    .A2(_07656_));
 sg13g2_a22oi_1 _26928_ (.Y(_07783_),
    .B1(_07782_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07645_),
    .A1(_05934_));
 sg13g2_nor2_1 _26929_ (.A(_07753_),
    .B(_07783_),
    .Y(_01096_));
 sg13g2_o21ai_1 _26930_ (.B1(_07642_),
    .Y(_07784_),
    .A1(_05940_),
    .A2(net152));
 sg13g2_a22oi_1 _26931_ (.Y(_07785_),
    .B1(_07784_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07778_),
    .A1(_07680_));
 sg13g2_nor2_1 _26932_ (.A(_07753_),
    .B(_07785_),
    .Y(_01097_));
 sg13g2_buf_1 _26933_ (.A(_06799_),
    .X(_07786_));
 sg13g2_o21ai_1 _26934_ (.B1(_07642_),
    .Y(_07787_),
    .A1(_05945_),
    .A2(net152));
 sg13g2_a22oi_1 _26935_ (.Y(_07788_),
    .B1(_07787_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07645_),
    .A1(_05945_));
 sg13g2_nor2_1 _26936_ (.A(_07786_),
    .B(_07788_),
    .Y(_01098_));
 sg13g2_nor2_1 _26937_ (.A(_07693_),
    .B(_07722_),
    .Y(_07789_));
 sg13g2_o21ai_1 _26938_ (.B1(_07642_),
    .Y(_07790_),
    .A1(net150),
    .A2(_07789_));
 sg13g2_a22oi_1 _26939_ (.Y(_07791_),
    .B1(_07790_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07778_),
    .A1(_07690_));
 sg13g2_nor2_1 _26940_ (.A(net651),
    .B(_07791_),
    .Y(_01099_));
 sg13g2_and2_1 _26941_ (.A(_07654_),
    .B(_07701_),
    .X(_07792_));
 sg13g2_buf_1 _26942_ (.A(_07792_),
    .X(_07793_));
 sg13g2_o21ai_1 _26943_ (.B1(_07642_),
    .Y(_07794_),
    .A1(net172),
    .A2(_07793_));
 sg13g2_a22oi_1 _26944_ (.Y(_07795_),
    .B1(_07794_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07793_),
    .A1(_07645_));
 sg13g2_nor2_1 _26945_ (.A(net651),
    .B(_07795_),
    .Y(_01100_));
 sg13g2_a21oi_1 _26946_ (.A1(_08332_),
    .A2(_00235_),
    .Y(_07796_),
    .B1(_00237_));
 sg13g2_nand2_1 _26947_ (.Y(_07797_),
    .A(_05733_),
    .B(_07796_));
 sg13g2_a21oi_1 _26948_ (.A1(_05731_),
    .A2(_07797_),
    .Y(_07798_),
    .B1(net288));
 sg13g2_nand2_1 _26949_ (.Y(_07799_),
    .A(_05731_),
    .B(_07798_));
 sg13g2_buf_1 _26950_ (.A(_07799_),
    .X(_07800_));
 sg13g2_inv_1 _26951_ (.Y(_07801_),
    .A(_03312_));
 sg13g2_nor3_1 _26952_ (.A(_07801_),
    .B(_10597_),
    .C(_05728_),
    .Y(_07802_));
 sg13g2_nor2b_1 _26953_ (.A(_07802_),
    .B_N(_07798_),
    .Y(_07803_));
 sg13g2_buf_2 _26954_ (.A(_07803_),
    .X(_07804_));
 sg13g2_o21ai_1 _26955_ (.B1(_07804_),
    .Y(_07805_),
    .A1(_07633_),
    .A2(net169));
 sg13g2_nor2_1 _26956_ (.A(_03527_),
    .B(_07799_),
    .Y(_07806_));
 sg13g2_buf_2 _26957_ (.A(_07806_),
    .X(_07807_));
 sg13g2_buf_1 _26958_ (.A(_07807_),
    .X(_07808_));
 sg13g2_a22oi_1 _26959_ (.Y(_07809_),
    .B1(net124),
    .B2(_07633_),
    .A2(_07805_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26960_ (.A(net651),
    .B(_07809_),
    .Y(_01101_));
 sg13g2_nor2b_1 _26961_ (.A(net169),
    .B_N(_07654_),
    .Y(_07810_));
 sg13g2_buf_1 _26962_ (.A(net169),
    .X(_07811_));
 sg13g2_buf_1 _26963_ (.A(_07804_),
    .X(_07812_));
 sg13g2_o21ai_1 _26964_ (.B1(net148),
    .Y(_07813_),
    .A1(_05799_),
    .A2(_07811_));
 sg13g2_a22oi_1 _26965_ (.Y(_07814_),
    .B1(_07813_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07810_),
    .A1(_07649_));
 sg13g2_nor2_1 _26966_ (.A(net651),
    .B(_07814_),
    .Y(_01102_));
 sg13g2_o21ai_1 _26967_ (.B1(net148),
    .Y(_07815_),
    .A1(_05805_),
    .A2(net149));
 sg13g2_a22oi_1 _26968_ (.Y(_07816_),
    .B1(_07815_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(net124),
    .A1(_05805_));
 sg13g2_nor2_1 _26969_ (.A(net651),
    .B(_07816_),
    .Y(_01103_));
 sg13g2_o21ai_1 _26970_ (.B1(net148),
    .Y(_07817_),
    .A1(_07671_),
    .A2(net149));
 sg13g2_a22oi_1 _26971_ (.Y(_07818_),
    .B1(_07817_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07810_),
    .A1(_07664_));
 sg13g2_nor2_1 _26972_ (.A(net651),
    .B(_07818_),
    .Y(_01104_));
 sg13g2_o21ai_1 _26973_ (.B1(_07812_),
    .Y(_07819_),
    .A1(_07676_),
    .A2(net149));
 sg13g2_a22oi_1 _26974_ (.Y(_07820_),
    .B1(_07819_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(_07808_),
    .A1(_07676_));
 sg13g2_nor2_1 _26975_ (.A(net651),
    .B(_07820_),
    .Y(_01105_));
 sg13g2_o21ai_1 _26976_ (.B1(net148),
    .Y(_07821_),
    .A1(_07681_),
    .A2(net149));
 sg13g2_a22oi_1 _26977_ (.Y(_07822_),
    .B1(_07821_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07810_),
    .A1(_07680_));
 sg13g2_nor2_1 _26978_ (.A(net651),
    .B(_07822_),
    .Y(_01106_));
 sg13g2_o21ai_1 _26979_ (.B1(net148),
    .Y(_07823_),
    .A1(_07685_),
    .A2(net149));
 sg13g2_a22oi_1 _26980_ (.Y(_07824_),
    .B1(_07823_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(_07808_),
    .A1(_07685_));
 sg13g2_nor2_1 _26981_ (.A(_07786_),
    .B(_07824_),
    .Y(_01107_));
 sg13g2_buf_1 _26982_ (.A(_06799_),
    .X(_07825_));
 sg13g2_a21oi_1 _26983_ (.A1(_03312_),
    .A2(_10488_),
    .Y(_07826_),
    .B1(_05731_));
 sg13g2_nor2b_1 _26984_ (.A(_07826_),
    .B_N(_07798_),
    .Y(_07827_));
 sg13g2_buf_2 _26985_ (.A(_07827_),
    .X(_07828_));
 sg13g2_buf_1 _26986_ (.A(_07828_),
    .X(_07829_));
 sg13g2_o21ai_1 _26987_ (.B1(net147),
    .Y(_07830_),
    .A1(_07694_),
    .A2(net149));
 sg13g2_a22oi_1 _26988_ (.Y(_07831_),
    .B1(_07830_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07810_),
    .A1(_07690_));
 sg13g2_nor2_1 _26989_ (.A(_07825_),
    .B(_07831_),
    .Y(_01108_));
 sg13g2_o21ai_1 _26990_ (.B1(_07829_),
    .Y(_07832_),
    .A1(_07710_),
    .A2(net149));
 sg13g2_a22oi_1 _26991_ (.Y(_07833_),
    .B1(_07832_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net124),
    .A1(_07710_));
 sg13g2_nor2_1 _26992_ (.A(_07825_),
    .B(_07833_),
    .Y(_01109_));
 sg13g2_nor2b_1 _26993_ (.A(net169),
    .B_N(_07708_),
    .Y(_07834_));
 sg13g2_o21ai_1 _26994_ (.B1(net147),
    .Y(_07835_),
    .A1(_05848_),
    .A2(net149));
 sg13g2_a22oi_1 _26995_ (.Y(_07836_),
    .B1(_07835_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07834_),
    .A1(_07649_));
 sg13g2_nor2_1 _26996_ (.A(net650),
    .B(_07836_),
    .Y(_01110_));
 sg13g2_buf_1 _26997_ (.A(net169),
    .X(_07837_));
 sg13g2_o21ai_1 _26998_ (.B1(net147),
    .Y(_07838_),
    .A1(_05855_),
    .A2(net146));
 sg13g2_a22oi_1 _26999_ (.Y(_07839_),
    .B1(_07838_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net124),
    .A1(_05855_));
 sg13g2_nor2_1 _27000_ (.A(net650),
    .B(_07839_),
    .Y(_01111_));
 sg13g2_o21ai_1 _27001_ (.B1(net148),
    .Y(_07840_),
    .A1(_07723_),
    .A2(_07837_));
 sg13g2_a22oi_1 _27002_ (.Y(_07841_),
    .B1(_07840_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net124),
    .A1(_07723_));
 sg13g2_nor2_1 _27003_ (.A(net650),
    .B(_07841_),
    .Y(_01112_));
 sg13g2_o21ai_1 _27004_ (.B1(net147),
    .Y(_07842_),
    .A1(_07726_),
    .A2(net146));
 sg13g2_a22oi_1 _27005_ (.Y(_07843_),
    .B1(_07842_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07834_),
    .A1(_07664_));
 sg13g2_nor2_1 _27006_ (.A(net650),
    .B(_07843_),
    .Y(_01113_));
 sg13g2_o21ai_1 _27007_ (.B1(_07829_),
    .Y(_07844_),
    .A1(_07730_),
    .A2(net146));
 sg13g2_a22oi_1 _27008_ (.Y(_07845_),
    .B1(_07844_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net124),
    .A1(_07730_));
 sg13g2_nor2_1 _27009_ (.A(net650),
    .B(_07845_),
    .Y(_01114_));
 sg13g2_o21ai_1 _27010_ (.B1(net147),
    .Y(_07846_),
    .A1(_07733_),
    .A2(net146));
 sg13g2_a22oi_1 _27011_ (.Y(_07847_),
    .B1(_07846_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07834_),
    .A1(_07680_));
 sg13g2_nor2_1 _27012_ (.A(net650),
    .B(_07847_),
    .Y(_01115_));
 sg13g2_o21ai_1 _27013_ (.B1(net147),
    .Y(_07848_),
    .A1(_07736_),
    .A2(_07837_));
 sg13g2_a22oi_1 _27014_ (.Y(_07849_),
    .B1(_07848_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net124),
    .A1(_07736_));
 sg13g2_nor2_1 _27015_ (.A(net650),
    .B(_07849_),
    .Y(_01116_));
 sg13g2_o21ai_1 _27016_ (.B1(net147),
    .Y(_07850_),
    .A1(_07740_),
    .A2(net146));
 sg13g2_a22oi_1 _27017_ (.Y(_07851_),
    .B1(_07850_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07834_),
    .A1(_07690_));
 sg13g2_nor2_1 _27018_ (.A(net650),
    .B(_07851_),
    .Y(_01117_));
 sg13g2_buf_1 _27019_ (.A(_06799_),
    .X(_07852_));
 sg13g2_o21ai_1 _27020_ (.B1(net147),
    .Y(_07853_),
    .A1(_07747_),
    .A2(net146));
 sg13g2_a22oi_1 _27021_ (.Y(_07854_),
    .B1(_07853_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net124),
    .A1(_07747_));
 sg13g2_nor2_1 _27022_ (.A(net649),
    .B(_07854_),
    .Y(_01118_));
 sg13g2_nor2b_1 _27023_ (.A(net169),
    .B_N(_07745_),
    .Y(_07855_));
 sg13g2_o21ai_1 _27024_ (.B1(_07828_),
    .Y(_07856_),
    .A1(_05895_),
    .A2(net146));
 sg13g2_a22oi_1 _27025_ (.Y(_07857_),
    .B1(_07856_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07855_),
    .A1(_07649_));
 sg13g2_nor2_1 _27026_ (.A(net649),
    .B(_07857_),
    .Y(_01119_));
 sg13g2_o21ai_1 _27027_ (.B1(_07828_),
    .Y(_07858_),
    .A1(_05900_),
    .A2(net146));
 sg13g2_a22oi_1 _27028_ (.Y(_07859_),
    .B1(_07858_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07807_),
    .A1(_05900_));
 sg13g2_nor2_1 _27029_ (.A(net649),
    .B(_07859_),
    .Y(_01120_));
 sg13g2_buf_1 _27030_ (.A(net169),
    .X(_07860_));
 sg13g2_o21ai_1 _27031_ (.B1(_07828_),
    .Y(_07861_),
    .A1(_07756_),
    .A2(net145));
 sg13g2_a22oi_1 _27032_ (.Y(_07862_),
    .B1(_07861_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07855_),
    .A1(_07664_));
 sg13g2_nor2_1 _27033_ (.A(net649),
    .B(_07862_),
    .Y(_01121_));
 sg13g2_o21ai_1 _27034_ (.B1(_07828_),
    .Y(_07863_),
    .A1(_07760_),
    .A2(net145));
 sg13g2_a22oi_1 _27035_ (.Y(_07864_),
    .B1(_07863_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07807_),
    .A1(_07760_));
 sg13g2_nor2_1 _27036_ (.A(net649),
    .B(_07864_),
    .Y(_01122_));
 sg13g2_inv_1 _27037_ (.Y(_07865_),
    .A(_07811_));
 sg13g2_o21ai_1 _27038_ (.B1(net148),
    .Y(_07866_),
    .A1(_07763_),
    .A2(net145));
 sg13g2_a22oi_1 _27039_ (.Y(_07867_),
    .B1(_07866_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07865_),
    .A1(_07765_));
 sg13g2_nor2_1 _27040_ (.A(_07852_),
    .B(_07867_),
    .Y(_01123_));
 sg13g2_o21ai_1 _27041_ (.B1(_07828_),
    .Y(_07868_),
    .A1(_07768_),
    .A2(net145));
 sg13g2_a22oi_1 _27042_ (.Y(_07869_),
    .B1(_07868_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07855_),
    .A1(_07680_));
 sg13g2_nor2_1 _27043_ (.A(net649),
    .B(_07869_),
    .Y(_01124_));
 sg13g2_o21ai_1 _27044_ (.B1(_07828_),
    .Y(_07870_),
    .A1(_07772_),
    .A2(net145));
 sg13g2_a22oi_1 _27045_ (.Y(_07871_),
    .B1(_07870_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07807_),
    .A1(_07772_));
 sg13g2_nor2_1 _27046_ (.A(net649),
    .B(_07871_),
    .Y(_01125_));
 sg13g2_o21ai_1 _27047_ (.B1(net148),
    .Y(_07872_),
    .A1(_07775_),
    .A2(_07860_));
 sg13g2_a22oi_1 _27048_ (.Y(_07873_),
    .B1(_07872_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07807_),
    .A1(_07775_));
 sg13g2_nor2_1 _27049_ (.A(_07852_),
    .B(_07873_),
    .Y(_01126_));
 sg13g2_nor2_1 _27050_ (.A(_07722_),
    .B(net169),
    .Y(_07874_));
 sg13g2_o21ai_1 _27051_ (.B1(_07812_),
    .Y(_07875_),
    .A1(_07779_),
    .A2(_07860_));
 sg13g2_a22oi_1 _27052_ (.Y(_07876_),
    .B1(_07875_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07874_),
    .A1(_07664_));
 sg13g2_nor2_1 _27053_ (.A(net649),
    .B(_07876_),
    .Y(_01127_));
 sg13g2_buf_2 _27054_ (.A(_06799_),
    .X(_07877_));
 sg13g2_o21ai_1 _27055_ (.B1(_07804_),
    .Y(_07878_),
    .A1(_05934_),
    .A2(net145));
 sg13g2_a22oi_1 _27056_ (.Y(_07879_),
    .B1(_07878_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07807_),
    .A1(_05934_));
 sg13g2_nor2_1 _27057_ (.A(net648),
    .B(_07879_),
    .Y(_01128_));
 sg13g2_o21ai_1 _27058_ (.B1(_07804_),
    .Y(_07880_),
    .A1(_05940_),
    .A2(net145));
 sg13g2_a22oi_1 _27059_ (.Y(_07881_),
    .B1(_07880_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07874_),
    .A1(_07680_));
 sg13g2_nor2_1 _27060_ (.A(net648),
    .B(_07881_),
    .Y(_01129_));
 sg13g2_o21ai_1 _27061_ (.B1(_07804_),
    .Y(_07882_),
    .A1(_05945_),
    .A2(net145));
 sg13g2_a22oi_1 _27062_ (.Y(_07883_),
    .B1(_07882_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07807_),
    .A1(_05945_));
 sg13g2_nor2_1 _27063_ (.A(net648),
    .B(_07883_),
    .Y(_01130_));
 sg13g2_o21ai_1 _27064_ (.B1(_07804_),
    .Y(_07884_),
    .A1(_07789_),
    .A2(_07800_));
 sg13g2_a22oi_1 _27065_ (.Y(_07885_),
    .B1(_07884_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07874_),
    .A1(_07690_));
 sg13g2_nor2_1 _27066_ (.A(_07877_),
    .B(_07885_),
    .Y(_01131_));
 sg13g2_o21ai_1 _27067_ (.B1(_07804_),
    .Y(_07886_),
    .A1(_07793_),
    .A2(_07800_));
 sg13g2_a22oi_1 _27068_ (.Y(_07887_),
    .B1(_07886_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07807_),
    .A1(_07793_));
 sg13g2_nor2_1 _27069_ (.A(_07877_),
    .B(_07887_),
    .Y(_01132_));
 sg13g2_inv_1 _27070_ (.Y(_07888_),
    .A(net390));
 sg13g2_nor2_1 _27071_ (.A(_07888_),
    .B(net129),
    .Y(_07889_));
 sg13g2_buf_2 _27072_ (.A(_07889_),
    .X(_07890_));
 sg13g2_nand2_1 _27073_ (.Y(_07891_),
    .A(net865),
    .B(_07890_));
 sg13g2_or2_1 _27074_ (.X(_07892_),
    .B(_06369_),
    .A(_07888_));
 sg13g2_buf_2 _27075_ (.A(_07892_),
    .X(_07893_));
 sg13g2_nand2_1 _27076_ (.Y(_07894_),
    .A(\cpu.gpio.r_enable_in[0] ),
    .B(_07893_));
 sg13g2_buf_1 _27077_ (.A(_06799_),
    .X(_07895_));
 sg13g2_a21oi_1 _27078_ (.A1(_07891_),
    .A2(_07894_),
    .Y(_01933_),
    .B1(net647));
 sg13g2_nand2_1 _27079_ (.Y(_07896_),
    .A(_10051_),
    .B(_07890_));
 sg13g2_nand2_1 _27080_ (.Y(_07897_),
    .A(_09093_),
    .B(_07893_));
 sg13g2_a21oi_1 _27081_ (.A1(_07896_),
    .A2(_07897_),
    .Y(_01934_),
    .B1(net647));
 sg13g2_nand2_1 _27082_ (.Y(_07898_),
    .A(_10057_),
    .B(_07890_));
 sg13g2_nand2_1 _27083_ (.Y(_07899_),
    .A(_09088_),
    .B(_07893_));
 sg13g2_a21oi_1 _27084_ (.A1(_07898_),
    .A2(_07899_),
    .Y(_01935_),
    .B1(_07895_));
 sg13g2_nand2_1 _27085_ (.Y(_07900_),
    .A(net1044),
    .B(_07890_));
 sg13g2_nand2_1 _27086_ (.Y(_07901_),
    .A(_09111_),
    .B(_07893_));
 sg13g2_a21oi_1 _27087_ (.A1(_07900_),
    .A2(_07901_),
    .Y(_01936_),
    .B1(net647));
 sg13g2_nand2_1 _27088_ (.Y(_07902_),
    .A(_10014_),
    .B(_07890_));
 sg13g2_nand2_1 _27089_ (.Y(_07903_),
    .A(_09090_),
    .B(_07893_));
 sg13g2_a21oi_1 _27090_ (.A1(_07902_),
    .A2(_07903_),
    .Y(_01937_),
    .B1(_07895_));
 sg13g2_nand2_1 _27091_ (.Y(_07904_),
    .A(_10020_),
    .B(_07890_));
 sg13g2_nand2_1 _27092_ (.Y(_07905_),
    .A(_09113_),
    .B(_07893_));
 sg13g2_a21oi_1 _27093_ (.A1(_07904_),
    .A2(_07905_),
    .Y(_01938_),
    .B1(net647));
 sg13g2_nand2_1 _27094_ (.Y(_07906_),
    .A(net1119),
    .B(_07890_));
 sg13g2_nand2_1 _27095_ (.Y(_07907_),
    .A(_09099_),
    .B(_07893_));
 sg13g2_a21oi_1 _27096_ (.A1(_07906_),
    .A2(_07907_),
    .Y(_01939_),
    .B1(net647));
 sg13g2_nand2_1 _27097_ (.Y(_07908_),
    .A(net1118),
    .B(_07890_));
 sg13g2_nand2_1 _27098_ (.Y(_07909_),
    .A(_09108_),
    .B(_07893_));
 sg13g2_a21oi_1 _27099_ (.A1(_07908_),
    .A2(_07909_),
    .Y(_01940_),
    .B1(net647));
 sg13g2_nor3_1 _27100_ (.A(_11843_),
    .B(_04855_),
    .C(_06369_),
    .Y(_07910_));
 sg13g2_buf_2 _27101_ (.A(_07910_),
    .X(_07911_));
 sg13g2_nand2_1 _27102_ (.Y(_07912_),
    .A(_10014_),
    .B(_07911_));
 sg13g2_nand2b_1 _27103_ (.Y(_07913_),
    .B(_09103_),
    .A_N(_07911_));
 sg13g2_a21oi_1 _27104_ (.A1(_07912_),
    .A2(_07913_),
    .Y(_01941_),
    .B1(net647));
 sg13g2_nand2_1 _27105_ (.Y(_07914_),
    .A(_10020_),
    .B(_07911_));
 sg13g2_nand2b_1 _27106_ (.Y(_07915_),
    .B(_09105_),
    .A_N(_07911_));
 sg13g2_a21oi_1 _27107_ (.A1(_07914_),
    .A2(_07915_),
    .Y(_01942_),
    .B1(net647));
 sg13g2_nand2_1 _27108_ (.Y(_07916_),
    .A(net1119),
    .B(_07911_));
 sg13g2_nand2b_1 _27109_ (.Y(_07917_),
    .B(\cpu.gpio.r_enable_io[6] ),
    .A_N(_07911_));
 sg13g2_buf_1 _27110_ (.A(net798),
    .X(_07918_));
 sg13g2_a21oi_1 _27111_ (.A1(_07916_),
    .A2(_07917_),
    .Y(_01943_),
    .B1(net646));
 sg13g2_nand2_1 _27112_ (.Y(_07919_),
    .A(net1118),
    .B(_07911_));
 sg13g2_nand2b_1 _27113_ (.Y(_07920_),
    .B(_09095_),
    .A_N(_07911_));
 sg13g2_a21oi_1 _27114_ (.A1(_07919_),
    .A2(_07920_),
    .Y(_01944_),
    .B1(_07918_));
 sg13g2_nand2_2 _27115_ (.Y(_07921_),
    .A(_04817_),
    .B(_04977_));
 sg13g2_nor2_1 _27116_ (.A(net129),
    .B(_07921_),
    .Y(_07922_));
 sg13g2_nand2_1 _27117_ (.Y(_07923_),
    .A(net1043),
    .B(_07922_));
 sg13g2_buf_1 _27118_ (.A(net129),
    .X(_07924_));
 sg13g2_o21ai_1 _27119_ (.B1(net8),
    .Y(_07925_),
    .A1(net109),
    .A2(_07921_));
 sg13g2_a21oi_1 _27120_ (.A1(_07923_),
    .A2(_07925_),
    .Y(_01945_),
    .B1(net646));
 sg13g2_nand2_1 _27121_ (.Y(_07926_),
    .A(net1042),
    .B(_07922_));
 sg13g2_o21ai_1 _27122_ (.B1(net9),
    .Y(_07927_),
    .A1(net109),
    .A2(_07921_));
 sg13g2_a21oi_1 _27123_ (.A1(_07926_),
    .A2(_07927_),
    .Y(_01946_),
    .B1(net646));
 sg13g2_nand2_1 _27124_ (.Y(_07928_),
    .A(net1119),
    .B(_07922_));
 sg13g2_o21ai_1 _27125_ (.B1(net10),
    .Y(_07929_),
    .A1(net109),
    .A2(_07921_));
 sg13g2_a21oi_1 _27126_ (.A1(_07928_),
    .A2(_07929_),
    .Y(_01947_),
    .B1(net646));
 sg13g2_nand2_1 _27127_ (.Y(_07930_),
    .A(net1118),
    .B(_07922_));
 sg13g2_o21ai_1 _27128_ (.B1(net11),
    .Y(_07931_),
    .A1(net129),
    .A2(_07921_));
 sg13g2_a21oi_1 _27129_ (.A1(_07930_),
    .A2(_07931_),
    .Y(_01948_),
    .B1(net646));
 sg13g2_nor2_1 _27130_ (.A(net386),
    .B(net129),
    .Y(_07932_));
 sg13g2_nand2_1 _27131_ (.Y(_07933_),
    .A(net865),
    .B(_07932_));
 sg13g2_o21ai_1 _27132_ (.B1(_04824_),
    .Y(_07934_),
    .A1(net386),
    .A2(net109));
 sg13g2_nand3_1 _27133_ (.B(_07933_),
    .C(_07934_),
    .A(net715),
    .Y(_01994_));
 sg13g2_nand2_1 _27134_ (.Y(_07935_),
    .A(net1040),
    .B(_07932_));
 sg13g2_buf_1 _27135_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07936_));
 sg13g2_o21ai_1 _27136_ (.B1(_07936_),
    .Y(_07937_),
    .A1(net386),
    .A2(net109));
 sg13g2_a21oi_1 _27137_ (.A1(_07935_),
    .A2(_07937_),
    .Y(_01995_),
    .B1(net646));
 sg13g2_nand2_1 _27138_ (.Y(_07938_),
    .A(net898),
    .B(_07932_));
 sg13g2_o21ai_1 _27139_ (.B1(\cpu.gpio.r_src_o[6][2] ),
    .Y(_07939_),
    .A1(net386),
    .A2(net109));
 sg13g2_a21oi_1 _27140_ (.A1(_07938_),
    .A2(_07939_),
    .Y(_01996_),
    .B1(net646));
 sg13g2_nand2_1 _27141_ (.Y(_07940_),
    .A(net1044),
    .B(_07932_));
 sg13g2_o21ai_1 _27142_ (.B1(\cpu.gpio.r_src_o[6][3] ),
    .Y(_07941_),
    .A1(_05015_),
    .A2(net109));
 sg13g2_a21oi_1 _27143_ (.A1(_07940_),
    .A2(_07941_),
    .Y(_01997_),
    .B1(net646));
 sg13g2_nor2_1 _27144_ (.A(_05274_),
    .B(net129),
    .Y(_07942_));
 sg13g2_nand2_1 _27145_ (.Y(_07943_),
    .A(net865),
    .B(_07942_));
 sg13g2_o21ai_1 _27146_ (.B1(_04830_),
    .Y(_07944_),
    .A1(_05274_),
    .A2(net109));
 sg13g2_a21oi_1 _27147_ (.A1(_07943_),
    .A2(_07944_),
    .Y(_02002_),
    .B1(_07918_));
 sg13g2_nand2_1 _27148_ (.Y(_07945_),
    .A(net1046),
    .B(_07942_));
 sg13g2_o21ai_1 _27149_ (.B1(\cpu.gpio.r_uart_rx_src[1] ),
    .Y(_07946_),
    .A1(_05274_),
    .A2(_07924_));
 sg13g2_buf_1 _27150_ (.A(_09232_),
    .X(_07947_));
 sg13g2_a21oi_1 _27151_ (.A1(_07945_),
    .A2(_07946_),
    .Y(_02003_),
    .B1(net645));
 sg13g2_nand2_1 _27152_ (.Y(_07948_),
    .A(net898),
    .B(_07942_));
 sg13g2_o21ai_1 _27153_ (.B1(\cpu.gpio.r_uart_rx_src[2] ),
    .Y(_07949_),
    .A1(_05274_),
    .A2(_07924_));
 sg13g2_a21oi_1 _27154_ (.A1(_07948_),
    .A2(_07949_),
    .Y(_02004_),
    .B1(_07947_));
 sg13g2_and2_1 _27155_ (.A(\cpu.i_wstrobe_d ),
    .B(_00312_),
    .X(_02261_));
 sg13g2_nor2_1 _27156_ (.A(_06425_),
    .B(_06438_),
    .Y(_07950_));
 sg13g2_nor2_1 _27157_ (.A(_06452_),
    .B(_07950_),
    .Y(_02262_));
 sg13g2_xor2_1 _27158_ (.B(_06453_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_07951_));
 sg13g2_nor2_1 _27159_ (.A(_06452_),
    .B(_07951_),
    .Y(_02263_));
 sg13g2_nand4_1 _27160_ (.B(_09995_),
    .C(net128),
    .A(net669),
    .Y(_07952_),
    .D(_04845_));
 sg13g2_nor2_1 _27161_ (.A(net609),
    .B(_07952_),
    .Y(_07953_));
 sg13g2_a21oi_1 _27162_ (.A1(\cpu.intr.r_clock ),
    .A2(_07952_),
    .Y(_07954_),
    .B1(_07953_));
 sg13g2_xnor2_1 _27163_ (.Y(_07955_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10079_));
 sg13g2_xnor2_1 _27164_ (.Y(_07956_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10126_));
 sg13g2_xnor2_1 _27165_ (.Y(_07957_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10120_));
 sg13g2_xnor2_1 _27166_ (.Y(_07958_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05477_));
 sg13g2_nand4_1 _27167_ (.B(_07956_),
    .C(_07957_),
    .A(_07955_),
    .Y(_07959_),
    .D(_07958_));
 sg13g2_xnor2_1 _27168_ (.Y(_07960_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10083_));
 sg13g2_xnor2_1 _27169_ (.Y(_07961_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10131_));
 sg13g2_xnor2_1 _27170_ (.Y(_07962_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10052_));
 sg13g2_xnor2_1 _27171_ (.Y(_07963_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05676_));
 sg13g2_nand4_1 _27172_ (.B(_07961_),
    .C(_07962_),
    .A(_07960_),
    .Y(_07964_),
    .D(_07963_));
 sg13g2_xnor2_1 _27173_ (.Y(_07965_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05184_));
 sg13g2_xnor2_1 _27174_ (.Y(_07966_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05295_));
 sg13g2_xnor2_1 _27175_ (.Y(_07967_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05665_));
 sg13g2_xnor2_1 _27176_ (.Y(_07968_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10095_));
 sg13g2_nand4_1 _27177_ (.B(_07966_),
    .C(_07967_),
    .A(_07965_),
    .Y(_07969_),
    .D(_07968_));
 sg13g2_xnor2_1 _27178_ (.Y(_07970_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10073_));
 sg13g2_xnor2_1 _27179_ (.Y(_07971_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10063_));
 sg13g2_xnor2_1 _27180_ (.Y(_07972_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05158_));
 sg13g2_xnor2_1 _27181_ (.Y(_07973_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10114_));
 sg13g2_nand4_1 _27182_ (.B(_07971_),
    .C(_07972_),
    .A(_07970_),
    .Y(_07974_),
    .D(_07973_));
 sg13g2_nor4_1 _27183_ (.A(_07959_),
    .B(_07964_),
    .C(_07969_),
    .D(_07974_),
    .Y(_07975_));
 sg13g2_xnor2_1 _27184_ (.Y(_07976_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10088_));
 sg13g2_xnor2_1 _27185_ (.Y(_07977_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05526_));
 sg13g2_xnor2_1 _27186_ (.Y(_07978_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04897_));
 sg13g2_xnor2_1 _27187_ (.Y(_07979_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10053_));
 sg13g2_nand4_1 _27188_ (.B(_07977_),
    .C(_07978_),
    .A(_07976_),
    .Y(_07980_),
    .D(_07979_));
 sg13g2_xnor2_1 _27189_ (.Y(_07981_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05008_));
 sg13g2_xnor2_1 _27190_ (.Y(_07982_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10101_));
 sg13g2_xnor2_1 _27191_ (.Y(_07983_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10106_));
 sg13g2_xnor2_1 _27192_ (.Y(_07984_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05133_));
 sg13g2_nand4_1 _27193_ (.B(_07982_),
    .C(_07983_),
    .A(_07981_),
    .Y(_07985_),
    .D(_07984_));
 sg13g2_xnor2_1 _27194_ (.Y(_07986_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(\cpu.intr.r_clock_count[31] ));
 sg13g2_xnor2_1 _27195_ (.Y(_07987_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10058_));
 sg13g2_xnor2_1 _27196_ (.Y(_07988_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10068_));
 sg13g2_xnor2_1 _27197_ (.Y(_07989_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05615_));
 sg13g2_nand4_1 _27198_ (.B(_07987_),
    .C(_07988_),
    .A(_07986_),
    .Y(_07990_),
    .D(_07989_));
 sg13g2_xnor2_1 _27199_ (.Y(_07991_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_04983_));
 sg13g2_xnor2_1 _27200_ (.Y(_07992_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05411_));
 sg13g2_xnor2_1 _27201_ (.Y(_07993_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05105_));
 sg13g2_xnor2_1 _27202_ (.Y(_07994_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05366_));
 sg13g2_nand4_1 _27203_ (.B(_07992_),
    .C(_07993_),
    .A(_07991_),
    .Y(_07995_),
    .D(_07994_));
 sg13g2_nor4_1 _27204_ (.A(_07980_),
    .B(_07985_),
    .C(_07990_),
    .D(_07995_),
    .Y(_07996_));
 sg13g2_nand2_1 _27205_ (.Y(_07997_),
    .A(_07975_),
    .B(_07996_));
 sg13g2_a21oi_1 _27206_ (.A1(_07954_),
    .A2(_07997_),
    .Y(_02424_),
    .B1(net645));
 sg13g2_and2_1 _27207_ (.A(net128),
    .B(net389),
    .X(_07998_));
 sg13g2_buf_1 _27208_ (.A(_07998_),
    .X(_07999_));
 sg13g2_nand2_1 _27209_ (.Y(_08000_),
    .A(net1047),
    .B(_07999_));
 sg13g2_nand2_1 _27210_ (.Y(_08001_),
    .A(net128),
    .B(net389));
 sg13g2_buf_1 _27211_ (.A(_08001_),
    .X(_08002_));
 sg13g2_nand2_1 _27212_ (.Y(_08003_),
    .A(_09129_),
    .B(_08002_));
 sg13g2_a21oi_1 _27213_ (.A1(_08000_),
    .A2(_08003_),
    .Y(_02473_),
    .B1(net645));
 sg13g2_nand2_1 _27214_ (.Y(_08004_),
    .A(net1046),
    .B(_07999_));
 sg13g2_nand2_1 _27215_ (.Y(_08005_),
    .A(_09124_),
    .B(_08002_));
 sg13g2_a21oi_1 _27216_ (.A1(_08004_),
    .A2(_08005_),
    .Y(_02474_),
    .B1(net645));
 sg13g2_nand2_1 _27217_ (.Y(_08006_),
    .A(net898),
    .B(_07999_));
 sg13g2_nand2_1 _27218_ (.Y(_08007_),
    .A(_09125_),
    .B(_08002_));
 sg13g2_a21oi_1 _27219_ (.A1(_08006_),
    .A2(_08007_),
    .Y(_02475_),
    .B1(net645));
 sg13g2_nand2_1 _27220_ (.Y(_08008_),
    .A(net1044),
    .B(_07999_));
 sg13g2_nand2_1 _27221_ (.Y(_08009_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_08002_));
 sg13g2_a21oi_1 _27222_ (.A1(_08008_),
    .A2(_08009_),
    .Y(_02476_),
    .B1(net645));
 sg13g2_nand2_1 _27223_ (.Y(_08010_),
    .A(net1043),
    .B(_07999_));
 sg13g2_nand2_1 _27224_ (.Y(_08011_),
    .A(_09118_),
    .B(_08002_));
 sg13g2_a21oi_1 _27225_ (.A1(_08010_),
    .A2(_08011_),
    .Y(_02477_),
    .B1(net645));
 sg13g2_nand2_1 _27226_ (.Y(_08012_),
    .A(net1042),
    .B(_07999_));
 sg13g2_nand2_1 _27227_ (.Y(_08013_),
    .A(_09122_),
    .B(_08002_));
 sg13g2_a21oi_1 _27228_ (.A1(_08012_),
    .A2(_08013_),
    .Y(_02478_),
    .B1(net645));
 sg13g2_nand3_1 _27229_ (.B(_06722_),
    .C(_04918_),
    .A(net1045),
    .Y(_08014_));
 sg13g2_nand3_1 _27230_ (.B(_06722_),
    .C(net427),
    .A(_10001_),
    .Y(_08015_));
 sg13g2_nand2_1 _27231_ (.Y(_08016_),
    .A(_09940_),
    .B(_08015_));
 sg13g2_a21oi_1 _27232_ (.A1(\cpu.intr.r_timer ),
    .A2(_08014_),
    .Y(_08017_),
    .B1(_08016_));
 sg13g2_nor2_1 _27233_ (.A(net648),
    .B(_08017_),
    .Y(_02479_));
 sg13g2_nand4_1 _27234_ (.B(_09826_),
    .C(_06886_),
    .A(_09777_),
    .Y(_08018_),
    .D(_06850_));
 sg13g2_buf_1 _27235_ (.A(_08018_),
    .X(_08019_));
 sg13g2_a21o_1 _27236_ (.A2(_09818_),
    .A1(_09800_),
    .B1(_08019_),
    .X(_08020_));
 sg13g2_o21ai_1 _27237_ (.B1(net802),
    .Y(_08021_),
    .A1(_06885_),
    .A2(_08019_));
 sg13g2_a21o_1 _27238_ (.A2(_08020_),
    .A1(net20),
    .B1(_08021_),
    .X(_02509_));
 sg13g2_nand3b_1 _27239_ (.B(\cpu.qspi.r_state[0] ),
    .C(_09779_),
    .Y(_08022_),
    .A_N(_09800_));
 sg13g2_a21o_1 _27240_ (.A2(_08022_),
    .A1(_06885_),
    .B1(_08019_),
    .X(_08023_));
 sg13g2_nand2_1 _27241_ (.Y(_08024_),
    .A(_09800_),
    .B(_06885_));
 sg13g2_nor2_1 _27242_ (.A(_09814_),
    .B(_08024_),
    .Y(_08025_));
 sg13g2_o21ai_1 _27243_ (.B1(net21),
    .Y(_08026_),
    .A1(_08019_),
    .A2(_08025_));
 sg13g2_nand3_1 _27244_ (.B(_08023_),
    .C(_08026_),
    .A(net715),
    .Y(_02510_));
 sg13g2_nor2b_1 _27245_ (.A(_09808_),
    .B_N(_09800_),
    .Y(_08027_));
 sg13g2_buf_1 _27246_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_08028_));
 sg13g2_o21ai_1 _27247_ (.B1(_08028_),
    .Y(_08029_),
    .A1(_08019_),
    .A2(_08027_));
 sg13g2_nand2b_1 _27248_ (.Y(_02511_),
    .B(_08029_),
    .A_N(_08021_));
 sg13g2_inv_1 _27249_ (.Y(_08030_),
    .A(\cpu.qspi.r_state[0] ));
 sg13g2_nand2_1 _27250_ (.Y(_08031_),
    .A(_08030_),
    .B(_06740_));
 sg13g2_nor3_1 _27251_ (.A(_09788_),
    .B(_09827_),
    .C(_08031_),
    .Y(_08032_));
 sg13g2_inv_1 _27252_ (.Y(_08033_),
    .A(_06739_));
 sg13g2_nor3_1 _27253_ (.A(_09842_),
    .B(_08033_),
    .C(_06746_),
    .Y(_08034_));
 sg13g2_nand2_1 _27254_ (.Y(_08035_),
    .A(_09822_),
    .B(_08034_));
 sg13g2_nor2_1 _27255_ (.A(_09795_),
    .B(_08035_),
    .Y(_08036_));
 sg13g2_a21oi_1 _27256_ (.A1(_08032_),
    .A2(_08036_),
    .Y(_08037_),
    .B1(_09779_));
 sg13g2_nor2_1 _27257_ (.A(net648),
    .B(_08037_),
    .Y(_02512_));
 sg13g2_nand2_1 _27258_ (.Y(_08038_),
    .A(_10033_),
    .B(_06781_));
 sg13g2_nand2_1 _27259_ (.Y(_08039_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06784_));
 sg13g2_a21oi_1 _27260_ (.A1(_08038_),
    .A2(_08039_),
    .Y(_02513_),
    .B1(_07947_));
 sg13g2_a21oi_1 _27261_ (.A1(net534),
    .A2(_04893_),
    .Y(_08040_),
    .B1(net972));
 sg13g2_nor2b_1 _27262_ (.A(_06779_),
    .B_N(_08040_),
    .Y(_08041_));
 sg13g2_inv_1 _27263_ (.Y(_08042_),
    .A(_07248_));
 sg13g2_a22oi_1 _27264_ (.Y(_08043_),
    .B1(_08041_),
    .B2(_08042_),
    .A2(_06795_),
    .A1(\cpu.qspi.r_mask[1] ));
 sg13g2_nand2_1 _27265_ (.Y(_02514_),
    .A(net694),
    .B(_08043_));
 sg13g2_nor2_1 _27266_ (.A(_07248_),
    .B(_06809_),
    .Y(_08044_));
 sg13g2_a21oi_1 _27267_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06809_),
    .Y(_08045_),
    .B1(_08044_));
 sg13g2_nor2_1 _27268_ (.A(net648),
    .B(_08045_),
    .Y(_02515_));
 sg13g2_nand2_1 _27269_ (.Y(_08046_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06784_));
 sg13g2_nand2_1 _27270_ (.Y(_08047_),
    .A(_10078_),
    .B(_06781_));
 sg13g2_nand3_1 _27271_ (.B(_08046_),
    .C(_08047_),
    .A(net715),
    .Y(_02516_));
 sg13g2_a22oi_1 _27272_ (.Y(_08048_),
    .B1(_08041_),
    .B2(_07243_),
    .A2(_06795_),
    .A1(\cpu.qspi.r_quad[1] ));
 sg13g2_nor2_1 _27273_ (.A(net648),
    .B(_08048_),
    .Y(_02517_));
 sg13g2_nand2_1 _27274_ (.Y(_08049_),
    .A(_00166_),
    .B(_06806_));
 sg13g2_o21ai_1 _27275_ (.B1(_08049_),
    .Y(_08050_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06806_));
 sg13g2_nand2_1 _27276_ (.Y(_02518_),
    .A(net694),
    .B(_08050_));
 sg13g2_nor2_1 _27277_ (.A(_04819_),
    .B(_06779_),
    .Y(_08051_));
 sg13g2_nand2_1 _27278_ (.Y(_08052_),
    .A(net865),
    .B(_08051_));
 sg13g2_o21ai_1 _27279_ (.B1(\cpu.qspi.r_rom_mode[0] ),
    .Y(_08053_),
    .A1(_04819_),
    .A2(_06779_));
 sg13g2_nand3_1 _27280_ (.B(_08052_),
    .C(_08053_),
    .A(net715),
    .Y(_02531_));
 sg13g2_nand2_1 _27281_ (.Y(_08054_),
    .A(net1040),
    .B(_08051_));
 sg13g2_o21ai_1 _27282_ (.B1(_09803_),
    .Y(_08055_),
    .A1(_04819_),
    .A2(_06779_));
 sg13g2_nand3_1 _27283_ (.B(_08054_),
    .C(_08055_),
    .A(net715),
    .Y(_02532_));
 sg13g2_nand3_1 _27284_ (.B(_09777_),
    .C(_08034_),
    .A(_11799_),
    .Y(_08056_));
 sg13g2_a21oi_1 _27285_ (.A1(_11778_),
    .A2(_06883_),
    .Y(_08057_),
    .B1(_08056_));
 sg13g2_nand2b_1 _27286_ (.Y(_08058_),
    .B(net4),
    .A_N(_08057_));
 sg13g2_nand2_1 _27287_ (.Y(_08059_),
    .A(_09829_),
    .B(_08032_));
 sg13g2_nand3_1 _27288_ (.B(_08030_),
    .C(_08059_),
    .A(_11777_),
    .Y(_08060_));
 sg13g2_nand2_1 _27289_ (.Y(_08061_),
    .A(_08057_),
    .B(_08060_));
 sg13g2_buf_1 _27290_ (.A(net798),
    .X(_08062_));
 sg13g2_a21oi_1 _27291_ (.A1(_08058_),
    .A2(_08061_),
    .Y(_02533_),
    .B1(net644));
 sg13g2_nand2b_1 _27292_ (.Y(_08063_),
    .B(net7),
    .A_N(_08057_));
 sg13g2_o21ai_1 _27293_ (.B1(_11777_),
    .Y(_08064_),
    .A1(_09821_),
    .A2(_08059_));
 sg13g2_nand2_1 _27294_ (.Y(_08065_),
    .A(_08057_),
    .B(_08064_));
 sg13g2_a21oi_1 _27295_ (.A1(_08063_),
    .A2(_08065_),
    .Y(_02534_),
    .B1(net644));
 sg13g2_nor3_1 _27296_ (.A(net1055),
    .B(net1127),
    .C(_09239_),
    .Y(_08066_));
 sg13g2_nor3_1 _27297_ (.A(_09235_),
    .B(_09255_),
    .C(_08066_),
    .Y(_08067_));
 sg13g2_buf_2 _27298_ (.A(_08067_),
    .X(_08068_));
 sg13g2_nand3_1 _27299_ (.B(net1055),
    .C(_08068_),
    .A(_09175_),
    .Y(_08069_));
 sg13g2_o21ai_1 _27300_ (.B1(_08069_),
    .Y(_08070_),
    .A1(_09175_),
    .A2(_08068_));
 sg13g2_nand2_1 _27301_ (.Y(_02540_),
    .A(net694),
    .B(_08070_));
 sg13g2_nand2_1 _27302_ (.Y(_08071_),
    .A(_09175_),
    .B(_11806_));
 sg13g2_a21oi_1 _27303_ (.A1(_08068_),
    .A2(_08071_),
    .Y(_08072_),
    .B1(_09176_));
 sg13g2_inv_1 _27304_ (.Y(_08073_),
    .A(_09175_));
 sg13g2_and4_1 _27305_ (.A(_08073_),
    .B(_09176_),
    .C(_11806_),
    .D(_08068_),
    .X(_08074_));
 sg13g2_o21ai_1 _27306_ (.B1(net694),
    .Y(_02541_),
    .A1(_08072_),
    .A2(_08074_));
 sg13g2_nor2_1 _27307_ (.A(_09175_),
    .B(_09176_),
    .Y(_08075_));
 sg13g2_or2_1 _27308_ (.X(_08076_),
    .B(_08075_),
    .A(_00207_));
 sg13g2_a21oi_1 _27309_ (.A1(_08068_),
    .A2(_08076_),
    .Y(_08077_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27310_ (.A(\cpu.spi.r_bits[2] ),
    .B(_11806_),
    .C(_08075_),
    .D(_08068_),
    .X(_08078_));
 sg13g2_o21ai_1 _27311_ (.B1(net694),
    .Y(_02542_),
    .A1(_08077_),
    .A2(_08078_));
 sg13g2_buf_1 _27312_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08079_));
 sg13g2_inv_1 _27313_ (.Y(_08080_),
    .A(_08079_));
 sg13g2_nor2b_1 _27314_ (.A(_09220_),
    .B_N(_09158_),
    .Y(_08081_));
 sg13g2_or2_1 _27315_ (.X(_08082_),
    .B(_09236_),
    .A(net1127));
 sg13g2_buf_1 _27316_ (.A(_08082_),
    .X(_08083_));
 sg13g2_nand2_1 _27317_ (.Y(_08084_),
    .A(_09210_),
    .B(_08083_));
 sg13g2_nor3_1 _27318_ (.A(net1125),
    .B(_09209_),
    .C(_08083_),
    .Y(_08085_));
 sg13g2_a21oi_1 _27319_ (.A1(net1020),
    .A2(net875),
    .Y(_08086_),
    .B1(_09225_));
 sg13g2_nor3_1 _27320_ (.A(_00259_),
    .B(_08085_),
    .C(_08086_),
    .Y(_08087_));
 sg13g2_a21oi_1 _27321_ (.A1(_00259_),
    .A2(_08084_),
    .Y(_08088_),
    .B1(_08087_));
 sg13g2_o21ai_1 _27322_ (.B1(_08088_),
    .Y(_08089_),
    .A1(_07006_),
    .A2(_08081_));
 sg13g2_buf_1 _27323_ (.A(_08089_),
    .X(_08090_));
 sg13g2_nor3_1 _27324_ (.A(_11810_),
    .B(net875),
    .C(_08090_),
    .Y(_08091_));
 sg13g2_inv_1 _27325_ (.Y(_08092_),
    .A(_08090_));
 sg13g2_a21oi_1 _27326_ (.A1(_08083_),
    .A2(_08092_),
    .Y(_08093_),
    .B1(net798));
 sg13g2_o21ai_1 _27327_ (.B1(_08093_),
    .Y(_02575_),
    .A1(_08080_),
    .A2(_08091_));
 sg13g2_nand2_1 _27328_ (.Y(_08094_),
    .A(_11824_),
    .B(net875));
 sg13g2_buf_1 _27329_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08095_));
 sg13g2_o21ai_1 _27330_ (.B1(_08095_),
    .Y(_08096_),
    .A1(_08090_),
    .A2(_08094_));
 sg13g2_nand2_1 _27331_ (.Y(_02576_),
    .A(_08093_),
    .B(_08096_));
 sg13g2_buf_1 _27332_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08097_));
 sg13g2_inv_1 _27333_ (.Y(_08098_),
    .A(_08097_));
 sg13g2_nor3_1 _27334_ (.A(_11824_),
    .B(net875),
    .C(_08090_),
    .Y(_08099_));
 sg13g2_o21ai_1 _27335_ (.B1(_08093_),
    .Y(_02577_),
    .A1(_08098_),
    .A2(_08099_));
 sg13g2_nand2_1 _27336_ (.Y(_08100_),
    .A(_09198_),
    .B(net410));
 sg13g2_nor3_1 _27337_ (.A(_07006_),
    .B(_09158_),
    .C(_09219_),
    .Y(_08101_));
 sg13g2_a21oi_1 _27338_ (.A1(_09173_),
    .A2(_08100_),
    .Y(_08102_),
    .B1(_08101_));
 sg13g2_nand2_1 _27339_ (.Y(_08103_),
    .A(_07215_),
    .B(_08102_));
 sg13g2_o21ai_1 _27340_ (.B1(_09121_),
    .Y(_08104_),
    .A1(_07216_),
    .A2(_08103_));
 sg13g2_nand3_1 _27341_ (.B(_07215_),
    .C(_08102_),
    .A(net1055),
    .Y(_08105_));
 sg13g2_a21oi_1 _27342_ (.A1(_08104_),
    .A2(_08105_),
    .Y(_02586_),
    .B1(net644));
 sg13g2_nand2b_1 _27343_ (.Y(_08106_),
    .B(_09225_),
    .A_N(\cpu.spi.r_ready ));
 sg13g2_nor3_1 _27344_ (.A(net1055),
    .B(_09239_),
    .C(_08083_),
    .Y(_08107_));
 sg13g2_nor2_1 _27345_ (.A(_08103_),
    .B(_08107_),
    .Y(_08108_));
 sg13g2_nand3b_1 _27346_ (.B(_09172_),
    .C(_08108_),
    .Y(_08109_),
    .A_N(_09236_));
 sg13g2_a21oi_1 _27347_ (.A1(_08106_),
    .A2(_08109_),
    .Y(_08110_),
    .B1(net1055));
 sg13g2_nor2_1 _27348_ (.A(\cpu.spi.r_ready ),
    .B(_08108_),
    .Y(_08111_));
 sg13g2_o21ai_1 _27349_ (.B1(net694),
    .Y(_02601_),
    .A1(_08110_),
    .A2(_08111_));
 sg13g2_nand2_1 _27350_ (.Y(_08112_),
    .A(_09215_),
    .B(_08068_));
 sg13g2_nand2_1 _27351_ (.Y(_08113_),
    .A(\cpu.spi.r_searching ),
    .B(_08112_));
 sg13g2_a21oi_1 _27352_ (.A1(_09085_),
    .A2(_09144_),
    .Y(_08114_),
    .B1(_07006_));
 sg13g2_nand3_1 _27353_ (.B(_08068_),
    .C(_08114_),
    .A(_09215_),
    .Y(_08115_));
 sg13g2_a21oi_1 _27354_ (.A1(_08113_),
    .A2(_08115_),
    .Y(_02602_),
    .B1(net644));
 sg13g2_and2_1 _27355_ (.A(net427),
    .B(_07322_),
    .X(_08116_));
 sg13g2_buf_2 _27356_ (.A(_08116_),
    .X(_08117_));
 sg13g2_nand2_1 _27357_ (.Y(_08118_),
    .A(net865),
    .B(_08117_));
 sg13g2_nand2_1 _27358_ (.Y(_08119_),
    .A(net427),
    .B(_07322_));
 sg13g2_buf_2 _27359_ (.A(_08119_),
    .X(_08120_));
 sg13g2_nand2_1 _27360_ (.Y(_08121_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08120_));
 sg13g2_nand3_1 _27361_ (.B(_08118_),
    .C(_08121_),
    .A(net715),
    .Y(_02624_));
 sg13g2_and2_1 _27362_ (.A(_04918_),
    .B(_07322_),
    .X(_08122_));
 sg13g2_buf_2 _27363_ (.A(_08122_),
    .X(_08123_));
 sg13g2_nand2_1 _27364_ (.Y(_08124_),
    .A(net898),
    .B(_08123_));
 sg13g2_nand2b_1 _27365_ (.Y(_08125_),
    .B(_09891_),
    .A_N(_08123_));
 sg13g2_a21oi_1 _27366_ (.A1(_08124_),
    .A2(_08125_),
    .Y(_02625_),
    .B1(net644));
 sg13g2_nand2_1 _27367_ (.Y(_08126_),
    .A(net1044),
    .B(_08123_));
 sg13g2_nand2b_1 _27368_ (.Y(_08127_),
    .B(\cpu.uart.r_div_value[11] ),
    .A_N(_08123_));
 sg13g2_a21oi_1 _27369_ (.A1(_08126_),
    .A2(_08127_),
    .Y(_02626_),
    .B1(net644));
 sg13g2_nand2_1 _27370_ (.Y(_08128_),
    .A(net1046),
    .B(_08117_));
 sg13g2_nand2_1 _27371_ (.Y(_08129_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27372_ (.A1(_08128_),
    .A2(_08129_),
    .Y(_02627_),
    .B1(net644));
 sg13g2_nand2_1 _27373_ (.Y(_08130_),
    .A(net1045),
    .B(_08117_));
 sg13g2_nand2_1 _27374_ (.Y(_08131_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27375_ (.A1(_08130_),
    .A2(_08131_),
    .Y(_02628_),
    .B1(net644));
 sg13g2_nand2_1 _27376_ (.Y(_08132_),
    .A(_10008_),
    .B(_08117_));
 sg13g2_nand2_1 _27377_ (.Y(_08133_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27378_ (.A1(_08132_),
    .A2(_08133_),
    .Y(_02629_),
    .B1(_08062_));
 sg13g2_nand2_1 _27379_ (.Y(_08134_),
    .A(net1043),
    .B(_08117_));
 sg13g2_nand2_1 _27380_ (.Y(_08135_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27381_ (.A1(_08134_),
    .A2(_08135_),
    .Y(_02630_),
    .B1(_08062_));
 sg13g2_nand2_1 _27382_ (.Y(_08136_),
    .A(net1042),
    .B(_08117_));
 sg13g2_nand2_1 _27383_ (.Y(_08137_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27384_ (.A1(_08136_),
    .A2(_08137_),
    .Y(_02631_),
    .B1(net655));
 sg13g2_nand2_1 _27385_ (.Y(_08138_),
    .A(net1119),
    .B(_08117_));
 sg13g2_nand2_1 _27386_ (.Y(_08139_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27387_ (.A1(_08138_),
    .A2(_08139_),
    .Y(_02632_),
    .B1(net655));
 sg13g2_nand2_1 _27388_ (.Y(_08140_),
    .A(net1118),
    .B(_08117_));
 sg13g2_nand2_1 _27389_ (.Y(_08141_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08120_));
 sg13g2_a21oi_1 _27390_ (.A1(_08140_),
    .A2(_08141_),
    .Y(_02633_),
    .B1(net655));
 sg13g2_nand2_1 _27391_ (.Y(_08142_),
    .A(net1047),
    .B(_08123_));
 sg13g2_nand2b_1 _27392_ (.Y(_08143_),
    .B(\cpu.uart.r_div_value[8] ),
    .A_N(_08123_));
 sg13g2_a21oi_1 _27393_ (.A1(_08142_),
    .A2(_08143_),
    .Y(_02634_),
    .B1(net655));
 sg13g2_nand2_1 _27394_ (.Y(_08144_),
    .A(net1046),
    .B(_08123_));
 sg13g2_nand2b_1 _27395_ (.Y(_08145_),
    .B(\cpu.uart.r_div_value[9] ),
    .A_N(_08123_));
 sg13g2_a21oi_1 _27396_ (.A1(_08144_),
    .A2(_08145_),
    .Y(_02635_),
    .B1(net655));
 sg13g2_nand3_1 _27397_ (.B(_04891_),
    .C(_07322_),
    .A(net1046),
    .Y(_08146_));
 sg13g2_nand3_1 _27398_ (.B(_08337_),
    .C(_07320_),
    .A(_11843_),
    .Y(_08147_));
 sg13g2_or4_1 _27399_ (.A(net1058),
    .B(_09145_),
    .C(net781),
    .D(_08147_),
    .X(_08148_));
 sg13g2_nand4_1 _27400_ (.B(net802),
    .C(_08146_),
    .A(_09128_),
    .Y(_08149_),
    .D(_08148_));
 sg13g2_nand2b_1 _27401_ (.Y(_02659_),
    .B(_08149_),
    .A_N(net173));
 sg13g2_and2_1 _27402_ (.A(net472),
    .B(_07322_),
    .X(_08150_));
 sg13g2_buf_1 _27403_ (.A(_08150_),
    .X(_08151_));
 sg13g2_mux2_1 _27404_ (.A0(\cpu.uart.r_r_invert ),
    .A1(_09996_),
    .S(_08151_),
    .X(_08152_));
 sg13g2_and2_1 _27405_ (.A(net682),
    .B(_08152_),
    .X(_02660_));
 sg13g2_a21oi_1 _27406_ (.A1(_07305_),
    .A2(_09869_),
    .Y(_08153_),
    .B1(net1085));
 sg13g2_a21oi_1 _27407_ (.A1(_07306_),
    .A2(_09869_),
    .Y(_08154_),
    .B1(_07380_));
 sg13g2_a221oi_1 _27408_ (.B2(_08153_),
    .C1(_08154_),
    .B1(_07304_),
    .A1(net939),
    .Y(_08155_),
    .A2(_07299_));
 sg13g2_a21oi_1 _27409_ (.A1(_07297_),
    .A2(_08155_),
    .Y(_08156_),
    .B1(_07377_));
 sg13g2_buf_2 _27410_ (.A(_08156_),
    .X(_08157_));
 sg13g2_o21ai_1 _27411_ (.B1(_08157_),
    .Y(_08158_),
    .A1(net939),
    .A2(_07380_));
 sg13g2_xnor2_1 _27412_ (.Y(_08159_),
    .A(_07306_),
    .B(_08158_));
 sg13g2_nor2_1 _27413_ (.A(net648),
    .B(_08159_),
    .Y(_02663_));
 sg13g2_o21ai_1 _27414_ (.B1(_08157_),
    .Y(_08160_),
    .A1(_07305_),
    .A2(net940));
 sg13g2_nand2_1 _27415_ (.Y(_08161_),
    .A(net1084),
    .B(_08160_));
 sg13g2_nand2b_1 _27416_ (.Y(_08162_),
    .B(net939),
    .A_N(net940));
 sg13g2_o21ai_1 _27417_ (.B1(_08162_),
    .Y(_08163_),
    .A1(net939),
    .A2(_07379_));
 sg13g2_nand3_1 _27418_ (.B(_08157_),
    .C(_08163_),
    .A(_07378_),
    .Y(_08164_));
 sg13g2_a21oi_1 _27419_ (.A1(_08161_),
    .A2(_08164_),
    .Y(_02664_),
    .B1(net655));
 sg13g2_nand2_1 _27420_ (.Y(_08165_),
    .A(_07305_),
    .B(net1084));
 sg13g2_nor3_1 _27421_ (.A(net939),
    .B(net940),
    .C(_08165_),
    .Y(_08166_));
 sg13g2_o21ai_1 _27422_ (.B1(_08157_),
    .Y(_08167_),
    .A1(net940),
    .A2(_07388_));
 sg13g2_a22oi_1 _27423_ (.Y(_08168_),
    .B1(_08167_),
    .B2(net939),
    .A2(_08166_),
    .A1(_08157_));
 sg13g2_nor2_1 _27424_ (.A(net712),
    .B(_08168_),
    .Y(_02665_));
 sg13g2_a21oi_1 _27425_ (.A1(_07388_),
    .A2(_08157_),
    .Y(_08169_),
    .B1(_07300_));
 sg13g2_nor2b_1 _27426_ (.A(_07303_),
    .B_N(net1084),
    .Y(_08170_));
 sg13g2_a21oi_1 _27427_ (.A1(_08157_),
    .A2(_08170_),
    .Y(_08171_),
    .B1(_06799_));
 sg13g2_nor2b_1 _27428_ (.A(_08169_),
    .B_N(_08171_),
    .Y(_02666_));
 sg13g2_nand2b_1 _27429_ (.Y(_08172_),
    .B(_07334_),
    .A_N(_09127_));
 sg13g2_nor2_1 _27430_ (.A(net937),
    .B(_07399_),
    .Y(_08173_));
 sg13g2_a21oi_1 _27431_ (.A1(_09987_),
    .A2(_04891_),
    .Y(_08174_),
    .B1(net430));
 sg13g2_o21ai_1 _27432_ (.B1(net595),
    .Y(_08175_),
    .A1(_00204_),
    .A2(net534));
 sg13g2_nand3_1 _27433_ (.B(_07420_),
    .C(_08175_),
    .A(_09362_),
    .Y(_08176_));
 sg13g2_o21ai_1 _27434_ (.B1(_08176_),
    .Y(_08177_),
    .A1(_07399_),
    .A2(_08174_));
 sg13g2_nand2_1 _27435_ (.Y(_08178_),
    .A(_07322_),
    .B(_08177_));
 sg13g2_a22oi_1 _27436_ (.Y(_08179_),
    .B1(_08178_),
    .B2(_09127_),
    .A2(_08173_),
    .A1(_08172_));
 sg13g2_nor2_1 _27437_ (.A(net712),
    .B(_08179_),
    .Y(_02668_));
 sg13g2_nand2_1 _27438_ (.Y(_08180_),
    .A(net1047),
    .B(_08151_));
 sg13g2_nand2b_1 _27439_ (.Y(_08181_),
    .B(\cpu.uart.r_x_invert ),
    .A_N(_08151_));
 sg13g2_a21oi_1 _27440_ (.A1(_08180_),
    .A2(_08181_),
    .Y(_02669_),
    .B1(net655));
 sg13g2_and2_1 _27441_ (.A(_07325_),
    .B(_07401_),
    .X(_08182_));
 sg13g2_o21ai_1 _27442_ (.B1(_08182_),
    .Y(_08183_),
    .A1(_07334_),
    .A2(_07409_));
 sg13g2_and3_1 _27443_ (.X(_08184_),
    .A(_07424_),
    .B(_07319_),
    .C(_07323_));
 sg13g2_a21oi_1 _27444_ (.A1(net936),
    .A2(_07425_),
    .Y(_08185_),
    .B1(_08184_));
 sg13g2_o21ai_1 _27445_ (.B1(_07414_),
    .Y(_08186_),
    .A1(_07338_),
    .A2(_08185_));
 sg13g2_buf_1 _27446_ (.A(_08186_),
    .X(_08187_));
 sg13g2_a21oi_1 _27447_ (.A1(_07323_),
    .A2(_07420_),
    .Y(_08188_),
    .B1(_08187_));
 sg13g2_mux2_1 _27448_ (.A0(net937),
    .A1(_08183_),
    .S(_08188_),
    .X(_08189_));
 sg13g2_and2_1 _27449_ (.A(net682),
    .B(_08189_),
    .X(_02672_));
 sg13g2_a21oi_1 _27450_ (.A1(net938),
    .A2(_07329_),
    .Y(_08190_),
    .B1(_07325_));
 sg13g2_o21ai_1 _27451_ (.B1(net1083),
    .Y(_08191_),
    .A1(_08187_),
    .A2(_08190_));
 sg13g2_inv_1 _27452_ (.Y(_08192_),
    .A(_08187_));
 sg13g2_nand3_1 _27453_ (.B(_08192_),
    .C(_08182_),
    .A(_07337_),
    .Y(_08193_));
 sg13g2_a21oi_1 _27454_ (.A1(_08191_),
    .A2(_08193_),
    .Y(_02673_),
    .B1(net655));
 sg13g2_a21oi_1 _27455_ (.A1(_07319_),
    .A2(_08192_),
    .Y(_08194_),
    .B1(net936));
 sg13g2_nand2b_1 _27456_ (.Y(_08195_),
    .B(_07334_),
    .A_N(_07409_));
 sg13g2_nand3_1 _27457_ (.B(_08192_),
    .C(_08195_),
    .A(_07315_),
    .Y(_08196_));
 sg13g2_nand3_1 _27458_ (.B(_07319_),
    .C(_07414_),
    .A(net936),
    .Y(_08197_));
 sg13g2_nand3_1 _27459_ (.B(_08196_),
    .C(_08197_),
    .A(net802),
    .Y(_08198_));
 sg13g2_nor2_1 _27460_ (.A(_08194_),
    .B(_08198_),
    .Y(_02674_));
 sg13g2_a21oi_1 _27461_ (.A1(_07319_),
    .A2(_08195_),
    .Y(_08199_),
    .B1(_07329_));
 sg13g2_o21ai_1 _27462_ (.B1(_07315_),
    .Y(_08200_),
    .A1(_08187_),
    .A2(_08199_));
 sg13g2_a21oi_1 _27463_ (.A1(_08197_),
    .A2(_08200_),
    .Y(_02675_),
    .B1(_07534_));
 sg13g2_nand2_1 _27464_ (.Y(\cpu.ex.genblk3.c_supmode ),
    .A(_07594_),
    .B(_07597_));
 sg13g2_nor2_1 _27465_ (.A(_08035_),
    .B(_08059_),
    .Y(_08201_));
 sg13g2_a22oi_1 _27466_ (.Y(_08202_),
    .B1(_09794_),
    .B2(_08201_),
    .A2(net626),
    .A1(_09790_));
 sg13g2_inv_1 _27467_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08202_));
 sg13g2_nor4_1 _27468_ (.A(_09788_),
    .B(_09778_),
    .C(net626),
    .D(_08031_),
    .Y(_08203_));
 sg13g2_a22oi_1 _27469_ (.Y(_08204_),
    .B1(_08036_),
    .B2(_08203_),
    .A2(net626),
    .A1(_09787_));
 sg13g2_nor2_1 _27470_ (.A(net830),
    .B(_08204_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27471_ (.A(_08282_),
    .B(_08204_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27472_ (.S0(_04830_),
    .A0(_09107_),
    .A1(_09094_),
    .A2(_09089_),
    .A3(_09112_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08205_));
 sg13g2_mux4_1 _27473_ (.S0(_04830_),
    .A0(_09091_),
    .A1(_09114_),
    .A2(_09100_),
    .A3(_09109_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08206_));
 sg13g2_mux2_1 _27474_ (.A0(_08205_),
    .A1(_08206_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27475_ (.S0(_04812_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_05269_),
    .X(_08207_));
 sg13g2_mux4_1 _27476_ (.S0(_04812_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_05269_),
    .X(_08208_));
 sg13g2_nor2b_1 _27477_ (.A(_05351_),
    .B_N(_08208_),
    .Y(_08209_));
 sg13g2_a21oi_1 _27478_ (.A1(_05351_),
    .A2(_08207_),
    .Y(_08210_),
    .B1(_08209_));
 sg13g2_nand2b_1 _27479_ (.Y(_08211_),
    .B(net1078),
    .A_N(_04812_));
 sg13g2_nand3_1 _27480_ (.B(_05269_),
    .C(net1081),
    .A(_04812_),
    .Y(_08212_));
 sg13g2_o21ai_1 _27481_ (.B1(_08212_),
    .Y(_08213_),
    .A1(_05269_),
    .A2(_08211_));
 sg13g2_nand3_1 _27482_ (.B(_00161_),
    .C(_08213_),
    .A(_05389_),
    .Y(_08214_));
 sg13g2_o21ai_1 _27483_ (.B1(_08214_),
    .Y(net16),
    .A1(_05389_),
    .A2(_08210_));
 sg13g2_mux4_1 _27484_ (.S0(_05504_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_05538_),
    .X(_08215_));
 sg13g2_mux4_1 _27485_ (.S0(_05504_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_05538_),
    .X(_08216_));
 sg13g2_nor2b_1 _27486_ (.A(_05630_),
    .B_N(_08216_),
    .Y(_08217_));
 sg13g2_a21oi_1 _27487_ (.A1(_05630_),
    .A2(_08215_),
    .Y(_08218_),
    .B1(_08217_));
 sg13g2_nand2b_1 _27488_ (.Y(_08219_),
    .B(net1078),
    .A_N(_05504_));
 sg13g2_nand3_1 _27489_ (.B(_05538_),
    .C(net1081),
    .A(_05504_),
    .Y(_08220_));
 sg13g2_o21ai_1 _27490_ (.B1(_08220_),
    .Y(_08221_),
    .A1(_05538_),
    .A2(_08219_));
 sg13g2_nand3_1 _27491_ (.B(_00160_),
    .C(_08221_),
    .A(_05018_),
    .Y(_08222_));
 sg13g2_o21ai_1 _27492_ (.B1(_08222_),
    .Y(net17),
    .A1(_05018_),
    .A2(_08218_));
 sg13g2_mux4_1 _27493_ (.S0(_04813_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_06398_),
    .X(_08223_));
 sg13g2_mux4_1 _27494_ (.S0(_04813_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(_07406_),
    .A2(net1101),
    .A3(net1102),
    .S1(_06398_),
    .X(_08224_));
 sg13g2_nor2b_1 _27495_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08224_),
    .Y(_08225_));
 sg13g2_a21oi_1 _27496_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08223_),
    .Y(_08226_),
    .B1(_08225_));
 sg13g2_nand2b_1 _27497_ (.Y(_08227_),
    .B(net1078),
    .A_N(_04813_));
 sg13g2_nand3_1 _27498_ (.B(net1081),
    .C(_06398_),
    .A(_04813_),
    .Y(_08228_));
 sg13g2_o21ai_1 _27499_ (.B1(_08228_),
    .Y(_08229_),
    .A1(_06398_),
    .A2(_08227_));
 sg13g2_nand3_1 _27500_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08229_),
    .A(_00094_),
    .Y(_08230_));
 sg13g2_o21ai_1 _27501_ (.B1(_08230_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08226_));
 sg13g2_mux4_1 _27502_ (.S0(_05505_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_06399_),
    .X(_08231_));
 sg13g2_mux4_1 _27503_ (.S0(_05505_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_06399_),
    .X(_08232_));
 sg13g2_nor2b_1 _27504_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08232_),
    .Y(_08233_));
 sg13g2_a21oi_1 _27505_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08231_),
    .Y(_08234_),
    .B1(_08233_));
 sg13g2_nand2b_1 _27506_ (.Y(_08235_),
    .B(net1078),
    .A_N(_05505_));
 sg13g2_nand3_1 _27507_ (.B(_06399_),
    .C(net1081),
    .A(_05505_),
    .Y(_08236_));
 sg13g2_o21ai_1 _27508_ (.B1(_08236_),
    .Y(_08237_),
    .A1(_06399_),
    .A2(_08235_));
 sg13g2_nand3_1 _27509_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08237_),
    .A(_00131_),
    .Y(_08238_));
 sg13g2_o21ai_1 _27510_ (.B1(_08238_),
    .Y(net19),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08234_));
 sg13g2_xor2_1 _27511_ (.B(clknet_leaf_76_clk),
    .A(\cpu.r_clk_invert ),
    .X(net22));
 sg13g2_mux4_1 _27512_ (.S0(_05498_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_06402_),
    .X(_08239_));
 sg13g2_mux4_1 _27513_ (.S0(_05498_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_06402_),
    .X(_08240_));
 sg13g2_nor2b_1 _27514_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08240_),
    .Y(_08241_));
 sg13g2_a21oi_1 _27515_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08239_),
    .Y(_08242_),
    .B1(_08241_));
 sg13g2_nand2b_1 _27516_ (.Y(_08243_),
    .B(net1078),
    .A_N(_05498_));
 sg13g2_nand3_1 _27517_ (.B(net1081),
    .C(_06402_),
    .A(_05498_),
    .Y(_08244_));
 sg13g2_o21ai_1 _27518_ (.B1(_08244_),
    .Y(_08245_),
    .A1(_06402_),
    .A2(_08243_));
 sg13g2_nand3_1 _27519_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08245_),
    .A(_00134_),
    .Y(_08246_));
 sg13g2_o21ai_1 _27520_ (.B1(_08246_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08242_));
 sg13g2_mux4_1 _27521_ (.S0(_04816_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_06407_),
    .X(_08247_));
 sg13g2_mux4_1 _27522_ (.S0(_04816_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_06407_),
    .X(_08248_));
 sg13g2_nor2b_1 _27523_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08248_),
    .Y(_08249_));
 sg13g2_a21oi_1 _27524_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08247_),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_nand2b_1 _27525_ (.Y(_08251_),
    .B(net1078),
    .A_N(_04816_));
 sg13g2_nand3_1 _27526_ (.B(net1081),
    .C(_06407_),
    .A(_04816_),
    .Y(_08252_));
 sg13g2_o21ai_1 _27527_ (.B1(_08252_),
    .Y(_08253_),
    .A1(_06407_),
    .A2(_08251_));
 sg13g2_nand3_1 _27528_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08253_),
    .A(_00096_),
    .Y(_08254_));
 sg13g2_o21ai_1 _27529_ (.B1(_08254_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08250_));
 sg13g2_mux4_1 _27530_ (.S0(_05503_),
    .A0(net1103),
    .A1(net1104),
    .A2(net1080),
    .A3(net1079),
    .S1(_06409_),
    .X(_08255_));
 sg13g2_mux4_1 _27531_ (.S0(_05503_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1082),
    .A2(net1101),
    .A3(net1102),
    .S1(_06409_),
    .X(_08256_));
 sg13g2_nor2b_1 _27532_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08256_),
    .Y(_08257_));
 sg13g2_a21oi_1 _27533_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08255_),
    .Y(_08258_),
    .B1(_08257_));
 sg13g2_nand2b_1 _27534_ (.Y(_08259_),
    .B(net1078),
    .A_N(_05503_));
 sg13g2_nand3_1 _27535_ (.B(net1081),
    .C(_06409_),
    .A(_05503_),
    .Y(_08260_));
 sg13g2_o21ai_1 _27536_ (.B1(_08260_),
    .Y(_08261_),
    .A1(_06409_),
    .A2(_08259_));
 sg13g2_nand3_1 _27537_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08261_),
    .A(_00133_),
    .Y(_08262_));
 sg13g2_o21ai_1 _27538_ (.B1(_08262_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08258_));
 sg13g2_mux4_1 _27539_ (.S0(_04824_),
    .A0(net1103),
    .A1(_11851_),
    .A2(net1080),
    .A3(_08095_),
    .S1(_07936_),
    .X(_08263_));
 sg13g2_mux4_1 _27540_ (.S0(_04824_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1082),
    .A2(_11877_),
    .A3(_11860_),
    .S1(_07936_),
    .X(_08264_));
 sg13g2_nor2b_1 _27541_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08264_),
    .Y(_08265_));
 sg13g2_a21oi_1 _27542_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08263_),
    .Y(_08266_),
    .B1(_08265_));
 sg13g2_nand2b_1 _27543_ (.Y(_08267_),
    .B(net1078),
    .A_N(_04824_));
 sg13g2_nand3_1 _27544_ (.B(_08028_),
    .C(_07936_),
    .A(_04824_),
    .Y(_08268_));
 sg13g2_o21ai_1 _27545_ (.B1(_08268_),
    .Y(_08269_),
    .A1(_07936_),
    .A2(_08267_));
 sg13g2_nand3_1 _27546_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08269_),
    .A(_00095_),
    .Y(_08270_));
 sg13g2_o21ai_1 _27547_ (.B1(_08270_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08266_));
 sg13g2_mux4_1 _27548_ (.S0(_05500_),
    .A0(_11858_),
    .A1(net1104),
    .A2(_08079_),
    .A3(net1079),
    .S1(_06414_),
    .X(_08271_));
 sg13g2_mux4_1 _27549_ (.S0(_05500_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1082),
    .A2(_11877_),
    .A3(_11860_),
    .S1(_06414_),
    .X(_08272_));
 sg13g2_nor2b_1 _27550_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08272_),
    .Y(_08273_));
 sg13g2_a21oi_1 _27551_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08271_),
    .Y(_08274_),
    .B1(_08273_));
 sg13g2_nand2b_1 _27552_ (.Y(_08275_),
    .B(_08097_),
    .A_N(_05500_));
 sg13g2_nand3_1 _27553_ (.B(net1081),
    .C(_06414_),
    .A(_05500_),
    .Y(_08276_));
 sg13g2_o21ai_1 _27554_ (.B1(_08276_),
    .Y(_08277_),
    .A1(_06414_),
    .A2(_08275_));
 sg13g2_nand3_1 _27555_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08277_),
    .A(_00132_),
    .Y(_08278_));
 sg13g2_o21ai_1 _27556_ (.B1(_08278_),
    .Y(net27),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08274_));
 sg13g2_dfrbp_1 _27557_ (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1138),
    .D(_00313_),
    .Q_N(_14891_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27558_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1139),
    .D(_00314_),
    .Q_N(_14890_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27559_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1140),
    .D(_00315_),
    .Q_N(_14889_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27560_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1141),
    .D(_00316_),
    .Q_N(_14888_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27561_ (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1142),
    .D(_00317_),
    .Q_N(_14887_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27563_ (.A(net7),
    .X(net5));
 sg13g2_buf_1 _27564_ (.A(net7),
    .X(net6));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1143),
    .D(_00318_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1144),
    .D(_00319_),
    .Q_N(_00091_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1145),
    .D(_00320_),
    .Q_N(_00101_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1146),
    .D(_00321_),
    .Q_N(_00111_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1147),
    .D(_00322_),
    .Q_N(_00117_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1148),
    .D(_00323_),
    .Q_N(_00128_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1149),
    .D(_00324_),
    .Q_N(_00139_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1150),
    .D(_00325_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1151),
    .D(_00326_),
    .Q_N(_00299_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1152),
    .D(_00327_),
    .Q_N(_00309_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1153),
    .D(_00328_),
    .Q_N(_00099_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1154),
    .D(_00329_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1155),
    .D(_00330_),
    .Q_N(_00109_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1156),
    .D(_00331_),
    .Q_N(_00115_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1157),
    .D(_00332_),
    .Q_N(_00126_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1158),
    .D(_00333_),
    .Q_N(_00137_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1159),
    .D(_00334_),
    .Q_N(_00295_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1160),
    .D(_00335_),
    .Q_N(_00300_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1161),
    .D(_00336_),
    .Q_N(_00310_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1162),
    .D(_00337_),
    .Q_N(_00100_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1163),
    .D(_00338_),
    .Q_N(_00110_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1164),
    .D(_00339_),
    .Q_N(_00116_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1165),
    .D(_00340_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1166),
    .D(_00341_),
    .Q_N(_00127_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1167),
    .D(_00342_),
    .Q_N(_00138_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1168),
    .D(_00343_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1169),
    .D(_00344_),
    .Q_N(_00108_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1170),
    .D(_00345_),
    .Q_N(_00114_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1171),
    .D(_00346_),
    .Q_N(_00125_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1172),
    .D(_00347_),
    .Q_N(_00136_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1173),
    .D(_00348_),
    .Q_N(_00296_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1174),
    .D(_00349_),
    .Q_N(_00301_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1175),
    .D(_00350_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1176),
    .D(_00351_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1177),
    .D(_00352_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1178),
    .D(_00353_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1179),
    .D(_00354_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1180),
    .D(_00355_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1181),
    .D(_00356_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1182),
    .D(_00357_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1183),
    .D(_00358_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1184),
    .D(_00359_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1185),
    .D(_00360_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1186),
    .D(_00361_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1187),
    .D(_00362_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1188),
    .D(_00363_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1189),
    .D(_00364_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1190),
    .D(_00365_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1191),
    .D(_00366_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1192),
    .D(_00367_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1193),
    .D(_00368_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1194),
    .D(_00369_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1195),
    .D(_00370_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1196),
    .D(_00371_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1197),
    .D(_00372_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1198),
    .D(_00373_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1199),
    .D(_00374_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1200),
    .D(_00375_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1201),
    .D(_00376_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1202),
    .D(_00377_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1203),
    .D(_00378_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1204),
    .D(_00379_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1205),
    .D(_00380_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1206),
    .D(_00381_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1207),
    .D(_00382_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1208),
    .D(_00383_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1209),
    .D(_00384_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1210),
    .D(_00385_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1211),
    .D(_00386_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1212),
    .D(_00387_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1213),
    .D(_00388_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1214),
    .D(_00389_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1215),
    .D(_00390_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1216),
    .D(_00391_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1217),
    .D(_00392_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1218),
    .D(_00393_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1219),
    .D(_00394_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1220),
    .D(_00395_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1221),
    .D(_00396_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1222),
    .D(_00397_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1223),
    .D(_00398_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1224),
    .D(_00399_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1225),
    .D(_00400_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1226),
    .D(_00401_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1227),
    .D(_00402_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1228),
    .D(_00403_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1229),
    .D(_00404_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1230),
    .D(_00405_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1231),
    .D(_00406_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1232),
    .D(_00407_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1233),
    .D(_00408_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1234),
    .D(_00409_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1235),
    .D(_00410_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1236),
    .D(_00411_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1237),
    .D(_00412_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1238),
    .D(_00413_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1239),
    .D(_00414_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1240),
    .D(_00415_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1241),
    .D(_00416_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1242),
    .D(_00417_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1243),
    .D(_00418_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1244),
    .D(_00419_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1245),
    .D(_00420_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1246),
    .D(_00421_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1247),
    .D(_00422_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1248),
    .D(_00423_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1249),
    .D(_00424_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1250),
    .D(_00425_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1251),
    .D(_00426_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1252),
    .D(_00427_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1253),
    .D(_00428_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1254),
    .D(_00429_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1255),
    .D(_00430_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1256),
    .D(_00431_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1257),
    .D(_00432_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1258),
    .D(_00433_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1259),
    .D(_00434_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1260),
    .D(_00435_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1261),
    .D(_00436_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1262),
    .D(_00437_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1263),
    .D(_00438_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1264),
    .D(_00439_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1265),
    .D(_00440_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1266),
    .D(_00441_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1267),
    .D(_00442_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1268),
    .D(_00443_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1269),
    .D(_00444_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1270),
    .D(_00445_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1271),
    .D(_00446_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1272),
    .D(_00447_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1273),
    .D(_00448_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1274),
    .D(_00449_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1275),
    .D(_00450_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1276),
    .D(_00451_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1277),
    .D(_00452_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1278),
    .D(_00453_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1279),
    .D(_00454_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1280),
    .D(_00455_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1281),
    .D(_00456_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1282),
    .D(_00457_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1283),
    .D(_00458_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1284),
    .D(_00459_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1285),
    .D(_00460_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1286),
    .D(_00461_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1287),
    .D(_00462_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1288),
    .D(_00463_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1289),
    .D(_00464_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1290),
    .D(_00465_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1291),
    .D(_00466_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1292),
    .D(_00467_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1293),
    .D(_00468_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1294),
    .D(_00469_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1295),
    .D(_00470_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1296),
    .D(_00471_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1297),
    .D(_00472_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1298),
    .D(_00473_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1299),
    .D(_00474_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1300),
    .D(_00475_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1301),
    .D(_00476_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1302),
    .D(_00477_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1303),
    .D(_00478_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1304),
    .D(_00479_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1305),
    .D(_00480_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1306),
    .D(_00481_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1307),
    .D(_00482_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1308),
    .D(_00483_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1309),
    .D(_00484_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1310),
    .D(_00485_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1311),
    .D(_00486_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1312),
    .D(_00487_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1313),
    .D(_00488_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1314),
    .D(_00489_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1315),
    .D(_00490_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1316),
    .D(_00491_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1317),
    .D(_00492_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1318),
    .D(_00493_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1319),
    .D(_00494_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1320),
    .D(_00495_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1321),
    .D(_00496_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1322),
    .D(_00497_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1323),
    .D(_00498_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1324),
    .D(_00499_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1325),
    .D(_00500_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1326),
    .D(_00501_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1327),
    .D(_00502_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1328),
    .D(_00503_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1329),
    .D(_00504_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1330),
    .D(_00505_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1331),
    .D(_00506_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1332),
    .D(_00507_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1333),
    .D(_00508_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1334),
    .D(_00509_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1335),
    .D(_00510_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1336),
    .D(_00511_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1337),
    .D(_00512_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1338),
    .D(_00513_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1339),
    .D(_00514_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1340),
    .D(_00515_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1341),
    .D(_00516_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1342),
    .D(_00517_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1343),
    .D(_00518_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1344),
    .D(_00519_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1345),
    .D(_00520_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1346),
    .D(_00521_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1347),
    .D(_00522_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1348),
    .D(_00523_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1349),
    .D(_00524_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1350),
    .D(_00525_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1351),
    .D(_00526_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1352),
    .D(_00527_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1353),
    .D(_00528_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1354),
    .D(_00529_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1355),
    .D(_00530_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1356),
    .D(_00531_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1357),
    .D(_00532_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1358),
    .D(_00533_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1359),
    .D(_00534_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1360),
    .D(_00535_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1361),
    .D(_00536_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1362),
    .D(_00537_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1363),
    .D(_00538_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1364),
    .D(_00539_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1365),
    .D(_00540_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1366),
    .D(_00541_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1367),
    .D(_00542_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1368),
    .D(_00543_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1369),
    .D(_00544_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1370),
    .D(_00545_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1371),
    .D(_00546_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1372),
    .D(_00547_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1373),
    .D(_00548_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1374),
    .D(_00549_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1375),
    .D(_00550_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1376),
    .D(_00551_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1377),
    .D(_00552_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1378),
    .D(_00553_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1379),
    .D(_00554_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1380),
    .D(_00555_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1381),
    .D(_00556_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1382),
    .D(_00557_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1383),
    .D(_00558_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1384),
    .D(_00559_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1385),
    .D(_00560_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1386),
    .D(_00561_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1387),
    .D(_00562_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1388),
    .D(_00563_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1389),
    .D(_00564_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1390),
    .D(_00565_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1391),
    .D(_00566_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1392),
    .D(_00567_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1393),
    .D(_00568_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1394),
    .D(_00569_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1395),
    .D(_00570_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1396),
    .D(_00571_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1397),
    .D(_00572_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1398),
    .D(_00573_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1399),
    .D(_00574_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1400),
    .D(_00575_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1401),
    .D(_00576_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1402),
    .D(_00577_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1403),
    .D(_00578_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1404),
    .D(_00579_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1405),
    .D(_00580_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1406),
    .D(_00581_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1407),
    .D(_00582_),
    .Q_N(_00311_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1408),
    .D(_00583_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1409),
    .D(_00584_),
    .Q_N(_00257_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1410),
    .D(_00585_),
    .Q_N(_00210_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1411),
    .D(_00586_),
    .Q_N(_00226_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1412),
    .D(_00587_),
    .Q_N(_00227_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1413),
    .D(_00588_),
    .Q_N(_00228_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1414),
    .D(_00589_),
    .Q_N(_00229_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1415),
    .D(_00590_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1416),
    .D(_00591_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1417),
    .D(_00592_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1418),
    .D(_00593_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1419),
    .D(_00594_),
    .Q_N(_00231_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1420),
    .D(_00595_),
    .Q_N(_00212_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1421),
    .D(_00596_),
    .Q_N(_00214_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1422),
    .D(_00597_),
    .Q_N(_00216_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1423),
    .D(_00598_),
    .Q_N(_00218_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1424),
    .D(_00599_),
    .Q_N(_00220_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1425),
    .D(_00600_),
    .Q_N(_00222_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1426),
    .D(_00601_),
    .Q_N(_00223_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1427),
    .D(_00602_),
    .Q_N(_00224_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1428),
    .D(_00603_),
    .Q_N(_00225_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1429),
    .D(_00604_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1430),
    .D(_00605_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1431),
    .D(_00606_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1432),
    .D(_00607_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1433),
    .D(_00608_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1434),
    .D(_00609_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1435),
    .D(_00610_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1436),
    .D(_00611_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1437),
    .D(_00612_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1438),
    .D(_00613_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1439),
    .D(_00614_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1440),
    .D(_00615_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1441),
    .D(_00616_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1442),
    .D(_00617_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1443),
    .D(_00618_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1444),
    .D(_00619_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1445),
    .D(_00620_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1446),
    .D(_00621_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1447),
    .D(_00622_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1448),
    .D(_00623_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1449),
    .D(_00624_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1450),
    .D(_00625_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1451),
    .D(_00626_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1452),
    .D(_00627_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1453),
    .D(_00628_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1454),
    .D(_00629_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1455),
    .D(_00630_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1456),
    .D(_00631_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1457),
    .D(_00632_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1458),
    .D(_00633_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1459),
    .D(_00634_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1460),
    .D(_00635_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1461),
    .D(_00636_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1462),
    .D(_00637_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1463),
    .D(_00638_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1464),
    .D(_00639_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1465),
    .D(_00640_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1466),
    .D(_00641_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1467),
    .D(_00642_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1468),
    .D(_00643_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1469),
    .D(_00644_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1470),
    .D(_00645_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1471),
    .D(_00646_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1472),
    .D(_00647_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1473),
    .D(_00648_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1474),
    .D(_00649_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1475),
    .D(_00650_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1476),
    .D(_00651_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1477),
    .D(_00652_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1478),
    .D(_00653_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1479),
    .D(_00654_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1480),
    .D(_00655_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1481),
    .D(_00656_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1482),
    .D(_00657_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1483),
    .D(_00658_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1484),
    .D(_00659_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1485),
    .D(_00660_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1486),
    .D(_00661_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1487),
    .D(_00662_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1488),
    .D(_00663_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1489),
    .D(_00664_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1490),
    .D(_00665_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1491),
    .D(_00666_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1492),
    .D(_00667_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1493),
    .D(_00668_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1494),
    .D(_00669_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1495),
    .D(_00670_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1496),
    .D(_00671_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1497),
    .D(_00672_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1498),
    .D(_00673_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1499),
    .D(_00674_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1500),
    .D(_00675_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1501),
    .D(_00676_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1502),
    .D(_00677_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1503),
    .D(_00678_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1504),
    .D(_00679_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1505),
    .D(_00680_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1506),
    .D(_00681_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1507),
    .D(_00682_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1508),
    .D(_00683_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1509),
    .D(_00684_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1510),
    .D(_00685_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1511),
    .D(_00686_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1512),
    .D(_00687_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1513),
    .D(_00688_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1514),
    .D(_00689_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1515),
    .D(_00690_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1516),
    .D(_00691_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1517),
    .D(_00692_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1518),
    .D(_00693_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1519),
    .D(_00694_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1520),
    .D(_00695_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1521),
    .D(_00696_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1522),
    .D(_00697_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1523),
    .D(_00698_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1524),
    .D(_00699_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1525),
    .D(_00700_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1526),
    .D(_00701_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1527),
    .D(_00702_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1528),
    .D(_00703_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1529),
    .D(_00704_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1530),
    .D(_00705_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1531),
    .D(_00706_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1532),
    .D(_00707_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1533),
    .D(_00708_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1534),
    .D(_00709_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1535),
    .D(_00710_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1536),
    .D(_00711_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1537),
    .D(_00712_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1538),
    .D(_00713_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1539),
    .D(_00714_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1540),
    .D(_00715_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1541),
    .D(_00716_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1542),
    .D(_00717_),
    .Q_N(_14532_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1543),
    .D(_00718_),
    .Q_N(_14531_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1544),
    .D(_00719_),
    .Q_N(_14530_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1545),
    .D(_00720_),
    .Q_N(_14529_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1546),
    .D(_00721_),
    .Q_N(_14528_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1547),
    .D(_00722_),
    .Q_N(_14527_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1548),
    .D(_00723_),
    .Q_N(_14526_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1549),
    .D(_00724_),
    .Q_N(_14525_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1550),
    .D(_00725_),
    .Q_N(_14524_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1551),
    .D(_00726_),
    .Q_N(_14523_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1552),
    .D(_00727_),
    .Q_N(_14522_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1553),
    .D(_00728_),
    .Q_N(_14521_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1554),
    .D(_00729_),
    .Q_N(_14520_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1555),
    .D(_00730_),
    .Q_N(_14519_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1556),
    .D(_00731_),
    .Q_N(_14518_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1557),
    .D(_00732_),
    .Q_N(_14517_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1558),
    .D(_00733_),
    .Q_N(_14516_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1559),
    .D(_00734_),
    .Q_N(_14515_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1560),
    .D(_00735_),
    .Q_N(_14514_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1561),
    .D(_00736_),
    .Q_N(_14513_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1562),
    .D(_00737_),
    .Q_N(_14512_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1563),
    .D(_00738_),
    .Q_N(_14511_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1564),
    .D(_00739_),
    .Q_N(_14510_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1565),
    .D(_00740_),
    .Q_N(_14509_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1566),
    .D(_00741_),
    .Q_N(_14508_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1567),
    .D(_00742_),
    .Q_N(_14507_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1568),
    .D(_00743_),
    .Q_N(_14506_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1569),
    .D(_00744_),
    .Q_N(_14505_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1570),
    .D(_00745_),
    .Q_N(_14504_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1571),
    .D(_00746_),
    .Q_N(_14503_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1572),
    .D(_00747_),
    .Q_N(_14502_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1573),
    .D(_00748_),
    .Q_N(_00254_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1574),
    .D(_00749_),
    .Q_N(_14501_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1575),
    .D(_00750_),
    .Q_N(_14500_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1576),
    .D(_00751_),
    .Q_N(_14499_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1577),
    .D(_00752_),
    .Q_N(_14498_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1578),
    .D(_00753_),
    .Q_N(_14497_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1579),
    .D(_00754_),
    .Q_N(_14496_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1580),
    .D(_00755_),
    .Q_N(_14495_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1581),
    .D(_00756_),
    .Q_N(_14494_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1582),
    .D(_00757_),
    .Q_N(_14493_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1583),
    .D(_00758_),
    .Q_N(_14492_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1584),
    .D(_00759_),
    .Q_N(_14491_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1585),
    .D(_00760_),
    .Q_N(_14490_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1586),
    .D(_00761_),
    .Q_N(_14489_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1587),
    .D(_00762_),
    .Q_N(_14488_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1588),
    .D(_00763_),
    .Q_N(_14487_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1589),
    .D(_00764_),
    .Q_N(_14486_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1590),
    .D(_00765_),
    .Q_N(_14485_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1591),
    .D(_00766_),
    .Q_N(_14484_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1592),
    .D(_00767_),
    .Q_N(_14483_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1593),
    .D(_00768_),
    .Q_N(_14482_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1594),
    .D(_00769_),
    .Q_N(_14481_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1595),
    .D(_00770_),
    .Q_N(_00238_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1596),
    .D(_00771_),
    .Q_N(_14480_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1597),
    .D(_00772_),
    .Q_N(_14479_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1598),
    .D(_00773_),
    .Q_N(_14892_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1599),
    .D(_00011_),
    .Q_N(_14893_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1600),
    .D(_00012_),
    .Q_N(_14894_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1601),
    .D(_00013_),
    .Q_N(_14895_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1602),
    .D(_00014_),
    .Q_N(_14896_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1603),
    .D(_00015_),
    .Q_N(_14897_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1604),
    .D(_00016_),
    .Q_N(_14898_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1605),
    .D(_00017_),
    .Q_N(_14899_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1606),
    .D(_00018_),
    .Q_N(_14900_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1607),
    .D(_00019_),
    .Q_N(_14901_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1608),
    .D(_00020_),
    .Q_N(_14478_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1609),
    .D(_00774_),
    .Q_N(_14477_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1610),
    .D(_00775_),
    .Q_N(_14476_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1611),
    .D(_00776_),
    .Q_N(_14475_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1612),
    .D(_00777_),
    .Q_N(_14902_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1613),
    .D(_00052_),
    .Q_N(_14474_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1614),
    .D(_00778_),
    .Q_N(_14473_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1615),
    .D(_00779_),
    .Q_N(_14472_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1616),
    .D(_00780_),
    .Q_N(_14471_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1617),
    .D(_00781_),
    .Q_N(_14470_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1618),
    .D(_00782_),
    .Q_N(_14469_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1619),
    .D(_00783_),
    .Q_N(_14468_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1620),
    .D(_00784_),
    .Q_N(_14467_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1621),
    .D(_00785_),
    .Q_N(_14466_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1622),
    .D(_00786_),
    .Q_N(_14465_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1623),
    .D(_00787_),
    .Q_N(_00294_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1624),
    .D(_00788_),
    .Q_N(_14464_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1625),
    .D(_00789_),
    .Q_N(_00255_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1626),
    .D(_00790_),
    .Q_N(_14463_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1627),
    .D(_00791_),
    .Q_N(_14462_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1628),
    .D(_00792_),
    .Q_N(_00174_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1629),
    .D(_00793_),
    .Q_N(_14903_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1630),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00175_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1631),
    .D(_00794_),
    .Q_N(_14461_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1632),
    .D(_00795_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1633),
    .D(_00796_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1634),
    .D(_00797_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1635),
    .D(_00798_),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1636),
    .D(_00799_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1637),
    .D(_00800_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1638),
    .D(_00801_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1639),
    .D(_00802_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1640),
    .D(_00803_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1641),
    .D(_00804_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1642),
    .D(_00805_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1643),
    .D(_00806_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1644),
    .D(_00807_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1645),
    .D(_00808_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1646),
    .D(_00809_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1647),
    .D(_00810_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1648),
    .D(_00811_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1649),
    .D(_00812_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1650),
    .D(_00813_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1651),
    .D(_00814_),
    .Q_N(_14441_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1652),
    .D(_00815_),
    .Q_N(_14440_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1653),
    .D(_00816_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1654),
    .D(_00817_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1655),
    .D(_00818_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1656),
    .D(_00819_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1657),
    .D(_00820_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1658),
    .D(_00821_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1659),
    .D(_00822_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1660),
    .D(_00823_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1661),
    .D(_00824_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1662),
    .D(_00825_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1663),
    .D(_00826_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1664),
    .D(_00827_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1665),
    .D(_00828_),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1666),
    .D(_00829_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1667),
    .D(_00830_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1668),
    .D(_00831_),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1669),
    .D(_00832_),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1670),
    .D(_00833_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1671),
    .D(_00834_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1672),
    .D(_00835_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1673),
    .D(_00836_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1674),
    .D(_00837_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1675),
    .D(_00838_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1676),
    .D(_00839_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1677),
    .D(_00840_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1678),
    .D(_00841_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1679),
    .D(_00842_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1680),
    .D(_00843_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1681),
    .D(_00844_),
    .Q_N(_14411_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1682),
    .D(_00845_),
    .Q_N(_14410_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1683),
    .D(_00846_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1684),
    .D(_00847_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1685),
    .D(_00848_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1686),
    .D(_00849_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1687),
    .D(_00850_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1688),
    .D(_00851_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1689),
    .D(_00852_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1690),
    .D(_00853_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1691),
    .D(_00854_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1692),
    .D(_00855_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1693),
    .D(_00856_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1694),
    .D(_00857_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1695),
    .D(_00858_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1696),
    .D(_00859_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1697),
    .D(_00860_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1698),
    .D(_00861_),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1699),
    .D(_00862_),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1700),
    .D(_00863_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1701),
    .D(_00864_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1702),
    .D(_00865_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1703),
    .D(_00866_),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1704),
    .D(_00867_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1705),
    .D(_00868_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1706),
    .D(_00869_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1707),
    .D(_00870_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1708),
    .D(_00871_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1709),
    .D(_00872_),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1710),
    .D(_00873_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1711),
    .D(_00874_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1712),
    .D(_00875_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1713),
    .D(_00876_),
    .Q_N(_00248_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1714),
    .D(_00877_),
    .Q_N(_00249_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1715),
    .D(_00878_),
    .Q_N(_00250_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1716),
    .D(_00879_),
    .Q_N(_00251_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1717),
    .D(_00880_),
    .Q_N(_00252_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1718),
    .D(_00881_),
    .Q_N(_00253_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1719),
    .D(_00882_),
    .Q_N(_00239_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1720),
    .D(_00883_),
    .Q_N(_00240_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1721),
    .D(_00884_),
    .Q_N(_00241_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1722),
    .D(_00885_),
    .Q_N(_00242_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1723),
    .D(_00886_),
    .Q_N(_00243_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1724),
    .D(_00887_),
    .Q_N(_00244_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1725),
    .D(_00888_),
    .Q_N(_00245_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1726),
    .D(_00889_),
    .Q_N(_00246_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1727),
    .D(_00890_),
    .Q_N(_00247_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1728),
    .D(_00891_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1729),
    .D(_00892_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1730),
    .D(_00893_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1731),
    .D(_00894_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1732),
    .D(_00895_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1733),
    .D(_00896_),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1734),
    .D(_00897_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1735),
    .D(_00898_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1736),
    .D(_00899_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1737),
    .D(_00900_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1738),
    .D(_00901_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1739),
    .D(_00902_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1740),
    .D(_00903_),
    .Q_N(_14367_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1741),
    .D(_00904_),
    .Q_N(_14366_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1742),
    .D(_00905_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1743),
    .D(_00906_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1744),
    .D(_00907_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1745),
    .D(_00908_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1746),
    .D(_00909_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1747),
    .D(_00910_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1748),
    .D(_00911_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1749),
    .D(_00912_),
    .Q_N(_14358_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1750),
    .D(_00913_),
    .Q_N(_14357_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1751),
    .D(_00914_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1752),
    .D(_00915_),
    .Q_N(_14355_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1753),
    .D(_00916_),
    .Q_N(_14354_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1754),
    .D(_00917_),
    .Q_N(_14353_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1755),
    .D(_00918_),
    .Q_N(_14352_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1756),
    .D(_00919_),
    .Q_N(_14351_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1757),
    .D(_00920_),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1758),
    .D(_00921_),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1759),
    .D(_00922_),
    .Q_N(_14904_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1760),
    .D(_00053_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net1761),
    .D(_00923_),
    .Q_N(_14905_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1762),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1763),
    .D(_00924_),
    .Q_N(_14346_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1764),
    .D(_00925_),
    .Q_N(_14345_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1765),
    .D(_00926_),
    .Q_N(_14344_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1766),
    .D(_00927_),
    .Q_N(_14343_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1767),
    .D(_00928_),
    .Q_N(_14342_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1768),
    .D(_00929_),
    .Q_N(_14341_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1769),
    .D(_00930_),
    .Q_N(_14340_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1770),
    .D(_00931_),
    .Q_N(_14339_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1771),
    .D(_00932_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1772),
    .D(_00933_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1773),
    .D(_00934_),
    .Q_N(_14336_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1774),
    .D(_00935_),
    .Q_N(_14335_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1775),
    .D(_00936_),
    .Q_N(_14334_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1776),
    .D(_00937_),
    .Q_N(_14333_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1777),
    .D(_00938_),
    .Q_N(_14332_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1778),
    .D(_00939_),
    .Q_N(_00171_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1779),
    .D(_00940_),
    .Q_N(_14331_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1780),
    .D(_00941_),
    .Q_N(_14330_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1781),
    .D(_00942_),
    .Q_N(_14329_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1782),
    .D(_00943_),
    .Q_N(_00179_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1783),
    .D(_00944_),
    .Q_N(_14328_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1784),
    .D(_00945_),
    .Q_N(_14327_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1785),
    .D(_00946_),
    .Q_N(_14326_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1786),
    .D(_00947_),
    .Q_N(_14325_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1787),
    .D(_00948_),
    .Q_N(_14324_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1788),
    .D(_00949_),
    .Q_N(_14323_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1789),
    .D(_00950_),
    .Q_N(_14322_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1790),
    .D(_00951_),
    .Q_N(_14321_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1791),
    .D(_00952_),
    .Q_N(_14320_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1792),
    .D(_00953_),
    .Q_N(_14319_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1793),
    .D(_00954_),
    .Q_N(_14318_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1794),
    .D(_00955_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1795),
    .D(_00956_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1796),
    .D(_00957_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1797),
    .D(_00958_),
    .Q_N(_14906_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1798),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_14907_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1799),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_14908_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1800),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_14909_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1801),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_14910_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1802),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_14911_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1803),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00147_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1804),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1805),
    .D(_00959_),
    .Q_N(_00293_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1806),
    .D(_00960_),
    .Q_N(_00292_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1807),
    .D(_00961_),
    .Q_N(_00291_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1808),
    .D(_00962_),
    .Q_N(_00290_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1809),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1810),
    .D(_00963_),
    .Q_N(_00289_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1811),
    .D(_00964_),
    .Q_N(_00288_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1812),
    .D(_00965_),
    .Q_N(_00287_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1813),
    .D(_00966_),
    .Q_N(_00286_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1814),
    .D(_00967_),
    .Q_N(_00285_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1815),
    .D(_00968_),
    .Q_N(_00284_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1816),
    .D(_00969_),
    .Q_N(_00283_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1817),
    .D(_00970_),
    .Q_N(_00282_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1818),
    .D(_00971_),
    .Q_N(_00281_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1819),
    .D(_00972_),
    .Q_N(_00280_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1820),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_14312_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1821),
    .D(_00973_),
    .Q_N(_00279_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1822),
    .D(_00974_),
    .Q_N(_14912_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1823),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_14913_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1824),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_14914_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1825),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_14915_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1826),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_14916_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1827),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_14917_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1828),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_14918_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1829),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_14919_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1830),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14920_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1831),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14921_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1832),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14922_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1833),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14923_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1834),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00181_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1835),
    .D(_00975_),
    .Q_N(_00182_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1836),
    .D(_00976_),
    .Q_N(_00273_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1837),
    .D(_00977_),
    .Q_N(_00272_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1838),
    .D(_00978_),
    .Q_N(_00178_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1839),
    .D(_00979_),
    .Q_N(_00177_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1840),
    .D(_00980_),
    .Q_N(_00176_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1841),
    .D(_00981_),
    .Q_N(_00271_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1842),
    .D(_00982_),
    .Q_N(_00173_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1843),
    .D(_00983_),
    .Q_N(_00172_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1844),
    .D(_00984_),
    .Q_N(_00278_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1845),
    .D(_00985_),
    .Q_N(_00277_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1846),
    .D(_00986_),
    .Q_N(_00276_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1847),
    .D(_00987_),
    .Q_N(_00270_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1848),
    .D(_00988_),
    .Q_N(_00275_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1849),
    .D(_00989_),
    .Q_N(_00274_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1850),
    .D(_00990_),
    .Q_N(_14311_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1851),
    .D(_00991_),
    .Q_N(_00180_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1852),
    .D(_00992_),
    .Q_N(_14310_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1853),
    .D(_00993_),
    .Q_N(_14309_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1854),
    .D(_00994_),
    .Q_N(_14308_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1855),
    .D(_00995_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1856),
    .D(_00996_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1857),
    .D(_00997_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1858),
    .D(_00998_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1859),
    .D(_00999_),
    .Q_N(_14303_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1860),
    .D(_01000_),
    .Q_N(_14302_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1861),
    .D(_01001_),
    .Q_N(_14301_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1862),
    .D(_01002_),
    .Q_N(_14300_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1863),
    .D(_01003_),
    .Q_N(_14299_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1864),
    .D(_01004_),
    .Q_N(_14298_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1865),
    .D(_01005_),
    .Q_N(_14297_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1866),
    .D(_01006_),
    .Q_N(_14296_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1867),
    .D(_01007_),
    .Q_N(_14295_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1868),
    .D(_01008_),
    .Q_N(_14294_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1869),
    .D(_01009_),
    .Q_N(_14293_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1870),
    .D(_01010_),
    .Q_N(_14292_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1871),
    .D(_01011_),
    .Q_N(_14291_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1872),
    .D(_01012_),
    .Q_N(_14290_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1873),
    .D(_01013_),
    .Q_N(_14289_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1874),
    .D(_01014_),
    .Q_N(_14288_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1875),
    .D(_01015_),
    .Q_N(_14287_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1876),
    .D(_01016_),
    .Q_N(_14286_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1877),
    .D(_01017_),
    .Q_N(_14285_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1878),
    .D(_01018_),
    .Q_N(_14284_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1879),
    .D(_01019_),
    .Q_N(_14283_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1880),
    .D(_01020_),
    .Q_N(_14282_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1881),
    .D(_01021_),
    .Q_N(_14281_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1882),
    .D(_01022_),
    .Q_N(_14280_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1883),
    .D(_01023_),
    .Q_N(_00237_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1884),
    .D(_01024_),
    .Q_N(_00219_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1885),
    .D(_01025_),
    .Q_N(_00221_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1886),
    .D(_01026_),
    .Q_N(_14279_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1887),
    .D(_01027_),
    .Q_N(_14278_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1888),
    .D(_01028_),
    .Q_N(_14277_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1889),
    .D(_01029_),
    .Q_N(_14276_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1890),
    .D(_01030_),
    .Q_N(_00256_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1891),
    .D(_01031_),
    .Q_N(_14275_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1892),
    .D(_01032_),
    .Q_N(_00203_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1893),
    .D(_01033_),
    .Q_N(_00208_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1894),
    .D(_01034_),
    .Q_N(_00209_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1895),
    .D(_01035_),
    .Q_N(_00211_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1896),
    .D(_01036_),
    .Q_N(_00213_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1897),
    .D(_01037_),
    .Q_N(_00215_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1898),
    .D(_01038_),
    .Q_N(_00217_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1899),
    .D(_01039_),
    .Q_N(_14274_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1900),
    .D(_01040_),
    .Q_N(_14273_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1901),
    .D(_01041_),
    .Q_N(_14272_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1902),
    .D(_01042_),
    .Q_N(_14271_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1903),
    .D(_01043_),
    .Q_N(_14924_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1904),
    .D(_00054_),
    .Q_N(_00236_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1905),
    .D(_01044_),
    .Q_N(_00204_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1906),
    .D(_01045_),
    .Q_N(_14270_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1907),
    .D(_01046_),
    .Q_N(_14269_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1908),
    .D(_01047_),
    .Q_N(_14268_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1909),
    .D(_01048_),
    .Q_N(_14267_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1910),
    .D(_01049_),
    .Q_N(_14266_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1911),
    .D(_01050_),
    .Q_N(_14265_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1912),
    .D(_01051_),
    .Q_N(_00162_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1913),
    .D(_01052_),
    .Q_N(_00163_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1914),
    .D(_01053_),
    .Q_N(_00268_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1915),
    .D(_01054_),
    .Q_N(_00164_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net1916),
    .D(_01055_),
    .Q_N(_00165_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1917),
    .D(_01056_),
    .Q_N(_00166_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1918),
    .D(_01057_),
    .Q_N(_00262_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1919),
    .D(_01058_),
    .Q_N(_14264_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1920),
    .D(_01059_),
    .Q_N(_14263_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1921),
    .D(_01060_),
    .Q_N(_14262_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1922),
    .D(_01061_),
    .Q_N(_14261_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1923),
    .D(_01062_),
    .Q_N(_00269_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1924),
    .D(_01063_),
    .Q_N(_14260_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1925),
    .D(_01064_),
    .Q_N(_00170_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1926),
    .D(_01065_),
    .Q_N(_14259_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1927),
    .D(_01066_),
    .Q_N(_00235_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1928),
    .D(_01067_),
    .Q_N(_14258_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1929),
    .D(_01068_),
    .Q_N(_14257_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1930),
    .D(_01069_),
    .Q_N(_14256_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1931),
    .D(_01070_),
    .Q_N(_14255_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1932),
    .D(_01071_),
    .Q_N(_14254_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1933),
    .D(_01072_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1934),
    .D(_01073_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1935),
    .D(_01074_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1936),
    .D(_01075_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1937),
    .D(_01076_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1938),
    .D(_01077_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1939),
    .D(_01078_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1940),
    .D(_01079_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1941),
    .D(_01080_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1942),
    .D(_01081_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1943),
    .D(_01082_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1944),
    .D(_01083_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1945),
    .D(_01084_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1946),
    .D(_01085_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1947),
    .D(_01086_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1948),
    .D(_01087_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1949),
    .D(_01088_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1950),
    .D(_01089_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1951),
    .D(_01090_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1952),
    .D(_01091_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1953),
    .D(_01092_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1954),
    .D(_01093_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1955),
    .D(_01094_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1956),
    .D(_01095_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1957),
    .D(_01096_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1958),
    .D(_01097_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1959),
    .D(_01098_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1960),
    .D(_01099_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1961),
    .D(_01100_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1962),
    .D(_01101_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1963),
    .D(_01102_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1964),
    .D(_01103_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1965),
    .D(_01104_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1966),
    .D(_01105_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1967),
    .D(_01106_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1968),
    .D(_01107_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1969),
    .D(_01108_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1970),
    .D(_01109_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1971),
    .D(_01110_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1972),
    .D(_01111_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1973),
    .D(_01112_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1974),
    .D(_01113_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1975),
    .D(_01114_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1976),
    .D(_01115_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1977),
    .D(_01116_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1978),
    .D(_01117_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1979),
    .D(_01118_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1980),
    .D(_01119_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1981),
    .D(_01120_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1982),
    .D(_01121_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1983),
    .D(_01122_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1984),
    .D(_01123_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1985),
    .D(_01124_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1986),
    .D(_01125_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1987),
    .D(_01126_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1988),
    .D(_01127_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1989),
    .D(_01128_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1990),
    .D(_01129_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1991),
    .D(_01130_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1992),
    .D(_01131_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1993),
    .D(_01132_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1994),
    .D(_01133_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1995),
    .D(_01134_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1996),
    .D(_01135_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1997),
    .D(_01136_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1998),
    .D(_01137_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1999),
    .D(_01138_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2000),
    .D(_01139_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2001),
    .D(_01140_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2002),
    .D(_01141_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2003),
    .D(_01142_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2004),
    .D(_01143_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2005),
    .D(_01144_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2006),
    .D(_01145_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2007),
    .D(_01146_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2008),
    .D(_01147_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2009),
    .D(_01148_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2010),
    .D(_01149_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net2011),
    .D(_01150_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2012),
    .D(_01151_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2013),
    .D(_01152_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2014),
    .D(_01153_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2015),
    .D(_01154_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2016),
    .D(_01155_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2017),
    .D(_01156_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2018),
    .D(_01157_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2019),
    .D(_01158_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2020),
    .D(_01159_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2021),
    .D(_01160_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2022),
    .D(_01161_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2023),
    .D(_01162_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2024),
    .D(_01163_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2025),
    .D(_01164_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2026),
    .D(_01165_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2027),
    .D(_01166_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2028),
    .D(_01167_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2029),
    .D(_01168_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2030),
    .D(_01169_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2031),
    .D(_01170_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2032),
    .D(_01171_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2033),
    .D(_01172_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2034),
    .D(_01173_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2035),
    .D(_01174_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2036),
    .D(_01175_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2037),
    .D(_01176_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2038),
    .D(_01177_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2039),
    .D(_01178_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2040),
    .D(_01179_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2041),
    .D(_01180_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2042),
    .D(_01181_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2043),
    .D(_01182_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2044),
    .D(_01183_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2045),
    .D(_01184_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2046),
    .D(_01185_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2047),
    .D(_01186_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2048),
    .D(_01187_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2049),
    .D(_01188_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2050),
    .D(_01189_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2051),
    .D(_01190_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2052),
    .D(_01191_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2053),
    .D(_01192_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2054),
    .D(_01193_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2055),
    .D(_01194_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2056),
    .D(_01195_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2057),
    .D(_01196_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2058),
    .D(_01197_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2059),
    .D(_01198_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2060),
    .D(_01199_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2061),
    .D(_01200_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2062),
    .D(_01201_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2063),
    .D(_01202_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2064),
    .D(_01203_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2065),
    .D(_01204_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2066),
    .D(_01205_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2067),
    .D(_01206_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2068),
    .D(_01207_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2069),
    .D(_01208_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2070),
    .D(_01209_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2071),
    .D(_01210_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2072),
    .D(_01211_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2073),
    .D(_01212_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2074),
    .D(_01213_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2075),
    .D(_01214_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2076),
    .D(_01215_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2077),
    .D(_01216_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2078),
    .D(_01217_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2079),
    .D(_01218_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2080),
    .D(_01219_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2081),
    .D(_01220_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2082),
    .D(_01221_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2083),
    .D(_01222_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2084),
    .D(_01223_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2085),
    .D(_01224_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2086),
    .D(_01225_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2087),
    .D(_01226_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2088),
    .D(_01227_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2089),
    .D(_01228_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net2090),
    .D(_01229_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2091),
    .D(_01230_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2092),
    .D(_01231_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2093),
    .D(_01232_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2094),
    .D(_01233_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2095),
    .D(_01234_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2096),
    .D(_01235_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2097),
    .D(_01236_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2098),
    .D(_01237_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2099),
    .D(_01238_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2100),
    .D(_01239_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2101),
    .D(_01240_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2102),
    .D(_01241_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2103),
    .D(_01242_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2104),
    .D(_01243_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2105),
    .D(_01244_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2106),
    .D(_01245_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2107),
    .D(_01246_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2108),
    .D(_01247_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2109),
    .D(_01248_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2110),
    .D(_01249_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2111),
    .D(_01250_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2112),
    .D(_01251_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2113),
    .D(_01252_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2114),
    .D(_01253_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2115),
    .D(_01254_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2116),
    .D(_01255_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2117),
    .D(_01256_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2118),
    .D(_01257_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2119),
    .D(_01258_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2120),
    .D(_01259_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2121),
    .D(_01260_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2122),
    .D(_01261_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2123),
    .D(_01262_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2124),
    .D(_01263_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2125),
    .D(_01264_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2126),
    .D(_01265_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2127),
    .D(_01266_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2128),
    .D(_01267_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2129),
    .D(_01268_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2130),
    .D(_01269_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2131),
    .D(_01270_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2132),
    .D(_01271_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2133),
    .D(_01272_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2134),
    .D(_01273_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2135),
    .D(_01274_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2136),
    .D(_01275_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2137),
    .D(_01276_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2138),
    .D(_01277_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2139),
    .D(_01278_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2140),
    .D(_01279_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2141),
    .D(_01280_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2142),
    .D(_01281_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2143),
    .D(_01282_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2144),
    .D(_01283_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2145),
    .D(_01284_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2146),
    .D(_01285_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2147),
    .D(_01286_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2148),
    .D(_01287_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2149),
    .D(_01288_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2150),
    .D(_01289_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2151),
    .D(_01290_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2152),
    .D(_01291_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2153),
    .D(_01292_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2154),
    .D(_01293_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2155),
    .D(_01294_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2156),
    .D(_01295_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2157),
    .D(_01296_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2158),
    .D(_01297_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2159),
    .D(_01298_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2160),
    .D(_01299_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2161),
    .D(_01300_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2162),
    .D(_01301_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2163),
    .D(_01302_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2164),
    .D(_01303_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2165),
    .D(_01304_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2166),
    .D(_01305_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2167),
    .D(_01306_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2168),
    .D(_01307_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2169),
    .D(_01308_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2170),
    .D(_01309_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2171),
    .D(_01310_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2172),
    .D(_01311_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2173),
    .D(_01312_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2174),
    .D(_01313_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2175),
    .D(_01314_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2176),
    .D(_01315_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2177),
    .D(_01316_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2178),
    .D(_01317_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2179),
    .D(_01318_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2180),
    .D(_01319_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2181),
    .D(_01320_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2182),
    .D(_01321_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2183),
    .D(_01322_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2184),
    .D(_01323_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2185),
    .D(_01324_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2186),
    .D(_01325_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2187),
    .D(_01326_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2188),
    .D(_01327_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2189),
    .D(_01328_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2190),
    .D(_01329_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2191),
    .D(_01330_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2192),
    .D(_01331_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2193),
    .D(_01332_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2194),
    .D(_01333_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2195),
    .D(_01334_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2196),
    .D(_01335_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2197),
    .D(_01336_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2198),
    .D(_01337_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2199),
    .D(_01338_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2200),
    .D(_01339_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2201),
    .D(_01340_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2202),
    .D(_01341_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2203),
    .D(_01342_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2204),
    .D(_01343_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2205),
    .D(_01344_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2206),
    .D(_01345_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2207),
    .D(_01346_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2208),
    .D(_01347_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2209),
    .D(_01348_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2210),
    .D(_01349_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2211),
    .D(_01350_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2212),
    .D(_01351_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2213),
    .D(_01352_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2214),
    .D(_01353_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2215),
    .D(_01354_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2216),
    .D(_01355_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2217),
    .D(_01356_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2218),
    .D(_01357_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2219),
    .D(_01358_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2220),
    .D(_01359_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2221),
    .D(_01360_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2222),
    .D(_01361_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2223),
    .D(_01362_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2224),
    .D(_01363_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2225),
    .D(_01364_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2226),
    .D(_01365_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2227),
    .D(_01366_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2228),
    .D(_01367_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2229),
    .D(_01368_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2230),
    .D(_01369_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2231),
    .D(_01370_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2232),
    .D(_01371_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2233),
    .D(_01372_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2234),
    .D(_01373_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2235),
    .D(_01374_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2236),
    .D(_01375_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2237),
    .D(_01376_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2238),
    .D(_01377_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2239),
    .D(_01378_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2240),
    .D(_01379_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2241),
    .D(_01380_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2242),
    .D(_01381_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2243),
    .D(_01382_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2244),
    .D(_01383_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2245),
    .D(_01384_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2246),
    .D(_01385_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2247),
    .D(_01386_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2248),
    .D(_01387_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2249),
    .D(_01388_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2250),
    .D(_01389_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2251),
    .D(_01390_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2252),
    .D(_01391_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2253),
    .D(_01392_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2254),
    .D(_01393_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2255),
    .D(_01394_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2256),
    .D(_01395_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2257),
    .D(_01396_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2258),
    .D(_01397_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2259),
    .D(_01398_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2260),
    .D(_01399_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2261),
    .D(_01400_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2262),
    .D(_01401_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net2263),
    .D(_01402_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2264),
    .D(_01403_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2265),
    .D(_01404_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2266),
    .D(_01405_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2267),
    .D(_01406_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2268),
    .D(_01407_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2269),
    .D(_01408_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2270),
    .D(_01409_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2271),
    .D(_01410_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2272),
    .D(_01411_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2273),
    .D(_01412_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2274),
    .D(_01413_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2275),
    .D(_01414_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2276),
    .D(_01415_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2277),
    .D(_01416_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2278),
    .D(_01417_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2279),
    .D(_01418_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2280),
    .D(_01419_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2281),
    .D(_01420_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2282),
    .D(_01421_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2283),
    .D(_01422_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2284),
    .D(_01423_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2285),
    .D(_01424_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2286),
    .D(_01425_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2287),
    .D(_01426_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2288),
    .D(_01427_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2289),
    .D(_01428_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2290),
    .D(_01429_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2291),
    .D(_01430_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2292),
    .D(_01431_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2293),
    .D(_01432_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2294),
    .D(_01433_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2295),
    .D(_01434_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2296),
    .D(_01435_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2297),
    .D(_01436_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2298),
    .D(_01437_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2299),
    .D(_01438_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2300),
    .D(_01439_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2301),
    .D(_01440_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net2302),
    .D(_01441_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2303),
    .D(_01442_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2304),
    .D(_01443_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2305),
    .D(_01444_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2306),
    .D(_01445_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2307),
    .D(_01446_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2308),
    .D(_01447_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2309),
    .D(_01448_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2310),
    .D(_01449_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2311),
    .D(_01450_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2312),
    .D(_01451_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2313),
    .D(_01452_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2314),
    .D(_01453_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2315),
    .D(_01454_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2316),
    .D(_01455_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2317),
    .D(_01456_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2318),
    .D(_01457_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2319),
    .D(_01458_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2320),
    .D(_01459_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2321),
    .D(_01460_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2322),
    .D(_01461_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2323),
    .D(_01462_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net2324),
    .D(_01463_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net2325),
    .D(_01464_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2326),
    .D(_01465_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2327),
    .D(_01466_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2328),
    .D(_01467_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2329),
    .D(_01468_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2330),
    .D(_01469_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2331),
    .D(_01470_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2332),
    .D(_01471_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2333),
    .D(_01472_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2334),
    .D(_01473_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2335),
    .D(_01474_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net2336),
    .D(_01475_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2337),
    .D(_01476_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2338),
    .D(_01477_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2339),
    .D(_01478_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2340),
    .D(_01479_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2341),
    .D(_01480_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net2342),
    .D(_01481_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2343),
    .D(_01482_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2344),
    .D(_01483_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2345),
    .D(_01484_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2346),
    .D(_01485_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2347),
    .D(_01486_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net2348),
    .D(_01487_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net2349),
    .D(_01488_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2350),
    .D(_01489_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2351),
    .D(_01490_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2352),
    .D(_01491_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2353),
    .D(_01492_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2354),
    .D(_01493_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2355),
    .D(_01494_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2356),
    .D(_01495_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net2357),
    .D(_01496_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2358),
    .D(_01497_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2359),
    .D(_01498_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net2360),
    .D(_01499_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2361),
    .D(_01500_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2362),
    .D(_01501_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2363),
    .D(_01502_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2364),
    .D(_01503_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2365),
    .D(_01504_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net2366),
    .D(_01505_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2367),
    .D(_01506_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2368),
    .D(_01507_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2369),
    .D(_01508_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net2370),
    .D(_01509_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net2371),
    .D(_01510_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net2372),
    .D(_01511_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net2373),
    .D(_01512_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2374),
    .D(_01513_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2375),
    .D(_01514_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2376),
    .D(_01515_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2377),
    .D(_01516_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2378),
    .D(_01517_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2379),
    .D(_01518_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2380),
    .D(_01519_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2381),
    .D(_01520_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2382),
    .D(_01521_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2383),
    .D(_01522_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2384),
    .D(_01523_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2385),
    .D(_01524_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2386),
    .D(_01525_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2387),
    .D(_01526_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2388),
    .D(_01527_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2389),
    .D(_01528_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net2390),
    .D(_01529_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2391),
    .D(_01530_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2392),
    .D(_01531_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2393),
    .D(_01532_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2394),
    .D(_01533_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2395),
    .D(_01534_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2396),
    .D(_01535_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2397),
    .D(_01536_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2398),
    .D(_01537_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2399),
    .D(_01538_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2400),
    .D(_01539_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2401),
    .D(_01540_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2402),
    .D(_01541_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2403),
    .D(_01542_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2404),
    .D(_01543_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2405),
    .D(_01544_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2406),
    .D(_01545_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2407),
    .D(_01546_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2408),
    .D(_01547_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2409),
    .D(_01548_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2410),
    .D(_01549_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2411),
    .D(_01550_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2412),
    .D(_01551_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net2413),
    .D(_01552_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2414),
    .D(_01553_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2415),
    .D(_01554_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2416),
    .D(_01555_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2417),
    .D(_01556_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2418),
    .D(_01557_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2419),
    .D(_01558_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2420),
    .D(_01559_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2421),
    .D(_01560_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2422),
    .D(_01561_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2423),
    .D(_01562_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2424),
    .D(_01563_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2425),
    .D(_01564_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2426),
    .D(_01565_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2427),
    .D(_01566_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2428),
    .D(_01567_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2429),
    .D(_01568_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2430),
    .D(_01569_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2431),
    .D(_01570_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2432),
    .D(_01571_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2433),
    .D(_01572_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2434),
    .D(_01573_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2435),
    .D(_01574_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2436),
    .D(_01575_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2437),
    .D(_01576_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2438),
    .D(_01577_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2439),
    .D(_01578_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2440),
    .D(_01579_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2441),
    .D(_01580_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2442),
    .D(_01581_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2443),
    .D(_01582_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2444),
    .D(_01583_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2445),
    .D(_01584_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2446),
    .D(_01585_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2447),
    .D(_01586_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2448),
    .D(_01587_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2449),
    .D(_01588_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2450),
    .D(_01589_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2451),
    .D(_01590_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net2452),
    .D(_01591_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2453),
    .D(_01592_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2454),
    .D(_01593_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2455),
    .D(_01594_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2456),
    .D(_01595_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2457),
    .D(_01596_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2458),
    .D(_01597_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2459),
    .D(_01598_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2460),
    .D(_01599_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2461),
    .D(_01600_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2462),
    .D(_01601_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2463),
    .D(_01602_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2464),
    .D(_01603_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2465),
    .D(_01604_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2466),
    .D(_01605_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2467),
    .D(_01606_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2468),
    .D(_01607_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2469),
    .D(_01608_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2470),
    .D(_01609_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2471),
    .D(_01610_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2472),
    .D(_01611_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2473),
    .D(_01612_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2474),
    .D(_01613_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2475),
    .D(_01614_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2476),
    .D(_01615_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2477),
    .D(_01616_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2478),
    .D(_01617_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2479),
    .D(_01618_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2480),
    .D(_01619_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2481),
    .D(_01620_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2482),
    .D(_01621_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2483),
    .D(_01622_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2484),
    .D(_01623_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2485),
    .D(_01624_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2486),
    .D(_01625_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2487),
    .D(_01626_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2488),
    .D(_01627_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2489),
    .D(_01628_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2490),
    .D(_01629_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2491),
    .D(_01630_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2492),
    .D(_01631_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2493),
    .D(_01632_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2494),
    .D(_01633_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2495),
    .D(_01634_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2496),
    .D(_01635_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2497),
    .D(_01636_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2498),
    .D(_01637_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2499),
    .D(_01638_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2500),
    .D(_01639_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2501),
    .D(_01640_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2502),
    .D(_01641_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2503),
    .D(_01642_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2504),
    .D(_01643_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2505),
    .D(_01644_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2506),
    .D(_01645_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2507),
    .D(_01646_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2508),
    .D(_01647_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2509),
    .D(_01648_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2510),
    .D(_01649_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2511),
    .D(_01650_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2512),
    .D(_01651_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2513),
    .D(_01652_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2514),
    .D(_01653_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2515),
    .D(_01654_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2516),
    .D(_01655_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2517),
    .D(_01656_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2518),
    .D(_01657_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2519),
    .D(_01658_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2520),
    .D(_01659_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2521),
    .D(_01660_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2522),
    .D(_01661_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2523),
    .D(_01662_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2524),
    .D(_01663_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2525),
    .D(_01664_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2526),
    .D(_01665_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2527),
    .D(_01666_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2528),
    .D(_01667_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2529),
    .D(_01668_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2530),
    .D(_01669_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2531),
    .D(_01670_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2532),
    .D(_01671_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2533),
    .D(_01672_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2534),
    .D(_01673_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2535),
    .D(_01674_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2536),
    .D(_01675_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2537),
    .D(_01676_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2538),
    .D(_01677_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2539),
    .D(_01678_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2540),
    .D(_01679_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2541),
    .D(_01680_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2542),
    .D(_01681_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2543),
    .D(_01682_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2544),
    .D(_01683_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2545),
    .D(_01684_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2546),
    .D(_01685_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2547),
    .D(_01686_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2548),
    .D(_01687_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2549),
    .D(_01688_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2550),
    .D(_01689_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2551),
    .D(_01690_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2552),
    .D(_01691_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2553),
    .D(_01692_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2554),
    .D(_01693_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2555),
    .D(_01694_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2556),
    .D(_01695_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2557),
    .D(_01696_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2558),
    .D(_01697_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2559),
    .D(_01698_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2560),
    .D(_01699_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2561),
    .D(_01700_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2562),
    .D(_01701_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2563),
    .D(_01702_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2564),
    .D(_01703_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2565),
    .D(_01704_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2566),
    .D(_01705_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2567),
    .D(_01706_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2568),
    .D(_01707_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2569),
    .D(_01708_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2570),
    .D(_01709_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2571),
    .D(_01710_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2572),
    .D(_01711_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2573),
    .D(_01712_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2574),
    .D(_01713_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2575),
    .D(_01714_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2576),
    .D(_01715_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2577),
    .D(_01716_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2578),
    .D(_01717_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2579),
    .D(_01718_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2580),
    .D(_01719_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2581),
    .D(_01720_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2582),
    .D(_01721_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2583),
    .D(_01722_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2584),
    .D(_01723_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2585),
    .D(_01724_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2586),
    .D(_01725_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2587),
    .D(_01726_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2588),
    .D(_01727_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2589),
    .D(_01728_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2590),
    .D(_01729_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2591),
    .D(_01730_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2592),
    .D(_01731_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2593),
    .D(_01732_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2594),
    .D(_01733_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2595),
    .D(_01734_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2596),
    .D(_01735_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2597),
    .D(_01736_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2598),
    .D(_01737_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2599),
    .D(_01738_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2600),
    .D(_01739_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2601),
    .D(_01740_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2602),
    .D(_01741_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2603),
    .D(_01742_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2604),
    .D(_01743_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2605),
    .D(_01744_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2606),
    .D(_01745_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2607),
    .D(_01746_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2608),
    .D(_01747_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2609),
    .D(_01748_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2610),
    .D(_01749_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2611),
    .D(_01750_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2612),
    .D(_01751_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2613),
    .D(_01752_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2614),
    .D(_01753_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2615),
    .D(_01754_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2616),
    .D(_01755_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2617),
    .D(_01756_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2618),
    .D(_01757_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2619),
    .D(_01758_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2620),
    .D(_01759_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2621),
    .D(_01760_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2622),
    .D(_01761_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2623),
    .D(_01762_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2624),
    .D(_01763_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2625),
    .D(_01764_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2626),
    .D(_01765_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2627),
    .D(_01766_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2628),
    .D(_01767_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2629),
    .D(_01768_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2630),
    .D(_01769_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2631),
    .D(_01770_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2632),
    .D(_01771_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2633),
    .D(_01772_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2634),
    .D(_01773_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2635),
    .D(_01774_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2636),
    .D(_01775_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2637),
    .D(_01776_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2638),
    .D(_01777_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2639),
    .D(_01778_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2640),
    .D(_01779_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2641),
    .D(_01780_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2642),
    .D(_01781_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2643),
    .D(_01782_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2644),
    .D(_01783_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2645),
    .D(_01784_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2646),
    .D(_01785_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2647),
    .D(_01786_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2648),
    .D(_01787_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2649),
    .D(_01788_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2650),
    .D(_01789_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2651),
    .D(_01790_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2652),
    .D(_01791_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2653),
    .D(_01792_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2654),
    .D(_01793_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2655),
    .D(_01794_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2656),
    .D(_01795_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2657),
    .D(_01796_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2658),
    .D(_01797_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2659),
    .D(_01798_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2660),
    .D(_01799_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2661),
    .D(_01800_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2662),
    .D(_01801_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2663),
    .D(_01802_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2664),
    .D(_01803_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2665),
    .D(_01804_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2666),
    .D(_01805_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2667),
    .D(_01806_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2668),
    .D(_01807_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2669),
    .D(_01808_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2670),
    .D(_01809_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2671),
    .D(_01810_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2672),
    .D(_01811_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2673),
    .D(_01812_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2674),
    .D(_01813_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2675),
    .D(_01814_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2676),
    .D(_01815_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2677),
    .D(_01816_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2678),
    .D(_01817_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2679),
    .D(_01818_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2680),
    .D(_01819_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2681),
    .D(_01820_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2682),
    .D(_01821_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2683),
    .D(_01822_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2684),
    .D(_01823_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2685),
    .D(_01824_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2686),
    .D(_01825_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2687),
    .D(_01826_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2688),
    .D(_01827_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2689),
    .D(_01828_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2690),
    .D(_01829_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2691),
    .D(_01830_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2692),
    .D(_01831_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2693),
    .D(_01832_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2694),
    .D(_01833_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2695),
    .D(_01834_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2696),
    .D(_01835_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2697),
    .D(_01836_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2698),
    .D(_01837_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2699),
    .D(_01838_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2700),
    .D(_01839_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2701),
    .D(_01840_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2702),
    .D(_01841_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2703),
    .D(_01842_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2704),
    .D(_01843_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2705),
    .D(_01844_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2706),
    .D(_01845_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2707),
    .D(_01846_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2708),
    .D(_01847_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2709),
    .D(_01848_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2710),
    .D(_01849_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2711),
    .D(_01850_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2712),
    .D(_01851_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2713),
    .D(_01852_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2714),
    .D(_01853_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2715),
    .D(_01854_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2716),
    .D(_01855_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2717),
    .D(_01856_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2718),
    .D(_01857_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2719),
    .D(_01858_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2720),
    .D(_01859_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net2721),
    .D(_01860_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2722),
    .D(_01861_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2723),
    .D(_01862_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2724),
    .D(_01863_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2725),
    .D(_01864_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2726),
    .D(_01865_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2727),
    .D(_01866_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2728),
    .D(_01867_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2729),
    .D(_01868_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2730),
    .D(_01869_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2731),
    .D(_01870_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2732),
    .D(_01871_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2733),
    .D(_01872_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2734),
    .D(_01873_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2735),
    .D(_01874_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net2736),
    .D(_01875_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2737),
    .D(_01876_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2738),
    .D(_01877_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2739),
    .D(_01878_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2740),
    .D(_01879_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2741),
    .D(_01880_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2742),
    .D(_01881_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2743),
    .D(_01882_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2744),
    .D(_01883_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2745),
    .D(_01884_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2746),
    .D(_01885_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2747),
    .D(_01886_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2748),
    .D(_01887_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2749),
    .D(_01888_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net2750),
    .D(_01889_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2751),
    .D(_01890_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net2752),
    .D(_01891_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net2753),
    .D(_01892_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2754),
    .D(_01893_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2755),
    .D(_01894_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2756),
    .D(_01895_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2757),
    .D(_01896_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net2758),
    .D(_01897_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net2759),
    .D(_01898_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2760),
    .D(_01899_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net2761),
    .D(_01900_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net2762),
    .D(_01901_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2763),
    .D(_01902_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2764),
    .D(_01903_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2765),
    .D(_01904_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2766),
    .D(_01905_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2767),
    .D(_01906_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2768),
    .D(_01907_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2769),
    .D(_01908_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net2770),
    .D(_01909_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2771),
    .D(_01910_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2772),
    .D(_01911_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2773),
    .D(_01912_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2774),
    .D(_01913_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2775),
    .D(_01914_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2776),
    .D(_01915_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2777),
    .D(_01916_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2778),
    .D(_01917_),
    .Q_N(_13408_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2779),
    .D(_01918_),
    .Q_N(_13407_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2780),
    .D(_01919_),
    .Q_N(_13406_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2781),
    .D(_01920_),
    .Q_N(_13405_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2782),
    .D(_01921_),
    .Q_N(_13404_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2783),
    .D(_01922_),
    .Q_N(_13403_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2784),
    .D(_01923_),
    .Q_N(_13402_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2785),
    .D(_01924_),
    .Q_N(_13401_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2786),
    .D(_01925_),
    .Q_N(_13400_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2787),
    .D(_01926_),
    .Q_N(_13399_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2788),
    .D(_01927_),
    .Q_N(_13398_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2789),
    .D(_01928_),
    .Q_N(_13397_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2790),
    .D(_01929_),
    .Q_N(_13396_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net2791),
    .D(_01930_),
    .Q_N(_13395_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2792),
    .D(_01931_),
    .Q_N(_13394_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2793),
    .D(_01932_),
    .Q_N(_13393_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2794),
    .D(_01933_),
    .Q_N(_13392_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2795),
    .D(_01934_),
    .Q_N(_13391_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2796),
    .D(_01935_),
    .Q_N(_13390_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2797),
    .D(_01936_),
    .Q_N(_13389_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2798),
    .D(_01937_),
    .Q_N(_13388_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2799),
    .D(_01938_),
    .Q_N(_13387_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2800),
    .D(_01939_),
    .Q_N(_13386_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2801),
    .D(_01940_),
    .Q_N(_13385_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2802),
    .D(_01941_),
    .Q_N(_13384_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2803),
    .D(_01942_),
    .Q_N(_13383_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2804),
    .D(_01943_),
    .Q_N(_13382_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2805),
    .D(_01944_),
    .Q_N(_13381_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2806),
    .D(_01945_),
    .Q_N(_13380_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2807),
    .D(_01946_),
    .Q_N(_13379_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2808),
    .D(_01947_),
    .Q_N(_13378_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2809),
    .D(_01948_),
    .Q_N(_13377_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2810),
    .D(_01949_),
    .Q_N(_13376_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2811),
    .D(_01950_),
    .Q_N(_13375_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2812),
    .D(_01951_),
    .Q_N(_13374_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2813),
    .D(_01952_),
    .Q_N(_13373_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2814),
    .D(_01953_),
    .Q_N(_13372_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2815),
    .D(_01954_),
    .Q_N(_13371_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2816),
    .D(_01955_),
    .Q_N(_13370_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2817),
    .D(_01956_),
    .Q_N(_13369_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2818),
    .D(_01957_),
    .Q_N(_13368_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2819),
    .D(_01958_),
    .Q_N(_13367_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2820),
    .D(_01959_),
    .Q_N(_00308_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2821),
    .D(_01960_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2822),
    .D(_01961_),
    .Q_N(_00107_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2823),
    .D(_01962_),
    .Q_N(_13366_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2824),
    .D(_01963_),
    .Q_N(_00124_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2825),
    .D(_01964_),
    .Q_N(_00135_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2826),
    .D(_01965_),
    .Q_N(_00146_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2827),
    .D(_01966_),
    .Q_N(_13365_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2828),
    .D(_01967_),
    .Q_N(_13364_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2829),
    .D(_01968_),
    .Q_N(_00161_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2830),
    .D(_01969_),
    .Q_N(_13363_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2831),
    .D(_01970_),
    .Q_N(_13362_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2832),
    .D(_01971_),
    .Q_N(_13361_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2833),
    .D(_01972_),
    .Q_N(_00160_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2834),
    .D(_01973_),
    .Q_N(_13360_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2835),
    .D(_01974_),
    .Q_N(_13359_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2836),
    .D(_01975_),
    .Q_N(_00304_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2837),
    .D(_01976_),
    .Q_N(_00094_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2838),
    .D(_01977_),
    .Q_N(_00104_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2839),
    .D(_01978_),
    .Q_N(_13358_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2840),
    .D(_01979_),
    .Q_N(_00120_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2841),
    .D(_01980_),
    .Q_N(_00131_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2842),
    .D(_01981_),
    .Q_N(_00142_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2843),
    .D(_01982_),
    .Q_N(_13357_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2844),
    .D(_01983_),
    .Q_N(_00123_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2845),
    .D(_01984_),
    .Q_N(_00134_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2846),
    .D(_01985_),
    .Q_N(_00145_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2847),
    .D(_01986_),
    .Q_N(_13356_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2848),
    .D(_01987_),
    .Q_N(_00306_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2849),
    .D(_01988_),
    .Q_N(_00096_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2850),
    .D(_01989_),
    .Q_N(_00106_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2851),
    .D(_01990_),
    .Q_N(_13355_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2852),
    .D(_01991_),
    .Q_N(_00122_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2853),
    .D(_01992_),
    .Q_N(_00133_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2854),
    .D(_01993_),
    .Q_N(_00144_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2855),
    .D(_01994_),
    .Q_N(_13354_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2856),
    .D(_01995_),
    .Q_N(_00305_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2857),
    .D(_01996_),
    .Q_N(_00095_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2858),
    .D(_01997_),
    .Q_N(_00105_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2859),
    .D(_01998_),
    .Q_N(_13353_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2860),
    .D(_01999_),
    .Q_N(_00121_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2861),
    .D(_02000_),
    .Q_N(_00132_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2862),
    .D(_02001_),
    .Q_N(_00143_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2863),
    .D(_02002_),
    .Q_N(_13352_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2864),
    .D(_02003_),
    .Q_N(_00307_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2865),
    .D(_02004_),
    .Q_N(_00097_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2866),
    .D(_02005_),
    .Q_N(_13351_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net2867),
    .D(_02006_),
    .Q_N(_00189_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2868),
    .D(_02007_),
    .Q_N(_00191_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2869),
    .D(_02008_),
    .Q_N(_00187_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2870),
    .D(_02009_),
    .Q_N(_00193_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2871),
    .D(_02010_),
    .Q_N(_00195_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2872),
    .D(_02011_),
    .Q_N(_00197_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2873),
    .D(_02012_),
    .Q_N(_13350_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2874),
    .D(_02013_),
    .Q_N(_00200_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2875),
    .D(_02014_),
    .Q_N(_00151_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2876),
    .D(_02015_),
    .Q_N(_00153_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2877),
    .D(_02016_),
    .Q_N(_00199_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2878),
    .D(_02017_),
    .Q_N(_00155_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2879),
    .D(_02018_),
    .Q_N(_00184_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2880),
    .D(_02019_),
    .Q_N(_00186_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2881),
    .D(_02020_),
    .Q_N(_00149_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2882),
    .D(_02021_),
    .Q_N(_00157_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2883),
    .D(_02022_),
    .Q_N(_00159_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2884),
    .D(_02023_),
    .Q_N(_00190_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2885),
    .D(_02024_),
    .Q_N(_00192_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2886),
    .D(_02025_),
    .Q_N(_00188_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2887),
    .D(_02026_),
    .Q_N(_00194_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2888),
    .D(_02027_),
    .Q_N(_00150_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2889),
    .D(_02028_),
    .Q_N(_00196_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2890),
    .D(_02029_),
    .Q_N(_00198_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2891),
    .D(_02030_),
    .Q_N(_00152_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2892),
    .D(_02031_),
    .Q_N(_00154_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2893),
    .D(_02032_),
    .Q_N(_00183_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2894),
    .D(_02033_),
    .Q_N(_00185_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2895),
    .D(_02034_),
    .Q_N(_00148_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net2896),
    .D(_02035_),
    .Q_N(_00156_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2897),
    .D(_02036_),
    .Q_N(_00158_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2898),
    .D(_02037_),
    .Q_N(_13349_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2899),
    .D(_02038_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2900),
    .D(_02039_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2901),
    .D(_02040_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2902),
    .D(_02041_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2903),
    .D(_02042_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2904),
    .D(_02043_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2905),
    .D(_02044_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2906),
    .D(_02045_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2907),
    .D(_02046_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2908),
    .D(_02047_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2909),
    .D(_02048_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2910),
    .D(_02049_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2911),
    .D(_02050_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2912),
    .D(_02051_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2913),
    .D(_02052_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2914),
    .D(_02053_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2915),
    .D(_02054_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2916),
    .D(_02055_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2917),
    .D(_02056_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2918),
    .D(_02057_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2919),
    .D(_02058_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2920),
    .D(_02059_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2921),
    .D(_02060_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2922),
    .D(_02061_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2923),
    .D(_02062_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2924),
    .D(_02063_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2925),
    .D(_02064_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2926),
    .D(_02065_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2927),
    .D(_02066_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2928),
    .D(_02067_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2929),
    .D(_02068_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2930),
    .D(_02069_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2931),
    .D(_02070_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2932),
    .D(_02071_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2933),
    .D(_02072_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2934),
    .D(_02073_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2935),
    .D(_02074_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2936),
    .D(_02075_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2937),
    .D(_02076_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2938),
    .D(_02077_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2939),
    .D(_02078_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2940),
    .D(_02079_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2941),
    .D(_02080_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2942),
    .D(_02081_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2943),
    .D(_02082_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2944),
    .D(_02083_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2945),
    .D(_02084_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2946),
    .D(_02085_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2947),
    .D(_02086_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2948),
    .D(_02087_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2949),
    .D(_02088_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2950),
    .D(_02089_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2951),
    .D(_02090_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2952),
    .D(_02091_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2953),
    .D(_02092_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2954),
    .D(_02093_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2955),
    .D(_02094_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2956),
    .D(_02095_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2957),
    .D(_02096_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2958),
    .D(_02097_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2959),
    .D(_02098_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2960),
    .D(_02099_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2961),
    .D(_02100_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2962),
    .D(_02101_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2963),
    .D(_02102_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net2964),
    .D(_02103_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2965),
    .D(_02104_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2966),
    .D(_02105_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2967),
    .D(_02106_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2968),
    .D(_02107_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2969),
    .D(_02108_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2970),
    .D(_02109_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2971),
    .D(_02110_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2972),
    .D(_02111_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2973),
    .D(_02112_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2974),
    .D(_02113_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2975),
    .D(_02114_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2976),
    .D(_02115_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2977),
    .D(_02116_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2978),
    .D(_02117_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2979),
    .D(_02118_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2980),
    .D(_02119_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2981),
    .D(_02120_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2982),
    .D(_02121_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2983),
    .D(_02122_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2984),
    .D(_02123_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2985),
    .D(_02124_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2986),
    .D(_02125_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2987),
    .D(_02126_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2988),
    .D(_02127_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2989),
    .D(_02128_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2990),
    .D(_02129_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2991),
    .D(_02130_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2992),
    .D(_02131_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net2993),
    .D(_02132_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2994),
    .D(_02133_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net2995),
    .D(_02134_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net2996),
    .D(_02135_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2997),
    .D(_02136_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2998),
    .D(_02137_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2999),
    .D(_02138_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3000),
    .D(_02139_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net3001),
    .D(_02140_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3002),
    .D(_02141_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3003),
    .D(_02142_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net3004),
    .D(_02143_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3005),
    .D(_02144_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3006),
    .D(_02145_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3007),
    .D(_02146_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3008),
    .D(_02147_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3009),
    .D(_02148_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3010),
    .D(_02149_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3011),
    .D(_02150_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3012),
    .D(_02151_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3013),
    .D(_02152_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3014),
    .D(_02153_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3015),
    .D(_02154_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3016),
    .D(_02155_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3017),
    .D(_02156_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3018),
    .D(_02157_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3019),
    .D(_02158_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3020),
    .D(_02159_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3021),
    .D(_02160_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3022),
    .D(_02161_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3023),
    .D(_02162_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3024),
    .D(_02163_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3025),
    .D(_02164_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3026),
    .D(_02165_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3027),
    .D(_02166_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3028),
    .D(_02167_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3029),
    .D(_02168_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3030),
    .D(_02169_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3031),
    .D(_02170_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3032),
    .D(_02171_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net3033),
    .D(_02172_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3034),
    .D(_02173_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3035),
    .D(_02174_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3036),
    .D(_02175_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3037),
    .D(_02176_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3038),
    .D(_02177_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3039),
    .D(_02178_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3040),
    .D(_02179_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3041),
    .D(_02180_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3042),
    .D(_02181_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3043),
    .D(_02182_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3044),
    .D(_02183_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3045),
    .D(_02184_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3046),
    .D(_02185_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3047),
    .D(_02186_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net3048),
    .D(_02187_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3049),
    .D(_02188_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3050),
    .D(_02189_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3051),
    .D(_02190_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3052),
    .D(_02191_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3053),
    .D(_02192_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3054),
    .D(_02193_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3055),
    .D(_02194_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3056),
    .D(_02195_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3057),
    .D(_02196_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3058),
    .D(_02197_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3059),
    .D(_02198_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3060),
    .D(_02199_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3061),
    .D(_02200_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3062),
    .D(_02201_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3063),
    .D(_02202_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3064),
    .D(_02203_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3065),
    .D(_02204_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net3066),
    .D(_02205_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3067),
    .D(_02206_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3068),
    .D(_02207_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3069),
    .D(_02208_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3070),
    .D(_02209_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3071),
    .D(_02210_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3072),
    .D(_02211_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3073),
    .D(_02212_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3074),
    .D(_02213_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3075),
    .D(_02214_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3076),
    .D(_02215_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3077),
    .D(_02216_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3078),
    .D(_02217_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3079),
    .D(_02218_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3080),
    .D(_02219_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3081),
    .D(_02220_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net3082),
    .D(_02221_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3083),
    .D(_02222_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3084),
    .D(_02223_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3085),
    .D(_02224_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net3086),
    .D(_02225_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3087),
    .D(_02226_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3088),
    .D(_02227_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3089),
    .D(_02228_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3090),
    .D(_02229_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3091),
    .D(_02230_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3092),
    .D(_02231_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3093),
    .D(_02232_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3094),
    .D(_02233_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net3095),
    .D(_02234_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3096),
    .D(_02235_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net3097),
    .D(_02236_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net3098),
    .D(_02237_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3099),
    .D(_02238_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net3100),
    .D(_02239_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3101),
    .D(_02240_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net3102),
    .D(_02241_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3103),
    .D(_02242_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3104),
    .D(_02243_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net3105),
    .D(_02244_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3106),
    .D(_02245_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3107),
    .D(_02246_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net3108),
    .D(_02247_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3109),
    .D(_02248_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3110),
    .D(_02249_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3111),
    .D(_02250_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net3112),
    .D(_02251_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net3113),
    .D(_02252_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net3114),
    .D(_02253_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net3115),
    .D(_02254_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net3116),
    .D(_02255_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net3117),
    .D(_02256_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3118),
    .D(_02257_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net3119),
    .D(_02258_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3120),
    .D(_02259_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3121),
    .D(_02260_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3122),
    .D(_02261_),
    .Q_N(_00312_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3123),
    .D(_02262_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net3124),
    .D(_02263_),
    .Q_N(_00234_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3125),
    .D(_02264_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net3126),
    .D(_02265_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3127),
    .D(_02266_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3128),
    .D(_02267_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3129),
    .D(_02268_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3130),
    .D(_02269_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3131),
    .D(_02270_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3132),
    .D(_02271_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3133),
    .D(_02272_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3134),
    .D(_02273_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3135),
    .D(_02274_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3136),
    .D(_02275_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3137),
    .D(_02276_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3138),
    .D(_02277_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3139),
    .D(_02278_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3140),
    .D(_02279_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3141),
    .D(_02280_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3142),
    .D(_02281_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3143),
    .D(_02282_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3144),
    .D(_02283_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3145),
    .D(_02284_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3146),
    .D(_02285_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3147),
    .D(_02286_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3148),
    .D(_02287_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3149),
    .D(_02288_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3150),
    .D(_02289_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3151),
    .D(_02290_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3152),
    .D(_02291_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3153),
    .D(_02292_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3154),
    .D(_02293_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3155),
    .D(_02294_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3156),
    .D(_02295_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3157),
    .D(_02296_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3158),
    .D(_02297_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3159),
    .D(_02298_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3160),
    .D(_02299_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3161),
    .D(_02300_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3162),
    .D(_02301_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3163),
    .D(_02302_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3164),
    .D(_02303_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3165),
    .D(_02304_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3166),
    .D(_02305_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3167),
    .D(_02306_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3168),
    .D(_02307_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3169),
    .D(_02308_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3170),
    .D(_02309_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3171),
    .D(_02310_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3172),
    .D(_02311_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3173),
    .D(_02312_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3174),
    .D(_02313_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3175),
    .D(_02314_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3176),
    .D(_02315_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3177),
    .D(_02316_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3178),
    .D(_02317_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3179),
    .D(_02318_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3180),
    .D(_02319_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3181),
    .D(_02320_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3182),
    .D(_02321_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3183),
    .D(_02322_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3184),
    .D(_02323_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3185),
    .D(_02324_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3186),
    .D(_02325_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3187),
    .D(_02326_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3188),
    .D(_02327_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3189),
    .D(_02328_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3190),
    .D(_02329_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3191),
    .D(_02330_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3192),
    .D(_02331_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3193),
    .D(_02332_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3194),
    .D(_02333_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3195),
    .D(_02334_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3196),
    .D(_02335_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3197),
    .D(_02336_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3198),
    .D(_02337_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3199),
    .D(_02338_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3200),
    .D(_02339_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3201),
    .D(_02340_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3202),
    .D(_02341_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3203),
    .D(_02342_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3204),
    .D(_02343_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3205),
    .D(_02344_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3206),
    .D(_02345_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3207),
    .D(_02346_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3208),
    .D(_02347_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3209),
    .D(_02348_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3210),
    .D(_02349_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3211),
    .D(_02350_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3212),
    .D(_02351_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3213),
    .D(_02352_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3214),
    .D(_02353_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3215),
    .D(_02354_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3216),
    .D(_02355_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3217),
    .D(_02356_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3218),
    .D(_02357_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3219),
    .D(_02358_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3220),
    .D(_02359_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3221),
    .D(_02360_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3222),
    .D(_02361_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3223),
    .D(_02362_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3224),
    .D(_02363_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3225),
    .D(_02364_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3226),
    .D(_02365_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3227),
    .D(_02366_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3228),
    .D(_02367_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3229),
    .D(_02368_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3230),
    .D(_02369_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3231),
    .D(_02370_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3232),
    .D(_02371_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3233),
    .D(_02372_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3234),
    .D(_02373_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3235),
    .D(_02374_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3236),
    .D(_02375_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3237),
    .D(_02376_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3238),
    .D(_02377_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3239),
    .D(_02378_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3240),
    .D(_02379_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3241),
    .D(_02380_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3242),
    .D(_02381_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3243),
    .D(_02382_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3244),
    .D(_02383_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3245),
    .D(_02384_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3246),
    .D(_02385_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3247),
    .D(_02386_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3248),
    .D(_02387_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3249),
    .D(_02388_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3250),
    .D(_02389_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3251),
    .D(_02390_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3252),
    .D(_02391_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3253),
    .D(_02392_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3254),
    .D(_02393_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3255),
    .D(_02394_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3256),
    .D(_02395_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3257),
    .D(_02396_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3258),
    .D(_02397_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3259),
    .D(_02398_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3260),
    .D(_02399_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3261),
    .D(_02400_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3262),
    .D(_02401_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3263),
    .D(_02402_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3264),
    .D(_02403_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3265),
    .D(_02404_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3266),
    .D(_02405_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3267),
    .D(_02406_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3268),
    .D(_02407_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3269),
    .D(_02408_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3270),
    .D(_02409_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3271),
    .D(_02410_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3272),
    .D(_02411_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3273),
    .D(_02412_),
    .Q_N(_12976_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3274),
    .D(_02413_),
    .Q_N(_12975_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3275),
    .D(_02414_),
    .Q_N(_12974_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3276),
    .D(_02415_),
    .Q_N(_12973_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3277),
    .D(_02416_),
    .Q_N(_12972_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3278),
    .D(_02417_),
    .Q_N(_12971_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3279),
    .D(_02418_),
    .Q_N(_12970_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net3280),
    .D(_02419_),
    .Q_N(_12969_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3281),
    .D(_02420_),
    .Q_N(_12968_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3282),
    .D(_02421_),
    .Q_N(_12967_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3283),
    .D(_02422_),
    .Q_N(_12966_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3284),
    .D(_02423_),
    .Q_N(_12965_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3285),
    .D(_02424_),
    .Q_N(_12964_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3286),
    .D(_02425_),
    .Q_N(_12963_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3287),
    .D(_02426_),
    .Q_N(_12962_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3288),
    .D(_02427_),
    .Q_N(_12961_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3289),
    .D(_02428_),
    .Q_N(_12960_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3290),
    .D(_02429_),
    .Q_N(_12959_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3291),
    .D(_02430_),
    .Q_N(_12958_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3292),
    .D(_02431_),
    .Q_N(_12957_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3293),
    .D(_02432_),
    .Q_N(_12956_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3294),
    .D(_02433_),
    .Q_N(_12955_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3295),
    .D(_02434_),
    .Q_N(_12954_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3296),
    .D(_02435_),
    .Q_N(_12953_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3297),
    .D(_02436_),
    .Q_N(_12952_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3298),
    .D(_02437_),
    .Q_N(_12951_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3299),
    .D(_02438_),
    .Q_N(_12950_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3300),
    .D(_02439_),
    .Q_N(_12949_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3301),
    .D(_02440_),
    .Q_N(_12948_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3302),
    .D(_02441_),
    .Q_N(_12947_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3303),
    .D(_02442_),
    .Q_N(_12946_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3304),
    .D(_02443_),
    .Q_N(_12945_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3305),
    .D(_02444_),
    .Q_N(_12944_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3306),
    .D(_02445_),
    .Q_N(_12943_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3307),
    .D(_02446_),
    .Q_N(_12942_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3308),
    .D(_02447_),
    .Q_N(_12941_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3309),
    .D(_02448_),
    .Q_N(_12940_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3310),
    .D(_02449_),
    .Q_N(_12939_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3311),
    .D(_02450_),
    .Q_N(_12938_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3312),
    .D(_02451_),
    .Q_N(_12937_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3313),
    .D(_02452_),
    .Q_N(_12936_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3314),
    .D(_02453_),
    .Q_N(_12935_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3315),
    .D(_02454_),
    .Q_N(_12934_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3316),
    .D(_02455_),
    .Q_N(_12933_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3317),
    .D(_02456_),
    .Q_N(_14925_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3318),
    .D(_00036_),
    .Q_N(_00267_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3319),
    .D(_00037_),
    .Q_N(_14926_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3320),
    .D(_00038_),
    .Q_N(_14927_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3321),
    .D(_00039_),
    .Q_N(_14928_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3322),
    .D(_00040_),
    .Q_N(_14929_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3323),
    .D(_00041_),
    .Q_N(_14930_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3324),
    .D(_00042_),
    .Q_N(_12932_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3325),
    .D(_02457_),
    .Q_N(_12931_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3326),
    .D(_02458_),
    .Q_N(_12930_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3327),
    .D(_02459_),
    .Q_N(_12929_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3328),
    .D(_02460_),
    .Q_N(_14931_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3329),
    .D(_00043_),
    .Q_N(_12928_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3330),
    .D(_02461_),
    .Q_N(_12927_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3331),
    .D(_02462_),
    .Q_N(_12926_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3332),
    .D(_02463_),
    .Q_N(_12925_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3333),
    .D(_02464_),
    .Q_N(_12924_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3334),
    .D(_02465_),
    .Q_N(_12923_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3335),
    .D(_02466_),
    .Q_N(_12922_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3336),
    .D(_02467_),
    .Q_N(_12921_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3337),
    .D(_02468_),
    .Q_N(_12920_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3338),
    .D(_02469_),
    .Q_N(_12919_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3339),
    .D(_02470_),
    .Q_N(_14932_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3340),
    .D(_00044_),
    .Q_N(_12918_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3341),
    .D(_02471_),
    .Q_N(_12917_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3342),
    .D(_02472_),
    .Q_N(_14933_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3343),
    .D(_00045_),
    .Q_N(_14934_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3344),
    .D(_00046_),
    .Q_N(_14935_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3345),
    .D(_00047_),
    .Q_N(_14936_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3346),
    .D(_00048_),
    .Q_N(_14937_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3347),
    .D(_00049_),
    .Q_N(_14938_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3348),
    .D(_00050_),
    .Q_N(_14939_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3349),
    .D(_00051_),
    .Q_N(_12916_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3350),
    .D(_02473_),
    .Q_N(_12915_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3351),
    .D(_02474_),
    .Q_N(_12914_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3352),
    .D(_02475_),
    .Q_N(_12913_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3353),
    .D(_02476_),
    .Q_N(_12912_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3354),
    .D(_02477_),
    .Q_N(_12911_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3355),
    .D(_02478_),
    .Q_N(_12910_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3356),
    .D(_02479_),
    .Q_N(_14940_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3357),
    .D(_00055_),
    .Q_N(_00266_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3358),
    .D(_00056_),
    .Q_N(_14941_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3359),
    .D(_00057_),
    .Q_N(_14942_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3360),
    .D(_00058_),
    .Q_N(_14943_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3361),
    .D(_00059_),
    .Q_N(_14944_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3362),
    .D(_00060_),
    .Q_N(_14945_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3363),
    .D(_00061_),
    .Q_N(_14946_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3364),
    .D(_00062_),
    .Q_N(_14947_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3365),
    .D(_00063_),
    .Q_N(_14948_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3366),
    .D(_00064_),
    .Q_N(_14949_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3367),
    .D(_00065_),
    .Q_N(_14950_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3368),
    .D(_00066_),
    .Q_N(_14951_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3369),
    .D(_00067_),
    .Q_N(_14952_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3370),
    .D(_00068_),
    .Q_N(_14953_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3371),
    .D(_00069_),
    .Q_N(_14954_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3372),
    .D(_00070_),
    .Q_N(_14955_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3373),
    .D(_00071_),
    .Q_N(_14956_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3374),
    .D(_00072_),
    .Q_N(_14957_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3375),
    .D(_00073_),
    .Q_N(_14958_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3376),
    .D(_00074_),
    .Q_N(_14959_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3377),
    .D(_00075_),
    .Q_N(_14960_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3378),
    .D(_00076_),
    .Q_N(_14961_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3379),
    .D(_00077_),
    .Q_N(_14962_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3380),
    .D(_00078_),
    .Q_N(_12909_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3381),
    .D(_02480_),
    .Q_N(_12908_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3382),
    .D(_02481_),
    .Q_N(_12907_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3383),
    .D(_02482_),
    .Q_N(_12906_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3384),
    .D(_02483_),
    .Q_N(_12905_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3385),
    .D(_02484_),
    .Q_N(_12904_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3386),
    .D(_02485_),
    .Q_N(_12903_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3387),
    .D(_02486_),
    .Q_N(_12902_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3388),
    .D(_02487_),
    .Q_N(_12901_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3389),
    .D(_02488_),
    .Q_N(_12900_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3390),
    .D(_02489_),
    .Q_N(_12899_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3391),
    .D(_02490_),
    .Q_N(_12898_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3392),
    .D(_02491_),
    .Q_N(_12897_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3393),
    .D(_02492_),
    .Q_N(_12896_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3394),
    .D(_02493_),
    .Q_N(_12895_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3395),
    .D(_02494_),
    .Q_N(_12894_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3396),
    .D(_02495_),
    .Q_N(_12893_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3397),
    .D(_02496_),
    .Q_N(_12892_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3398),
    .D(_02497_),
    .Q_N(_12891_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3399),
    .D(_02498_),
    .Q_N(_12890_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3400),
    .D(_02499_),
    .Q_N(_12889_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3401),
    .D(_02500_),
    .Q_N(_12888_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3402),
    .D(_02501_),
    .Q_N(_12887_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3403),
    .D(_02502_),
    .Q_N(_12886_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3404),
    .D(_02503_),
    .Q_N(_12885_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3405),
    .D(_02504_),
    .Q_N(_00168_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3406),
    .D(_02505_),
    .Q_N(_12884_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3407),
    .D(_02506_),
    .Q_N(_00167_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3408),
    .D(_02507_),
    .Q_N(_12883_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3409),
    .D(_02508_),
    .Q_N(_00232_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3410),
    .D(_02509_),
    .Q_N(_12882_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3411),
    .D(_02510_),
    .Q_N(_12881_),
    .Q(net21));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3412),
    .D(_02511_),
    .Q_N(_12880_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3413),
    .D(_02512_),
    .Q_N(_12879_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3414),
    .D(_02513_),
    .Q_N(_12878_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3415),
    .D(_02514_),
    .Q_N(_12877_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3416),
    .D(_02515_),
    .Q_N(_12876_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3417),
    .D(_02516_),
    .Q_N(_12875_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3418),
    .D(_02517_),
    .Q_N(_12874_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3419),
    .D(_02518_),
    .Q_N(_12873_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3420),
    .D(_02519_),
    .Q_N(_12872_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3421),
    .D(_02520_),
    .Q_N(_12871_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3422),
    .D(_02521_),
    .Q_N(_12870_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3423),
    .D(_02522_),
    .Q_N(_12869_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3424),
    .D(_02523_),
    .Q_N(_12868_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3425),
    .D(_02524_),
    .Q_N(_12867_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3426),
    .D(_02525_),
    .Q_N(_12866_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3427),
    .D(_02526_),
    .Q_N(_12865_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3428),
    .D(_02527_),
    .Q_N(_12864_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3429),
    .D(_02528_),
    .Q_N(_12863_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3430),
    .D(_02529_),
    .Q_N(_12862_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3431),
    .D(_02530_),
    .Q_N(_12861_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3432),
    .D(_02531_),
    .Q_N(_12860_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3433),
    .D(_02532_),
    .Q_N(_14963_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net3434),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14964_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3435),
    .D(_00021_),
    .Q_N(_00258_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3436),
    .D(_00008_),
    .Q_N(_14965_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3437),
    .D(_00022_),
    .Q_N(_14966_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3438),
    .D(_00023_),
    .Q_N(_14967_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3439),
    .D(_00009_),
    .Q_N(_14968_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3440),
    .D(_00024_),
    .Q_N(_14969_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net3441),
    .D(_00010_),
    .Q_N(_14970_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3442),
    .D(_00025_),
    .Q_N(_14971_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3443),
    .D(_00026_),
    .Q_N(_14972_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3444),
    .D(_00001_),
    .Q_N(_14973_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3445),
    .D(_00027_),
    .Q_N(_14974_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3446),
    .D(_00002_),
    .Q_N(_14975_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3447),
    .D(_00028_),
    .Q_N(_14976_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3448),
    .D(_00003_),
    .Q_N(_14977_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3449),
    .D(_00004_),
    .Q_N(_14978_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3450),
    .D(_00005_),
    .Q_N(_14979_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3451),
    .D(_00006_),
    .Q_N(_00169_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3452),
    .D(_00007_),
    .Q_N(_12859_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3453),
    .D(_02533_),
    .Q_N(_12858_),
    .Q(net4));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3454),
    .D(_02534_),
    .Q_N(_12857_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3455),
    .D(_02535_),
    .Q_N(_12856_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3456),
    .D(_02536_),
    .Q_N(_12855_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3457),
    .D(_02537_),
    .Q_N(_12854_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3458),
    .D(_02538_),
    .Q_N(_14980_),
    .Q(net15));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net3459),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14981_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net3460),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00233_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3461),
    .D(_02539_),
    .Q_N(_12853_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3462),
    .D(_02540_),
    .Q_N(_12852_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3463),
    .D(_02541_),
    .Q_N(_12851_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3464),
    .D(_02542_),
    .Q_N(_12850_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3465),
    .D(_02543_),
    .Q_N(_00298_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3466),
    .D(_02544_),
    .Q_N(_00303_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3467),
    .D(_02545_),
    .Q_N(_00093_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3468),
    .D(_02546_),
    .Q_N(_00103_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3469),
    .D(_02547_),
    .Q_N(_00113_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3470),
    .D(_02548_),
    .Q_N(_00119_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3471),
    .D(_02549_),
    .Q_N(_00130_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3472),
    .D(_02550_),
    .Q_N(_00141_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3473),
    .D(_02551_),
    .Q_N(_00297_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3474),
    .D(_02552_),
    .Q_N(_00302_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3475),
    .D(_02553_),
    .Q_N(_00092_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3476),
    .D(_02554_),
    .Q_N(_00102_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3477),
    .D(_02555_),
    .Q_N(_00112_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3478),
    .D(_02556_),
    .Q_N(_00118_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3479),
    .D(_02557_),
    .Q_N(_00129_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3480),
    .D(_02558_),
    .Q_N(_00140_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3481),
    .D(_02559_),
    .Q_N(_12849_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3482),
    .D(_02560_),
    .Q_N(_12848_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3483),
    .D(_02561_),
    .Q_N(_12847_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3484),
    .D(_02562_),
    .Q_N(_12846_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3485),
    .D(_02563_),
    .Q_N(_12845_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3486),
    .D(_02564_),
    .Q_N(_12844_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3487),
    .D(_02565_),
    .Q_N(_12843_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3488),
    .D(_02566_),
    .Q_N(_12842_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3489),
    .D(_02567_),
    .Q_N(_12841_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3490),
    .D(_02568_),
    .Q_N(_12840_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3491),
    .D(_02569_),
    .Q_N(_12839_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3492),
    .D(_02570_),
    .Q_N(_12838_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3493),
    .D(_02571_),
    .Q_N(_12837_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3494),
    .D(_02572_),
    .Q_N(_12836_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3495),
    .D(_02573_),
    .Q_N(_12835_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3496),
    .D(_02574_),
    .Q_N(_12834_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3497),
    .D(_02575_),
    .Q_N(_12833_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3498),
    .D(_02576_),
    .Q_N(_12832_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3499),
    .D(_02577_),
    .Q_N(_12831_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3500),
    .D(_02578_),
    .Q_N(_12830_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3501),
    .D(_02579_),
    .Q_N(_12829_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3502),
    .D(_02580_),
    .Q_N(_12828_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3503),
    .D(_02581_),
    .Q_N(_12827_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3504),
    .D(_02582_),
    .Q_N(_12826_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3505),
    .D(_02583_),
    .Q_N(_12825_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3506),
    .D(_02584_),
    .Q_N(_12824_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3507),
    .D(_02585_),
    .Q_N(_00202_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3508),
    .D(_02586_),
    .Q_N(_12823_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3509),
    .D(_02587_),
    .Q_N(_00205_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3510),
    .D(_02588_),
    .Q_N(_12822_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3511),
    .D(_02589_),
    .Q_N(_12821_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3512),
    .D(_02590_),
    .Q_N(_12820_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3513),
    .D(_02591_),
    .Q_N(_12819_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3514),
    .D(_02592_),
    .Q_N(_12818_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3515),
    .D(_02593_),
    .Q_N(_12817_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3516),
    .D(_02594_),
    .Q_N(_12816_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3517),
    .D(_02595_),
    .Q_N(_12815_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3518),
    .D(_02596_),
    .Q_N(_12814_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3519),
    .D(_02597_),
    .Q_N(_12813_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3520),
    .D(_02598_),
    .Q_N(_12812_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3521),
    .D(_02599_),
    .Q_N(_12811_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3522),
    .D(_02600_),
    .Q_N(_12810_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3523),
    .D(_02601_),
    .Q_N(_12809_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3524),
    .D(_02602_),
    .Q_N(_00201_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3525),
    .D(_02603_),
    .Q_N(_12808_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3526),
    .D(_02604_),
    .Q_N(_12807_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3527),
    .D(_02605_),
    .Q_N(_00263_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3528),
    .D(_02606_),
    .Q_N(_00264_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net3529),
    .D(_02607_),
    .Q_N(_14982_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3530),
    .D(_00029_),
    .Q_N(_14983_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3531),
    .D(_00030_),
    .Q_N(_00206_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3532),
    .D(_00031_),
    .Q_N(_14984_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3533),
    .D(_00032_),
    .Q_N(_14985_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3534),
    .D(_00033_),
    .Q_N(_00259_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3535),
    .D(_00034_),
    .Q_N(_14986_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3536),
    .D(_00035_),
    .Q_N(_00207_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3537),
    .D(_02608_),
    .Q_N(_12806_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3538),
    .D(_02609_),
    .Q_N(_12805_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3539),
    .D(_02610_),
    .Q_N(_12804_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3540),
    .D(_02611_),
    .Q_N(_12803_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3541),
    .D(_02612_),
    .Q_N(_12802_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3542),
    .D(_02613_),
    .Q_N(_12801_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3543),
    .D(_02614_),
    .Q_N(_12800_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3544),
    .D(_02615_),
    .Q_N(_12799_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3545),
    .D(_02616_),
    .Q_N(_00265_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3546),
    .D(_02617_),
    .Q_N(_12798_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3547),
    .D(_02618_),
    .Q_N(_12797_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3548),
    .D(_02619_),
    .Q_N(_12796_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3549),
    .D(_02620_),
    .Q_N(_12795_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3550),
    .D(_02621_),
    .Q_N(_12794_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3551),
    .D(_02622_),
    .Q_N(_12793_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3552),
    .D(_02623_),
    .Q_N(_14987_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3553),
    .D(_00079_),
    .Q_N(_00260_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3554),
    .D(_00080_),
    .Q_N(_14988_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3555),
    .D(_00081_),
    .Q_N(_14989_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3556),
    .D(_00082_),
    .Q_N(_14990_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3557),
    .D(_00083_),
    .Q_N(_14991_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3558),
    .D(_00084_),
    .Q_N(_14992_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3559),
    .D(_00085_),
    .Q_N(_14993_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3560),
    .D(_00086_),
    .Q_N(_14994_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3561),
    .D(_00087_),
    .Q_N(_14995_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3562),
    .D(_00088_),
    .Q_N(_14996_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3563),
    .D(_00089_),
    .Q_N(_14997_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3564),
    .D(_00090_),
    .Q_N(_12792_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3565),
    .D(_02624_),
    .Q_N(_12791_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3566),
    .D(_02625_),
    .Q_N(_12790_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3567),
    .D(_02626_),
    .Q_N(_12789_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3568),
    .D(_02627_),
    .Q_N(_12788_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3569),
    .D(_02628_),
    .Q_N(_12787_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3570),
    .D(_02629_),
    .Q_N(_12786_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3571),
    .D(_02630_),
    .Q_N(_12785_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3572),
    .D(_02631_),
    .Q_N(_12784_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3573),
    .D(_02632_),
    .Q_N(_12783_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3574),
    .D(_02633_),
    .Q_N(_12782_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3575),
    .D(_02634_),
    .Q_N(_12781_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3576),
    .D(_02635_),
    .Q_N(_12780_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3577),
    .D(_02636_),
    .Q_N(_12779_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3578),
    .D(_02637_),
    .Q_N(_12778_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3579),
    .D(_02638_),
    .Q_N(_12777_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3580),
    .D(_02639_),
    .Q_N(_12776_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3581),
    .D(_02640_),
    .Q_N(_12775_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3582),
    .D(_02641_),
    .Q_N(_12774_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3583),
    .D(_02642_),
    .Q_N(_12773_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3584),
    .D(_02643_),
    .Q_N(_12772_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3585),
    .D(_02644_),
    .Q_N(_12771_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3586),
    .D(_02645_),
    .Q_N(_12770_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3587),
    .D(_02646_),
    .Q_N(_12769_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3588),
    .D(_02647_),
    .Q_N(_12768_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3589),
    .D(_02648_),
    .Q_N(_12767_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3590),
    .D(_02649_),
    .Q_N(_12766_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3591),
    .D(_02650_),
    .Q_N(_12765_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3592),
    .D(_02651_),
    .Q_N(_12764_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3593),
    .D(_02652_),
    .Q_N(_12763_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3594),
    .D(_02653_),
    .Q_N(_12762_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3595),
    .D(_02654_),
    .Q_N(_12761_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3596),
    .D(_02655_),
    .Q_N(_12760_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3597),
    .D(_02656_),
    .Q_N(_12759_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3598),
    .D(_02657_),
    .Q_N(_12758_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3599),
    .D(_02658_),
    .Q_N(_14998_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3600),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12757_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3601),
    .D(_02659_),
    .Q_N(_12756_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3602),
    .D(_02660_),
    .Q_N(_12755_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3603),
    .D(_02661_),
    .Q_N(_12754_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3604),
    .D(_02662_),
    .Q_N(_12753_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3605),
    .D(_02663_),
    .Q_N(_12752_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3606),
    .D(_02664_),
    .Q_N(_12751_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3607),
    .D(_02665_),
    .Q_N(_12750_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3608),
    .D(_02666_),
    .Q_N(_12749_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3609),
    .D(_02667_),
    .Q_N(_12748_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3610),
    .D(_02668_),
    .Q_N(_12747_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3611),
    .D(_02669_),
    .Q_N(_00261_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3612),
    .D(_02670_),
    .Q_N(_12746_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3613),
    .D(_02671_),
    .Q_N(_12745_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3614),
    .D(_02672_),
    .Q_N(_12744_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3615),
    .D(_02673_),
    .Q_N(_12743_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3616),
    .D(_02674_),
    .Q_N(_12742_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3617),
    .D(_02675_),
    .Q_N(_14999_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3618),
    .D(_00000_),
    .Q_N(_12741_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[5]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[0]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[1]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[2]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[3]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[4]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[5]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[6]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_oe[7]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[0]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[1]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[2]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[3]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[4]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[5]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[6]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_out[7]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[0]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[1]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[2]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[3]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[4]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[5]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[6]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout28 (.A(_11364_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_06742_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_07344_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_07017_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_07263_),
    .X(net32));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(_07219_));
 sg13g2_buf_2 fanout34 (.A(_04971_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_03992_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02827_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02799_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02773_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02765_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02710_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02676_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_12716_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_12708_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_12653_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12619_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12593_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12584_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12506_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12480_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12472_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12418_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12388_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12363_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12355_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12298_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12264_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12238_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12230_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12173_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_12140_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12112_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_12102_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_11979_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_11923_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_11902_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_06406_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06392_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_06383_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_05691_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_05689_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_05176_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_04961_));
 sg13g2_buf_2 fanout73 (.A(_04750_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_03703_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_03561_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_12539_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_12038_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_11579_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_10724_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_06731_));
 sg13g2_buf_4 fanout81 (.X(net81),
    .A(_06725_));
 sg13g2_buf_2 fanout82 (.A(_05155_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04187_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03837_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_11439_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_11406_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_11369_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_09221_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_07447_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_07002_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_06844_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_06821_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_04070_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_03979_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_03096_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_11368_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_11336_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_10111_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_10100_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_10055_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_10048_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_09955_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_09944_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_09943_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_09836_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_09220_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_09062_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_08855_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_07924_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_07442_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_04069_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_03866_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_03862_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_03853_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_03843_),
    .X(net115));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(_03258_));
 sg13g2_buf_2 fanout117 (.A(_03146_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_11240_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_10040_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_09837_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_09067_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_08856_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_08854_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_07808_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_07646_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_07436_),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_06728_));
 sg13g2_buf_2 fanout128 (.A(_06722_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_06369_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_04224_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_04213_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04189_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04061_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04053_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04046_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04043_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_03968_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_03895_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_03852_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_03242_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_11709_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_11707_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_09989_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_09980_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_07860_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_07837_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_07829_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_07812_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_07811_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_07737_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_07665_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_07656_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_07435_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_04065_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_04063_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_04057_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_04039_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_03924_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_03910_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_03899_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_03897_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_03893_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_03891_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_03872_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_03857_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_03838_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_02996_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_10292_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_07800_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_07698_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_07657_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_07639_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_07313_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03921_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_03909_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_03902_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_03896_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_03890_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_03885_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_03881_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_03877_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_03856_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_03847_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_03202_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_03144_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_03128_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_03015_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_02999_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_02995_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_02982_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_11600_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_11536_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_10879_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_10690_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_09852_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_09063_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_09054_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_09044_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_08989_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_04050_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_03839_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_03585_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_03222_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_03129_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_03098_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_03097_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_03071_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_03017_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_03007_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_11763_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_11695_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_11562_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_11452_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_11447_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_11030_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_10635_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_10426_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_09872_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_09064_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_09056_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_08933_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_04080_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_04054_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_03613_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_03124_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_03006_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_02994_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_11566_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_11522_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_11514_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_11454_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_11451_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_11432_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11421_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_11359_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_11243_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_10937_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_10914_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_10796_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_10717_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_10634_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_10483_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_10329_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_09871_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_06630_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_06597_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_06595_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_06594_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_06520_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_06355_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_06354_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_06298_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_06297_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_06185_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_06184_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_06070_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_06069_),
    .X(net257));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(_05954_));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(_05932_));
 sg13g2_buf_4 fanout260 (.X(net260),
    .A(_05915_));
 sg13g2_buf_4 fanout261 (.X(net261),
    .A(_05910_));
 sg13g2_buf_4 fanout262 (.X(net262),
    .A(_05892_));
 sg13g2_buf_4 fanout263 (.X(net263),
    .A(_05872_));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(_05869_));
 sg13g2_buf_4 fanout265 (.X(net265),
    .A(_05863_));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_05844_));
 sg13g2_buf_4 fanout267 (.X(net267),
    .A(_05822_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_05814_));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_05790_));
 sg13g2_buf_2 fanout270 (.A(_05206_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_03563_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_03559_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_03001_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_02993_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_11609_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_11497_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_11367_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_11253_),
    .X(net278));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(_10795_));
 sg13g2_buf_2 fanout280 (.A(_10761_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_10659_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_10601_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_10547_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_10456_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_10390_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_10364_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_09070_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_08405_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_06631_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_06616_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_06614_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_06613_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_06519_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_06343_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_06342_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_06286_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_06285_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_06274_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_06273_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_06262_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_06261_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_06250_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_06249_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_06238_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06237_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06225_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06224_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06169_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06168_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06156_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06155_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06144_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06143_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_06132_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_06131_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_06121_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_06120_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_06109_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06108_),
    .X(net319));
 sg13g2_buf_2 fanout320 (.A(_06056_),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(_06055_),
    .X(net321));
 sg13g2_buf_2 fanout322 (.A(_06039_),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(_06038_),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(_06026_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(_06025_),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(_06013_),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(_06012_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_06000_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_05999_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_05963_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05962_),
    .X(net331));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_05951_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_05948_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_05943_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_05937_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_05928_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_05925_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05922_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_05919_));
 sg13g2_buf_4 fanout340 (.X(net340),
    .A(_05903_));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(_05898_));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(_05889_));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_05884_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_05876_));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(_05858_));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(_05851_));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_05840_));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(_05834_));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(_05831_));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(_05808_));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(_05802_));
 sg13g2_buf_2 fanout352 (.A(_03981_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_03053_),
    .X(net353));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(_02939_));
 sg13g2_buf_2 fanout355 (.A(_02937_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_02914_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_02912_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_10658_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_10567_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_09211_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_08507_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_08439_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_06670_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_06668_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_06667_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_06574_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_06457_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_06331_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_06330_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_06320_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_06319_),
    .X(net371));
 sg13g2_buf_2 fanout372 (.A(_06309_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_06308_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_06211_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_06210_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_06198_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_06197_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_06096_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_06095_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_06083_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_06082_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_05988_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_05987_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_05977_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_05976_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_05015_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_04982_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_04906_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_04891_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_04849_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_04401_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_03729_),
    .X(net392));
 sg13g2_buf_4 fanout393 (.X(net393),
    .A(_02981_));
 sg13g2_buf_4 fanout394 (.X(net394),
    .A(_02980_));
 sg13g2_buf_4 fanout395 (.X(net395),
    .A(_02964_));
 sg13g2_buf_2 fanout396 (.A(_02963_),
    .X(net396));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_02940_));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(_02915_));
 sg13g2_buf_2 fanout399 (.A(_12176_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_12030_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_11425_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_11419_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_11292_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_09804_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_09661_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_09636_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_09590_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_09566_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_09307_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_09210_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_08841_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_08819_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_08798_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_08581_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_08547_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_06689_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_06687_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_06686_),
    .X(net418));
 sg13g2_buf_2 fanout419 (.A(_06651_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_06649_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_06648_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_06575_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_06456_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_06366_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_06365_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_06364_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_05285_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_05035_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_04974_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_04909_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_04896_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_04708_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_04706_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_03483_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_03475_),
    .X(net435));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(_02976_));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(_02973_));
 sg13g2_buf_2 fanout438 (.A(_02962_),
    .X(net438));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(_02961_));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_02960_));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(_02957_));
 sg13g2_buf_2 fanout442 (.A(_02904_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_02829_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_11424_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_11418_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_10727_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_10045_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_09532_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_09385_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_09275_),
    .X(net450));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(_08996_));
 sg13g2_buf_2 fanout452 (.A(_08776_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_08752_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_08728_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_08706_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_08549_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_08474_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_08455_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_08402_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_07018_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_06708_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_06706_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_06705_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_06035_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_05974_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_05905_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_05853_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_05828_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_05793_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_05779_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_05696_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_04821_),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_04787_));
 sg13g2_buf_2 fanout474 (.A(_04766_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_04758_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_04705_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_03479_),
    .X(net477));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(_02977_));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(_02974_));
 sg13g2_buf_4 fanout480 (.X(net480),
    .A(_02958_));
 sg13g2_buf_2 fanout481 (.A(_02903_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_02896_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_02892_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_02889_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_02762_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_02712_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_12655_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_12421_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_12300_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_12097_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_12068_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_12064_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_12057_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_12053_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_12046_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_12042_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_12034_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_11937_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_11417_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_11316_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_10251_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_10044_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_10036_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_09278_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_09274_),
    .X(net505));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(_09243_));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(_09166_));
 sg13g2_buf_2 fanout508 (.A(_08730_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_08653_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_08601_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_08556_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_08551_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_08548_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_08488_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_08482_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_08473_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_08454_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_07557_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_06235_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_06221_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_06214_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_06208_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_06200_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_06189_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_06106_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_06093_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_06086_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_06080_),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_06072_),
    .X(net529));
 sg13g2_buf_2 fanout530 (.A(_06060_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_05973_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_04981_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_04914_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_04806_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_04782_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_04757_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_04755_),
    .X(net537));
 sg13g2_buf_2 fanout538 (.A(_04709_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_04699_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_04696_),
    .X(net540));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_04695_));
 sg13g2_buf_2 fanout542 (.A(_03553_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_03545_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_03539_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_03537_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_03535_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_03520_),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_03519_));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(_03515_));
 sg13g2_buf_4 fanout550 (.X(net550),
    .A(_03482_));
 sg13g2_buf_4 fanout551 (.X(net551),
    .A(_03478_));
 sg13g2_buf_2 fanout552 (.A(_03473_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_03468_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_03466_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_03462_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_02979_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_02938_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_02911_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_02907_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_02902_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_02900_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_02895_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_02891_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_02888_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_12469_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_12352_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_11906_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_11467_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_10250_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(_10238_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_10035_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_09593_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_09267_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_09242_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_09165_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_08625_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_08564_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_08550_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_08487_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_08481_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_08472_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_08453_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_07348_),
    .X(net583));
 sg13g2_buf_2 fanout584 (.A(_07220_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_07019_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_05912_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_05904_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_05893_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_05860_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_05852_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_05841_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_05792_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_04979_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_04977_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_04893_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_04777_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_04753_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_04698_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_03544_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_03536_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_03527_),
    .X(net601));
 sg13g2_buf_4 fanout602 (.X(net602),
    .A(_03525_));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(_03512_));
 sg13g2_buf_2 fanout604 (.A(_03500_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_03499_),
    .X(net605));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_03494_));
 sg13g2_buf_4 fanout607 (.X(net607),
    .A(_03489_));
 sg13g2_buf_2 fanout608 (.A(_03477_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_03472_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_03467_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_03465_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_03461_),
    .X(net612));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(_02910_));
 sg13g2_buf_2 fanout614 (.A(_02906_),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(_02899_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_02894_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_11889_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_11378_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_10941_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_10875_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_10838_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_10224_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_10213_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_10166_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_10148_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_09792_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_09678_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_09487_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_09478_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_09426_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_09336_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_09331_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_09241_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_09164_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_08902_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_08563_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_08559_),
    .X(net637));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(_08511_));
 sg13g2_buf_2 fanout639 (.A(_08486_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_08480_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_08471_),
    .X(net641));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(_08465_));
 sg13g2_buf_2 fanout643 (.A(_08452_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_08062_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_07947_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_07918_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_07895_),
    .X(net647));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(_07877_));
 sg13g2_buf_2 fanout649 (.A(_07852_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_07825_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_07786_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_07753_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_07713_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_07621_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_07534_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_07009_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_06800_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_06173_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_06043_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_05916_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_05864_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_05803_),
    .X(net662));
 sg13g2_buf_2 fanout663 (.A(_05002_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_04965_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_04958_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_04885_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_04776_),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_04734_));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_03541_));
 sg13g2_buf_2 fanout670 (.A(_03531_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_03530_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_03526_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_03471_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_03469_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_02920_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_02909_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_12705_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_12227_),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_11879_));
 sg13g2_buf_2 fanout680 (.A(_11839_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_11835_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_11776_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_10886_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_10842_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_10226_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_10220_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_10196_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_10190_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_10179_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_10176_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_10147_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_09910_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_09904_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_09830_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_09575_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_09563_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_09484_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_09483_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_09481_),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_09479_));
 sg13g2_buf_8 fanout701 (.A(_09465_),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(_09462_),
    .X(net702));
 sg13g2_buf_4 fanout703 (.X(net703),
    .A(_09439_));
 sg13g2_buf_8 fanout704 (.A(_09427_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_09322_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_09314_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_09298_),
    .X(net707));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(_09294_));
 sg13g2_buf_8 fanout709 (.A(_09284_),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(_09265_),
    .X(net710));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_09254_));
 sg13g2_buf_2 fanout712 (.A(_09233_),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(_09163_));
 sg13g2_buf_4 fanout714 (.X(net714),
    .A(_09142_));
 sg13g2_buf_2 fanout715 (.A(_09084_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_08778_),
    .X(net716));
 sg13g2_buf_4 fanout717 (.X(net717),
    .A(_08608_));
 sg13g2_buf_8 fanout718 (.A(_08540_),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(_08536_),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(_08529_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_08516_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_08510_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_08464_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_08461_));
 sg13g2_buf_8 fanout725 (.A(_08418_),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(_08411_),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_08408_));
 sg13g2_buf_2 fanout728 (.A(_06191_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_06180_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_06178_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_06176_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_06062_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_06050_),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(_06048_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_06046_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_05911_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_05859_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_05795_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_05791_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_04964_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_03529_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_03507_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_03506_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_03470_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_02948_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_02946_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_02933_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_02929_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_02926_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_02923_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_02919_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_12648_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_12645_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_12581_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_12025_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_12019_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_11843_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_11838_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_10892_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_10887_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_10850_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_10847_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_10819_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_10816_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_10813_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_10434_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_10429_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_10306_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_10301_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_10229_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_10219_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_10210_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_10207_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_10202_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_10195_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_10189_),
    .X(net776));
 sg13g2_buf_4 fanout777 (.X(net777),
    .A(_10178_));
 sg13g2_buf_2 fanout778 (.A(_10175_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_09903_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_09902_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_09594_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_09537_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_09492_),
    .X(net783));
 sg13g2_buf_4 fanout784 (.X(net784),
    .A(_09466_));
 sg13g2_buf_4 fanout785 (.X(net785),
    .A(_09461_));
 sg13g2_buf_4 fanout786 (.X(net786),
    .A(_09440_));
 sg13g2_buf_4 fanout787 (.X(net787),
    .A(_09432_));
 sg13g2_buf_4 fanout788 (.X(net788),
    .A(_09428_));
 sg13g2_buf_2 fanout789 (.A(_09387_),
    .X(net789));
 sg13g2_buf_4 fanout790 (.X(net790),
    .A(_09351_));
 sg13g2_buf_8 fanout791 (.A(_09343_),
    .X(net791));
 sg13g2_buf_4 fanout792 (.X(net792),
    .A(_09301_));
 sg13g2_buf_4 fanout793 (.X(net793),
    .A(_09293_));
 sg13g2_buf_4 fanout794 (.X(net794),
    .A(_09287_));
 sg13g2_buf_4 fanout795 (.X(net795),
    .A(_09283_));
 sg13g2_buf_2 fanout796 (.A(_09253_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_09246_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_09232_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_09162_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(_09157_),
    .X(net800));
 sg13g2_buf_2 fanout801 (.A(_09141_),
    .X(net801));
 sg13g2_buf_2 fanout802 (.A(_09083_),
    .X(net802));
 sg13g2_buf_2 fanout803 (.A(_08991_),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(_08692_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_08670_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_08607_),
    .X(net806));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(_08541_));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_08537_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_08534_));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_08531_));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(_08528_));
 sg13g2_buf_2 fanout812 (.A(_08517_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_08515_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_08509_),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_08463_));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(_08460_));
 sg13g2_buf_2 fanout817 (.A(_08458_),
    .X(net817));
 sg13g2_buf_4 fanout818 (.X(net818),
    .A(_08432_));
 sg13g2_buf_2 fanout819 (.A(_08428_),
    .X(net819));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(_08424_));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(_08422_));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(_08416_));
 sg13g2_buf_4 fanout823 (.X(net823),
    .A(_08414_));
 sg13g2_buf_4 fanout824 (.X(net824),
    .A(_08410_));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_08407_));
 sg13g2_buf_2 fanout826 (.A(_08311_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_07225_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_06843_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_06825_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_06818_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_06539_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_06517_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_06500_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_06472_),
    .X(net834));
 sg13g2_buf_2 fanout835 (.A(_06436_),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_06385_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_06381_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_06234_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_06105_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_05972_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_05878_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_05877_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_05873_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_05824_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_05823_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_05815_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_05760_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_05756_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_03509_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_03508_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_03502_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_03495_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_03455_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_03011_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_02956_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_02954_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_02952_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_02950_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_02947_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_02945_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_02932_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_02928_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_02925_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_02922_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_02804_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_12631_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_12399_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_12282_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_12269_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_11997_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_11994_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_11990_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_11855_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_11834_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_11827_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_11810_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_11414_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_10894_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_10863_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_10852_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_10835_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_10812_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_10809_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_10806_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_10802_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_10801_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_10540_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_10299_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_10281_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_10243_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_10218_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_10194_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_10186_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_10185_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_10177_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_10174_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_10151_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_10057_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_10049_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_09997_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_09901_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_09769_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_09454_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_09446_),
    .X(net904));
 sg13g2_buf_4 fanout905 (.X(net905),
    .A(_09435_));
 sg13g2_buf_2 fanout906 (.A(_09431_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_09371_),
    .X(net907));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(_09352_));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(_09344_));
 sg13g2_buf_2 fanout910 (.A(_09319_),
    .X(net910));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(_09295_));
 sg13g2_buf_4 fanout912 (.X(net912),
    .A(_09290_));
 sg13g2_buf_2 fanout913 (.A(_09286_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_09251_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_09245_),
    .X(net915));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(_09231_));
 sg13g2_buf_2 fanout917 (.A(_09161_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09140_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_09082_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_08897_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_08868_),
    .X(net921));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(_08695_));
 sg13g2_buf_4 fanout923 (.X(net923),
    .A(_08654_));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(_08530_));
 sg13g2_buf_2 fanout925 (.A(_08514_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_08477_),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_08462_));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(_08459_));
 sg13g2_buf_2 fanout929 (.A(_08457_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_08431_),
    .X(net930));
 sg13g2_buf_4 fanout931 (.X(net931),
    .A(_08427_));
 sg13g2_buf_2 fanout932 (.A(_08423_),
    .X(net932));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(_08421_));
 sg13g2_buf_4 fanout934 (.X(net934),
    .A(_08413_));
 sg13g2_buf_2 fanout935 (.A(_08281_),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_07329_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_07325_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_07315_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_07303_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_07300_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_06817_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_06557_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_06556_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_06555_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_06553_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_06541_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_06537_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_06533_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_06516_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_06514_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_06512_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_06502_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_06499_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_06497_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_06476_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_06470_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_06464_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_06442_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_06429_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_06417_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_05881_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_05880_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_05879_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_05827_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_05826_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_05825_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_05772_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_05755_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_05747_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_05740_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_04817_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_04778_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_04688_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_04648_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_04589_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_04562_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_04534_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_04033_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_03969_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_03463_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_03454_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_03424_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_03010_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_02953_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_02951_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_02949_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_02877_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_02779_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_12551_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_12500_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_12425_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_12419_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_12411_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_12409_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_12324_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_12271_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_12247_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_12203_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_12129_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_12093_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_12089_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_12086_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_12082_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_12078_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_12015_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_12011_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_11980_),
    .X(net1007));
 sg13g2_buf_4 fanout1008 (.X(net1008),
    .A(_11960_));
 sg13g2_buf_2 fanout1009 (.A(_11947_),
    .X(net1009));
 sg13g2_buf_4 fanout1010 (.X(net1010),
    .A(_11941_));
 sg13g2_buf_4 fanout1011 (.X(net1011),
    .A(_11926_));
 sg13g2_buf_2 fanout1012 (.A(_11919_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_11910_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_11909_),
    .X(net1014));
 sg13g2_buf_4 fanout1015 (.X(net1015),
    .A(_11905_));
 sg13g2_buf_2 fanout1016 (.A(_11833_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_11817_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_11816_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_11814_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_11809_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_11646_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_11530_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_11261_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_10808_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_10805_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_10798_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_10797_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_10324_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_10295_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_10242_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_10182_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_10181_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_10173_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_10168_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_10167_),
    .X(net1035));
 sg13g2_buf_4 fanout1036 (.X(net1036),
    .A(_10158_));
 sg13g2_buf_2 fanout1037 (.A(_10144_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_10078_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_10062_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_10051_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_10034_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_10020_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_10014_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_10008_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_10002_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_09996_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_09988_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_09848_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_09453_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_09309_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_09250_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_09244_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_09230_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_09217_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_09174_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_09160_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_09155_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_09151_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_09139_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_09074_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_09049_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_08858_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_08643_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_08615_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_08525_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_08450_),
    .X(net1066));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(_08446_));
 sg13g2_buf_2 fanout1068 (.A(_08443_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_08412_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_08409_),
    .X(net1070));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(_08388_));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(_08377_));
 sg13g2_buf_2 fanout1073 (.A(_08299_),
    .X(net1073));
 sg13g2_buf_4 fanout1074 (.X(net1074),
    .A(_08296_));
 sg13g2_buf_8 fanout1075 (.A(_08294_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_08291_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_08280_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_08097_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_08095_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_08079_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_08028_),
    .X(net1081));
 sg13g2_buf_2 fanout1082 (.A(_07406_),
    .X(net1082));
 sg13g2_buf_2 fanout1083 (.A(_07316_),
    .X(net1083));
 sg13g2_buf_2 fanout1084 (.A(_07301_),
    .X(net1084));
 sg13g2_buf_2 fanout1085 (.A(_07299_),
    .X(net1085));
 sg13g2_buf_2 fanout1086 (.A(_05734_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_02692_),
    .X(net1087));
 sg13g2_buf_2 fanout1088 (.A(_02686_),
    .X(net1088));
 sg13g2_buf_2 fanout1089 (.A(_02677_),
    .X(net1089));
 sg13g2_buf_2 fanout1090 (.A(_12607_),
    .X(net1090));
 sg13g2_buf_2 fanout1091 (.A(_12585_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_12452_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_12020_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_11998_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_11959_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_11940_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_11925_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_11907_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_11904_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_11881_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_11877_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_11860_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_11858_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_11851_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_11678_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_11675_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_11618_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_11495_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_11344_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_11275_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_10785_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_10781_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_10516_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_10160_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_10149_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_10142_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_10138_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_10033_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_10027_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_09907_),
    .X(net1120));
 sg13g2_buf_1 fanout1121 (.A(_09847_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_09801_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_09317_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_09277_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_09223_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_09216_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_09171_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_09143_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_09138_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_09066_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_08364_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_08341_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_08336_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_08332_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_08320_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_08289_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_08283_),
    .X(net1137));
 sg13g2_tiehi _27557__1138 (.L_HI(net1138));
 sg13g2_tiehi _27558__1139 (.L_HI(net1139));
 sg13g2_tiehi _27559__1140 (.L_HI(net1140));
 sg13g2_tiehi _27560__1141 (.L_HI(net1141));
 sg13g2_tiehi _27561__1142 (.L_HI(net1142));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1143  (.L_HI(net1143));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1144  (.L_HI(net1144));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1145  (.L_HI(net1145));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1146  (.L_HI(net1146));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1147  (.L_HI(net1147));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1148  (.L_HI(net1148));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1149  (.L_HI(net1149));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1150  (.L_HI(net1150));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1151  (.L_HI(net1151));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1152  (.L_HI(net1152));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1153  (.L_HI(net1153));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1154  (.L_HI(net1154));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1155  (.L_HI(net1155));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1156  (.L_HI(net1156));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1157  (.L_HI(net1157));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1158  (.L_HI(net1158));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1159  (.L_HI(net1159));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1160  (.L_HI(net1160));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1161  (.L_HI(net1161));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1162  (.L_HI(net1162));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1163  (.L_HI(net1163));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1164  (.L_HI(net1164));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1165  (.L_HI(net1165));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1166  (.L_HI(net1166));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1167  (.L_HI(net1167));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1168  (.L_HI(net1168));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1169  (.L_HI(net1169));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1170  (.L_HI(net1170));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1171  (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_DFFE_PP__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_DFFE_PP__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_DFFE_PP__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_DFFE_PP__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_DFFE_PP__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_DFFE_PP__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_DFFE_PP__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_DFFE_PP__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_DFFE_PP__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_DFFE_PP__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_DFFE_PP__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_DFFE_PP__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_DFFE_PP__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_DFFE_PP__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_DFFE_PP__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_DFFE_PP__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_DFFE_PP__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_DFFE_PP__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_DFFE_PP__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_DFFE_PP__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_DFFE_PP__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_DFFE_PP__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_DFFE_PP__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.spi.r_count[0]$_DFFE_PP__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.spi.r_count[1]$_DFFE_PP__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.spi.r_count[2]$_DFFE_PP__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_count[3]$_DFFE_PP__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_count[4]$_DFFE_PP__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_count[5]$_DFFE_PP__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_count[6]$_DFFE_PP__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_count[7]$_DFFE_PP__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_DFFE_PP__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_DFFE_PP__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_DFFE_PP__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_src[0]$_DFFE_PP__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_src[1]$_DFFE_PP__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_src[2]$_DFFE_PP__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3614  (.L_HI(net3614));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3615  (.L_HI(net3615));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3616  (.L_HI(net3616));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3617  (.L_HI(net3617));
 sg13g2_tiehi \r_reset$_DFF_P__3618  (.L_HI(net3618));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_63__leaf_clk));
 sg13g2_inv_4 clkload7 (.A(clknet_leaf_255_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_leaf_256_clk));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_262_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_263_clk));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_123_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_124_clk));
 sg13g2_buf_16 clkload13 (.A(clknet_leaf_125_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_121_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00203_));
 sg13g2_antennanp ANTENNA_2 (.A(_00203_));
 sg13g2_antennanp ANTENNA_3 (.A(_00209_));
 sg13g2_antennanp ANTENNA_4 (.A(_00784_));
 sg13g2_antennanp ANTENNA_5 (.A(_00923_));
 sg13g2_antennanp ANTENNA_6 (.A(_01032_));
 sg13g2_antennanp ANTENNA_7 (.A(_01034_));
 sg13g2_antennanp ANTENNA_8 (.A(_01034_));
 sg13g2_antennanp ANTENNA_9 (.A(_02779_));
 sg13g2_antennanp ANTENNA_10 (.A(_02779_));
 sg13g2_antennanp ANTENNA_11 (.A(_02779_));
 sg13g2_antennanp ANTENNA_12 (.A(_02779_));
 sg13g2_antennanp ANTENNA_13 (.A(_02910_));
 sg13g2_antennanp ANTENNA_14 (.A(_02910_));
 sg13g2_antennanp ANTENNA_15 (.A(_02910_));
 sg13g2_antennanp ANTENNA_16 (.A(_02910_));
 sg13g2_antennanp ANTENNA_17 (.A(_02910_));
 sg13g2_antennanp ANTENNA_18 (.A(_02910_));
 sg13g2_antennanp ANTENNA_19 (.A(_02910_));
 sg13g2_antennanp ANTENNA_20 (.A(_02910_));
 sg13g2_antennanp ANTENNA_21 (.A(_02910_));
 sg13g2_antennanp ANTENNA_22 (.A(_02932_));
 sg13g2_antennanp ANTENNA_23 (.A(_02932_));
 sg13g2_antennanp ANTENNA_24 (.A(_02932_));
 sg13g2_antennanp ANTENNA_25 (.A(_02955_));
 sg13g2_antennanp ANTENNA_26 (.A(_02955_));
 sg13g2_antennanp ANTENNA_27 (.A(_02955_));
 sg13g2_antennanp ANTENNA_28 (.A(_02955_));
 sg13g2_antennanp ANTENNA_29 (.A(_02955_));
 sg13g2_antennanp ANTENNA_30 (.A(_02955_));
 sg13g2_antennanp ANTENNA_31 (.A(_02955_));
 sg13g2_antennanp ANTENNA_32 (.A(_02955_));
 sg13g2_antennanp ANTENNA_33 (.A(_02955_));
 sg13g2_antennanp ANTENNA_34 (.A(_02955_));
 sg13g2_antennanp ANTENNA_35 (.A(_02955_));
 sg13g2_antennanp ANTENNA_36 (.A(_02955_));
 sg13g2_antennanp ANTENNA_37 (.A(_02955_));
 sg13g2_antennanp ANTENNA_38 (.A(_02955_));
 sg13g2_antennanp ANTENNA_39 (.A(_03053_));
 sg13g2_antennanp ANTENNA_40 (.A(_03053_));
 sg13g2_antennanp ANTENNA_41 (.A(_03053_));
 sg13g2_antennanp ANTENNA_42 (.A(_03053_));
 sg13g2_antennanp ANTENNA_43 (.A(_03478_));
 sg13g2_antennanp ANTENNA_44 (.A(_03478_));
 sg13g2_antennanp ANTENNA_45 (.A(_03478_));
 sg13g2_antennanp ANTENNA_46 (.A(_03478_));
 sg13g2_antennanp ANTENNA_47 (.A(_03478_));
 sg13g2_antennanp ANTENNA_48 (.A(_03478_));
 sg13g2_antennanp ANTENNA_49 (.A(_03478_));
 sg13g2_antennanp ANTENNA_50 (.A(_03478_));
 sg13g2_antennanp ANTENNA_51 (.A(_03478_));
 sg13g2_antennanp ANTENNA_52 (.A(_03527_));
 sg13g2_antennanp ANTENNA_53 (.A(_03527_));
 sg13g2_antennanp ANTENNA_54 (.A(_03527_));
 sg13g2_antennanp ANTENNA_55 (.A(_04734_));
 sg13g2_antennanp ANTENNA_56 (.A(_04734_));
 sg13g2_antennanp ANTENNA_57 (.A(_04734_));
 sg13g2_antennanp ANTENNA_58 (.A(_04734_));
 sg13g2_antennanp ANTENNA_59 (.A(_04751_));
 sg13g2_antennanp ANTENNA_60 (.A(_04775_));
 sg13g2_antennanp ANTENNA_61 (.A(_04778_));
 sg13g2_antennanp ANTENNA_62 (.A(_04778_));
 sg13g2_antennanp ANTENNA_63 (.A(_04778_));
 sg13g2_antennanp ANTENNA_64 (.A(_04927_));
 sg13g2_antennanp ANTENNA_65 (.A(_04985_));
 sg13g2_antennanp ANTENNA_66 (.A(_04985_));
 sg13g2_antennanp ANTENNA_67 (.A(_05003_));
 sg13g2_antennanp ANTENNA_68 (.A(_05126_));
 sg13g2_antennanp ANTENNA_69 (.A(_05149_));
 sg13g2_antennanp ANTENNA_70 (.A(_05160_));
 sg13g2_antennanp ANTENNA_71 (.A(_05174_));
 sg13g2_antennanp ANTENNA_72 (.A(_05215_));
 sg13g2_antennanp ANTENNA_73 (.A(_05309_));
 sg13g2_antennanp ANTENNA_74 (.A(_05446_));
 sg13g2_antennanp ANTENNA_75 (.A(_05583_));
 sg13g2_antennanp ANTENNA_76 (.A(_05597_));
 sg13g2_antennanp ANTENNA_77 (.A(_05653_));
 sg13g2_antennanp ANTENNA_78 (.A(_05667_));
 sg13g2_antennanp ANTENNA_79 (.A(_05669_));
 sg13g2_antennanp ANTENNA_80 (.A(_05680_));
 sg13g2_antennanp ANTENNA_81 (.A(_05700_));
 sg13g2_antennanp ANTENNA_82 (.A(_05706_));
 sg13g2_antennanp ANTENNA_83 (.A(_05712_));
 sg13g2_antennanp ANTENNA_84 (.A(_05724_));
 sg13g2_antennanp ANTENNA_85 (.A(_05895_));
 sg13g2_antennanp ANTENNA_86 (.A(_05895_));
 sg13g2_antennanp ANTENNA_87 (.A(_05895_));
 sg13g2_antennanp ANTENNA_88 (.A(_05895_));
 sg13g2_antennanp ANTENNA_89 (.A(_05895_));
 sg13g2_antennanp ANTENNA_90 (.A(_05900_));
 sg13g2_antennanp ANTENNA_91 (.A(_05900_));
 sg13g2_antennanp ANTENNA_92 (.A(_05900_));
 sg13g2_antennanp ANTENNA_93 (.A(_05900_));
 sg13g2_antennanp ANTENNA_94 (.A(_05900_));
 sg13g2_antennanp ANTENNA_95 (.A(_05900_));
 sg13g2_antennanp ANTENNA_96 (.A(_05900_));
 sg13g2_antennanp ANTENNA_97 (.A(_05955_));
 sg13g2_antennanp ANTENNA_98 (.A(_06556_));
 sg13g2_antennanp ANTENNA_99 (.A(_06556_));
 sg13g2_antennanp ANTENNA_100 (.A(_06556_));
 sg13g2_antennanp ANTENNA_101 (.A(_06556_));
 sg13g2_antennanp ANTENNA_102 (.A(_06556_));
 sg13g2_antennanp ANTENNA_103 (.A(_06556_));
 sg13g2_antennanp ANTENNA_104 (.A(_06556_));
 sg13g2_antennanp ANTENNA_105 (.A(_06556_));
 sg13g2_antennanp ANTENNA_106 (.A(_07576_));
 sg13g2_antennanp ANTENNA_107 (.A(_07576_));
 sg13g2_antennanp ANTENNA_108 (.A(_07877_));
 sg13g2_antennanp ANTENNA_109 (.A(_07877_));
 sg13g2_antennanp ANTENNA_110 (.A(_07877_));
 sg13g2_antennanp ANTENNA_111 (.A(_08204_));
 sg13g2_antennanp ANTENNA_112 (.A(_08204_));
 sg13g2_antennanp ANTENNA_113 (.A(_08328_));
 sg13g2_antennanp ANTENNA_114 (.A(_08328_));
 sg13g2_antennanp ANTENNA_115 (.A(_08408_));
 sg13g2_antennanp ANTENNA_116 (.A(_08408_));
 sg13g2_antennanp ANTENNA_117 (.A(_08408_));
 sg13g2_antennanp ANTENNA_118 (.A(_08408_));
 sg13g2_antennanp ANTENNA_119 (.A(_08439_));
 sg13g2_antennanp ANTENNA_120 (.A(_08439_));
 sg13g2_antennanp ANTENNA_121 (.A(_08439_));
 sg13g2_antennanp ANTENNA_122 (.A(_08439_));
 sg13g2_antennanp ANTENNA_123 (.A(_08439_));
 sg13g2_antennanp ANTENNA_124 (.A(_08439_));
 sg13g2_antennanp ANTENNA_125 (.A(_08444_));
 sg13g2_antennanp ANTENNA_126 (.A(_08444_));
 sg13g2_antennanp ANTENNA_127 (.A(_08444_));
 sg13g2_antennanp ANTENNA_128 (.A(_08444_));
 sg13g2_antennanp ANTENNA_129 (.A(_08444_));
 sg13g2_antennanp ANTENNA_130 (.A(_08444_));
 sg13g2_antennanp ANTENNA_131 (.A(_08444_));
 sg13g2_antennanp ANTENNA_132 (.A(_08444_));
 sg13g2_antennanp ANTENNA_133 (.A(_08444_));
 sg13g2_antennanp ANTENNA_134 (.A(_08449_));
 sg13g2_antennanp ANTENNA_135 (.A(_08449_));
 sg13g2_antennanp ANTENNA_136 (.A(_08449_));
 sg13g2_antennanp ANTENNA_137 (.A(_08449_));
 sg13g2_antennanp ANTENNA_138 (.A(_08449_));
 sg13g2_antennanp ANTENNA_139 (.A(_08449_));
 sg13g2_antennanp ANTENNA_140 (.A(_08449_));
 sg13g2_antennanp ANTENNA_141 (.A(_08449_));
 sg13g2_antennanp ANTENNA_142 (.A(_08449_));
 sg13g2_antennanp ANTENNA_143 (.A(_08449_));
 sg13g2_antennanp ANTENNA_144 (.A(_08507_));
 sg13g2_antennanp ANTENNA_145 (.A(_08507_));
 sg13g2_antennanp ANTENNA_146 (.A(_08507_));
 sg13g2_antennanp ANTENNA_147 (.A(_08680_));
 sg13g2_antennanp ANTENNA_148 (.A(_08680_));
 sg13g2_antennanp ANTENNA_149 (.A(_08680_));
 sg13g2_antennanp ANTENNA_150 (.A(_08680_));
 sg13g2_antennanp ANTENNA_151 (.A(_08680_));
 sg13g2_antennanp ANTENNA_152 (.A(_08706_));
 sg13g2_antennanp ANTENNA_153 (.A(_08706_));
 sg13g2_antennanp ANTENNA_154 (.A(_08706_));
 sg13g2_antennanp ANTENNA_155 (.A(_08706_));
 sg13g2_antennanp ANTENNA_156 (.A(_08706_));
 sg13g2_antennanp ANTENNA_157 (.A(_08706_));
 sg13g2_antennanp ANTENNA_158 (.A(_08752_));
 sg13g2_antennanp ANTENNA_159 (.A(_08752_));
 sg13g2_antennanp ANTENNA_160 (.A(_08752_));
 sg13g2_antennanp ANTENNA_161 (.A(_08776_));
 sg13g2_antennanp ANTENNA_162 (.A(_08776_));
 sg13g2_antennanp ANTENNA_163 (.A(_08776_));
 sg13g2_antennanp ANTENNA_164 (.A(_08798_));
 sg13g2_antennanp ANTENNA_165 (.A(_08798_));
 sg13g2_antennanp ANTENNA_166 (.A(_08798_));
 sg13g2_antennanp ANTENNA_167 (.A(_08818_));
 sg13g2_antennanp ANTENNA_168 (.A(_08840_));
 sg13g2_antennanp ANTENNA_169 (.A(_08840_));
 sg13g2_antennanp ANTENNA_170 (.A(_08851_));
 sg13g2_antennanp ANTENNA_171 (.A(_08851_));
 sg13g2_antennanp ANTENNA_172 (.A(_08851_));
 sg13g2_antennanp ANTENNA_173 (.A(_08851_));
 sg13g2_antennanp ANTENNA_174 (.A(_09080_));
 sg13g2_antennanp ANTENNA_175 (.A(_09080_));
 sg13g2_antennanp ANTENNA_176 (.A(_09084_));
 sg13g2_antennanp ANTENNA_177 (.A(_09084_));
 sg13g2_antennanp ANTENNA_178 (.A(_09084_));
 sg13g2_antennanp ANTENNA_179 (.A(_09084_));
 sg13g2_antennanp ANTENNA_180 (.A(_09084_));
 sg13g2_antennanp ANTENNA_181 (.A(_09084_));
 sg13g2_antennanp ANTENNA_182 (.A(_09084_));
 sg13g2_antennanp ANTENNA_183 (.A(_09084_));
 sg13g2_antennanp ANTENNA_184 (.A(_09084_));
 sg13g2_antennanp ANTENNA_185 (.A(_09131_));
 sg13g2_antennanp ANTENNA_186 (.A(_09131_));
 sg13g2_antennanp ANTENNA_187 (.A(_09131_));
 sg13g2_antennanp ANTENNA_188 (.A(_09131_));
 sg13g2_antennanp ANTENNA_189 (.A(_09140_));
 sg13g2_antennanp ANTENNA_190 (.A(_09140_));
 sg13g2_antennanp ANTENNA_191 (.A(_09140_));
 sg13g2_antennanp ANTENNA_192 (.A(_09140_));
 sg13g2_antennanp ANTENNA_193 (.A(_09140_));
 sg13g2_antennanp ANTENNA_194 (.A(_09141_));
 sg13g2_antennanp ANTENNA_195 (.A(_09141_));
 sg13g2_antennanp ANTENNA_196 (.A(_09141_));
 sg13g2_antennanp ANTENNA_197 (.A(_09141_));
 sg13g2_antennanp ANTENNA_198 (.A(_09141_));
 sg13g2_antennanp ANTENNA_199 (.A(_09149_));
 sg13g2_antennanp ANTENNA_200 (.A(_09149_));
 sg13g2_antennanp ANTENNA_201 (.A(_09149_));
 sg13g2_antennanp ANTENNA_202 (.A(_09149_));
 sg13g2_antennanp ANTENNA_203 (.A(_09149_));
 sg13g2_antennanp ANTENNA_204 (.A(_09149_));
 sg13g2_antennanp ANTENNA_205 (.A(_09150_));
 sg13g2_antennanp ANTENNA_206 (.A(_09150_));
 sg13g2_antennanp ANTENNA_207 (.A(_09150_));
 sg13g2_antennanp ANTENNA_208 (.A(_09150_));
 sg13g2_antennanp ANTENNA_209 (.A(_09151_));
 sg13g2_antennanp ANTENNA_210 (.A(_09151_));
 sg13g2_antennanp ANTENNA_211 (.A(_09151_));
 sg13g2_antennanp ANTENNA_212 (.A(_09151_));
 sg13g2_antennanp ANTENNA_213 (.A(_09162_));
 sg13g2_antennanp ANTENNA_214 (.A(_09162_));
 sg13g2_antennanp ANTENNA_215 (.A(_09162_));
 sg13g2_antennanp ANTENNA_216 (.A(_09163_));
 sg13g2_antennanp ANTENNA_217 (.A(_09163_));
 sg13g2_antennanp ANTENNA_218 (.A(_09163_));
 sg13g2_antennanp ANTENNA_219 (.A(_09230_));
 sg13g2_antennanp ANTENNA_220 (.A(_09230_));
 sg13g2_antennanp ANTENNA_221 (.A(_09230_));
 sg13g2_antennanp ANTENNA_222 (.A(_09230_));
 sg13g2_antennanp ANTENNA_223 (.A(_09230_));
 sg13g2_antennanp ANTENNA_224 (.A(_09253_));
 sg13g2_antennanp ANTENNA_225 (.A(_09253_));
 sg13g2_antennanp ANTENNA_226 (.A(_09253_));
 sg13g2_antennanp ANTENNA_227 (.A(_09253_));
 sg13g2_antennanp ANTENNA_228 (.A(_09253_));
 sg13g2_antennanp ANTENNA_229 (.A(_09253_));
 sg13g2_antennanp ANTENNA_230 (.A(_09253_));
 sg13g2_antennanp ANTENNA_231 (.A(_09253_));
 sg13g2_antennanp ANTENNA_232 (.A(_09253_));
 sg13g2_antennanp ANTENNA_233 (.A(_09253_));
 sg13g2_antennanp ANTENNA_234 (.A(_09254_));
 sg13g2_antennanp ANTENNA_235 (.A(_09254_));
 sg13g2_antennanp ANTENNA_236 (.A(_09254_));
 sg13g2_antennanp ANTENNA_237 (.A(_09254_));
 sg13g2_antennanp ANTENNA_238 (.A(_09306_));
 sg13g2_antennanp ANTENNA_239 (.A(_09395_));
 sg13g2_antennanp ANTENNA_240 (.A(_09395_));
 sg13g2_antennanp ANTENNA_241 (.A(_09395_));
 sg13g2_antennanp ANTENNA_242 (.A(_09395_));
 sg13g2_antennanp ANTENNA_243 (.A(_09395_));
 sg13g2_antennanp ANTENNA_244 (.A(_09395_));
 sg13g2_antennanp ANTENNA_245 (.A(_09395_));
 sg13g2_antennanp ANTENNA_246 (.A(_09395_));
 sg13g2_antennanp ANTENNA_247 (.A(_09395_));
 sg13g2_antennanp ANTENNA_248 (.A(_09395_));
 sg13g2_antennanp ANTENNA_249 (.A(_09395_));
 sg13g2_antennanp ANTENNA_250 (.A(_09395_));
 sg13g2_antennanp ANTENNA_251 (.A(_09395_));
 sg13g2_antennanp ANTENNA_252 (.A(_09420_));
 sg13g2_antennanp ANTENNA_253 (.A(_09420_));
 sg13g2_antennanp ANTENNA_254 (.A(_09420_));
 sg13g2_antennanp ANTENNA_255 (.A(_09420_));
 sg13g2_antennanp ANTENNA_256 (.A(_09426_));
 sg13g2_antennanp ANTENNA_257 (.A(_09426_));
 sg13g2_antennanp ANTENNA_258 (.A(_09426_));
 sg13g2_antennanp ANTENNA_259 (.A(_09426_));
 sg13g2_antennanp ANTENNA_260 (.A(_09436_));
 sg13g2_antennanp ANTENNA_261 (.A(_09437_));
 sg13g2_antennanp ANTENNA_262 (.A(_09437_));
 sg13g2_antennanp ANTENNA_263 (.A(_09445_));
 sg13g2_antennanp ANTENNA_264 (.A(_09498_));
 sg13g2_antennanp ANTENNA_265 (.A(_09499_));
 sg13g2_antennanp ANTENNA_266 (.A(_09499_));
 sg13g2_antennanp ANTENNA_267 (.A(_09505_));
 sg13g2_antennanp ANTENNA_268 (.A(_09531_));
 sg13g2_antennanp ANTENNA_269 (.A(_09587_));
 sg13g2_antennanp ANTENNA_270 (.A(_09615_));
 sg13g2_antennanp ANTENNA_271 (.A(_09660_));
 sg13g2_antennanp ANTENNA_272 (.A(_09660_));
 sg13g2_antennanp ANTENNA_273 (.A(_09660_));
 sg13g2_antennanp ANTENNA_274 (.A(_09660_));
 sg13g2_antennanp ANTENNA_275 (.A(_09907_));
 sg13g2_antennanp ANTENNA_276 (.A(_09907_));
 sg13g2_antennanp ANTENNA_277 (.A(_09907_));
 sg13g2_antennanp ANTENNA_278 (.A(_09907_));
 sg13g2_antennanp ANTENNA_279 (.A(_10042_));
 sg13g2_antennanp ANTENNA_280 (.A(_10042_));
 sg13g2_antennanp ANTENNA_281 (.A(_10042_));
 sg13g2_antennanp ANTENNA_282 (.A(_10042_));
 sg13g2_antennanp ANTENNA_283 (.A(_10042_));
 sg13g2_antennanp ANTENNA_284 (.A(_10113_));
 sg13g2_antennanp ANTENNA_285 (.A(_10113_));
 sg13g2_antennanp ANTENNA_286 (.A(_10113_));
 sg13g2_antennanp ANTENNA_287 (.A(_10113_));
 sg13g2_antennanp ANTENNA_288 (.A(_10113_));
 sg13g2_antennanp ANTENNA_289 (.A(_10113_));
 sg13g2_antennanp ANTENNA_290 (.A(_10113_));
 sg13g2_antennanp ANTENNA_291 (.A(_10113_));
 sg13g2_antennanp ANTENNA_292 (.A(_10113_));
 sg13g2_antennanp ANTENNA_293 (.A(_10113_));
 sg13g2_antennanp ANTENNA_294 (.A(_10113_));
 sg13g2_antennanp ANTENNA_295 (.A(_10113_));
 sg13g2_antennanp ANTENNA_296 (.A(_10113_));
 sg13g2_antennanp ANTENNA_297 (.A(_10113_));
 sg13g2_antennanp ANTENNA_298 (.A(_10113_));
 sg13g2_antennanp ANTENNA_299 (.A(_10113_));
 sg13g2_antennanp ANTENNA_300 (.A(_10113_));
 sg13g2_antennanp ANTENNA_301 (.A(_10113_));
 sg13g2_antennanp ANTENNA_302 (.A(_10113_));
 sg13g2_antennanp ANTENNA_303 (.A(_10113_));
 sg13g2_antennanp ANTENNA_304 (.A(_10119_));
 sg13g2_antennanp ANTENNA_305 (.A(_10119_));
 sg13g2_antennanp ANTENNA_306 (.A(_10119_));
 sg13g2_antennanp ANTENNA_307 (.A(_10119_));
 sg13g2_antennanp ANTENNA_308 (.A(_10119_));
 sg13g2_antennanp ANTENNA_309 (.A(_10119_));
 sg13g2_antennanp ANTENNA_310 (.A(_10119_));
 sg13g2_antennanp ANTENNA_311 (.A(_10119_));
 sg13g2_antennanp ANTENNA_312 (.A(_10297_));
 sg13g2_antennanp ANTENNA_313 (.A(_10297_));
 sg13g2_antennanp ANTENNA_314 (.A(_10297_));
 sg13g2_antennanp ANTENNA_315 (.A(_10297_));
 sg13g2_antennanp ANTENNA_316 (.A(_10297_));
 sg13g2_antennanp ANTENNA_317 (.A(_10297_));
 sg13g2_antennanp ANTENNA_318 (.A(_10297_));
 sg13g2_antennanp ANTENNA_319 (.A(_10297_));
 sg13g2_antennanp ANTENNA_320 (.A(_10297_));
 sg13g2_antennanp ANTENNA_321 (.A(_10297_));
 sg13g2_antennanp ANTENNA_322 (.A(_10330_));
 sg13g2_antennanp ANTENNA_323 (.A(_10330_));
 sg13g2_antennanp ANTENNA_324 (.A(_10330_));
 sg13g2_antennanp ANTENNA_325 (.A(_10330_));
 sg13g2_antennanp ANTENNA_326 (.A(_10330_));
 sg13g2_antennanp ANTENNA_327 (.A(_10330_));
 sg13g2_antennanp ANTENNA_328 (.A(_10330_));
 sg13g2_antennanp ANTENNA_329 (.A(_10330_));
 sg13g2_antennanp ANTENNA_330 (.A(_10330_));
 sg13g2_antennanp ANTENNA_331 (.A(_10368_));
 sg13g2_antennanp ANTENNA_332 (.A(_10368_));
 sg13g2_antennanp ANTENNA_333 (.A(_10368_));
 sg13g2_antennanp ANTENNA_334 (.A(_10368_));
 sg13g2_antennanp ANTENNA_335 (.A(_10368_));
 sg13g2_antennanp ANTENNA_336 (.A(_10368_));
 sg13g2_antennanp ANTENNA_337 (.A(_10368_));
 sg13g2_antennanp ANTENNA_338 (.A(_10368_));
 sg13g2_antennanp ANTENNA_339 (.A(_10368_));
 sg13g2_antennanp ANTENNA_340 (.A(_10368_));
 sg13g2_antennanp ANTENNA_341 (.A(_10368_));
 sg13g2_antennanp ANTENNA_342 (.A(_10368_));
 sg13g2_antennanp ANTENNA_343 (.A(_10368_));
 sg13g2_antennanp ANTENNA_344 (.A(_10458_));
 sg13g2_antennanp ANTENNA_345 (.A(_10458_));
 sg13g2_antennanp ANTENNA_346 (.A(_10458_));
 sg13g2_antennanp ANTENNA_347 (.A(_10458_));
 sg13g2_antennanp ANTENNA_348 (.A(_10458_));
 sg13g2_antennanp ANTENNA_349 (.A(_10458_));
 sg13g2_antennanp ANTENNA_350 (.A(_10458_));
 sg13g2_antennanp ANTENNA_351 (.A(_10458_));
 sg13g2_antennanp ANTENNA_352 (.A(_10458_));
 sg13g2_antennanp ANTENNA_353 (.A(_10458_));
 sg13g2_antennanp ANTENNA_354 (.A(_10458_));
 sg13g2_antennanp ANTENNA_355 (.A(_10629_));
 sg13g2_antennanp ANTENNA_356 (.A(_10629_));
 sg13g2_antennanp ANTENNA_357 (.A(_10629_));
 sg13g2_antennanp ANTENNA_358 (.A(_10629_));
 sg13g2_antennanp ANTENNA_359 (.A(_10629_));
 sg13g2_antennanp ANTENNA_360 (.A(_10629_));
 sg13g2_antennanp ANTENNA_361 (.A(_10634_));
 sg13g2_antennanp ANTENNA_362 (.A(_10634_));
 sg13g2_antennanp ANTENNA_363 (.A(_10634_));
 sg13g2_antennanp ANTENNA_364 (.A(_10779_));
 sg13g2_antennanp ANTENNA_365 (.A(_11031_));
 sg13g2_antennanp ANTENNA_366 (.A(_11031_));
 sg13g2_antennanp ANTENNA_367 (.A(_11031_));
 sg13g2_antennanp ANTENNA_368 (.A(_11031_));
 sg13g2_antennanp ANTENNA_369 (.A(_11031_));
 sg13g2_antennanp ANTENNA_370 (.A(_11032_));
 sg13g2_antennanp ANTENNA_371 (.A(_11032_));
 sg13g2_antennanp ANTENNA_372 (.A(_11032_));
 sg13g2_antennanp ANTENNA_373 (.A(_11032_));
 sg13g2_antennanp ANTENNA_374 (.A(_11032_));
 sg13g2_antennanp ANTENNA_375 (.A(_11032_));
 sg13g2_antennanp ANTENNA_376 (.A(_11032_));
 sg13g2_antennanp ANTENNA_377 (.A(_11032_));
 sg13g2_antennanp ANTENNA_378 (.A(_11210_));
 sg13g2_antennanp ANTENNA_379 (.A(_11776_));
 sg13g2_antennanp ANTENNA_380 (.A(_11776_));
 sg13g2_antennanp ANTENNA_381 (.A(_11776_));
 sg13g2_antennanp ANTENNA_382 (.A(_11919_));
 sg13g2_antennanp ANTENNA_383 (.A(_11919_));
 sg13g2_antennanp ANTENNA_384 (.A(_11919_));
 sg13g2_antennanp ANTENNA_385 (.A(_11919_));
 sg13g2_antennanp ANTENNA_386 (.A(_11926_));
 sg13g2_antennanp ANTENNA_387 (.A(_11926_));
 sg13g2_antennanp ANTENNA_388 (.A(_11926_));
 sg13g2_antennanp ANTENNA_389 (.A(_11926_));
 sg13g2_antennanp ANTENNA_390 (.A(_11926_));
 sg13g2_antennanp ANTENNA_391 (.A(_11926_));
 sg13g2_antennanp ANTENNA_392 (.A(_11926_));
 sg13g2_antennanp ANTENNA_393 (.A(_11926_));
 sg13g2_antennanp ANTENNA_394 (.A(_11926_));
 sg13g2_antennanp ANTENNA_395 (.A(_11941_));
 sg13g2_antennanp ANTENNA_396 (.A(_11941_));
 sg13g2_antennanp ANTENNA_397 (.A(_11941_));
 sg13g2_antennanp ANTENNA_398 (.A(_11941_));
 sg13g2_antennanp ANTENNA_399 (.A(_11941_));
 sg13g2_antennanp ANTENNA_400 (.A(_11941_));
 sg13g2_antennanp ANTENNA_401 (.A(_11941_));
 sg13g2_antennanp ANTENNA_402 (.A(_11941_));
 sg13g2_antennanp ANTENNA_403 (.A(_11941_));
 sg13g2_antennanp ANTENNA_404 (.A(_11941_));
 sg13g2_antennanp ANTENNA_405 (.A(_11941_));
 sg13g2_antennanp ANTENNA_406 (.A(_11941_));
 sg13g2_antennanp ANTENNA_407 (.A(_11941_));
 sg13g2_antennanp ANTENNA_408 (.A(_11941_));
 sg13g2_antennanp ANTENNA_409 (.A(_11941_));
 sg13g2_antennanp ANTENNA_410 (.A(_11941_));
 sg13g2_antennanp ANTENNA_411 (.A(_11941_));
 sg13g2_antennanp ANTENNA_412 (.A(_11941_));
 sg13g2_antennanp ANTENNA_413 (.A(_11960_));
 sg13g2_antennanp ANTENNA_414 (.A(_11960_));
 sg13g2_antennanp ANTENNA_415 (.A(_11960_));
 sg13g2_antennanp ANTENNA_416 (.A(_11960_));
 sg13g2_antennanp ANTENNA_417 (.A(_11960_));
 sg13g2_antennanp ANTENNA_418 (.A(_11960_));
 sg13g2_antennanp ANTENNA_419 (.A(_11960_));
 sg13g2_antennanp ANTENNA_420 (.A(_11960_));
 sg13g2_antennanp ANTENNA_421 (.A(_11960_));
 sg13g2_antennanp ANTENNA_422 (.A(_12351_));
 sg13g2_antennanp ANTENNA_423 (.A(_12351_));
 sg13g2_antennanp ANTENNA_424 (.A(_12351_));
 sg13g2_antennanp ANTENNA_425 (.A(_12351_));
 sg13g2_antennanp ANTENNA_426 (.A(_12351_));
 sg13g2_antennanp ANTENNA_427 (.A(_12648_));
 sg13g2_antennanp ANTENNA_428 (.A(_12648_));
 sg13g2_antennanp ANTENNA_429 (.A(_12648_));
 sg13g2_antennanp ANTENNA_430 (.A(clk));
 sg13g2_antennanp ANTENNA_431 (.A(clk));
 sg13g2_antennanp ANTENNA_432 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_433 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_434 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_435 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_436 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_437 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_438 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_439 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_440 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_441 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_442 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_443 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_444 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_445 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_446 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_447 (.A(uio_in[0]));
 sg13g2_antennanp ANTENNA_448 (.A(net4));
 sg13g2_antennanp ANTENNA_449 (.A(net4));
 sg13g2_antennanp ANTENNA_450 (.A(net4));
 sg13g2_antennanp ANTENNA_451 (.A(net12));
 sg13g2_antennanp ANTENNA_452 (.A(net12));
 sg13g2_antennanp ANTENNA_453 (.A(net12));
 sg13g2_antennanp ANTENNA_454 (.A(net13));
 sg13g2_antennanp ANTENNA_455 (.A(net13));
 sg13g2_antennanp ANTENNA_456 (.A(net13));
 sg13g2_antennanp ANTENNA_457 (.A(net14));
 sg13g2_antennanp ANTENNA_458 (.A(net14));
 sg13g2_antennanp ANTENNA_459 (.A(net14));
 sg13g2_antennanp ANTENNA_460 (.A(net15));
 sg13g2_antennanp ANTENNA_461 (.A(net15));
 sg13g2_antennanp ANTENNA_462 (.A(net15));
 sg13g2_antennanp ANTENNA_463 (.A(net71));
 sg13g2_antennanp ANTENNA_464 (.A(net71));
 sg13g2_antennanp ANTENNA_465 (.A(net71));
 sg13g2_antennanp ANTENNA_466 (.A(net71));
 sg13g2_antennanp ANTENNA_467 (.A(net71));
 sg13g2_antennanp ANTENNA_468 (.A(net71));
 sg13g2_antennanp ANTENNA_469 (.A(net71));
 sg13g2_antennanp ANTENNA_470 (.A(net71));
 sg13g2_antennanp ANTENNA_471 (.A(net71));
 sg13g2_antennanp ANTENNA_472 (.A(net506));
 sg13g2_antennanp ANTENNA_473 (.A(net506));
 sg13g2_antennanp ANTENNA_474 (.A(net506));
 sg13g2_antennanp ANTENNA_475 (.A(net506));
 sg13g2_antennanp ANTENNA_476 (.A(net506));
 sg13g2_antennanp ANTENNA_477 (.A(net506));
 sg13g2_antennanp ANTENNA_478 (.A(net506));
 sg13g2_antennanp ANTENNA_479 (.A(net506));
 sg13g2_antennanp ANTENNA_480 (.A(net506));
 sg13g2_antennanp ANTENNA_481 (.A(net506));
 sg13g2_antennanp ANTENNA_482 (.A(net507));
 sg13g2_antennanp ANTENNA_483 (.A(net507));
 sg13g2_antennanp ANTENNA_484 (.A(net507));
 sg13g2_antennanp ANTENNA_485 (.A(net507));
 sg13g2_antennanp ANTENNA_486 (.A(net507));
 sg13g2_antennanp ANTENNA_487 (.A(net507));
 sg13g2_antennanp ANTENNA_488 (.A(net507));
 sg13g2_antennanp ANTENNA_489 (.A(net507));
 sg13g2_antennanp ANTENNA_490 (.A(net507));
 sg13g2_antennanp ANTENNA_491 (.A(net507));
 sg13g2_antennanp ANTENNA_492 (.A(net507));
 sg13g2_antennanp ANTENNA_493 (.A(net507));
 sg13g2_antennanp ANTENNA_494 (.A(net507));
 sg13g2_antennanp ANTENNA_495 (.A(net507));
 sg13g2_antennanp ANTENNA_496 (.A(net507));
 sg13g2_antennanp ANTENNA_497 (.A(net599));
 sg13g2_antennanp ANTENNA_498 (.A(net599));
 sg13g2_antennanp ANTENNA_499 (.A(net599));
 sg13g2_antennanp ANTENNA_500 (.A(net599));
 sg13g2_antennanp ANTENNA_501 (.A(net599));
 sg13g2_antennanp ANTENNA_502 (.A(net599));
 sg13g2_antennanp ANTENNA_503 (.A(net599));
 sg13g2_antennanp ANTENNA_504 (.A(net599));
 sg13g2_antennanp ANTENNA_505 (.A(net601));
 sg13g2_antennanp ANTENNA_506 (.A(net601));
 sg13g2_antennanp ANTENNA_507 (.A(net601));
 sg13g2_antennanp ANTENNA_508 (.A(net601));
 sg13g2_antennanp ANTENNA_509 (.A(net601));
 sg13g2_antennanp ANTENNA_510 (.A(net601));
 sg13g2_antennanp ANTENNA_511 (.A(net601));
 sg13g2_antennanp ANTENNA_512 (.A(net601));
 sg13g2_antennanp ANTENNA_513 (.A(net601));
 sg13g2_antennanp ANTENNA_514 (.A(net601));
 sg13g2_antennanp ANTENNA_515 (.A(net601));
 sg13g2_antennanp ANTENNA_516 (.A(net601));
 sg13g2_antennanp ANTENNA_517 (.A(net601));
 sg13g2_antennanp ANTENNA_518 (.A(net601));
 sg13g2_antennanp ANTENNA_519 (.A(net601));
 sg13g2_antennanp ANTENNA_520 (.A(net601));
 sg13g2_antennanp ANTENNA_521 (.A(net601));
 sg13g2_antennanp ANTENNA_522 (.A(net601));
 sg13g2_antennanp ANTENNA_523 (.A(net601));
 sg13g2_antennanp ANTENNA_524 (.A(net601));
 sg13g2_antennanp ANTENNA_525 (.A(net601));
 sg13g2_antennanp ANTENNA_526 (.A(net613));
 sg13g2_antennanp ANTENNA_527 (.A(net613));
 sg13g2_antennanp ANTENNA_528 (.A(net613));
 sg13g2_antennanp ANTENNA_529 (.A(net613));
 sg13g2_antennanp ANTENNA_530 (.A(net613));
 sg13g2_antennanp ANTENNA_531 (.A(net613));
 sg13g2_antennanp ANTENNA_532 (.A(net613));
 sg13g2_antennanp ANTENNA_533 (.A(net613));
 sg13g2_antennanp ANTENNA_534 (.A(net613));
 sg13g2_antennanp ANTENNA_535 (.A(net613));
 sg13g2_antennanp ANTENNA_536 (.A(net613));
 sg13g2_antennanp ANTENNA_537 (.A(net613));
 sg13g2_antennanp ANTENNA_538 (.A(net669));
 sg13g2_antennanp ANTENNA_539 (.A(net669));
 sg13g2_antennanp ANTENNA_540 (.A(net669));
 sg13g2_antennanp ANTENNA_541 (.A(net669));
 sg13g2_antennanp ANTENNA_542 (.A(net669));
 sg13g2_antennanp ANTENNA_543 (.A(net669));
 sg13g2_antennanp ANTENNA_544 (.A(net669));
 sg13g2_antennanp ANTENNA_545 (.A(net669));
 sg13g2_antennanp ANTENNA_546 (.A(net669));
 sg13g2_antennanp ANTENNA_547 (.A(net669));
 sg13g2_antennanp ANTENNA_548 (.A(net669));
 sg13g2_antennanp ANTENNA_549 (.A(net669));
 sg13g2_antennanp ANTENNA_550 (.A(net669));
 sg13g2_antennanp ANTENNA_551 (.A(net669));
 sg13g2_antennanp ANTENNA_552 (.A(net669));
 sg13g2_antennanp ANTENNA_553 (.A(net682));
 sg13g2_antennanp ANTENNA_554 (.A(net682));
 sg13g2_antennanp ANTENNA_555 (.A(net682));
 sg13g2_antennanp ANTENNA_556 (.A(net682));
 sg13g2_antennanp ANTENNA_557 (.A(net682));
 sg13g2_antennanp ANTENNA_558 (.A(net682));
 sg13g2_antennanp ANTENNA_559 (.A(net682));
 sg13g2_antennanp ANTENNA_560 (.A(net682));
 sg13g2_antennanp ANTENNA_561 (.A(net682));
 sg13g2_antennanp ANTENNA_562 (.A(net682));
 sg13g2_antennanp ANTENNA_563 (.A(net682));
 sg13g2_antennanp ANTENNA_564 (.A(net696));
 sg13g2_antennanp ANTENNA_565 (.A(net696));
 sg13g2_antennanp ANTENNA_566 (.A(net696));
 sg13g2_antennanp ANTENNA_567 (.A(net696));
 sg13g2_antennanp ANTENNA_568 (.A(net696));
 sg13g2_antennanp ANTENNA_569 (.A(net696));
 sg13g2_antennanp ANTENNA_570 (.A(net696));
 sg13g2_antennanp ANTENNA_571 (.A(net696));
 sg13g2_antennanp ANTENNA_572 (.A(net696));
 sg13g2_antennanp ANTENNA_573 (.A(net696));
 sg13g2_antennanp ANTENNA_574 (.A(net696));
 sg13g2_antennanp ANTENNA_575 (.A(net696));
 sg13g2_antennanp ANTENNA_576 (.A(net696));
 sg13g2_antennanp ANTENNA_577 (.A(net696));
 sg13g2_antennanp ANTENNA_578 (.A(net696));
 sg13g2_antennanp ANTENNA_579 (.A(net717));
 sg13g2_antennanp ANTENNA_580 (.A(net717));
 sg13g2_antennanp ANTENNA_581 (.A(net717));
 sg13g2_antennanp ANTENNA_582 (.A(net717));
 sg13g2_antennanp ANTENNA_583 (.A(net717));
 sg13g2_antennanp ANTENNA_584 (.A(net717));
 sg13g2_antennanp ANTENNA_585 (.A(net717));
 sg13g2_antennanp ANTENNA_586 (.A(net717));
 sg13g2_antennanp ANTENNA_587 (.A(net717));
 sg13g2_antennanp ANTENNA_588 (.A(net717));
 sg13g2_antennanp ANTENNA_589 (.A(net717));
 sg13g2_antennanp ANTENNA_590 (.A(net717));
 sg13g2_antennanp ANTENNA_591 (.A(net717));
 sg13g2_antennanp ANTENNA_592 (.A(net717));
 sg13g2_antennanp ANTENNA_593 (.A(net717));
 sg13g2_antennanp ANTENNA_594 (.A(net717));
 sg13g2_antennanp ANTENNA_595 (.A(net717));
 sg13g2_antennanp ANTENNA_596 (.A(net717));
 sg13g2_antennanp ANTENNA_597 (.A(net717));
 sg13g2_antennanp ANTENNA_598 (.A(net717));
 sg13g2_antennanp ANTENNA_599 (.A(net717));
 sg13g2_antennanp ANTENNA_600 (.A(net717));
 sg13g2_antennanp ANTENNA_601 (.A(net717));
 sg13g2_antennanp ANTENNA_602 (.A(net796));
 sg13g2_antennanp ANTENNA_603 (.A(net796));
 sg13g2_antennanp ANTENNA_604 (.A(net796));
 sg13g2_antennanp ANTENNA_605 (.A(net796));
 sg13g2_antennanp ANTENNA_606 (.A(net796));
 sg13g2_antennanp ANTENNA_607 (.A(net796));
 sg13g2_antennanp ANTENNA_608 (.A(net796));
 sg13g2_antennanp ANTENNA_609 (.A(net796));
 sg13g2_antennanp ANTENNA_610 (.A(net796));
 sg13g2_antennanp ANTENNA_611 (.A(net796));
 sg13g2_antennanp ANTENNA_612 (.A(net796));
 sg13g2_antennanp ANTENNA_613 (.A(net796));
 sg13g2_antennanp ANTENNA_614 (.A(net796));
 sg13g2_antennanp ANTENNA_615 (.A(net802));
 sg13g2_antennanp ANTENNA_616 (.A(net802));
 sg13g2_antennanp ANTENNA_617 (.A(net802));
 sg13g2_antennanp ANTENNA_618 (.A(net802));
 sg13g2_antennanp ANTENNA_619 (.A(net802));
 sg13g2_antennanp ANTENNA_620 (.A(net802));
 sg13g2_antennanp ANTENNA_621 (.A(net802));
 sg13g2_antennanp ANTENNA_622 (.A(net802));
 sg13g2_antennanp ANTENNA_623 (.A(net802));
 sg13g2_antennanp ANTENNA_624 (.A(net802));
 sg13g2_antennanp ANTENNA_625 (.A(net802));
 sg13g2_antennanp ANTENNA_626 (.A(net802));
 sg13g2_antennanp ANTENNA_627 (.A(net802));
 sg13g2_antennanp ANTENNA_628 (.A(net802));
 sg13g2_antennanp ANTENNA_629 (.A(net802));
 sg13g2_antennanp ANTENNA_630 (.A(net802));
 sg13g2_antennanp ANTENNA_631 (.A(net849));
 sg13g2_antennanp ANTENNA_632 (.A(net849));
 sg13g2_antennanp ANTENNA_633 (.A(net849));
 sg13g2_antennanp ANTENNA_634 (.A(net849));
 sg13g2_antennanp ANTENNA_635 (.A(net849));
 sg13g2_antennanp ANTENNA_636 (.A(net849));
 sg13g2_antennanp ANTENNA_637 (.A(net849));
 sg13g2_antennanp ANTENNA_638 (.A(net849));
 sg13g2_antennanp ANTENNA_639 (.A(net849));
 sg13g2_antennanp ANTENNA_640 (.A(net849));
 sg13g2_antennanp ANTENNA_641 (.A(net849));
 sg13g2_antennanp ANTENNA_642 (.A(net849));
 sg13g2_antennanp ANTENNA_643 (.A(net849));
 sg13g2_antennanp ANTENNA_644 (.A(net849));
 sg13g2_antennanp ANTENNA_645 (.A(net849));
 sg13g2_antennanp ANTENNA_646 (.A(net849));
 sg13g2_antennanp ANTENNA_647 (.A(net849));
 sg13g2_antennanp ANTENNA_648 (.A(net849));
 sg13g2_antennanp ANTENNA_649 (.A(net850));
 sg13g2_antennanp ANTENNA_650 (.A(net850));
 sg13g2_antennanp ANTENNA_651 (.A(net850));
 sg13g2_antennanp ANTENNA_652 (.A(net850));
 sg13g2_antennanp ANTENNA_653 (.A(net850));
 sg13g2_antennanp ANTENNA_654 (.A(net850));
 sg13g2_antennanp ANTENNA_655 (.A(net850));
 sg13g2_antennanp ANTENNA_656 (.A(net850));
 sg13g2_antennanp ANTENNA_657 (.A(net850));
 sg13g2_antennanp ANTENNA_658 (.A(net904));
 sg13g2_antennanp ANTENNA_659 (.A(net904));
 sg13g2_antennanp ANTENNA_660 (.A(net904));
 sg13g2_antennanp ANTENNA_661 (.A(net904));
 sg13g2_antennanp ANTENNA_662 (.A(net904));
 sg13g2_antennanp ANTENNA_663 (.A(net904));
 sg13g2_antennanp ANTENNA_664 (.A(net904));
 sg13g2_antennanp ANTENNA_665 (.A(net904));
 sg13g2_antennanp ANTENNA_666 (.A(net904));
 sg13g2_antennanp ANTENNA_667 (.A(net904));
 sg13g2_antennanp ANTENNA_668 (.A(net904));
 sg13g2_antennanp ANTENNA_669 (.A(net904));
 sg13g2_antennanp ANTENNA_670 (.A(net904));
 sg13g2_antennanp ANTENNA_671 (.A(net904));
 sg13g2_antennanp ANTENNA_672 (.A(net904));
 sg13g2_antennanp ANTENNA_673 (.A(net904));
 sg13g2_antennanp ANTENNA_674 (.A(net904));
 sg13g2_antennanp ANTENNA_675 (.A(net904));
 sg13g2_antennanp ANTENNA_676 (.A(net974));
 sg13g2_antennanp ANTENNA_677 (.A(net974));
 sg13g2_antennanp ANTENNA_678 (.A(net974));
 sg13g2_antennanp ANTENNA_679 (.A(net974));
 sg13g2_antennanp ANTENNA_680 (.A(net974));
 sg13g2_antennanp ANTENNA_681 (.A(net974));
 sg13g2_antennanp ANTENNA_682 (.A(net974));
 sg13g2_antennanp ANTENNA_683 (.A(net974));
 sg13g2_antennanp ANTENNA_684 (.A(net974));
 sg13g2_antennanp ANTENNA_685 (.A(net977));
 sg13g2_antennanp ANTENNA_686 (.A(net977));
 sg13g2_antennanp ANTENNA_687 (.A(net977));
 sg13g2_antennanp ANTENNA_688 (.A(net977));
 sg13g2_antennanp ANTENNA_689 (.A(net977));
 sg13g2_antennanp ANTENNA_690 (.A(net977));
 sg13g2_antennanp ANTENNA_691 (.A(net977));
 sg13g2_antennanp ANTENNA_692 (.A(net977));
 sg13g2_antennanp ANTENNA_693 (.A(net977));
 sg13g2_antennanp ANTENNA_694 (.A(net977));
 sg13g2_antennanp ANTENNA_695 (.A(net977));
 sg13g2_antennanp ANTENNA_696 (.A(net977));
 sg13g2_antennanp ANTENNA_697 (.A(net977));
 sg13g2_antennanp ANTENNA_698 (.A(net977));
 sg13g2_antennanp ANTENNA_699 (.A(net977));
 sg13g2_antennanp ANTENNA_700 (.A(net977));
 sg13g2_antennanp ANTENNA_701 (.A(net977));
 sg13g2_antennanp ANTENNA_702 (.A(net977));
 sg13g2_antennanp ANTENNA_703 (.A(net977));
 sg13g2_antennanp ANTENNA_704 (.A(net977));
 sg13g2_antennanp ANTENNA_705 (.A(net977));
 sg13g2_antennanp ANTENNA_706 (.A(net977));
 sg13g2_antennanp ANTENNA_707 (.A(net977));
 sg13g2_antennanp ANTENNA_708 (.A(net1008));
 sg13g2_antennanp ANTENNA_709 (.A(net1008));
 sg13g2_antennanp ANTENNA_710 (.A(net1008));
 sg13g2_antennanp ANTENNA_711 (.A(net1008));
 sg13g2_antennanp ANTENNA_712 (.A(net1008));
 sg13g2_antennanp ANTENNA_713 (.A(net1008));
 sg13g2_antennanp ANTENNA_714 (.A(net1008));
 sg13g2_antennanp ANTENNA_715 (.A(net1008));
 sg13g2_antennanp ANTENNA_716 (.A(net1008));
 sg13g2_antennanp ANTENNA_717 (.A(net1008));
 sg13g2_antennanp ANTENNA_718 (.A(net1008));
 sg13g2_antennanp ANTENNA_719 (.A(net1008));
 sg13g2_antennanp ANTENNA_720 (.A(net1008));
 sg13g2_antennanp ANTENNA_721 (.A(net1008));
 sg13g2_antennanp ANTENNA_722 (.A(net1008));
 sg13g2_antennanp ANTENNA_723 (.A(net1008));
 sg13g2_antennanp ANTENNA_724 (.A(net1008));
 sg13g2_antennanp ANTENNA_725 (.A(net1008));
 sg13g2_antennanp ANTENNA_726 (.A(net1008));
 sg13g2_antennanp ANTENNA_727 (.A(net1008));
 sg13g2_antennanp ANTENNA_728 (.A(net1008));
 sg13g2_antennanp ANTENNA_729 (.A(net1008));
 sg13g2_antennanp ANTENNA_730 (.A(net1008));
 sg13g2_antennanp ANTENNA_731 (.A(net1008));
 sg13g2_antennanp ANTENNA_732 (.A(net1008));
 sg13g2_antennanp ANTENNA_733 (.A(net1008));
 sg13g2_antennanp ANTENNA_734 (.A(net1008));
 sg13g2_antennanp ANTENNA_735 (.A(net1008));
 sg13g2_antennanp ANTENNA_736 (.A(net1008));
 sg13g2_antennanp ANTENNA_737 (.A(net1008));
 sg13g2_antennanp ANTENNA_738 (.A(net1008));
 sg13g2_antennanp ANTENNA_739 (.A(net1008));
 sg13g2_antennanp ANTENNA_740 (.A(net1008));
 sg13g2_antennanp ANTENNA_741 (.A(net1008));
 sg13g2_antennanp ANTENNA_742 (.A(net1008));
 sg13g2_antennanp ANTENNA_743 (.A(net1008));
 sg13g2_antennanp ANTENNA_744 (.A(net1010));
 sg13g2_antennanp ANTENNA_745 (.A(net1010));
 sg13g2_antennanp ANTENNA_746 (.A(net1010));
 sg13g2_antennanp ANTENNA_747 (.A(net1010));
 sg13g2_antennanp ANTENNA_748 (.A(net1010));
 sg13g2_antennanp ANTENNA_749 (.A(net1010));
 sg13g2_antennanp ANTENNA_750 (.A(net1010));
 sg13g2_antennanp ANTENNA_751 (.A(net1010));
 sg13g2_antennanp ANTENNA_752 (.A(net1012));
 sg13g2_antennanp ANTENNA_753 (.A(net1012));
 sg13g2_antennanp ANTENNA_754 (.A(net1012));
 sg13g2_antennanp ANTENNA_755 (.A(net1012));
 sg13g2_antennanp ANTENNA_756 (.A(net1012));
 sg13g2_antennanp ANTENNA_757 (.A(net1012));
 sg13g2_antennanp ANTENNA_758 (.A(net1012));
 sg13g2_antennanp ANTENNA_759 (.A(net1012));
 sg13g2_antennanp ANTENNA_760 (.A(net1012));
 sg13g2_antennanp ANTENNA_761 (.A(net1015));
 sg13g2_antennanp ANTENNA_762 (.A(net1015));
 sg13g2_antennanp ANTENNA_763 (.A(net1015));
 sg13g2_antennanp ANTENNA_764 (.A(net1015));
 sg13g2_antennanp ANTENNA_765 (.A(net1015));
 sg13g2_antennanp ANTENNA_766 (.A(net1015));
 sg13g2_antennanp ANTENNA_767 (.A(net1015));
 sg13g2_antennanp ANTENNA_768 (.A(net1015));
 sg13g2_antennanp ANTENNA_769 (.A(net1015));
 sg13g2_antennanp ANTENNA_770 (.A(net1015));
 sg13g2_antennanp ANTENNA_771 (.A(net1015));
 sg13g2_antennanp ANTENNA_772 (.A(net1015));
 sg13g2_antennanp ANTENNA_773 (.A(net1015));
 sg13g2_antennanp ANTENNA_774 (.A(net1015));
 sg13g2_antennanp ANTENNA_775 (.A(net1015));
 sg13g2_antennanp ANTENNA_776 (.A(net1015));
 sg13g2_antennanp ANTENNA_777 (.A(net1053));
 sg13g2_antennanp ANTENNA_778 (.A(net1053));
 sg13g2_antennanp ANTENNA_779 (.A(net1053));
 sg13g2_antennanp ANTENNA_780 (.A(net1053));
 sg13g2_antennanp ANTENNA_781 (.A(net1053));
 sg13g2_antennanp ANTENNA_782 (.A(net1053));
 sg13g2_antennanp ANTENNA_783 (.A(net1053));
 sg13g2_antennanp ANTENNA_784 (.A(net1053));
 sg13g2_antennanp ANTENNA_785 (.A(net1058));
 sg13g2_antennanp ANTENNA_786 (.A(net1058));
 sg13g2_antennanp ANTENNA_787 (.A(net1058));
 sg13g2_antennanp ANTENNA_788 (.A(net1058));
 sg13g2_antennanp ANTENNA_789 (.A(net1058));
 sg13g2_antennanp ANTENNA_790 (.A(net1058));
 sg13g2_antennanp ANTENNA_791 (.A(net1058));
 sg13g2_antennanp ANTENNA_792 (.A(net1058));
 sg13g2_antennanp ANTENNA_793 (.A(net1058));
 sg13g2_antennanp ANTENNA_794 (.A(net1058));
 sg13g2_antennanp ANTENNA_795 (.A(net1058));
 sg13g2_antennanp ANTENNA_796 (.A(net1058));
 sg13g2_antennanp ANTENNA_797 (.A(net1058));
 sg13g2_antennanp ANTENNA_798 (.A(net1058));
 sg13g2_antennanp ANTENNA_799 (.A(net1058));
 sg13g2_antennanp ANTENNA_800 (.A(net1058));
 sg13g2_antennanp ANTENNA_801 (.A(net1058));
 sg13g2_antennanp ANTENNA_802 (.A(net1058));
 sg13g2_antennanp ANTENNA_803 (.A(net1058));
 sg13g2_antennanp ANTENNA_804 (.A(net1058));
 sg13g2_antennanp ANTENNA_805 (.A(net1094));
 sg13g2_antennanp ANTENNA_806 (.A(net1094));
 sg13g2_antennanp ANTENNA_807 (.A(net1094));
 sg13g2_antennanp ANTENNA_808 (.A(net1094));
 sg13g2_antennanp ANTENNA_809 (.A(net1094));
 sg13g2_antennanp ANTENNA_810 (.A(net1094));
 sg13g2_antennanp ANTENNA_811 (.A(net1094));
 sg13g2_antennanp ANTENNA_812 (.A(net1094));
 sg13g2_antennanp ANTENNA_813 (.A(net1094));
 sg13g2_antennanp ANTENNA_814 (.A(_00203_));
 sg13g2_antennanp ANTENNA_815 (.A(_00203_));
 sg13g2_antennanp ANTENNA_816 (.A(_00209_));
 sg13g2_antennanp ANTENNA_817 (.A(_00784_));
 sg13g2_antennanp ANTENNA_818 (.A(_00784_));
 sg13g2_antennanp ANTENNA_819 (.A(_00923_));
 sg13g2_antennanp ANTENNA_820 (.A(_01032_));
 sg13g2_antennanp ANTENNA_821 (.A(_01034_));
 sg13g2_antennanp ANTENNA_822 (.A(_01034_));
 sg13g2_antennanp ANTENNA_823 (.A(_02779_));
 sg13g2_antennanp ANTENNA_824 (.A(_02779_));
 sg13g2_antennanp ANTENNA_825 (.A(_02779_));
 sg13g2_antennanp ANTENNA_826 (.A(_02779_));
 sg13g2_antennanp ANTENNA_827 (.A(_02910_));
 sg13g2_antennanp ANTENNA_828 (.A(_02910_));
 sg13g2_antennanp ANTENNA_829 (.A(_02910_));
 sg13g2_antennanp ANTENNA_830 (.A(_02910_));
 sg13g2_antennanp ANTENNA_831 (.A(_02910_));
 sg13g2_antennanp ANTENNA_832 (.A(_02910_));
 sg13g2_antennanp ANTENNA_833 (.A(_02910_));
 sg13g2_antennanp ANTENNA_834 (.A(_02910_));
 sg13g2_antennanp ANTENNA_835 (.A(_02910_));
 sg13g2_antennanp ANTENNA_836 (.A(_02955_));
 sg13g2_antennanp ANTENNA_837 (.A(_02955_));
 sg13g2_antennanp ANTENNA_838 (.A(_02955_));
 sg13g2_antennanp ANTENNA_839 (.A(_02955_));
 sg13g2_antennanp ANTENNA_840 (.A(_02955_));
 sg13g2_antennanp ANTENNA_841 (.A(_02955_));
 sg13g2_antennanp ANTENNA_842 (.A(_02955_));
 sg13g2_antennanp ANTENNA_843 (.A(_02955_));
 sg13g2_antennanp ANTENNA_844 (.A(_02955_));
 sg13g2_antennanp ANTENNA_845 (.A(_02955_));
 sg13g2_antennanp ANTENNA_846 (.A(_02955_));
 sg13g2_antennanp ANTENNA_847 (.A(_02955_));
 sg13g2_antennanp ANTENNA_848 (.A(_02955_));
 sg13g2_antennanp ANTENNA_849 (.A(_02955_));
 sg13g2_antennanp ANTENNA_850 (.A(_03053_));
 sg13g2_antennanp ANTENNA_851 (.A(_03053_));
 sg13g2_antennanp ANTENNA_852 (.A(_03053_));
 sg13g2_antennanp ANTENNA_853 (.A(_03053_));
 sg13g2_antennanp ANTENNA_854 (.A(_03478_));
 sg13g2_antennanp ANTENNA_855 (.A(_03478_));
 sg13g2_antennanp ANTENNA_856 (.A(_03478_));
 sg13g2_antennanp ANTENNA_857 (.A(_03478_));
 sg13g2_antennanp ANTENNA_858 (.A(_03527_));
 sg13g2_antennanp ANTENNA_859 (.A(_03527_));
 sg13g2_antennanp ANTENNA_860 (.A(_03527_));
 sg13g2_antennanp ANTENNA_861 (.A(_04734_));
 sg13g2_antennanp ANTENNA_862 (.A(_04734_));
 sg13g2_antennanp ANTENNA_863 (.A(_04734_));
 sg13g2_antennanp ANTENNA_864 (.A(_04734_));
 sg13g2_antennanp ANTENNA_865 (.A(_04751_));
 sg13g2_antennanp ANTENNA_866 (.A(_04775_));
 sg13g2_antennanp ANTENNA_867 (.A(_04778_));
 sg13g2_antennanp ANTENNA_868 (.A(_04778_));
 sg13g2_antennanp ANTENNA_869 (.A(_04778_));
 sg13g2_antennanp ANTENNA_870 (.A(_04927_));
 sg13g2_antennanp ANTENNA_871 (.A(_04985_));
 sg13g2_antennanp ANTENNA_872 (.A(_04985_));
 sg13g2_antennanp ANTENNA_873 (.A(_05003_));
 sg13g2_antennanp ANTENNA_874 (.A(_05090_));
 sg13g2_antennanp ANTENNA_875 (.A(_05090_));
 sg13g2_antennanp ANTENNA_876 (.A(_05090_));
 sg13g2_antennanp ANTENNA_877 (.A(_05126_));
 sg13g2_antennanp ANTENNA_878 (.A(_05149_));
 sg13g2_antennanp ANTENNA_879 (.A(_05160_));
 sg13g2_antennanp ANTENNA_880 (.A(_05174_));
 sg13g2_antennanp ANTENNA_881 (.A(_05201_));
 sg13g2_antennanp ANTENNA_882 (.A(_05215_));
 sg13g2_antennanp ANTENNA_883 (.A(_05309_));
 sg13g2_antennanp ANTENNA_884 (.A(_05583_));
 sg13g2_antennanp ANTENNA_885 (.A(_05653_));
 sg13g2_antennanp ANTENNA_886 (.A(_05667_));
 sg13g2_antennanp ANTENNA_887 (.A(_05669_));
 sg13g2_antennanp ANTENNA_888 (.A(_05680_));
 sg13g2_antennanp ANTENNA_889 (.A(_05700_));
 sg13g2_antennanp ANTENNA_890 (.A(_05700_));
 sg13g2_antennanp ANTENNA_891 (.A(_05706_));
 sg13g2_antennanp ANTENNA_892 (.A(_05706_));
 sg13g2_antennanp ANTENNA_893 (.A(_05712_));
 sg13g2_antennanp ANTENNA_894 (.A(_05724_));
 sg13g2_antennanp ANTENNA_895 (.A(_05724_));
 sg13g2_antennanp ANTENNA_896 (.A(_05895_));
 sg13g2_antennanp ANTENNA_897 (.A(_05895_));
 sg13g2_antennanp ANTENNA_898 (.A(_05895_));
 sg13g2_antennanp ANTENNA_899 (.A(_05895_));
 sg13g2_antennanp ANTENNA_900 (.A(_05895_));
 sg13g2_antennanp ANTENNA_901 (.A(_05900_));
 sg13g2_antennanp ANTENNA_902 (.A(_05900_));
 sg13g2_antennanp ANTENNA_903 (.A(_05900_));
 sg13g2_antennanp ANTENNA_904 (.A(_05900_));
 sg13g2_antennanp ANTENNA_905 (.A(_05900_));
 sg13g2_antennanp ANTENNA_906 (.A(_05900_));
 sg13g2_antennanp ANTENNA_907 (.A(_05900_));
 sg13g2_antennanp ANTENNA_908 (.A(_05955_));
 sg13g2_antennanp ANTENNA_909 (.A(_06556_));
 sg13g2_antennanp ANTENNA_910 (.A(_06556_));
 sg13g2_antennanp ANTENNA_911 (.A(_06556_));
 sg13g2_antennanp ANTENNA_912 (.A(_06556_));
 sg13g2_antennanp ANTENNA_913 (.A(_06556_));
 sg13g2_antennanp ANTENNA_914 (.A(_06556_));
 sg13g2_antennanp ANTENNA_915 (.A(_07576_));
 sg13g2_antennanp ANTENNA_916 (.A(_07576_));
 sg13g2_antennanp ANTENNA_917 (.A(_07877_));
 sg13g2_antennanp ANTENNA_918 (.A(_07877_));
 sg13g2_antennanp ANTENNA_919 (.A(_07877_));
 sg13g2_antennanp ANTENNA_920 (.A(_08204_));
 sg13g2_antennanp ANTENNA_921 (.A(_08204_));
 sg13g2_antennanp ANTENNA_922 (.A(_08299_));
 sg13g2_antennanp ANTENNA_923 (.A(_08299_));
 sg13g2_antennanp ANTENNA_924 (.A(_08299_));
 sg13g2_antennanp ANTENNA_925 (.A(_08327_));
 sg13g2_antennanp ANTENNA_926 (.A(_08327_));
 sg13g2_antennanp ANTENNA_927 (.A(_08327_));
 sg13g2_antennanp ANTENNA_928 (.A(_08328_));
 sg13g2_antennanp ANTENNA_929 (.A(_08328_));
 sg13g2_antennanp ANTENNA_930 (.A(_08328_));
 sg13g2_antennanp ANTENNA_931 (.A(_08408_));
 sg13g2_antennanp ANTENNA_932 (.A(_08408_));
 sg13g2_antennanp ANTENNA_933 (.A(_08408_));
 sg13g2_antennanp ANTENNA_934 (.A(_08408_));
 sg13g2_antennanp ANTENNA_935 (.A(_08408_));
 sg13g2_antennanp ANTENNA_936 (.A(_08439_));
 sg13g2_antennanp ANTENNA_937 (.A(_08439_));
 sg13g2_antennanp ANTENNA_938 (.A(_08439_));
 sg13g2_antennanp ANTENNA_939 (.A(_08439_));
 sg13g2_antennanp ANTENNA_940 (.A(_08439_));
 sg13g2_antennanp ANTENNA_941 (.A(_08439_));
 sg13g2_antennanp ANTENNA_942 (.A(_08507_));
 sg13g2_antennanp ANTENNA_943 (.A(_08507_));
 sg13g2_antennanp ANTENNA_944 (.A(_08507_));
 sg13g2_antennanp ANTENNA_945 (.A(_08507_));
 sg13g2_antennanp ANTENNA_946 (.A(_08507_));
 sg13g2_antennanp ANTENNA_947 (.A(_08507_));
 sg13g2_antennanp ANTENNA_948 (.A(_08680_));
 sg13g2_antennanp ANTENNA_949 (.A(_08680_));
 sg13g2_antennanp ANTENNA_950 (.A(_08680_));
 sg13g2_antennanp ANTENNA_951 (.A(_08680_));
 sg13g2_antennanp ANTENNA_952 (.A(_08680_));
 sg13g2_antennanp ANTENNA_953 (.A(_08706_));
 sg13g2_antennanp ANTENNA_954 (.A(_08706_));
 sg13g2_antennanp ANTENNA_955 (.A(_08706_));
 sg13g2_antennanp ANTENNA_956 (.A(_08706_));
 sg13g2_antennanp ANTENNA_957 (.A(_08706_));
 sg13g2_antennanp ANTENNA_958 (.A(_08706_));
 sg13g2_antennanp ANTENNA_959 (.A(_08706_));
 sg13g2_antennanp ANTENNA_960 (.A(_08706_));
 sg13g2_antennanp ANTENNA_961 (.A(_08706_));
 sg13g2_antennanp ANTENNA_962 (.A(_08752_));
 sg13g2_antennanp ANTENNA_963 (.A(_08752_));
 sg13g2_antennanp ANTENNA_964 (.A(_08752_));
 sg13g2_antennanp ANTENNA_965 (.A(_08776_));
 sg13g2_antennanp ANTENNA_966 (.A(_08776_));
 sg13g2_antennanp ANTENNA_967 (.A(_08776_));
 sg13g2_antennanp ANTENNA_968 (.A(_08798_));
 sg13g2_antennanp ANTENNA_969 (.A(_08798_));
 sg13g2_antennanp ANTENNA_970 (.A(_08798_));
 sg13g2_antennanp ANTENNA_971 (.A(_08818_));
 sg13g2_antennanp ANTENNA_972 (.A(_08840_));
 sg13g2_antennanp ANTENNA_973 (.A(_08851_));
 sg13g2_antennanp ANTENNA_974 (.A(_08851_));
 sg13g2_antennanp ANTENNA_975 (.A(_08851_));
 sg13g2_antennanp ANTENNA_976 (.A(_08851_));
 sg13g2_antennanp ANTENNA_977 (.A(_08851_));
 sg13g2_antennanp ANTENNA_978 (.A(_08851_));
 sg13g2_antennanp ANTENNA_979 (.A(_09084_));
 sg13g2_antennanp ANTENNA_980 (.A(_09084_));
 sg13g2_antennanp ANTENNA_981 (.A(_09084_));
 sg13g2_antennanp ANTENNA_982 (.A(_09131_));
 sg13g2_antennanp ANTENNA_983 (.A(_09131_));
 sg13g2_antennanp ANTENNA_984 (.A(_09131_));
 sg13g2_antennanp ANTENNA_985 (.A(_09131_));
 sg13g2_antennanp ANTENNA_986 (.A(_09141_));
 sg13g2_antennanp ANTENNA_987 (.A(_09141_));
 sg13g2_antennanp ANTENNA_988 (.A(_09141_));
 sg13g2_antennanp ANTENNA_989 (.A(_09141_));
 sg13g2_antennanp ANTENNA_990 (.A(_09141_));
 sg13g2_antennanp ANTENNA_991 (.A(_09141_));
 sg13g2_antennanp ANTENNA_992 (.A(_09149_));
 sg13g2_antennanp ANTENNA_993 (.A(_09149_));
 sg13g2_antennanp ANTENNA_994 (.A(_09149_));
 sg13g2_antennanp ANTENNA_995 (.A(_09149_));
 sg13g2_antennanp ANTENNA_996 (.A(_09149_));
 sg13g2_antennanp ANTENNA_997 (.A(_09149_));
 sg13g2_antennanp ANTENNA_998 (.A(_09150_));
 sg13g2_antennanp ANTENNA_999 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1000 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1001 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1002 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1003 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1004 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1005 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1006 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1007 (.A(_09162_));
 sg13g2_antennanp ANTENNA_1008 (.A(_09162_));
 sg13g2_antennanp ANTENNA_1009 (.A(_09162_));
 sg13g2_antennanp ANTENNA_1010 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1011 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1012 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1013 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1014 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1015 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1016 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1017 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1018 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1019 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1020 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1021 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1022 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1023 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1024 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1025 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1026 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1027 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1028 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1029 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1030 (.A(_09306_));
 sg13g2_antennanp ANTENNA_1031 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1032 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1033 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1034 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1035 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1036 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1037 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1038 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1039 (.A(_09436_));
 sg13g2_antennanp ANTENNA_1040 (.A(_09437_));
 sg13g2_antennanp ANTENNA_1041 (.A(_09437_));
 sg13g2_antennanp ANTENNA_1042 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1043 (.A(_09498_));
 sg13g2_antennanp ANTENNA_1044 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1045 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1046 (.A(_09505_));
 sg13g2_antennanp ANTENNA_1047 (.A(_09531_));
 sg13g2_antennanp ANTENNA_1048 (.A(_09587_));
 sg13g2_antennanp ANTENNA_1049 (.A(_09589_));
 sg13g2_antennanp ANTENNA_1050 (.A(_09615_));
 sg13g2_antennanp ANTENNA_1051 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1052 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1053 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1054 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1055 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1056 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1057 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1058 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1059 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1060 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1061 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1062 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1063 (.A(_10042_));
 sg13g2_antennanp ANTENNA_1064 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1065 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1066 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1067 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1068 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1069 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1070 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1071 (.A(_10113_));
 sg13g2_antennanp ANTENNA_1072 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1073 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1074 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1075 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1076 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1077 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1078 (.A(_10297_));
 sg13g2_antennanp ANTENNA_1079 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1080 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1081 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1082 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1083 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1084 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1085 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1086 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1087 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1088 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1089 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1090 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1091 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1092 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1093 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1094 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1095 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1096 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1097 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1098 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1099 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1100 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1101 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1102 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1103 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1104 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1105 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1106 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1107 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1108 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1109 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1110 (.A(_10779_));
 sg13g2_antennanp ANTENNA_1111 (.A(_11031_));
 sg13g2_antennanp ANTENNA_1112 (.A(_11031_));
 sg13g2_antennanp ANTENNA_1113 (.A(_11031_));
 sg13g2_antennanp ANTENNA_1114 (.A(_11031_));
 sg13g2_antennanp ANTENNA_1115 (.A(_11031_));
 sg13g2_antennanp ANTENNA_1116 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1117 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1118 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1119 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1120 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1121 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1122 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1123 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1124 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1125 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1126 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1127 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1128 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1129 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1130 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1131 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1132 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1133 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1134 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1135 (.A(_12648_));
 sg13g2_antennanp ANTENNA_1136 (.A(_12648_));
 sg13g2_antennanp ANTENNA_1137 (.A(_12648_));
 sg13g2_antennanp ANTENNA_1138 (.A(clk));
 sg13g2_antennanp ANTENNA_1139 (.A(clk));
 sg13g2_antennanp ANTENNA_1140 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1141 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1142 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1143 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1144 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1145 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1146 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1147 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1148 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1149 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1150 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1151 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1152 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1153 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1154 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1155 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1156 (.A(net4));
 sg13g2_antennanp ANTENNA_1157 (.A(net4));
 sg13g2_antennanp ANTENNA_1158 (.A(net4));
 sg13g2_antennanp ANTENNA_1159 (.A(net12));
 sg13g2_antennanp ANTENNA_1160 (.A(net12));
 sg13g2_antennanp ANTENNA_1161 (.A(net12));
 sg13g2_antennanp ANTENNA_1162 (.A(net13));
 sg13g2_antennanp ANTENNA_1163 (.A(net13));
 sg13g2_antennanp ANTENNA_1164 (.A(net13));
 sg13g2_antennanp ANTENNA_1165 (.A(net14));
 sg13g2_antennanp ANTENNA_1166 (.A(net14));
 sg13g2_antennanp ANTENNA_1167 (.A(net14));
 sg13g2_antennanp ANTENNA_1168 (.A(net15));
 sg13g2_antennanp ANTENNA_1169 (.A(net15));
 sg13g2_antennanp ANTENNA_1170 (.A(net15));
 sg13g2_antennanp ANTENNA_1171 (.A(net506));
 sg13g2_antennanp ANTENNA_1172 (.A(net506));
 sg13g2_antennanp ANTENNA_1173 (.A(net506));
 sg13g2_antennanp ANTENNA_1174 (.A(net506));
 sg13g2_antennanp ANTENNA_1175 (.A(net506));
 sg13g2_antennanp ANTENNA_1176 (.A(net506));
 sg13g2_antennanp ANTENNA_1177 (.A(net506));
 sg13g2_antennanp ANTENNA_1178 (.A(net506));
 sg13g2_antennanp ANTENNA_1179 (.A(net506));
 sg13g2_antennanp ANTENNA_1180 (.A(net506));
 sg13g2_antennanp ANTENNA_1181 (.A(net506));
 sg13g2_antennanp ANTENNA_1182 (.A(net506));
 sg13g2_antennanp ANTENNA_1183 (.A(net506));
 sg13g2_antennanp ANTENNA_1184 (.A(net506));
 sg13g2_antennanp ANTENNA_1185 (.A(net506));
 sg13g2_antennanp ANTENNA_1186 (.A(net506));
 sg13g2_antennanp ANTENNA_1187 (.A(net506));
 sg13g2_antennanp ANTENNA_1188 (.A(net506));
 sg13g2_antennanp ANTENNA_1189 (.A(net507));
 sg13g2_antennanp ANTENNA_1190 (.A(net507));
 sg13g2_antennanp ANTENNA_1191 (.A(net507));
 sg13g2_antennanp ANTENNA_1192 (.A(net507));
 sg13g2_antennanp ANTENNA_1193 (.A(net507));
 sg13g2_antennanp ANTENNA_1194 (.A(net507));
 sg13g2_antennanp ANTENNA_1195 (.A(net507));
 sg13g2_antennanp ANTENNA_1196 (.A(net507));
 sg13g2_antennanp ANTENNA_1197 (.A(net507));
 sg13g2_antennanp ANTENNA_1198 (.A(net507));
 sg13g2_antennanp ANTENNA_1199 (.A(net507));
 sg13g2_antennanp ANTENNA_1200 (.A(net507));
 sg13g2_antennanp ANTENNA_1201 (.A(net507));
 sg13g2_antennanp ANTENNA_1202 (.A(net507));
 sg13g2_antennanp ANTENNA_1203 (.A(net507));
 sg13g2_antennanp ANTENNA_1204 (.A(net507));
 sg13g2_antennanp ANTENNA_1205 (.A(net507));
 sg13g2_antennanp ANTENNA_1206 (.A(net507));
 sg13g2_antennanp ANTENNA_1207 (.A(net507));
 sg13g2_antennanp ANTENNA_1208 (.A(net507));
 sg13g2_antennanp ANTENNA_1209 (.A(net507));
 sg13g2_antennanp ANTENNA_1210 (.A(net507));
 sg13g2_antennanp ANTENNA_1211 (.A(net507));
 sg13g2_antennanp ANTENNA_1212 (.A(net551));
 sg13g2_antennanp ANTENNA_1213 (.A(net551));
 sg13g2_antennanp ANTENNA_1214 (.A(net551));
 sg13g2_antennanp ANTENNA_1215 (.A(net551));
 sg13g2_antennanp ANTENNA_1216 (.A(net551));
 sg13g2_antennanp ANTENNA_1217 (.A(net551));
 sg13g2_antennanp ANTENNA_1218 (.A(net551));
 sg13g2_antennanp ANTENNA_1219 (.A(net551));
 sg13g2_antennanp ANTENNA_1220 (.A(net551));
 sg13g2_antennanp ANTENNA_1221 (.A(net551));
 sg13g2_antennanp ANTENNA_1222 (.A(net551));
 sg13g2_antennanp ANTENNA_1223 (.A(net551));
 sg13g2_antennanp ANTENNA_1224 (.A(net551));
 sg13g2_antennanp ANTENNA_1225 (.A(net551));
 sg13g2_antennanp ANTENNA_1226 (.A(net551));
 sg13g2_antennanp ANTENNA_1227 (.A(net551));
 sg13g2_antennanp ANTENNA_1228 (.A(net551));
 sg13g2_antennanp ANTENNA_1229 (.A(net551));
 sg13g2_antennanp ANTENNA_1230 (.A(net551));
 sg13g2_antennanp ANTENNA_1231 (.A(net551));
 sg13g2_antennanp ANTENNA_1232 (.A(net551));
 sg13g2_antennanp ANTENNA_1233 (.A(net551));
 sg13g2_antennanp ANTENNA_1234 (.A(net551));
 sg13g2_antennanp ANTENNA_1235 (.A(net551));
 sg13g2_antennanp ANTENNA_1236 (.A(net599));
 sg13g2_antennanp ANTENNA_1237 (.A(net599));
 sg13g2_antennanp ANTENNA_1238 (.A(net599));
 sg13g2_antennanp ANTENNA_1239 (.A(net599));
 sg13g2_antennanp ANTENNA_1240 (.A(net599));
 sg13g2_antennanp ANTENNA_1241 (.A(net599));
 sg13g2_antennanp ANTENNA_1242 (.A(net599));
 sg13g2_antennanp ANTENNA_1243 (.A(net599));
 sg13g2_antennanp ANTENNA_1244 (.A(net610));
 sg13g2_antennanp ANTENNA_1245 (.A(net610));
 sg13g2_antennanp ANTENNA_1246 (.A(net610));
 sg13g2_antennanp ANTENNA_1247 (.A(net610));
 sg13g2_antennanp ANTENNA_1248 (.A(net610));
 sg13g2_antennanp ANTENNA_1249 (.A(net610));
 sg13g2_antennanp ANTENNA_1250 (.A(net610));
 sg13g2_antennanp ANTENNA_1251 (.A(net610));
 sg13g2_antennanp ANTENNA_1252 (.A(net610));
 sg13g2_antennanp ANTENNA_1253 (.A(net610));
 sg13g2_antennanp ANTENNA_1254 (.A(net610));
 sg13g2_antennanp ANTENNA_1255 (.A(net610));
 sg13g2_antennanp ANTENNA_1256 (.A(net610));
 sg13g2_antennanp ANTENNA_1257 (.A(net610));
 sg13g2_antennanp ANTENNA_1258 (.A(net610));
 sg13g2_antennanp ANTENNA_1259 (.A(net610));
 sg13g2_antennanp ANTENNA_1260 (.A(net610));
 sg13g2_antennanp ANTENNA_1261 (.A(net610));
 sg13g2_antennanp ANTENNA_1262 (.A(net610));
 sg13g2_antennanp ANTENNA_1263 (.A(net610));
 sg13g2_antennanp ANTENNA_1264 (.A(net613));
 sg13g2_antennanp ANTENNA_1265 (.A(net613));
 sg13g2_antennanp ANTENNA_1266 (.A(net613));
 sg13g2_antennanp ANTENNA_1267 (.A(net613));
 sg13g2_antennanp ANTENNA_1268 (.A(net613));
 sg13g2_antennanp ANTENNA_1269 (.A(net613));
 sg13g2_antennanp ANTENNA_1270 (.A(net613));
 sg13g2_antennanp ANTENNA_1271 (.A(net613));
 sg13g2_antennanp ANTENNA_1272 (.A(net613));
 sg13g2_antennanp ANTENNA_1273 (.A(net613));
 sg13g2_antennanp ANTENNA_1274 (.A(net613));
 sg13g2_antennanp ANTENNA_1275 (.A(net613));
 sg13g2_antennanp ANTENNA_1276 (.A(net613));
 sg13g2_antennanp ANTENNA_1277 (.A(net613));
 sg13g2_antennanp ANTENNA_1278 (.A(net613));
 sg13g2_antennanp ANTENNA_1279 (.A(net669));
 sg13g2_antennanp ANTENNA_1280 (.A(net669));
 sg13g2_antennanp ANTENNA_1281 (.A(net669));
 sg13g2_antennanp ANTENNA_1282 (.A(net669));
 sg13g2_antennanp ANTENNA_1283 (.A(net669));
 sg13g2_antennanp ANTENNA_1284 (.A(net669));
 sg13g2_antennanp ANTENNA_1285 (.A(net669));
 sg13g2_antennanp ANTENNA_1286 (.A(net669));
 sg13g2_antennanp ANTENNA_1287 (.A(net669));
 sg13g2_antennanp ANTENNA_1288 (.A(net669));
 sg13g2_antennanp ANTENNA_1289 (.A(net669));
 sg13g2_antennanp ANTENNA_1290 (.A(net669));
 sg13g2_antennanp ANTENNA_1291 (.A(net669));
 sg13g2_antennanp ANTENNA_1292 (.A(net669));
 sg13g2_antennanp ANTENNA_1293 (.A(net669));
 sg13g2_antennanp ANTENNA_1294 (.A(net669));
 sg13g2_antennanp ANTENNA_1295 (.A(net696));
 sg13g2_antennanp ANTENNA_1296 (.A(net696));
 sg13g2_antennanp ANTENNA_1297 (.A(net696));
 sg13g2_antennanp ANTENNA_1298 (.A(net696));
 sg13g2_antennanp ANTENNA_1299 (.A(net696));
 sg13g2_antennanp ANTENNA_1300 (.A(net696));
 sg13g2_antennanp ANTENNA_1301 (.A(net696));
 sg13g2_antennanp ANTENNA_1302 (.A(net696));
 sg13g2_antennanp ANTENNA_1303 (.A(net696));
 sg13g2_antennanp ANTENNA_1304 (.A(net717));
 sg13g2_antennanp ANTENNA_1305 (.A(net717));
 sg13g2_antennanp ANTENNA_1306 (.A(net717));
 sg13g2_antennanp ANTENNA_1307 (.A(net717));
 sg13g2_antennanp ANTENNA_1308 (.A(net717));
 sg13g2_antennanp ANTENNA_1309 (.A(net717));
 sg13g2_antennanp ANTENNA_1310 (.A(net717));
 sg13g2_antennanp ANTENNA_1311 (.A(net717));
 sg13g2_antennanp ANTENNA_1312 (.A(net717));
 sg13g2_antennanp ANTENNA_1313 (.A(net724));
 sg13g2_antennanp ANTENNA_1314 (.A(net724));
 sg13g2_antennanp ANTENNA_1315 (.A(net724));
 sg13g2_antennanp ANTENNA_1316 (.A(net724));
 sg13g2_antennanp ANTENNA_1317 (.A(net724));
 sg13g2_antennanp ANTENNA_1318 (.A(net724));
 sg13g2_antennanp ANTENNA_1319 (.A(net724));
 sg13g2_antennanp ANTENNA_1320 (.A(net724));
 sg13g2_antennanp ANTENNA_1321 (.A(net724));
 sg13g2_antennanp ANTENNA_1322 (.A(net724));
 sg13g2_antennanp ANTENNA_1323 (.A(net724));
 sg13g2_antennanp ANTENNA_1324 (.A(net724));
 sg13g2_antennanp ANTENNA_1325 (.A(net724));
 sg13g2_antennanp ANTENNA_1326 (.A(net724));
 sg13g2_antennanp ANTENNA_1327 (.A(net724));
 sg13g2_antennanp ANTENNA_1328 (.A(net724));
 sg13g2_antennanp ANTENNA_1329 (.A(net802));
 sg13g2_antennanp ANTENNA_1330 (.A(net802));
 sg13g2_antennanp ANTENNA_1331 (.A(net802));
 sg13g2_antennanp ANTENNA_1332 (.A(net802));
 sg13g2_antennanp ANTENNA_1333 (.A(net802));
 sg13g2_antennanp ANTENNA_1334 (.A(net802));
 sg13g2_antennanp ANTENNA_1335 (.A(net802));
 sg13g2_antennanp ANTENNA_1336 (.A(net802));
 sg13g2_antennanp ANTENNA_1337 (.A(net802));
 sg13g2_antennanp ANTENNA_1338 (.A(net850));
 sg13g2_antennanp ANTENNA_1339 (.A(net850));
 sg13g2_antennanp ANTENNA_1340 (.A(net850));
 sg13g2_antennanp ANTENNA_1341 (.A(net850));
 sg13g2_antennanp ANTENNA_1342 (.A(net850));
 sg13g2_antennanp ANTENNA_1343 (.A(net850));
 sg13g2_antennanp ANTENNA_1344 (.A(net850));
 sg13g2_antennanp ANTENNA_1345 (.A(net850));
 sg13g2_antennanp ANTENNA_1346 (.A(net850));
 sg13g2_antennanp ANTENNA_1347 (.A(net904));
 sg13g2_antennanp ANTENNA_1348 (.A(net904));
 sg13g2_antennanp ANTENNA_1349 (.A(net904));
 sg13g2_antennanp ANTENNA_1350 (.A(net904));
 sg13g2_antennanp ANTENNA_1351 (.A(net904));
 sg13g2_antennanp ANTENNA_1352 (.A(net904));
 sg13g2_antennanp ANTENNA_1353 (.A(net904));
 sg13g2_antennanp ANTENNA_1354 (.A(net904));
 sg13g2_antennanp ANTENNA_1355 (.A(net904));
 sg13g2_antennanp ANTENNA_1356 (.A(net974));
 sg13g2_antennanp ANTENNA_1357 (.A(net974));
 sg13g2_antennanp ANTENNA_1358 (.A(net974));
 sg13g2_antennanp ANTENNA_1359 (.A(net974));
 sg13g2_antennanp ANTENNA_1360 (.A(net974));
 sg13g2_antennanp ANTENNA_1361 (.A(net974));
 sg13g2_antennanp ANTENNA_1362 (.A(net974));
 sg13g2_antennanp ANTENNA_1363 (.A(net974));
 sg13g2_antennanp ANTENNA_1364 (.A(net974));
 sg13g2_antennanp ANTENNA_1365 (.A(net977));
 sg13g2_antennanp ANTENNA_1366 (.A(net977));
 sg13g2_antennanp ANTENNA_1367 (.A(net977));
 sg13g2_antennanp ANTENNA_1368 (.A(net977));
 sg13g2_antennanp ANTENNA_1369 (.A(net977));
 sg13g2_antennanp ANTENNA_1370 (.A(net977));
 sg13g2_antennanp ANTENNA_1371 (.A(net977));
 sg13g2_antennanp ANTENNA_1372 (.A(net977));
 sg13g2_antennanp ANTENNA_1373 (.A(net977));
 sg13g2_antennanp ANTENNA_1374 (.A(net1008));
 sg13g2_antennanp ANTENNA_1375 (.A(net1008));
 sg13g2_antennanp ANTENNA_1376 (.A(net1008));
 sg13g2_antennanp ANTENNA_1377 (.A(net1008));
 sg13g2_antennanp ANTENNA_1378 (.A(net1008));
 sg13g2_antennanp ANTENNA_1379 (.A(net1008));
 sg13g2_antennanp ANTENNA_1380 (.A(net1008));
 sg13g2_antennanp ANTENNA_1381 (.A(net1008));
 sg13g2_antennanp ANTENNA_1382 (.A(net1008));
 sg13g2_antennanp ANTENNA_1383 (.A(net1008));
 sg13g2_antennanp ANTENNA_1384 (.A(net1008));
 sg13g2_antennanp ANTENNA_1385 (.A(net1008));
 sg13g2_antennanp ANTENNA_1386 (.A(net1008));
 sg13g2_antennanp ANTENNA_1387 (.A(net1008));
 sg13g2_antennanp ANTENNA_1388 (.A(net1008));
 sg13g2_antennanp ANTENNA_1389 (.A(net1008));
 sg13g2_antennanp ANTENNA_1390 (.A(net1015));
 sg13g2_antennanp ANTENNA_1391 (.A(net1015));
 sg13g2_antennanp ANTENNA_1392 (.A(net1015));
 sg13g2_antennanp ANTENNA_1393 (.A(net1015));
 sg13g2_antennanp ANTENNA_1394 (.A(net1015));
 sg13g2_antennanp ANTENNA_1395 (.A(net1015));
 sg13g2_antennanp ANTENNA_1396 (.A(net1015));
 sg13g2_antennanp ANTENNA_1397 (.A(net1015));
 sg13g2_antennanp ANTENNA_1398 (.A(net1015));
 sg13g2_antennanp ANTENNA_1399 (.A(net1015));
 sg13g2_antennanp ANTENNA_1400 (.A(net1015));
 sg13g2_antennanp ANTENNA_1401 (.A(net1015));
 sg13g2_antennanp ANTENNA_1402 (.A(net1015));
 sg13g2_antennanp ANTENNA_1403 (.A(net1015));
 sg13g2_antennanp ANTENNA_1404 (.A(net1015));
 sg13g2_antennanp ANTENNA_1405 (.A(net1015));
 sg13g2_antennanp ANTENNA_1406 (.A(net1053));
 sg13g2_antennanp ANTENNA_1407 (.A(net1053));
 sg13g2_antennanp ANTENNA_1408 (.A(net1053));
 sg13g2_antennanp ANTENNA_1409 (.A(net1053));
 sg13g2_antennanp ANTENNA_1410 (.A(net1053));
 sg13g2_antennanp ANTENNA_1411 (.A(net1053));
 sg13g2_antennanp ANTENNA_1412 (.A(net1053));
 sg13g2_antennanp ANTENNA_1413 (.A(net1053));
 sg13g2_antennanp ANTENNA_1414 (.A(net1053));
 sg13g2_antennanp ANTENNA_1415 (.A(net1058));
 sg13g2_antennanp ANTENNA_1416 (.A(net1058));
 sg13g2_antennanp ANTENNA_1417 (.A(net1058));
 sg13g2_antennanp ANTENNA_1418 (.A(net1058));
 sg13g2_antennanp ANTENNA_1419 (.A(net1058));
 sg13g2_antennanp ANTENNA_1420 (.A(net1058));
 sg13g2_antennanp ANTENNA_1421 (.A(net1058));
 sg13g2_antennanp ANTENNA_1422 (.A(net1058));
 sg13g2_antennanp ANTENNA_1423 (.A(net1058));
 sg13g2_antennanp ANTENNA_1424 (.A(net1058));
 sg13g2_antennanp ANTENNA_1425 (.A(net1058));
 sg13g2_antennanp ANTENNA_1426 (.A(net1058));
 sg13g2_antennanp ANTENNA_1427 (.A(net1058));
 sg13g2_antennanp ANTENNA_1428 (.A(net1058));
 sg13g2_antennanp ANTENNA_1429 (.A(net1058));
 sg13g2_antennanp ANTENNA_1430 (.A(net1094));
 sg13g2_antennanp ANTENNA_1431 (.A(net1094));
 sg13g2_antennanp ANTENNA_1432 (.A(net1094));
 sg13g2_antennanp ANTENNA_1433 (.A(net1094));
 sg13g2_antennanp ANTENNA_1434 (.A(net1094));
 sg13g2_antennanp ANTENNA_1435 (.A(net1094));
 sg13g2_antennanp ANTENNA_1436 (.A(net1094));
 sg13g2_antennanp ANTENNA_1437 (.A(net1094));
 sg13g2_antennanp ANTENNA_1438 (.A(net1094));
 sg13g2_antennanp ANTENNA_1439 (.A(_00203_));
 sg13g2_antennanp ANTENNA_1440 (.A(_00203_));
 sg13g2_antennanp ANTENNA_1441 (.A(_00209_));
 sg13g2_antennanp ANTENNA_1442 (.A(_00209_));
 sg13g2_antennanp ANTENNA_1443 (.A(_00784_));
 sg13g2_antennanp ANTENNA_1444 (.A(_00784_));
 sg13g2_antennanp ANTENNA_1445 (.A(_00923_));
 sg13g2_antennanp ANTENNA_1446 (.A(_01034_));
 sg13g2_antennanp ANTENNA_1447 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1448 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1449 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1450 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1451 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1452 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1453 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1454 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1455 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1456 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1457 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1458 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1459 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1460 (.A(_03053_));
 sg13g2_antennanp ANTENNA_1461 (.A(_03053_));
 sg13g2_antennanp ANTENNA_1462 (.A(_03053_));
 sg13g2_antennanp ANTENNA_1463 (.A(_03053_));
 sg13g2_antennanp ANTENNA_1464 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1465 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1466 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1467 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1468 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1469 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1470 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1471 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1472 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1473 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1474 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1475 (.A(_04751_));
 sg13g2_antennanp ANTENNA_1476 (.A(_04775_));
 sg13g2_antennanp ANTENNA_1477 (.A(_04775_));
 sg13g2_antennanp ANTENNA_1478 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1479 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1480 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1481 (.A(_04985_));
 sg13g2_antennanp ANTENNA_1482 (.A(_04985_));
 sg13g2_antennanp ANTENNA_1483 (.A(_05003_));
 sg13g2_antennanp ANTENNA_1484 (.A(_05126_));
 sg13g2_antennanp ANTENNA_1485 (.A(_05149_));
 sg13g2_antennanp ANTENNA_1486 (.A(_05174_));
 sg13g2_antennanp ANTENNA_1487 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1488 (.A(_05215_));
 sg13g2_antennanp ANTENNA_1489 (.A(_05309_));
 sg13g2_antennanp ANTENNA_1490 (.A(_05583_));
 sg13g2_antennanp ANTENNA_1491 (.A(_05653_));
 sg13g2_antennanp ANTENNA_1492 (.A(_05667_));
 sg13g2_antennanp ANTENNA_1493 (.A(_05669_));
 sg13g2_antennanp ANTENNA_1494 (.A(_05680_));
 sg13g2_antennanp ANTENNA_1495 (.A(_05700_));
 sg13g2_antennanp ANTENNA_1496 (.A(_05706_));
 sg13g2_antennanp ANTENNA_1497 (.A(_05712_));
 sg13g2_antennanp ANTENNA_1498 (.A(_05724_));
 sg13g2_antennanp ANTENNA_1499 (.A(_05724_));
 sg13g2_antennanp ANTENNA_1500 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1501 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1502 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1503 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1504 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1505 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1506 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1507 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1508 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1509 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1510 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1511 (.A(_05900_));
 sg13g2_antennanp ANTENNA_1512 (.A(_05955_));
 sg13g2_antennanp ANTENNA_1513 (.A(_06556_));
 sg13g2_antennanp ANTENNA_1514 (.A(_06556_));
 sg13g2_antennanp ANTENNA_1515 (.A(_06556_));
 sg13g2_antennanp ANTENNA_1516 (.A(_06556_));
 sg13g2_antennanp ANTENNA_1517 (.A(_06818_));
 sg13g2_antennanp ANTENNA_1518 (.A(_06818_));
 sg13g2_antennanp ANTENNA_1519 (.A(_06818_));
 sg13g2_antennanp ANTENNA_1520 (.A(_06818_));
 sg13g2_antennanp ANTENNA_1521 (.A(_07576_));
 sg13g2_antennanp ANTENNA_1522 (.A(_07576_));
 sg13g2_antennanp ANTENNA_1523 (.A(_07877_));
 sg13g2_antennanp ANTENNA_1524 (.A(_07877_));
 sg13g2_antennanp ANTENNA_1525 (.A(_07877_));
 sg13g2_antennanp ANTENNA_1526 (.A(_08204_));
 sg13g2_antennanp ANTENNA_1527 (.A(_08204_));
 sg13g2_antennanp ANTENNA_1528 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1529 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1530 (.A(_08327_));
 sg13g2_antennanp ANTENNA_1531 (.A(_08408_));
 sg13g2_antennanp ANTENNA_1532 (.A(_08408_));
 sg13g2_antennanp ANTENNA_1533 (.A(_08408_));
 sg13g2_antennanp ANTENNA_1534 (.A(_08408_));
 sg13g2_antennanp ANTENNA_1535 (.A(_08408_));
 sg13g2_antennanp ANTENNA_1536 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1537 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1538 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1539 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1540 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1541 (.A(_08439_));
 sg13g2_antennanp ANTENNA_1542 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1543 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1544 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1545 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1546 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1547 (.A(_08507_));
 sg13g2_antennanp ANTENNA_1548 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1549 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1550 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1551 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1552 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1553 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1554 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1555 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1556 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1557 (.A(_08798_));
 sg13g2_antennanp ANTENNA_1558 (.A(_08798_));
 sg13g2_antennanp ANTENNA_1559 (.A(_08798_));
 sg13g2_antennanp ANTENNA_1560 (.A(_08818_));
 sg13g2_antennanp ANTENNA_1561 (.A(_08840_));
 sg13g2_antennanp ANTENNA_1562 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1563 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1564 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1565 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1566 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1567 (.A(_08851_));
 sg13g2_antennanp ANTENNA_1568 (.A(_09084_));
 sg13g2_antennanp ANTENNA_1569 (.A(_09084_));
 sg13g2_antennanp ANTENNA_1570 (.A(_09084_));
 sg13g2_antennanp ANTENNA_1571 (.A(_09131_));
 sg13g2_antennanp ANTENNA_1572 (.A(_09131_));
 sg13g2_antennanp ANTENNA_1573 (.A(_09131_));
 sg13g2_antennanp ANTENNA_1574 (.A(_09131_));
 sg13g2_antennanp ANTENNA_1575 (.A(_09140_));
 sg13g2_antennanp ANTENNA_1576 (.A(_09140_));
 sg13g2_antennanp ANTENNA_1577 (.A(_09140_));
 sg13g2_antennanp ANTENNA_1578 (.A(_09141_));
 sg13g2_antennanp ANTENNA_1579 (.A(_09141_));
 sg13g2_antennanp ANTENNA_1580 (.A(_09141_));
 sg13g2_antennanp ANTENNA_1581 (.A(_09141_));
 sg13g2_antennanp ANTENNA_1582 (.A(_09149_));
 sg13g2_antennanp ANTENNA_1583 (.A(_09149_));
 sg13g2_antennanp ANTENNA_1584 (.A(_09149_));
 sg13g2_antennanp ANTENNA_1585 (.A(_09149_));
 sg13g2_antennanp ANTENNA_1586 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1587 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1588 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1589 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1590 (.A(_09150_));
 sg13g2_antennanp ANTENNA_1591 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1592 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1593 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1594 (.A(_09151_));
 sg13g2_antennanp ANTENNA_1595 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1596 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1597 (.A(_09163_));
 sg13g2_antennanp ANTENNA_1598 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1599 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1600 (.A(_09230_));
 sg13g2_antennanp ANTENNA_1601 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1602 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1603 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1604 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1605 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1606 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1607 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1608 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1609 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1610 (.A(_09253_));
 sg13g2_antennanp ANTENNA_1611 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1612 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1613 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1614 (.A(_09254_));
 sg13g2_antennanp ANTENNA_1615 (.A(_09306_));
 sg13g2_antennanp ANTENNA_1616 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1617 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1618 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1619 (.A(_09420_));
 sg13g2_antennanp ANTENNA_1620 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1621 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1622 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1623 (.A(_09426_));
 sg13g2_antennanp ANTENNA_1624 (.A(_09436_));
 sg13g2_antennanp ANTENNA_1625 (.A(_09437_));
 sg13g2_antennanp ANTENNA_1626 (.A(_09437_));
 sg13g2_antennanp ANTENNA_1627 (.A(_09445_));
 sg13g2_antennanp ANTENNA_1628 (.A(_09498_));
 sg13g2_antennanp ANTENNA_1629 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1630 (.A(_09499_));
 sg13g2_antennanp ANTENNA_1631 (.A(_09505_));
 sg13g2_antennanp ANTENNA_1632 (.A(_09531_));
 sg13g2_antennanp ANTENNA_1633 (.A(_09587_));
 sg13g2_antennanp ANTENNA_1634 (.A(_09589_));
 sg13g2_antennanp ANTENNA_1635 (.A(_09589_));
 sg13g2_antennanp ANTENNA_1636 (.A(_09615_));
 sg13g2_antennanp ANTENNA_1637 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1638 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1639 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1640 (.A(_09660_));
 sg13g2_antennanp ANTENNA_1641 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1642 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1643 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1644 (.A(_09907_));
 sg13g2_antennanp ANTENNA_1645 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1646 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1647 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1648 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1649 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1650 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1651 (.A(_10330_));
 sg13g2_antennanp ANTENNA_1652 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1653 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1654 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1655 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1656 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1657 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1658 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1659 (.A(_10368_));
 sg13g2_antennanp ANTENNA_1660 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1661 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1662 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1663 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1664 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1665 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1666 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1667 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1668 (.A(_10458_));
 sg13g2_antennanp ANTENNA_1669 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1670 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1671 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1672 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1673 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1674 (.A(_10478_));
 sg13g2_antennanp ANTENNA_1675 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1676 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1677 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1678 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1679 (.A(_10629_));
 sg13g2_antennanp ANTENNA_1680 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1681 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1682 (.A(_10634_));
 sg13g2_antennanp ANTENNA_1683 (.A(_10779_));
 sg13g2_antennanp ANTENNA_1684 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1685 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1686 (.A(_11776_));
 sg13g2_antennanp ANTENNA_1687 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1688 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1689 (.A(_11919_));
 sg13g2_antennanp ANTENNA_1690 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1691 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1692 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1693 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1694 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1695 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1696 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1697 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1698 (.A(_11926_));
 sg13g2_antennanp ANTENNA_1699 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1700 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1701 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1702 (.A(_11960_));
 sg13g2_antennanp ANTENNA_1703 (.A(clk));
 sg13g2_antennanp ANTENNA_1704 (.A(clk));
 sg13g2_antennanp ANTENNA_1705 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1706 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1707 (.A(\cpu.ex.r_mult[29] ));
 sg13g2_antennanp ANTENNA_1708 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1709 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1710 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_1711 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1712 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1713 (.A(\cpu.ex.r_mult[31] ));
 sg13g2_antennanp ANTENNA_1714 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1715 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1716 (.A(net4));
 sg13g2_antennanp ANTENNA_1717 (.A(net4));
 sg13g2_antennanp ANTENNA_1718 (.A(net4));
 sg13g2_antennanp ANTENNA_1719 (.A(net12));
 sg13g2_antennanp ANTENNA_1720 (.A(net12));
 sg13g2_antennanp ANTENNA_1721 (.A(net12));
 sg13g2_antennanp ANTENNA_1722 (.A(net13));
 sg13g2_antennanp ANTENNA_1723 (.A(net13));
 sg13g2_antennanp ANTENNA_1724 (.A(net13));
 sg13g2_antennanp ANTENNA_1725 (.A(net14));
 sg13g2_antennanp ANTENNA_1726 (.A(net14));
 sg13g2_antennanp ANTENNA_1727 (.A(net14));
 sg13g2_antennanp ANTENNA_1728 (.A(net15));
 sg13g2_antennanp ANTENNA_1729 (.A(net15));
 sg13g2_antennanp ANTENNA_1730 (.A(net15));
 sg13g2_antennanp ANTENNA_1731 (.A(net506));
 sg13g2_antennanp ANTENNA_1732 (.A(net506));
 sg13g2_antennanp ANTENNA_1733 (.A(net506));
 sg13g2_antennanp ANTENNA_1734 (.A(net506));
 sg13g2_antennanp ANTENNA_1735 (.A(net506));
 sg13g2_antennanp ANTENNA_1736 (.A(net506));
 sg13g2_antennanp ANTENNA_1737 (.A(net506));
 sg13g2_antennanp ANTENNA_1738 (.A(net506));
 sg13g2_antennanp ANTENNA_1739 (.A(net506));
 sg13g2_antennanp ANTENNA_1740 (.A(net506));
 sg13g2_antennanp ANTENNA_1741 (.A(net506));
 sg13g2_antennanp ANTENNA_1742 (.A(net507));
 sg13g2_antennanp ANTENNA_1743 (.A(net507));
 sg13g2_antennanp ANTENNA_1744 (.A(net507));
 sg13g2_antennanp ANTENNA_1745 (.A(net507));
 sg13g2_antennanp ANTENNA_1746 (.A(net507));
 sg13g2_antennanp ANTENNA_1747 (.A(net507));
 sg13g2_antennanp ANTENNA_1748 (.A(net507));
 sg13g2_antennanp ANTENNA_1749 (.A(net507));
 sg13g2_antennanp ANTENNA_1750 (.A(net507));
 sg13g2_antennanp ANTENNA_1751 (.A(net507));
 sg13g2_antennanp ANTENNA_1752 (.A(net507));
 sg13g2_antennanp ANTENNA_1753 (.A(net507));
 sg13g2_antennanp ANTENNA_1754 (.A(net507));
 sg13g2_antennanp ANTENNA_1755 (.A(net507));
 sg13g2_antennanp ANTENNA_1756 (.A(net507));
 sg13g2_antennanp ANTENNA_1757 (.A(net507));
 sg13g2_antennanp ANTENNA_1758 (.A(net507));
 sg13g2_antennanp ANTENNA_1759 (.A(net507));
 sg13g2_antennanp ANTENNA_1760 (.A(net507));
 sg13g2_antennanp ANTENNA_1761 (.A(net599));
 sg13g2_antennanp ANTENNA_1762 (.A(net599));
 sg13g2_antennanp ANTENNA_1763 (.A(net599));
 sg13g2_antennanp ANTENNA_1764 (.A(net599));
 sg13g2_antennanp ANTENNA_1765 (.A(net599));
 sg13g2_antennanp ANTENNA_1766 (.A(net599));
 sg13g2_antennanp ANTENNA_1767 (.A(net599));
 sg13g2_antennanp ANTENNA_1768 (.A(net599));
 sg13g2_antennanp ANTENNA_1769 (.A(net610));
 sg13g2_antennanp ANTENNA_1770 (.A(net610));
 sg13g2_antennanp ANTENNA_1771 (.A(net610));
 sg13g2_antennanp ANTENNA_1772 (.A(net610));
 sg13g2_antennanp ANTENNA_1773 (.A(net610));
 sg13g2_antennanp ANTENNA_1774 (.A(net610));
 sg13g2_antennanp ANTENNA_1775 (.A(net610));
 sg13g2_antennanp ANTENNA_1776 (.A(net610));
 sg13g2_antennanp ANTENNA_1777 (.A(net610));
 sg13g2_antennanp ANTENNA_1778 (.A(net610));
 sg13g2_antennanp ANTENNA_1779 (.A(net610));
 sg13g2_antennanp ANTENNA_1780 (.A(net610));
 sg13g2_antennanp ANTENNA_1781 (.A(net610));
 sg13g2_antennanp ANTENNA_1782 (.A(net610));
 sg13g2_antennanp ANTENNA_1783 (.A(net610));
 sg13g2_antennanp ANTENNA_1784 (.A(net610));
 sg13g2_antennanp ANTENNA_1785 (.A(net610));
 sg13g2_antennanp ANTENNA_1786 (.A(net610));
 sg13g2_antennanp ANTENNA_1787 (.A(net610));
 sg13g2_antennanp ANTENNA_1788 (.A(net610));
 sg13g2_antennanp ANTENNA_1789 (.A(net613));
 sg13g2_antennanp ANTENNA_1790 (.A(net613));
 sg13g2_antennanp ANTENNA_1791 (.A(net613));
 sg13g2_antennanp ANTENNA_1792 (.A(net613));
 sg13g2_antennanp ANTENNA_1793 (.A(net613));
 sg13g2_antennanp ANTENNA_1794 (.A(net613));
 sg13g2_antennanp ANTENNA_1795 (.A(net613));
 sg13g2_antennanp ANTENNA_1796 (.A(net613));
 sg13g2_antennanp ANTENNA_1797 (.A(net613));
 sg13g2_antennanp ANTENNA_1798 (.A(net613));
 sg13g2_antennanp ANTENNA_1799 (.A(net613));
 sg13g2_antennanp ANTENNA_1800 (.A(net613));
 sg13g2_antennanp ANTENNA_1801 (.A(net613));
 sg13g2_antennanp ANTENNA_1802 (.A(net613));
 sg13g2_antennanp ANTENNA_1803 (.A(net613));
 sg13g2_antennanp ANTENNA_1804 (.A(net613));
 sg13g2_antennanp ANTENNA_1805 (.A(net696));
 sg13g2_antennanp ANTENNA_1806 (.A(net696));
 sg13g2_antennanp ANTENNA_1807 (.A(net696));
 sg13g2_antennanp ANTENNA_1808 (.A(net696));
 sg13g2_antennanp ANTENNA_1809 (.A(net696));
 sg13g2_antennanp ANTENNA_1810 (.A(net696));
 sg13g2_antennanp ANTENNA_1811 (.A(net696));
 sg13g2_antennanp ANTENNA_1812 (.A(net696));
 sg13g2_antennanp ANTENNA_1813 (.A(net696));
 sg13g2_antennanp ANTENNA_1814 (.A(net717));
 sg13g2_antennanp ANTENNA_1815 (.A(net717));
 sg13g2_antennanp ANTENNA_1816 (.A(net717));
 sg13g2_antennanp ANTENNA_1817 (.A(net717));
 sg13g2_antennanp ANTENNA_1818 (.A(net717));
 sg13g2_antennanp ANTENNA_1819 (.A(net717));
 sg13g2_antennanp ANTENNA_1820 (.A(net717));
 sg13g2_antennanp ANTENNA_1821 (.A(net717));
 sg13g2_antennanp ANTENNA_1822 (.A(net717));
 sg13g2_antennanp ANTENNA_1823 (.A(net724));
 sg13g2_antennanp ANTENNA_1824 (.A(net724));
 sg13g2_antennanp ANTENNA_1825 (.A(net724));
 sg13g2_antennanp ANTENNA_1826 (.A(net724));
 sg13g2_antennanp ANTENNA_1827 (.A(net724));
 sg13g2_antennanp ANTENNA_1828 (.A(net724));
 sg13g2_antennanp ANTENNA_1829 (.A(net724));
 sg13g2_antennanp ANTENNA_1830 (.A(net724));
 sg13g2_antennanp ANTENNA_1831 (.A(net724));
 sg13g2_antennanp ANTENNA_1832 (.A(net724));
 sg13g2_antennanp ANTENNA_1833 (.A(net724));
 sg13g2_antennanp ANTENNA_1834 (.A(net724));
 sg13g2_antennanp ANTENNA_1835 (.A(net724));
 sg13g2_antennanp ANTENNA_1836 (.A(net724));
 sg13g2_antennanp ANTENNA_1837 (.A(net724));
 sg13g2_antennanp ANTENNA_1838 (.A(net724));
 sg13g2_antennanp ANTENNA_1839 (.A(net802));
 sg13g2_antennanp ANTENNA_1840 (.A(net802));
 sg13g2_antennanp ANTENNA_1841 (.A(net802));
 sg13g2_antennanp ANTENNA_1842 (.A(net802));
 sg13g2_antennanp ANTENNA_1843 (.A(net802));
 sg13g2_antennanp ANTENNA_1844 (.A(net802));
 sg13g2_antennanp ANTENNA_1845 (.A(net802));
 sg13g2_antennanp ANTENNA_1846 (.A(net802));
 sg13g2_antennanp ANTENNA_1847 (.A(net802));
 sg13g2_antennanp ANTENNA_1848 (.A(net802));
 sg13g2_antennanp ANTENNA_1849 (.A(net802));
 sg13g2_antennanp ANTENNA_1850 (.A(net802));
 sg13g2_antennanp ANTENNA_1851 (.A(net802));
 sg13g2_antennanp ANTENNA_1852 (.A(net802));
 sg13g2_antennanp ANTENNA_1853 (.A(net802));
 sg13g2_antennanp ANTENNA_1854 (.A(net802));
 sg13g2_antennanp ANTENNA_1855 (.A(net850));
 sg13g2_antennanp ANTENNA_1856 (.A(net850));
 sg13g2_antennanp ANTENNA_1857 (.A(net850));
 sg13g2_antennanp ANTENNA_1858 (.A(net850));
 sg13g2_antennanp ANTENNA_1859 (.A(net850));
 sg13g2_antennanp ANTENNA_1860 (.A(net850));
 sg13g2_antennanp ANTENNA_1861 (.A(net850));
 sg13g2_antennanp ANTENNA_1862 (.A(net850));
 sg13g2_antennanp ANTENNA_1863 (.A(net850));
 sg13g2_antennanp ANTENNA_1864 (.A(net974));
 sg13g2_antennanp ANTENNA_1865 (.A(net974));
 sg13g2_antennanp ANTENNA_1866 (.A(net974));
 sg13g2_antennanp ANTENNA_1867 (.A(net974));
 sg13g2_antennanp ANTENNA_1868 (.A(net974));
 sg13g2_antennanp ANTENNA_1869 (.A(net974));
 sg13g2_antennanp ANTENNA_1870 (.A(net974));
 sg13g2_antennanp ANTENNA_1871 (.A(net974));
 sg13g2_antennanp ANTENNA_1872 (.A(net974));
 sg13g2_antennanp ANTENNA_1873 (.A(net977));
 sg13g2_antennanp ANTENNA_1874 (.A(net977));
 sg13g2_antennanp ANTENNA_1875 (.A(net977));
 sg13g2_antennanp ANTENNA_1876 (.A(net977));
 sg13g2_antennanp ANTENNA_1877 (.A(net977));
 sg13g2_antennanp ANTENNA_1878 (.A(net977));
 sg13g2_antennanp ANTENNA_1879 (.A(net977));
 sg13g2_antennanp ANTENNA_1880 (.A(net977));
 sg13g2_antennanp ANTENNA_1881 (.A(net977));
 sg13g2_antennanp ANTENNA_1882 (.A(net1008));
 sg13g2_antennanp ANTENNA_1883 (.A(net1008));
 sg13g2_antennanp ANTENNA_1884 (.A(net1008));
 sg13g2_antennanp ANTENNA_1885 (.A(net1008));
 sg13g2_antennanp ANTENNA_1886 (.A(net1008));
 sg13g2_antennanp ANTENNA_1887 (.A(net1008));
 sg13g2_antennanp ANTENNA_1888 (.A(net1008));
 sg13g2_antennanp ANTENNA_1889 (.A(net1008));
 sg13g2_antennanp ANTENNA_1890 (.A(net1008));
 sg13g2_antennanp ANTENNA_1891 (.A(net1008));
 sg13g2_antennanp ANTENNA_1892 (.A(net1008));
 sg13g2_antennanp ANTENNA_1893 (.A(net1008));
 sg13g2_antennanp ANTENNA_1894 (.A(net1008));
 sg13g2_antennanp ANTENNA_1895 (.A(net1008));
 sg13g2_antennanp ANTENNA_1896 (.A(net1008));
 sg13g2_antennanp ANTENNA_1897 (.A(net1008));
 sg13g2_antennanp ANTENNA_1898 (.A(net1012));
 sg13g2_antennanp ANTENNA_1899 (.A(net1012));
 sg13g2_antennanp ANTENNA_1900 (.A(net1012));
 sg13g2_antennanp ANTENNA_1901 (.A(net1012));
 sg13g2_antennanp ANTENNA_1902 (.A(net1012));
 sg13g2_antennanp ANTENNA_1903 (.A(net1012));
 sg13g2_antennanp ANTENNA_1904 (.A(net1012));
 sg13g2_antennanp ANTENNA_1905 (.A(net1012));
 sg13g2_antennanp ANTENNA_1906 (.A(net1012));
 sg13g2_antennanp ANTENNA_1907 (.A(net1053));
 sg13g2_antennanp ANTENNA_1908 (.A(net1053));
 sg13g2_antennanp ANTENNA_1909 (.A(net1053));
 sg13g2_antennanp ANTENNA_1910 (.A(net1053));
 sg13g2_antennanp ANTENNA_1911 (.A(net1053));
 sg13g2_antennanp ANTENNA_1912 (.A(net1053));
 sg13g2_antennanp ANTENNA_1913 (.A(net1053));
 sg13g2_antennanp ANTENNA_1914 (.A(net1053));
 sg13g2_antennanp ANTENNA_1915 (.A(net1053));
 sg13g2_antennanp ANTENNA_1916 (.A(net1058));
 sg13g2_antennanp ANTENNA_1917 (.A(net1058));
 sg13g2_antennanp ANTENNA_1918 (.A(net1058));
 sg13g2_antennanp ANTENNA_1919 (.A(net1058));
 sg13g2_antennanp ANTENNA_1920 (.A(net1058));
 sg13g2_antennanp ANTENNA_1921 (.A(net1058));
 sg13g2_antennanp ANTENNA_1922 (.A(net1058));
 sg13g2_antennanp ANTENNA_1923 (.A(net1058));
 sg13g2_antennanp ANTENNA_1924 (.A(net1058));
 sg13g2_antennanp ANTENNA_1925 (.A(net1058));
 sg13g2_antennanp ANTENNA_1926 (.A(net1058));
 sg13g2_antennanp ANTENNA_1927 (.A(net1058));
 sg13g2_antennanp ANTENNA_1928 (.A(net1058));
 sg13g2_antennanp ANTENNA_1929 (.A(net1058));
 sg13g2_antennanp ANTENNA_1930 (.A(net1058));
 sg13g2_antennanp ANTENNA_1931 (.A(_00203_));
 sg13g2_antennanp ANTENNA_1932 (.A(_00203_));
 sg13g2_antennanp ANTENNA_1933 (.A(_00209_));
 sg13g2_antennanp ANTENNA_1934 (.A(_00784_));
 sg13g2_antennanp ANTENNA_1935 (.A(_00784_));
 sg13g2_antennanp ANTENNA_1936 (.A(_00923_));
 sg13g2_antennanp ANTENNA_1937 (.A(_01034_));
 sg13g2_antennanp ANTENNA_1938 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1939 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1940 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1941 (.A(_02779_));
 sg13g2_antennanp ANTENNA_1942 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1943 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1944 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1945 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1946 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1947 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1948 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1949 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1950 (.A(_02910_));
 sg13g2_antennanp ANTENNA_1951 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1952 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1953 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1954 (.A(_03478_));
 sg13g2_antennanp ANTENNA_1955 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1956 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1957 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1958 (.A(_03527_));
 sg13g2_antennanp ANTENNA_1959 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1960 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1961 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1962 (.A(_04734_));
 sg13g2_antennanp ANTENNA_1963 (.A(_04751_));
 sg13g2_antennanp ANTENNA_1964 (.A(_04775_));
 sg13g2_antennanp ANTENNA_1965 (.A(_04775_));
 sg13g2_antennanp ANTENNA_1966 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1967 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1968 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1969 (.A(_04778_));
 sg13g2_antennanp ANTENNA_1970 (.A(_04927_));
 sg13g2_antennanp ANTENNA_1971 (.A(_04985_));
 sg13g2_antennanp ANTENNA_1972 (.A(_04985_));
 sg13g2_antennanp ANTENNA_1973 (.A(_05003_));
 sg13g2_antennanp ANTENNA_1974 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1975 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1976 (.A(_05090_));
 sg13g2_antennanp ANTENNA_1977 (.A(_05126_));
 sg13g2_antennanp ANTENNA_1978 (.A(_05149_));
 sg13g2_antennanp ANTENNA_1979 (.A(_05160_));
 sg13g2_antennanp ANTENNA_1980 (.A(_05174_));
 sg13g2_antennanp ANTENNA_1981 (.A(_05201_));
 sg13g2_antennanp ANTENNA_1982 (.A(_05215_));
 sg13g2_antennanp ANTENNA_1983 (.A(_05309_));
 sg13g2_antennanp ANTENNA_1984 (.A(_05583_));
 sg13g2_antennanp ANTENNA_1985 (.A(_05653_));
 sg13g2_antennanp ANTENNA_1986 (.A(_05667_));
 sg13g2_antennanp ANTENNA_1987 (.A(_05667_));
 sg13g2_antennanp ANTENNA_1988 (.A(_05669_));
 sg13g2_antennanp ANTENNA_1989 (.A(_05680_));
 sg13g2_antennanp ANTENNA_1990 (.A(_05706_));
 sg13g2_antennanp ANTENNA_1991 (.A(_05712_));
 sg13g2_antennanp ANTENNA_1992 (.A(_05724_));
 sg13g2_antennanp ANTENNA_1993 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1994 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1995 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1996 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1997 (.A(_05895_));
 sg13g2_antennanp ANTENNA_1998 (.A(_05955_));
 sg13g2_antennanp ANTENNA_1999 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2000 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2001 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2002 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2003 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2004 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2005 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2006 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2007 (.A(_07576_));
 sg13g2_antennanp ANTENNA_2008 (.A(_07576_));
 sg13g2_antennanp ANTENNA_2009 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2010 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2011 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2012 (.A(_08204_));
 sg13g2_antennanp ANTENNA_2013 (.A(_08204_));
 sg13g2_antennanp ANTENNA_2014 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2015 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2016 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2017 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2018 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2019 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2020 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2021 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2022 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2023 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2024 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2025 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2026 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2027 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2028 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2029 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2030 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2031 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2032 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2033 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2034 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2035 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2036 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2037 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2038 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2039 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2040 (.A(_08818_));
 sg13g2_antennanp ANTENNA_2041 (.A(_08840_));
 sg13g2_antennanp ANTENNA_2042 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2043 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2044 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2045 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2046 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2047 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2048 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2049 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2050 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2051 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2052 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2053 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2054 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2055 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2056 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2057 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2058 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2059 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2060 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2061 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2062 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2063 (.A(_09143_));
 sg13g2_antennanp ANTENNA_2064 (.A(_09143_));
 sg13g2_antennanp ANTENNA_2065 (.A(_09143_));
 sg13g2_antennanp ANTENNA_2066 (.A(_09143_));
 sg13g2_antennanp ANTENNA_2067 (.A(_09143_));
 sg13g2_antennanp ANTENNA_2068 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2069 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2070 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2071 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2072 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2073 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2074 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2075 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2076 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2077 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2078 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2079 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2080 (.A(_09151_));
 sg13g2_antennanp ANTENNA_2081 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2082 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2083 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2084 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2085 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2086 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2087 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2088 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2089 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2090 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2091 (.A(_09306_));
 sg13g2_antennanp ANTENNA_2092 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2093 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2094 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2095 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2096 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2097 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2098 (.A(_09436_));
 sg13g2_antennanp ANTENNA_2099 (.A(_09437_));
 sg13g2_antennanp ANTENNA_2100 (.A(_09437_));
 sg13g2_antennanp ANTENNA_2101 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2102 (.A(_09498_));
 sg13g2_antennanp ANTENNA_2103 (.A(_09499_));
 sg13g2_antennanp ANTENNA_2104 (.A(_09499_));
 sg13g2_antennanp ANTENNA_2105 (.A(_09505_));
 sg13g2_antennanp ANTENNA_2106 (.A(_09531_));
 sg13g2_antennanp ANTENNA_2107 (.A(_09587_));
 sg13g2_antennanp ANTENNA_2108 (.A(_09615_));
 sg13g2_antennanp ANTENNA_2109 (.A(_09660_));
 sg13g2_antennanp ANTENNA_2110 (.A(_09660_));
 sg13g2_antennanp ANTENNA_2111 (.A(_09660_));
 sg13g2_antennanp ANTENNA_2112 (.A(_09660_));
 sg13g2_antennanp ANTENNA_2113 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2114 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2115 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2116 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2117 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2118 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2119 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2120 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2121 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2122 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2123 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2124 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2125 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2126 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2127 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2128 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2129 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2130 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2131 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2132 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2133 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2134 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2135 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2136 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2137 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2138 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2139 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2140 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2141 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2142 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2143 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2144 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2145 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2146 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2147 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2148 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2149 (.A(_10629_));
 sg13g2_antennanp ANTENNA_2150 (.A(_10629_));
 sg13g2_antennanp ANTENNA_2151 (.A(_10629_));
 sg13g2_antennanp ANTENNA_2152 (.A(_10629_));
 sg13g2_antennanp ANTENNA_2153 (.A(_10629_));
 sg13g2_antennanp ANTENNA_2154 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2155 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2156 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2157 (.A(_11210_));
 sg13g2_antennanp ANTENNA_2158 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2159 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2160 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2161 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2162 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2163 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2164 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2165 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2166 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2167 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2168 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2169 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2170 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2171 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2172 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2173 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2174 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2175 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2176 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2177 (.A(clk));
 sg13g2_antennanp ANTENNA_2178 (.A(clk));
 sg13g2_antennanp ANTENNA_2179 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2180 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2181 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2182 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2183 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2184 (.A(net4));
 sg13g2_antennanp ANTENNA_2185 (.A(net4));
 sg13g2_antennanp ANTENNA_2186 (.A(net4));
 sg13g2_antennanp ANTENNA_2187 (.A(net12));
 sg13g2_antennanp ANTENNA_2188 (.A(net12));
 sg13g2_antennanp ANTENNA_2189 (.A(net12));
 sg13g2_antennanp ANTENNA_2190 (.A(net13));
 sg13g2_antennanp ANTENNA_2191 (.A(net13));
 sg13g2_antennanp ANTENNA_2192 (.A(net13));
 sg13g2_antennanp ANTENNA_2193 (.A(net14));
 sg13g2_antennanp ANTENNA_2194 (.A(net14));
 sg13g2_antennanp ANTENNA_2195 (.A(net14));
 sg13g2_antennanp ANTENNA_2196 (.A(net506));
 sg13g2_antennanp ANTENNA_2197 (.A(net506));
 sg13g2_antennanp ANTENNA_2198 (.A(net506));
 sg13g2_antennanp ANTENNA_2199 (.A(net506));
 sg13g2_antennanp ANTENNA_2200 (.A(net506));
 sg13g2_antennanp ANTENNA_2201 (.A(net506));
 sg13g2_antennanp ANTENNA_2202 (.A(net506));
 sg13g2_antennanp ANTENNA_2203 (.A(net506));
 sg13g2_antennanp ANTENNA_2204 (.A(net506));
 sg13g2_antennanp ANTENNA_2205 (.A(net506));
 sg13g2_antennanp ANTENNA_2206 (.A(net506));
 sg13g2_antennanp ANTENNA_2207 (.A(net507));
 sg13g2_antennanp ANTENNA_2208 (.A(net507));
 sg13g2_antennanp ANTENNA_2209 (.A(net507));
 sg13g2_antennanp ANTENNA_2210 (.A(net507));
 sg13g2_antennanp ANTENNA_2211 (.A(net507));
 sg13g2_antennanp ANTENNA_2212 (.A(net507));
 sg13g2_antennanp ANTENNA_2213 (.A(net507));
 sg13g2_antennanp ANTENNA_2214 (.A(net507));
 sg13g2_antennanp ANTENNA_2215 (.A(net507));
 sg13g2_antennanp ANTENNA_2216 (.A(net507));
 sg13g2_antennanp ANTENNA_2217 (.A(net507));
 sg13g2_antennanp ANTENNA_2218 (.A(net507));
 sg13g2_antennanp ANTENNA_2219 (.A(net507));
 sg13g2_antennanp ANTENNA_2220 (.A(net507));
 sg13g2_antennanp ANTENNA_2221 (.A(net507));
 sg13g2_antennanp ANTENNA_2222 (.A(net507));
 sg13g2_antennanp ANTENNA_2223 (.A(net507));
 sg13g2_antennanp ANTENNA_2224 (.A(net507));
 sg13g2_antennanp ANTENNA_2225 (.A(net507));
 sg13g2_antennanp ANTENNA_2226 (.A(net551));
 sg13g2_antennanp ANTENNA_2227 (.A(net551));
 sg13g2_antennanp ANTENNA_2228 (.A(net551));
 sg13g2_antennanp ANTENNA_2229 (.A(net551));
 sg13g2_antennanp ANTENNA_2230 (.A(net551));
 sg13g2_antennanp ANTENNA_2231 (.A(net551));
 sg13g2_antennanp ANTENNA_2232 (.A(net551));
 sg13g2_antennanp ANTENNA_2233 (.A(net551));
 sg13g2_antennanp ANTENNA_2234 (.A(net551));
 sg13g2_antennanp ANTENNA_2235 (.A(net551));
 sg13g2_antennanp ANTENNA_2236 (.A(net551));
 sg13g2_antennanp ANTENNA_2237 (.A(net551));
 sg13g2_antennanp ANTENNA_2238 (.A(net551));
 sg13g2_antennanp ANTENNA_2239 (.A(net551));
 sg13g2_antennanp ANTENNA_2240 (.A(net551));
 sg13g2_antennanp ANTENNA_2241 (.A(net551));
 sg13g2_antennanp ANTENNA_2242 (.A(net551));
 sg13g2_antennanp ANTENNA_2243 (.A(net551));
 sg13g2_antennanp ANTENNA_2244 (.A(net551));
 sg13g2_antennanp ANTENNA_2245 (.A(net551));
 sg13g2_antennanp ANTENNA_2246 (.A(net551));
 sg13g2_antennanp ANTENNA_2247 (.A(net551));
 sg13g2_antennanp ANTENNA_2248 (.A(net551));
 sg13g2_antennanp ANTENNA_2249 (.A(net551));
 sg13g2_antennanp ANTENNA_2250 (.A(net599));
 sg13g2_antennanp ANTENNA_2251 (.A(net599));
 sg13g2_antennanp ANTENNA_2252 (.A(net599));
 sg13g2_antennanp ANTENNA_2253 (.A(net599));
 sg13g2_antennanp ANTENNA_2254 (.A(net599));
 sg13g2_antennanp ANTENNA_2255 (.A(net599));
 sg13g2_antennanp ANTENNA_2256 (.A(net599));
 sg13g2_antennanp ANTENNA_2257 (.A(net599));
 sg13g2_antennanp ANTENNA_2258 (.A(net613));
 sg13g2_antennanp ANTENNA_2259 (.A(net613));
 sg13g2_antennanp ANTENNA_2260 (.A(net613));
 sg13g2_antennanp ANTENNA_2261 (.A(net613));
 sg13g2_antennanp ANTENNA_2262 (.A(net613));
 sg13g2_antennanp ANTENNA_2263 (.A(net613));
 sg13g2_antennanp ANTENNA_2264 (.A(net613));
 sg13g2_antennanp ANTENNA_2265 (.A(net613));
 sg13g2_antennanp ANTENNA_2266 (.A(net613));
 sg13g2_antennanp ANTENNA_2267 (.A(net613));
 sg13g2_antennanp ANTENNA_2268 (.A(net613));
 sg13g2_antennanp ANTENNA_2269 (.A(net613));
 sg13g2_antennanp ANTENNA_2270 (.A(net613));
 sg13g2_antennanp ANTENNA_2271 (.A(net613));
 sg13g2_antennanp ANTENNA_2272 (.A(net613));
 sg13g2_antennanp ANTENNA_2273 (.A(net682));
 sg13g2_antennanp ANTENNA_2274 (.A(net682));
 sg13g2_antennanp ANTENNA_2275 (.A(net682));
 sg13g2_antennanp ANTENNA_2276 (.A(net682));
 sg13g2_antennanp ANTENNA_2277 (.A(net682));
 sg13g2_antennanp ANTENNA_2278 (.A(net682));
 sg13g2_antennanp ANTENNA_2279 (.A(net682));
 sg13g2_antennanp ANTENNA_2280 (.A(net682));
 sg13g2_antennanp ANTENNA_2281 (.A(net682));
 sg13g2_antennanp ANTENNA_2282 (.A(net696));
 sg13g2_antennanp ANTENNA_2283 (.A(net696));
 sg13g2_antennanp ANTENNA_2284 (.A(net696));
 sg13g2_antennanp ANTENNA_2285 (.A(net696));
 sg13g2_antennanp ANTENNA_2286 (.A(net696));
 sg13g2_antennanp ANTENNA_2287 (.A(net696));
 sg13g2_antennanp ANTENNA_2288 (.A(net696));
 sg13g2_antennanp ANTENNA_2289 (.A(net696));
 sg13g2_antennanp ANTENNA_2290 (.A(net696));
 sg13g2_antennanp ANTENNA_2291 (.A(net802));
 sg13g2_antennanp ANTENNA_2292 (.A(net802));
 sg13g2_antennanp ANTENNA_2293 (.A(net802));
 sg13g2_antennanp ANTENNA_2294 (.A(net802));
 sg13g2_antennanp ANTENNA_2295 (.A(net802));
 sg13g2_antennanp ANTENNA_2296 (.A(net802));
 sg13g2_antennanp ANTENNA_2297 (.A(net802));
 sg13g2_antennanp ANTENNA_2298 (.A(net802));
 sg13g2_antennanp ANTENNA_2299 (.A(net802));
 sg13g2_antennanp ANTENNA_2300 (.A(net850));
 sg13g2_antennanp ANTENNA_2301 (.A(net850));
 sg13g2_antennanp ANTENNA_2302 (.A(net850));
 sg13g2_antennanp ANTENNA_2303 (.A(net850));
 sg13g2_antennanp ANTENNA_2304 (.A(net850));
 sg13g2_antennanp ANTENNA_2305 (.A(net850));
 sg13g2_antennanp ANTENNA_2306 (.A(net850));
 sg13g2_antennanp ANTENNA_2307 (.A(net850));
 sg13g2_antennanp ANTENNA_2308 (.A(net850));
 sg13g2_antennanp ANTENNA_2309 (.A(net974));
 sg13g2_antennanp ANTENNA_2310 (.A(net974));
 sg13g2_antennanp ANTENNA_2311 (.A(net974));
 sg13g2_antennanp ANTENNA_2312 (.A(net974));
 sg13g2_antennanp ANTENNA_2313 (.A(net974));
 sg13g2_antennanp ANTENNA_2314 (.A(net974));
 sg13g2_antennanp ANTENNA_2315 (.A(net974));
 sg13g2_antennanp ANTENNA_2316 (.A(net974));
 sg13g2_antennanp ANTENNA_2317 (.A(net974));
 sg13g2_antennanp ANTENNA_2318 (.A(net977));
 sg13g2_antennanp ANTENNA_2319 (.A(net977));
 sg13g2_antennanp ANTENNA_2320 (.A(net977));
 sg13g2_antennanp ANTENNA_2321 (.A(net977));
 sg13g2_antennanp ANTENNA_2322 (.A(net977));
 sg13g2_antennanp ANTENNA_2323 (.A(net977));
 sg13g2_antennanp ANTENNA_2324 (.A(net977));
 sg13g2_antennanp ANTENNA_2325 (.A(net977));
 sg13g2_antennanp ANTENNA_2326 (.A(net977));
 sg13g2_antennanp ANTENNA_2327 (.A(net1008));
 sg13g2_antennanp ANTENNA_2328 (.A(net1008));
 sg13g2_antennanp ANTENNA_2329 (.A(net1008));
 sg13g2_antennanp ANTENNA_2330 (.A(net1008));
 sg13g2_antennanp ANTENNA_2331 (.A(net1008));
 sg13g2_antennanp ANTENNA_2332 (.A(net1008));
 sg13g2_antennanp ANTENNA_2333 (.A(net1008));
 sg13g2_antennanp ANTENNA_2334 (.A(net1008));
 sg13g2_antennanp ANTENNA_2335 (.A(net1008));
 sg13g2_antennanp ANTENNA_2336 (.A(net1008));
 sg13g2_antennanp ANTENNA_2337 (.A(net1008));
 sg13g2_antennanp ANTENNA_2338 (.A(net1008));
 sg13g2_antennanp ANTENNA_2339 (.A(net1008));
 sg13g2_antennanp ANTENNA_2340 (.A(net1008));
 sg13g2_antennanp ANTENNA_2341 (.A(net1008));
 sg13g2_antennanp ANTENNA_2342 (.A(net1008));
 sg13g2_antennanp ANTENNA_2343 (.A(net1053));
 sg13g2_antennanp ANTENNA_2344 (.A(net1053));
 sg13g2_antennanp ANTENNA_2345 (.A(net1053));
 sg13g2_antennanp ANTENNA_2346 (.A(net1053));
 sg13g2_antennanp ANTENNA_2347 (.A(net1053));
 sg13g2_antennanp ANTENNA_2348 (.A(net1053));
 sg13g2_antennanp ANTENNA_2349 (.A(net1053));
 sg13g2_antennanp ANTENNA_2350 (.A(net1053));
 sg13g2_antennanp ANTENNA_2351 (.A(net1058));
 sg13g2_antennanp ANTENNA_2352 (.A(net1058));
 sg13g2_antennanp ANTENNA_2353 (.A(net1058));
 sg13g2_antennanp ANTENNA_2354 (.A(net1058));
 sg13g2_antennanp ANTENNA_2355 (.A(net1058));
 sg13g2_antennanp ANTENNA_2356 (.A(net1058));
 sg13g2_antennanp ANTENNA_2357 (.A(net1058));
 sg13g2_antennanp ANTENNA_2358 (.A(net1058));
 sg13g2_antennanp ANTENNA_2359 (.A(net1058));
 sg13g2_antennanp ANTENNA_2360 (.A(net1058));
 sg13g2_antennanp ANTENNA_2361 (.A(net1058));
 sg13g2_antennanp ANTENNA_2362 (.A(net1058));
 sg13g2_antennanp ANTENNA_2363 (.A(net1058));
 sg13g2_antennanp ANTENNA_2364 (.A(net1058));
 sg13g2_antennanp ANTENNA_2365 (.A(net1058));
 sg13g2_antennanp ANTENNA_2366 (.A(_00209_));
 sg13g2_antennanp ANTENNA_2367 (.A(_00209_));
 sg13g2_antennanp ANTENNA_2368 (.A(_00784_));
 sg13g2_antennanp ANTENNA_2369 (.A(_00784_));
 sg13g2_antennanp ANTENNA_2370 (.A(_00923_));
 sg13g2_antennanp ANTENNA_2371 (.A(_01034_));
 sg13g2_antennanp ANTENNA_2372 (.A(_02779_));
 sg13g2_antennanp ANTENNA_2373 (.A(_02779_));
 sg13g2_antennanp ANTENNA_2374 (.A(_02779_));
 sg13g2_antennanp ANTENNA_2375 (.A(_02779_));
 sg13g2_antennanp ANTENNA_2376 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2377 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2378 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2379 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2380 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2381 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2382 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2383 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2384 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2385 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2386 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2387 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2388 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2389 (.A(_02910_));
 sg13g2_antennanp ANTENNA_2390 (.A(_03478_));
 sg13g2_antennanp ANTENNA_2391 (.A(_03478_));
 sg13g2_antennanp ANTENNA_2392 (.A(_03478_));
 sg13g2_antennanp ANTENNA_2393 (.A(_03478_));
 sg13g2_antennanp ANTENNA_2394 (.A(_03527_));
 sg13g2_antennanp ANTENNA_2395 (.A(_03527_));
 sg13g2_antennanp ANTENNA_2396 (.A(_03527_));
 sg13g2_antennanp ANTENNA_2397 (.A(_03527_));
 sg13g2_antennanp ANTENNA_2398 (.A(_04734_));
 sg13g2_antennanp ANTENNA_2399 (.A(_04734_));
 sg13g2_antennanp ANTENNA_2400 (.A(_04734_));
 sg13g2_antennanp ANTENNA_2401 (.A(_04734_));
 sg13g2_antennanp ANTENNA_2402 (.A(_04751_));
 sg13g2_antennanp ANTENNA_2403 (.A(_04751_));
 sg13g2_antennanp ANTENNA_2404 (.A(_04775_));
 sg13g2_antennanp ANTENNA_2405 (.A(_04775_));
 sg13g2_antennanp ANTENNA_2406 (.A(_04778_));
 sg13g2_antennanp ANTENNA_2407 (.A(_04778_));
 sg13g2_antennanp ANTENNA_2408 (.A(_04778_));
 sg13g2_antennanp ANTENNA_2409 (.A(_04778_));
 sg13g2_antennanp ANTENNA_2410 (.A(_04927_));
 sg13g2_antennanp ANTENNA_2411 (.A(_04985_));
 sg13g2_antennanp ANTENNA_2412 (.A(_04985_));
 sg13g2_antennanp ANTENNA_2413 (.A(_05090_));
 sg13g2_antennanp ANTENNA_2414 (.A(_05090_));
 sg13g2_antennanp ANTENNA_2415 (.A(_05126_));
 sg13g2_antennanp ANTENNA_2416 (.A(_05149_));
 sg13g2_antennanp ANTENNA_2417 (.A(_05160_));
 sg13g2_antennanp ANTENNA_2418 (.A(_05174_));
 sg13g2_antennanp ANTENNA_2419 (.A(_05201_));
 sg13g2_antennanp ANTENNA_2420 (.A(_05215_));
 sg13g2_antennanp ANTENNA_2421 (.A(_05309_));
 sg13g2_antennanp ANTENNA_2422 (.A(_05583_));
 sg13g2_antennanp ANTENNA_2423 (.A(_05653_));
 sg13g2_antennanp ANTENNA_2424 (.A(_05667_));
 sg13g2_antennanp ANTENNA_2425 (.A(_05667_));
 sg13g2_antennanp ANTENNA_2426 (.A(_05669_));
 sg13g2_antennanp ANTENNA_2427 (.A(_05680_));
 sg13g2_antennanp ANTENNA_2428 (.A(_05700_));
 sg13g2_antennanp ANTENNA_2429 (.A(_05706_));
 sg13g2_antennanp ANTENNA_2430 (.A(_05712_));
 sg13g2_antennanp ANTENNA_2431 (.A(_05724_));
 sg13g2_antennanp ANTENNA_2432 (.A(_05895_));
 sg13g2_antennanp ANTENNA_2433 (.A(_05895_));
 sg13g2_antennanp ANTENNA_2434 (.A(_05895_));
 sg13g2_antennanp ANTENNA_2435 (.A(_05895_));
 sg13g2_antennanp ANTENNA_2436 (.A(_05895_));
 sg13g2_antennanp ANTENNA_2437 (.A(_05955_));
 sg13g2_antennanp ANTENNA_2438 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2439 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2440 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2441 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2442 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2443 (.A(_06556_));
 sg13g2_antennanp ANTENNA_2444 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2445 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2446 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2447 (.A(_06818_));
 sg13g2_antennanp ANTENNA_2448 (.A(_07576_));
 sg13g2_antennanp ANTENNA_2449 (.A(_07576_));
 sg13g2_antennanp ANTENNA_2450 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2451 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2452 (.A(_07877_));
 sg13g2_antennanp ANTENNA_2453 (.A(_08204_));
 sg13g2_antennanp ANTENNA_2454 (.A(_08204_));
 sg13g2_antennanp ANTENNA_2455 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2456 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2457 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2458 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2459 (.A(_08408_));
 sg13g2_antennanp ANTENNA_2460 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2461 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2462 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2463 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2464 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2465 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2466 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2467 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2468 (.A(_08439_));
 sg13g2_antennanp ANTENNA_2469 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2470 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2471 (.A(_08507_));
 sg13g2_antennanp ANTENNA_2472 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2473 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2474 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2475 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2476 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2477 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2478 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2479 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2480 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2481 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2482 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2483 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2484 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2485 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2486 (.A(_08798_));
 sg13g2_antennanp ANTENNA_2487 (.A(_08818_));
 sg13g2_antennanp ANTENNA_2488 (.A(_08840_));
 sg13g2_antennanp ANTENNA_2489 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2490 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2491 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2492 (.A(_08851_));
 sg13g2_antennanp ANTENNA_2493 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2494 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2495 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2496 (.A(_08868_));
 sg13g2_antennanp ANTENNA_2497 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2498 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2499 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2500 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2501 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2502 (.A(_09084_));
 sg13g2_antennanp ANTENNA_2503 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2504 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2505 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2506 (.A(_09131_));
 sg13g2_antennanp ANTENNA_2507 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2508 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2509 (.A(_09140_));
 sg13g2_antennanp ANTENNA_2510 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2511 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2512 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2513 (.A(_09141_));
 sg13g2_antennanp ANTENNA_2514 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2515 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2516 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2517 (.A(_09149_));
 sg13g2_antennanp ANTENNA_2518 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2519 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2520 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2521 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2522 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2523 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2524 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2525 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2526 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2527 (.A(_09150_));
 sg13g2_antennanp ANTENNA_2528 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2529 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2530 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2531 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2532 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2533 (.A(_09163_));
 sg13g2_antennanp ANTENNA_2534 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2535 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2536 (.A(_09230_));
 sg13g2_antennanp ANTENNA_2537 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2538 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2539 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2540 (.A(_09254_));
 sg13g2_antennanp ANTENNA_2541 (.A(_09306_));
 sg13g2_antennanp ANTENNA_2542 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2543 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2544 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2545 (.A(_09426_));
 sg13g2_antennanp ANTENNA_2546 (.A(_09436_));
 sg13g2_antennanp ANTENNA_2547 (.A(_09437_));
 sg13g2_antennanp ANTENNA_2548 (.A(_09437_));
 sg13g2_antennanp ANTENNA_2549 (.A(_09445_));
 sg13g2_antennanp ANTENNA_2550 (.A(_09498_));
 sg13g2_antennanp ANTENNA_2551 (.A(_09499_));
 sg13g2_antennanp ANTENNA_2552 (.A(_09499_));
 sg13g2_antennanp ANTENNA_2553 (.A(_09505_));
 sg13g2_antennanp ANTENNA_2554 (.A(_09531_));
 sg13g2_antennanp ANTENNA_2555 (.A(_09587_));
 sg13g2_antennanp ANTENNA_2556 (.A(_09615_));
 sg13g2_antennanp ANTENNA_2557 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2558 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2559 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2560 (.A(_09907_));
 sg13g2_antennanp ANTENNA_2561 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2562 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2563 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2564 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2565 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2566 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2567 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2568 (.A(_10113_));
 sg13g2_antennanp ANTENNA_2569 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2570 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2571 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2572 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2573 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2574 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2575 (.A(_10330_));
 sg13g2_antennanp ANTENNA_2576 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2577 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2578 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2579 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2580 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2581 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2582 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2583 (.A(_10368_));
 sg13g2_antennanp ANTENNA_2584 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2585 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2586 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2587 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2588 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2589 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2590 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2591 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2592 (.A(_10458_));
 sg13g2_antennanp ANTENNA_2593 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2594 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2595 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2596 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2597 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2598 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2599 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2600 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2601 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2602 (.A(_10478_));
 sg13g2_antennanp ANTENNA_2603 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2604 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2605 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2606 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2607 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2608 (.A(_10634_));
 sg13g2_antennanp ANTENNA_2609 (.A(_10779_));
 sg13g2_antennanp ANTENNA_2610 (.A(_11210_));
 sg13g2_antennanp ANTENNA_2611 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2612 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2613 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2614 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2615 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2616 (.A(_11776_));
 sg13g2_antennanp ANTENNA_2617 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2618 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2619 (.A(_11919_));
 sg13g2_antennanp ANTENNA_2620 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2621 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2622 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2623 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2624 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2625 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2626 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2627 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2628 (.A(_11926_));
 sg13g2_antennanp ANTENNA_2629 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2630 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2631 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2632 (.A(_11960_));
 sg13g2_antennanp ANTENNA_2633 (.A(clk));
 sg13g2_antennanp ANTENNA_2634 (.A(clk));
 sg13g2_antennanp ANTENNA_2635 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2636 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2637 (.A(\cpu.ex.r_mult[30] ));
 sg13g2_antennanp ANTENNA_2638 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2639 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2640 (.A(net4));
 sg13g2_antennanp ANTENNA_2641 (.A(net4));
 sg13g2_antennanp ANTENNA_2642 (.A(net4));
 sg13g2_antennanp ANTENNA_2643 (.A(net12));
 sg13g2_antennanp ANTENNA_2644 (.A(net12));
 sg13g2_antennanp ANTENNA_2645 (.A(net12));
 sg13g2_antennanp ANTENNA_2646 (.A(net13));
 sg13g2_antennanp ANTENNA_2647 (.A(net13));
 sg13g2_antennanp ANTENNA_2648 (.A(net13));
 sg13g2_antennanp ANTENNA_2649 (.A(net14));
 sg13g2_antennanp ANTENNA_2650 (.A(net14));
 sg13g2_antennanp ANTENNA_2651 (.A(net14));
 sg13g2_antennanp ANTENNA_2652 (.A(net506));
 sg13g2_antennanp ANTENNA_2653 (.A(net506));
 sg13g2_antennanp ANTENNA_2654 (.A(net506));
 sg13g2_antennanp ANTENNA_2655 (.A(net506));
 sg13g2_antennanp ANTENNA_2656 (.A(net506));
 sg13g2_antennanp ANTENNA_2657 (.A(net506));
 sg13g2_antennanp ANTENNA_2658 (.A(net506));
 sg13g2_antennanp ANTENNA_2659 (.A(net506));
 sg13g2_antennanp ANTENNA_2660 (.A(net507));
 sg13g2_antennanp ANTENNA_2661 (.A(net507));
 sg13g2_antennanp ANTENNA_2662 (.A(net507));
 sg13g2_antennanp ANTENNA_2663 (.A(net507));
 sg13g2_antennanp ANTENNA_2664 (.A(net507));
 sg13g2_antennanp ANTENNA_2665 (.A(net507));
 sg13g2_antennanp ANTENNA_2666 (.A(net507));
 sg13g2_antennanp ANTENNA_2667 (.A(net507));
 sg13g2_antennanp ANTENNA_2668 (.A(net507));
 sg13g2_antennanp ANTENNA_2669 (.A(net507));
 sg13g2_antennanp ANTENNA_2670 (.A(net507));
 sg13g2_antennanp ANTENNA_2671 (.A(net507));
 sg13g2_antennanp ANTENNA_2672 (.A(net507));
 sg13g2_antennanp ANTENNA_2673 (.A(net507));
 sg13g2_antennanp ANTENNA_2674 (.A(net507));
 sg13g2_antennanp ANTENNA_2675 (.A(net507));
 sg13g2_antennanp ANTENNA_2676 (.A(net507));
 sg13g2_antennanp ANTENNA_2677 (.A(net507));
 sg13g2_antennanp ANTENNA_2678 (.A(net507));
 sg13g2_antennanp ANTENNA_2679 (.A(net507));
 sg13g2_antennanp ANTENNA_2680 (.A(net507));
 sg13g2_antennanp ANTENNA_2681 (.A(net507));
 sg13g2_antennanp ANTENNA_2682 (.A(net507));
 sg13g2_antennanp ANTENNA_2683 (.A(net551));
 sg13g2_antennanp ANTENNA_2684 (.A(net551));
 sg13g2_antennanp ANTENNA_2685 (.A(net551));
 sg13g2_antennanp ANTENNA_2686 (.A(net551));
 sg13g2_antennanp ANTENNA_2687 (.A(net551));
 sg13g2_antennanp ANTENNA_2688 (.A(net551));
 sg13g2_antennanp ANTENNA_2689 (.A(net551));
 sg13g2_antennanp ANTENNA_2690 (.A(net551));
 sg13g2_antennanp ANTENNA_2691 (.A(net551));
 sg13g2_antennanp ANTENNA_2692 (.A(net551));
 sg13g2_antennanp ANTENNA_2693 (.A(net551));
 sg13g2_antennanp ANTENNA_2694 (.A(net551));
 sg13g2_antennanp ANTENNA_2695 (.A(net551));
 sg13g2_antennanp ANTENNA_2696 (.A(net551));
 sg13g2_antennanp ANTENNA_2697 (.A(net551));
 sg13g2_antennanp ANTENNA_2698 (.A(net551));
 sg13g2_antennanp ANTENNA_2699 (.A(net551));
 sg13g2_antennanp ANTENNA_2700 (.A(net551));
 sg13g2_antennanp ANTENNA_2701 (.A(net551));
 sg13g2_antennanp ANTENNA_2702 (.A(net551));
 sg13g2_antennanp ANTENNA_2703 (.A(net551));
 sg13g2_antennanp ANTENNA_2704 (.A(net551));
 sg13g2_antennanp ANTENNA_2705 (.A(net551));
 sg13g2_antennanp ANTENNA_2706 (.A(net551));
 sg13g2_antennanp ANTENNA_2707 (.A(net613));
 sg13g2_antennanp ANTENNA_2708 (.A(net613));
 sg13g2_antennanp ANTENNA_2709 (.A(net613));
 sg13g2_antennanp ANTENNA_2710 (.A(net613));
 sg13g2_antennanp ANTENNA_2711 (.A(net613));
 sg13g2_antennanp ANTENNA_2712 (.A(net613));
 sg13g2_antennanp ANTENNA_2713 (.A(net613));
 sg13g2_antennanp ANTENNA_2714 (.A(net613));
 sg13g2_antennanp ANTENNA_2715 (.A(net613));
 sg13g2_antennanp ANTENNA_2716 (.A(net613));
 sg13g2_antennanp ANTENNA_2717 (.A(net613));
 sg13g2_antennanp ANTENNA_2718 (.A(net613));
 sg13g2_antennanp ANTENNA_2719 (.A(net613));
 sg13g2_antennanp ANTENNA_2720 (.A(net613));
 sg13g2_antennanp ANTENNA_2721 (.A(net613));
 sg13g2_antennanp ANTENNA_2722 (.A(net682));
 sg13g2_antennanp ANTENNA_2723 (.A(net682));
 sg13g2_antennanp ANTENNA_2724 (.A(net682));
 sg13g2_antennanp ANTENNA_2725 (.A(net682));
 sg13g2_antennanp ANTENNA_2726 (.A(net682));
 sg13g2_antennanp ANTENNA_2727 (.A(net682));
 sg13g2_antennanp ANTENNA_2728 (.A(net682));
 sg13g2_antennanp ANTENNA_2729 (.A(net682));
 sg13g2_antennanp ANTENNA_2730 (.A(net682));
 sg13g2_antennanp ANTENNA_2731 (.A(net696));
 sg13g2_antennanp ANTENNA_2732 (.A(net696));
 sg13g2_antennanp ANTENNA_2733 (.A(net696));
 sg13g2_antennanp ANTENNA_2734 (.A(net696));
 sg13g2_antennanp ANTENNA_2735 (.A(net696));
 sg13g2_antennanp ANTENNA_2736 (.A(net696));
 sg13g2_antennanp ANTENNA_2737 (.A(net696));
 sg13g2_antennanp ANTENNA_2738 (.A(net696));
 sg13g2_antennanp ANTENNA_2739 (.A(net696));
 sg13g2_antennanp ANTENNA_2740 (.A(net802));
 sg13g2_antennanp ANTENNA_2741 (.A(net802));
 sg13g2_antennanp ANTENNA_2742 (.A(net802));
 sg13g2_antennanp ANTENNA_2743 (.A(net802));
 sg13g2_antennanp ANTENNA_2744 (.A(net802));
 sg13g2_antennanp ANTENNA_2745 (.A(net802));
 sg13g2_antennanp ANTENNA_2746 (.A(net802));
 sg13g2_antennanp ANTENNA_2747 (.A(net802));
 sg13g2_antennanp ANTENNA_2748 (.A(net802));
 sg13g2_antennanp ANTENNA_2749 (.A(net850));
 sg13g2_antennanp ANTENNA_2750 (.A(net850));
 sg13g2_antennanp ANTENNA_2751 (.A(net850));
 sg13g2_antennanp ANTENNA_2752 (.A(net850));
 sg13g2_antennanp ANTENNA_2753 (.A(net850));
 sg13g2_antennanp ANTENNA_2754 (.A(net850));
 sg13g2_antennanp ANTENNA_2755 (.A(net850));
 sg13g2_antennanp ANTENNA_2756 (.A(net850));
 sg13g2_antennanp ANTENNA_2757 (.A(net850));
 sg13g2_antennanp ANTENNA_2758 (.A(net977));
 sg13g2_antennanp ANTENNA_2759 (.A(net977));
 sg13g2_antennanp ANTENNA_2760 (.A(net977));
 sg13g2_antennanp ANTENNA_2761 (.A(net977));
 sg13g2_antennanp ANTENNA_2762 (.A(net977));
 sg13g2_antennanp ANTENNA_2763 (.A(net977));
 sg13g2_antennanp ANTENNA_2764 (.A(net977));
 sg13g2_antennanp ANTENNA_2765 (.A(net977));
 sg13g2_antennanp ANTENNA_2766 (.A(net977));
 sg13g2_antennanp ANTENNA_2767 (.A(net1008));
 sg13g2_antennanp ANTENNA_2768 (.A(net1008));
 sg13g2_antennanp ANTENNA_2769 (.A(net1008));
 sg13g2_antennanp ANTENNA_2770 (.A(net1008));
 sg13g2_antennanp ANTENNA_2771 (.A(net1008));
 sg13g2_antennanp ANTENNA_2772 (.A(net1008));
 sg13g2_antennanp ANTENNA_2773 (.A(net1008));
 sg13g2_antennanp ANTENNA_2774 (.A(net1008));
 sg13g2_antennanp ANTENNA_2775 (.A(net1008));
 sg13g2_antennanp ANTENNA_2776 (.A(net1008));
 sg13g2_antennanp ANTENNA_2777 (.A(net1008));
 sg13g2_antennanp ANTENNA_2778 (.A(net1008));
 sg13g2_antennanp ANTENNA_2779 (.A(net1008));
 sg13g2_antennanp ANTENNA_2780 (.A(net1008));
 sg13g2_antennanp ANTENNA_2781 (.A(net1008));
 sg13g2_antennanp ANTENNA_2782 (.A(net1008));
 sg13g2_antennanp ANTENNA_2783 (.A(net1008));
 sg13g2_antennanp ANTENNA_2784 (.A(net1008));
 sg13g2_antennanp ANTENNA_2785 (.A(net1008));
 sg13g2_antennanp ANTENNA_2786 (.A(net1008));
 sg13g2_antennanp ANTENNA_2787 (.A(net1008));
 sg13g2_antennanp ANTENNA_2788 (.A(net1008));
 sg13g2_antennanp ANTENNA_2789 (.A(net1008));
 sg13g2_antennanp ANTENNA_2790 (.A(net1008));
 sg13g2_antennanp ANTENNA_2791 (.A(net1015));
 sg13g2_antennanp ANTENNA_2792 (.A(net1015));
 sg13g2_antennanp ANTENNA_2793 (.A(net1015));
 sg13g2_antennanp ANTENNA_2794 (.A(net1015));
 sg13g2_antennanp ANTENNA_2795 (.A(net1015));
 sg13g2_antennanp ANTENNA_2796 (.A(net1015));
 sg13g2_antennanp ANTENNA_2797 (.A(net1015));
 sg13g2_antennanp ANTENNA_2798 (.A(net1015));
 sg13g2_antennanp ANTENNA_2799 (.A(net1015));
 sg13g2_antennanp ANTENNA_2800 (.A(net1015));
 sg13g2_antennanp ANTENNA_2801 (.A(net1015));
 sg13g2_antennanp ANTENNA_2802 (.A(net1015));
 sg13g2_antennanp ANTENNA_2803 (.A(net1015));
 sg13g2_antennanp ANTENNA_2804 (.A(net1015));
 sg13g2_antennanp ANTENNA_2805 (.A(net1015));
 sg13g2_antennanp ANTENNA_2806 (.A(net1015));
 sg13g2_antennanp ANTENNA_2807 (.A(net1053));
 sg13g2_antennanp ANTENNA_2808 (.A(net1053));
 sg13g2_antennanp ANTENNA_2809 (.A(net1053));
 sg13g2_antennanp ANTENNA_2810 (.A(net1053));
 sg13g2_antennanp ANTENNA_2811 (.A(net1053));
 sg13g2_antennanp ANTENNA_2812 (.A(net1053));
 sg13g2_antennanp ANTENNA_2813 (.A(net1053));
 sg13g2_antennanp ANTENNA_2814 (.A(net1053));
 sg13g2_antennanp ANTENNA_2815 (.A(net1053));
 sg13g2_antennanp ANTENNA_2816 (.A(net1058));
 sg13g2_antennanp ANTENNA_2817 (.A(net1058));
 sg13g2_antennanp ANTENNA_2818 (.A(net1058));
 sg13g2_antennanp ANTENNA_2819 (.A(net1058));
 sg13g2_antennanp ANTENNA_2820 (.A(net1058));
 sg13g2_antennanp ANTENNA_2821 (.A(net1058));
 sg13g2_antennanp ANTENNA_2822 (.A(net1058));
 sg13g2_antennanp ANTENNA_2823 (.A(net1058));
 sg13g2_antennanp ANTENNA_2824 (.A(net1058));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_4 FILLER_0_42 ();
 sg13g2_fill_2 FILLER_0_46 ();
 sg13g2_fill_2 FILLER_0_53 ();
 sg13g2_fill_2 FILLER_0_64 ();
 sg13g2_fill_1 FILLER_0_66 ();
 sg13g2_decap_8 FILLER_0_96 ();
 sg13g2_decap_8 FILLER_0_103 ();
 sg13g2_fill_2 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_138 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_decap_8 FILLER_0_213 ();
 sg13g2_decap_8 FILLER_0_220 ();
 sg13g2_fill_1 FILLER_0_227 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_fill_1 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_fill_2 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_4 FILLER_0_389 ();
 sg13g2_fill_2 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_decap_4 FILLER_0_432 ();
 sg13g2_decap_8 FILLER_0_440 ();
 sg13g2_fill_2 FILLER_0_473 ();
 sg13g2_fill_2 FILLER_0_479 ();
 sg13g2_fill_2 FILLER_0_507 ();
 sg13g2_fill_1 FILLER_0_509 ();
 sg13g2_decap_8 FILLER_0_514 ();
 sg13g2_decap_8 FILLER_0_521 ();
 sg13g2_decap_8 FILLER_0_528 ();
 sg13g2_decap_8 FILLER_0_535 ();
 sg13g2_decap_8 FILLER_0_542 ();
 sg13g2_decap_8 FILLER_0_549 ();
 sg13g2_decap_8 FILLER_0_556 ();
 sg13g2_fill_2 FILLER_0_563 ();
 sg13g2_decap_8 FILLER_0_612 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_4 FILLER_0_626 ();
 sg13g2_fill_1 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_fill_2 FILLER_0_671 ();
 sg13g2_fill_1 FILLER_0_673 ();
 sg13g2_fill_1 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_705 ();
 sg13g2_fill_2 FILLER_0_712 ();
 sg13g2_fill_1 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_719 ();
 sg13g2_decap_8 FILLER_0_726 ();
 sg13g2_decap_8 FILLER_0_733 ();
 sg13g2_decap_8 FILLER_0_740 ();
 sg13g2_fill_1 FILLER_0_747 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_fill_1 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_771 ();
 sg13g2_decap_8 FILLER_0_778 ();
 sg13g2_decap_8 FILLER_0_785 ();
 sg13g2_decap_8 FILLER_0_792 ();
 sg13g2_decap_8 FILLER_0_799 ();
 sg13g2_decap_8 FILLER_0_806 ();
 sg13g2_decap_8 FILLER_0_813 ();
 sg13g2_decap_8 FILLER_0_820 ();
 sg13g2_decap_8 FILLER_0_827 ();
 sg13g2_decap_8 FILLER_0_860 ();
 sg13g2_decap_4 FILLER_0_867 ();
 sg13g2_fill_1 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_905 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_4 FILLER_0_926 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_4 FILLER_0_1003 ();
 sg13g2_fill_2 FILLER_0_1007 ();
 sg13g2_decap_8 FILLER_0_1035 ();
 sg13g2_decap_8 FILLER_0_1042 ();
 sg13g2_decap_8 FILLER_0_1049 ();
 sg13g2_decap_4 FILLER_0_1056 ();
 sg13g2_fill_2 FILLER_0_1060 ();
 sg13g2_decap_8 FILLER_0_1092 ();
 sg13g2_decap_4 FILLER_0_1099 ();
 sg13g2_fill_1 FILLER_0_1103 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_fill_1 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1164 ();
 sg13g2_decap_8 FILLER_0_1171 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_decap_8 FILLER_0_1211 ();
 sg13g2_decap_8 FILLER_0_1218 ();
 sg13g2_decap_8 FILLER_0_1225 ();
 sg13g2_fill_1 FILLER_0_1232 ();
 sg13g2_decap_8 FILLER_0_1237 ();
 sg13g2_fill_2 FILLER_0_1244 ();
 sg13g2_decap_8 FILLER_0_1272 ();
 sg13g2_decap_8 FILLER_0_1279 ();
 sg13g2_decap_8 FILLER_0_1312 ();
 sg13g2_decap_4 FILLER_0_1319 ();
 sg13g2_fill_1 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1350 ();
 sg13g2_decap_8 FILLER_0_1357 ();
 sg13g2_decap_8 FILLER_0_1364 ();
 sg13g2_decap_8 FILLER_0_1371 ();
 sg13g2_decap_8 FILLER_0_1378 ();
 sg13g2_decap_8 FILLER_0_1385 ();
 sg13g2_decap_4 FILLER_0_1392 ();
 sg13g2_fill_1 FILLER_0_1396 ();
 sg13g2_decap_8 FILLER_0_1411 ();
 sg13g2_decap_8 FILLER_0_1418 ();
 sg13g2_decap_8 FILLER_0_1425 ();
 sg13g2_decap_8 FILLER_0_1436 ();
 sg13g2_decap_8 FILLER_0_1443 ();
 sg13g2_decap_8 FILLER_0_1450 ();
 sg13g2_decap_8 FILLER_0_1457 ();
 sg13g2_decap_8 FILLER_0_1464 ();
 sg13g2_decap_8 FILLER_0_1471 ();
 sg13g2_decap_8 FILLER_0_1478 ();
 sg13g2_fill_2 FILLER_0_1485 ();
 sg13g2_fill_1 FILLER_0_1487 ();
 sg13g2_decap_8 FILLER_0_1514 ();
 sg13g2_decap_8 FILLER_0_1521 ();
 sg13g2_decap_8 FILLER_0_1528 ();
 sg13g2_fill_2 FILLER_0_1535 ();
 sg13g2_fill_1 FILLER_0_1537 ();
 sg13g2_decap_8 FILLER_0_1546 ();
 sg13g2_decap_8 FILLER_0_1553 ();
 sg13g2_decap_8 FILLER_0_1560 ();
 sg13g2_fill_2 FILLER_0_1567 ();
 sg13g2_decap_8 FILLER_0_1599 ();
 sg13g2_decap_8 FILLER_0_1606 ();
 sg13g2_decap_8 FILLER_0_1613 ();
 sg13g2_decap_8 FILLER_0_1620 ();
 sg13g2_fill_1 FILLER_0_1627 ();
 sg13g2_decap_8 FILLER_0_1684 ();
 sg13g2_decap_8 FILLER_0_1691 ();
 sg13g2_decap_8 FILLER_0_1698 ();
 sg13g2_decap_8 FILLER_0_1705 ();
 sg13g2_decap_8 FILLER_0_1712 ();
 sg13g2_decap_8 FILLER_0_1719 ();
 sg13g2_fill_2 FILLER_0_1726 ();
 sg13g2_decap_4 FILLER_0_1767 ();
 sg13g2_fill_1 FILLER_0_1771 ();
 sg13g2_decap_8 FILLER_0_1802 ();
 sg13g2_decap_8 FILLER_0_1809 ();
 sg13g2_decap_4 FILLER_0_1816 ();
 sg13g2_decap_4 FILLER_0_1846 ();
 sg13g2_fill_1 FILLER_0_1850 ();
 sg13g2_decap_8 FILLER_0_1877 ();
 sg13g2_decap_4 FILLER_0_1884 ();
 sg13g2_fill_1 FILLER_0_1888 ();
 sg13g2_decap_8 FILLER_0_1915 ();
 sg13g2_decap_8 FILLER_0_1922 ();
 sg13g2_decap_8 FILLER_0_1929 ();
 sg13g2_fill_2 FILLER_0_1936 ();
 sg13g2_fill_1 FILLER_0_1938 ();
 sg13g2_decap_8 FILLER_0_1969 ();
 sg13g2_decap_8 FILLER_0_1976 ();
 sg13g2_fill_2 FILLER_0_1983 ();
 sg13g2_decap_8 FILLER_0_2011 ();
 sg13g2_fill_1 FILLER_0_2018 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_decap_8 FILLER_0_2037 ();
 sg13g2_fill_2 FILLER_0_2044 ();
 sg13g2_decap_8 FILLER_0_2054 ();
 sg13g2_fill_2 FILLER_0_2061 ();
 sg13g2_fill_2 FILLER_0_2084 ();
 sg13g2_fill_1 FILLER_0_2086 ();
 sg13g2_fill_1 FILLER_0_2097 ();
 sg13g2_decap_8 FILLER_0_2102 ();
 sg13g2_decap_8 FILLER_0_2109 ();
 sg13g2_decap_8 FILLER_0_2116 ();
 sg13g2_decap_8 FILLER_0_2123 ();
 sg13g2_decap_8 FILLER_0_2130 ();
 sg13g2_fill_2 FILLER_0_2137 ();
 sg13g2_decap_8 FILLER_0_2147 ();
 sg13g2_decap_8 FILLER_0_2154 ();
 sg13g2_decap_8 FILLER_0_2161 ();
 sg13g2_decap_8 FILLER_0_2168 ();
 sg13g2_fill_1 FILLER_0_2175 ();
 sg13g2_decap_8 FILLER_0_2180 ();
 sg13g2_decap_8 FILLER_0_2187 ();
 sg13g2_decap_8 FILLER_0_2194 ();
 sg13g2_decap_8 FILLER_0_2201 ();
 sg13g2_fill_2 FILLER_0_2208 ();
 sg13g2_decap_8 FILLER_0_2214 ();
 sg13g2_decap_8 FILLER_0_2221 ();
 sg13g2_fill_1 FILLER_0_2228 ();
 sg13g2_decap_8 FILLER_0_2233 ();
 sg13g2_decap_8 FILLER_0_2240 ();
 sg13g2_decap_8 FILLER_0_2247 ();
 sg13g2_decap_8 FILLER_0_2254 ();
 sg13g2_decap_8 FILLER_0_2261 ();
 sg13g2_decap_8 FILLER_0_2268 ();
 sg13g2_decap_8 FILLER_0_2275 ();
 sg13g2_decap_8 FILLER_0_2282 ();
 sg13g2_decap_8 FILLER_0_2289 ();
 sg13g2_decap_8 FILLER_0_2296 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_8 FILLER_0_2310 ();
 sg13g2_decap_8 FILLER_0_2317 ();
 sg13g2_decap_8 FILLER_0_2324 ();
 sg13g2_decap_8 FILLER_0_2331 ();
 sg13g2_decap_8 FILLER_0_2338 ();
 sg13g2_decap_8 FILLER_0_2345 ();
 sg13g2_decap_8 FILLER_0_2352 ();
 sg13g2_decap_8 FILLER_0_2359 ();
 sg13g2_decap_4 FILLER_0_2366 ();
 sg13g2_fill_1 FILLER_0_2370 ();
 sg13g2_decap_8 FILLER_0_2400 ();
 sg13g2_fill_2 FILLER_0_2407 ();
 sg13g2_fill_1 FILLER_0_2409 ();
 sg13g2_decap_8 FILLER_0_2424 ();
 sg13g2_decap_8 FILLER_0_2431 ();
 sg13g2_decap_8 FILLER_0_2438 ();
 sg13g2_decap_8 FILLER_0_2445 ();
 sg13g2_decap_8 FILLER_0_2452 ();
 sg13g2_decap_8 FILLER_0_2459 ();
 sg13g2_fill_2 FILLER_0_2466 ();
 sg13g2_fill_1 FILLER_0_2468 ();
 sg13g2_decap_8 FILLER_0_2473 ();
 sg13g2_decap_8 FILLER_0_2480 ();
 sg13g2_decap_8 FILLER_0_2487 ();
 sg13g2_decap_8 FILLER_0_2494 ();
 sg13g2_decap_8 FILLER_0_2501 ();
 sg13g2_decap_8 FILLER_0_2508 ();
 sg13g2_decap_8 FILLER_0_2515 ();
 sg13g2_decap_8 FILLER_0_2522 ();
 sg13g2_decap_8 FILLER_0_2529 ();
 sg13g2_decap_8 FILLER_0_2536 ();
 sg13g2_decap_8 FILLER_0_2543 ();
 sg13g2_decap_8 FILLER_0_2550 ();
 sg13g2_decap_8 FILLER_0_2557 ();
 sg13g2_decap_8 FILLER_0_2564 ();
 sg13g2_decap_8 FILLER_0_2571 ();
 sg13g2_decap_8 FILLER_0_2578 ();
 sg13g2_decap_8 FILLER_0_2585 ();
 sg13g2_decap_8 FILLER_0_2592 ();
 sg13g2_decap_8 FILLER_0_2599 ();
 sg13g2_decap_8 FILLER_0_2606 ();
 sg13g2_decap_8 FILLER_0_2613 ();
 sg13g2_decap_8 FILLER_0_2620 ();
 sg13g2_decap_8 FILLER_0_2627 ();
 sg13g2_decap_8 FILLER_0_2634 ();
 sg13g2_decap_8 FILLER_0_2641 ();
 sg13g2_decap_8 FILLER_0_2648 ();
 sg13g2_decap_8 FILLER_0_2655 ();
 sg13g2_decap_8 FILLER_0_2662 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_51 ();
 sg13g2_fill_1 FILLER_1_63 ();
 sg13g2_fill_2 FILLER_1_86 ();
 sg13g2_fill_1 FILLER_1_88 ();
 sg13g2_decap_4 FILLER_1_123 ();
 sg13g2_fill_2 FILLER_1_127 ();
 sg13g2_fill_2 FILLER_1_159 ();
 sg13g2_fill_1 FILLER_1_161 ();
 sg13g2_decap_4 FILLER_1_172 ();
 sg13g2_fill_2 FILLER_1_176 ();
 sg13g2_fill_2 FILLER_1_204 ();
 sg13g2_decap_4 FILLER_1_230 ();
 sg13g2_fill_2 FILLER_1_234 ();
 sg13g2_decap_4 FILLER_1_240 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_4 FILLER_1_277 ();
 sg13g2_fill_1 FILLER_1_337 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_fill_2 FILLER_1_364 ();
 sg13g2_fill_2 FILLER_1_418 ();
 sg13g2_fill_1 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_451 ();
 sg13g2_fill_1 FILLER_1_458 ();
 sg13g2_fill_2 FILLER_1_477 ();
 sg13g2_fill_2 FILLER_1_524 ();
 sg13g2_decap_4 FILLER_1_530 ();
 sg13g2_fill_1 FILLER_1_560 ();
 sg13g2_fill_1 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_622 ();
 sg13g2_decap_8 FILLER_1_629 ();
 sg13g2_decap_4 FILLER_1_636 ();
 sg13g2_fill_1 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_fill_1 FILLER_1_685 ();
 sg13g2_decap_4 FILLER_1_689 ();
 sg13g2_fill_2 FILLER_1_693 ();
 sg13g2_fill_1 FILLER_1_699 ();
 sg13g2_fill_2 FILLER_1_705 ();
 sg13g2_fill_1 FILLER_1_707 ();
 sg13g2_decap_4 FILLER_1_734 ();
 sg13g2_fill_2 FILLER_1_738 ();
 sg13g2_fill_2 FILLER_1_779 ();
 sg13g2_decap_4 FILLER_1_791 ();
 sg13g2_fill_2 FILLER_1_795 ();
 sg13g2_fill_2 FILLER_1_806 ();
 sg13g2_decap_8 FILLER_1_834 ();
 sg13g2_fill_1 FILLER_1_841 ();
 sg13g2_decap_4 FILLER_1_872 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_fill_2 FILLER_1_923 ();
 sg13g2_fill_2 FILLER_1_955 ();
 sg13g2_fill_1 FILLER_1_957 ();
 sg13g2_fill_2 FILLER_1_984 ();
 sg13g2_fill_1 FILLER_1_986 ();
 sg13g2_fill_2 FILLER_1_1013 ();
 sg13g2_fill_1 FILLER_1_1015 ();
 sg13g2_fill_1 FILLER_1_1020 ();
 sg13g2_fill_2 FILLER_1_1056 ();
 sg13g2_fill_1 FILLER_1_1058 ();
 sg13g2_fill_1 FILLER_1_1067 ();
 sg13g2_fill_2 FILLER_1_1073 ();
 sg13g2_fill_1 FILLER_1_1075 ();
 sg13g2_fill_2 FILLER_1_1102 ();
 sg13g2_fill_1 FILLER_1_1138 ();
 sg13g2_decap_4 FILLER_1_1173 ();
 sg13g2_decap_4 FILLER_1_1211 ();
 sg13g2_fill_1 FILLER_1_1215 ();
 sg13g2_decap_8 FILLER_1_1279 ();
 sg13g2_decap_4 FILLER_1_1286 ();
 sg13g2_fill_1 FILLER_1_1290 ();
 sg13g2_fill_2 FILLER_1_1317 ();
 sg13g2_fill_1 FILLER_1_1357 ();
 sg13g2_fill_2 FILLER_1_1384 ();
 sg13g2_fill_1 FILLER_1_1396 ();
 sg13g2_fill_2 FILLER_1_1423 ();
 sg13g2_decap_4 FILLER_1_1451 ();
 sg13g2_fill_1 FILLER_1_1455 ();
 sg13g2_fill_2 FILLER_1_1460 ();
 sg13g2_fill_2 FILLER_1_1488 ();
 sg13g2_fill_1 FILLER_1_1490 ();
 sg13g2_fill_2 FILLER_1_1517 ();
 sg13g2_fill_2 FILLER_1_1529 ();
 sg13g2_fill_1 FILLER_1_1531 ();
 sg13g2_fill_1 FILLER_1_1558 ();
 sg13g2_fill_2 FILLER_1_1585 ();
 sg13g2_decap_8 FILLER_1_1607 ();
 sg13g2_decap_8 FILLER_1_1614 ();
 sg13g2_fill_2 FILLER_1_1621 ();
 sg13g2_fill_2 FILLER_1_1627 ();
 sg13g2_decap_8 FILLER_1_1639 ();
 sg13g2_decap_8 FILLER_1_1646 ();
 sg13g2_fill_2 FILLER_1_1657 ();
 sg13g2_fill_1 FILLER_1_1659 ();
 sg13g2_decap_8 FILLER_1_1670 ();
 sg13g2_fill_1 FILLER_1_1677 ();
 sg13g2_decap_8 FILLER_1_1714 ();
 sg13g2_decap_4 FILLER_1_1721 ();
 sg13g2_fill_2 FILLER_1_1751 ();
 sg13g2_fill_1 FILLER_1_1753 ();
 sg13g2_decap_8 FILLER_1_1786 ();
 sg13g2_decap_8 FILLER_1_1793 ();
 sg13g2_decap_8 FILLER_1_1800 ();
 sg13g2_fill_2 FILLER_1_1807 ();
 sg13g2_fill_1 FILLER_1_1839 ();
 sg13g2_decap_8 FILLER_1_1873 ();
 sg13g2_decap_4 FILLER_1_1880 ();
 sg13g2_decap_4 FILLER_1_1920 ();
 sg13g2_fill_2 FILLER_1_1924 ();
 sg13g2_decap_8 FILLER_1_1962 ();
 sg13g2_decap_4 FILLER_1_1969 ();
 sg13g2_fill_1 FILLER_1_1999 ();
 sg13g2_fill_2 FILLER_1_2036 ();
 sg13g2_fill_1 FILLER_1_2038 ();
 sg13g2_decap_8 FILLER_1_2065 ();
 sg13g2_fill_1 FILLER_1_2072 ();
 sg13g2_fill_1 FILLER_1_2113 ();
 sg13g2_fill_2 FILLER_1_2118 ();
 sg13g2_fill_2 FILLER_1_2130 ();
 sg13g2_fill_2 FILLER_1_2158 ();
 sg13g2_decap_8 FILLER_1_2196 ();
 sg13g2_fill_2 FILLER_1_2229 ();
 sg13g2_fill_1 FILLER_1_2231 ();
 sg13g2_decap_4 FILLER_1_2245 ();
 sg13g2_fill_1 FILLER_1_2249 ();
 sg13g2_decap_8 FILLER_1_2280 ();
 sg13g2_decap_8 FILLER_1_2287 ();
 sg13g2_decap_8 FILLER_1_2294 ();
 sg13g2_decap_8 FILLER_1_2301 ();
 sg13g2_decap_8 FILLER_1_2308 ();
 sg13g2_decap_8 FILLER_1_2315 ();
 sg13g2_decap_8 FILLER_1_2322 ();
 sg13g2_decap_8 FILLER_1_2329 ();
 sg13g2_decap_8 FILLER_1_2336 ();
 sg13g2_fill_2 FILLER_1_2343 ();
 sg13g2_decap_8 FILLER_1_2349 ();
 sg13g2_decap_4 FILLER_1_2356 ();
 sg13g2_fill_1 FILLER_1_2360 ();
 sg13g2_decap_4 FILLER_1_2453 ();
 sg13g2_fill_1 FILLER_1_2457 ();
 sg13g2_decap_8 FILLER_1_2488 ();
 sg13g2_decap_8 FILLER_1_2495 ();
 sg13g2_decap_8 FILLER_1_2502 ();
 sg13g2_decap_8 FILLER_1_2509 ();
 sg13g2_decap_8 FILLER_1_2516 ();
 sg13g2_decap_8 FILLER_1_2523 ();
 sg13g2_decap_8 FILLER_1_2530 ();
 sg13g2_decap_8 FILLER_1_2537 ();
 sg13g2_decap_8 FILLER_1_2544 ();
 sg13g2_decap_8 FILLER_1_2551 ();
 sg13g2_decap_8 FILLER_1_2558 ();
 sg13g2_decap_8 FILLER_1_2565 ();
 sg13g2_decap_8 FILLER_1_2572 ();
 sg13g2_decap_8 FILLER_1_2579 ();
 sg13g2_decap_8 FILLER_1_2586 ();
 sg13g2_decap_8 FILLER_1_2593 ();
 sg13g2_decap_8 FILLER_1_2600 ();
 sg13g2_decap_8 FILLER_1_2607 ();
 sg13g2_decap_8 FILLER_1_2614 ();
 sg13g2_decap_8 FILLER_1_2621 ();
 sg13g2_decap_8 FILLER_1_2628 ();
 sg13g2_decap_8 FILLER_1_2635 ();
 sg13g2_decap_8 FILLER_1_2642 ();
 sg13g2_decap_8 FILLER_1_2649 ();
 sg13g2_decap_8 FILLER_1_2656 ();
 sg13g2_decap_8 FILLER_1_2663 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_11 ();
 sg13g2_fill_2 FILLER_2_15 ();
 sg13g2_fill_1 FILLER_2_17 ();
 sg13g2_fill_1 FILLER_2_25 ();
 sg13g2_fill_2 FILLER_2_71 ();
 sg13g2_fill_1 FILLER_2_73 ();
 sg13g2_fill_2 FILLER_2_103 ();
 sg13g2_decap_8 FILLER_2_115 ();
 sg13g2_fill_2 FILLER_2_122 ();
 sg13g2_fill_2 FILLER_2_170 ();
 sg13g2_decap_4 FILLER_2_208 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_fill_2 FILLER_2_348 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_fill_2 FILLER_2_365 ();
 sg13g2_fill_1 FILLER_2_371 ();
 sg13g2_fill_1 FILLER_2_376 ();
 sg13g2_fill_1 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_407 ();
 sg13g2_decap_4 FILLER_2_414 ();
 sg13g2_fill_2 FILLER_2_453 ();
 sg13g2_fill_1 FILLER_2_455 ();
 sg13g2_decap_4 FILLER_2_482 ();
 sg13g2_fill_1 FILLER_2_486 ();
 sg13g2_decap_4 FILLER_2_491 ();
 sg13g2_fill_1 FILLER_2_495 ();
 sg13g2_fill_1 FILLER_2_501 ();
 sg13g2_decap_4 FILLER_2_537 ();
 sg13g2_fill_2 FILLER_2_541 ();
 sg13g2_fill_2 FILLER_2_571 ();
 sg13g2_fill_2 FILLER_2_601 ();
 sg13g2_fill_1 FILLER_2_622 ();
 sg13g2_fill_2 FILLER_2_628 ();
 sg13g2_fill_1 FILLER_2_630 ();
 sg13g2_fill_2 FILLER_2_636 ();
 sg13g2_fill_2 FILLER_2_653 ();
 sg13g2_fill_1 FILLER_2_674 ();
 sg13g2_fill_1 FILLER_2_680 ();
 sg13g2_fill_1 FILLER_2_685 ();
 sg13g2_decap_4 FILLER_2_732 ();
 sg13g2_fill_1 FILLER_2_736 ();
 sg13g2_fill_1 FILLER_2_747 ();
 sg13g2_fill_2 FILLER_2_774 ();
 sg13g2_fill_1 FILLER_2_776 ();
 sg13g2_fill_2 FILLER_2_834 ();
 sg13g2_fill_1 FILLER_2_836 ();
 sg13g2_decap_4 FILLER_2_874 ();
 sg13g2_fill_1 FILLER_2_878 ();
 sg13g2_decap_8 FILLER_2_904 ();
 sg13g2_decap_8 FILLER_2_911 ();
 sg13g2_fill_2 FILLER_2_918 ();
 sg13g2_fill_1 FILLER_2_920 ();
 sg13g2_fill_1 FILLER_2_925 ();
 sg13g2_fill_2 FILLER_2_935 ();
 sg13g2_fill_1 FILLER_2_937 ();
 sg13g2_decap_4 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_993 ();
 sg13g2_decap_4 FILLER_2_1004 ();
 sg13g2_decap_4 FILLER_2_1012 ();
 sg13g2_fill_1 FILLER_2_1016 ();
 sg13g2_fill_2 FILLER_2_1052 ();
 sg13g2_fill_1 FILLER_2_1102 ();
 sg13g2_decap_4 FILLER_2_1125 ();
 sg13g2_fill_1 FILLER_2_1129 ();
 sg13g2_fill_1 FILLER_2_1158 ();
 sg13g2_fill_1 FILLER_2_1186 ();
 sg13g2_fill_1 FILLER_2_1192 ();
 sg13g2_fill_1 FILLER_2_1224 ();
 sg13g2_decap_4 FILLER_2_1272 ();
 sg13g2_fill_2 FILLER_2_1276 ();
 sg13g2_fill_2 FILLER_2_1288 ();
 sg13g2_fill_1 FILLER_2_1290 ();
 sg13g2_decap_8 FILLER_2_1321 ();
 sg13g2_fill_1 FILLER_2_1328 ();
 sg13g2_fill_2 FILLER_2_1343 ();
 sg13g2_fill_1 FILLER_2_1481 ();
 sg13g2_fill_2 FILLER_2_1506 ();
 sg13g2_fill_1 FILLER_2_1508 ();
 sg13g2_fill_1 FILLER_2_1571 ();
 sg13g2_fill_1 FILLER_2_1645 ();
 sg13g2_fill_2 FILLER_2_1672 ();
 sg13g2_fill_2 FILLER_2_1700 ();
 sg13g2_fill_2 FILLER_2_1706 ();
 sg13g2_fill_1 FILLER_2_1712 ();
 sg13g2_fill_1 FILLER_2_1743 ();
 sg13g2_decap_4 FILLER_2_1811 ();
 sg13g2_fill_2 FILLER_2_1823 ();
 sg13g2_fill_2 FILLER_2_1835 ();
 sg13g2_decap_8 FILLER_2_1869 ();
 sg13g2_decap_8 FILLER_2_1876 ();
 sg13g2_decap_8 FILLER_2_1883 ();
 sg13g2_fill_1 FILLER_2_1890 ();
 sg13g2_decap_4 FILLER_2_1899 ();
 sg13g2_fill_1 FILLER_2_1903 ();
 sg13g2_fill_2 FILLER_2_1914 ();
 sg13g2_fill_1 FILLER_2_1942 ();
 sg13g2_fill_1 FILLER_2_1983 ();
 sg13g2_fill_2 FILLER_2_1994 ();
 sg13g2_fill_1 FILLER_2_1996 ();
 sg13g2_fill_2 FILLER_2_2001 ();
 sg13g2_fill_1 FILLER_2_2003 ();
 sg13g2_fill_1 FILLER_2_2076 ();
 sg13g2_decap_4 FILLER_2_2199 ();
 sg13g2_fill_2 FILLER_2_2213 ();
 sg13g2_fill_1 FILLER_2_2215 ();
 sg13g2_decap_4 FILLER_2_2246 ();
 sg13g2_decap_8 FILLER_2_2312 ();
 sg13g2_decap_8 FILLER_2_2319 ();
 sg13g2_fill_2 FILLER_2_2326 ();
 sg13g2_fill_2 FILLER_2_2331 ();
 sg13g2_fill_1 FILLER_2_2333 ();
 sg13g2_decap_8 FILLER_2_2360 ();
 sg13g2_decap_4 FILLER_2_2367 ();
 sg13g2_fill_2 FILLER_2_2404 ();
 sg13g2_decap_8 FILLER_2_2484 ();
 sg13g2_fill_2 FILLER_2_2491 ();
 sg13g2_fill_1 FILLER_2_2493 ();
 sg13g2_decap_8 FILLER_2_2524 ();
 sg13g2_decap_8 FILLER_2_2531 ();
 sg13g2_decap_8 FILLER_2_2538 ();
 sg13g2_decap_8 FILLER_2_2545 ();
 sg13g2_decap_8 FILLER_2_2552 ();
 sg13g2_decap_8 FILLER_2_2559 ();
 sg13g2_decap_8 FILLER_2_2566 ();
 sg13g2_decap_8 FILLER_2_2573 ();
 sg13g2_decap_8 FILLER_2_2580 ();
 sg13g2_decap_8 FILLER_2_2587 ();
 sg13g2_decap_8 FILLER_2_2594 ();
 sg13g2_decap_8 FILLER_2_2601 ();
 sg13g2_decap_8 FILLER_2_2608 ();
 sg13g2_decap_8 FILLER_2_2615 ();
 sg13g2_decap_8 FILLER_2_2622 ();
 sg13g2_decap_8 FILLER_2_2629 ();
 sg13g2_decap_8 FILLER_2_2636 ();
 sg13g2_decap_8 FILLER_2_2643 ();
 sg13g2_decap_8 FILLER_2_2650 ();
 sg13g2_decap_8 FILLER_2_2657 ();
 sg13g2_decap_4 FILLER_2_2664 ();
 sg13g2_fill_2 FILLER_2_2668 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_61 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_1 FILLER_3_82 ();
 sg13g2_fill_1 FILLER_3_86 ();
 sg13g2_decap_8 FILLER_3_103 ();
 sg13g2_fill_1 FILLER_3_110 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_fill_2 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_fill_1 FILLER_3_282 ();
 sg13g2_decap_4 FILLER_3_287 ();
 sg13g2_fill_1 FILLER_3_291 ();
 sg13g2_decap_4 FILLER_3_302 ();
 sg13g2_fill_1 FILLER_3_306 ();
 sg13g2_fill_1 FILLER_3_358 ();
 sg13g2_fill_1 FILLER_3_364 ();
 sg13g2_fill_1 FILLER_3_380 ();
 sg13g2_fill_2 FILLER_3_416 ();
 sg13g2_fill_1 FILLER_3_418 ();
 sg13g2_fill_1 FILLER_3_433 ();
 sg13g2_fill_1 FILLER_3_438 ();
 sg13g2_fill_1 FILLER_3_458 ();
 sg13g2_fill_1 FILLER_3_463 ();
 sg13g2_fill_1 FILLER_3_474 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_fill_2 FILLER_3_487 ();
 sg13g2_fill_2 FILLER_3_494 ();
 sg13g2_decap_4 FILLER_3_501 ();
 sg13g2_fill_2 FILLER_3_515 ();
 sg13g2_fill_1 FILLER_3_517 ();
 sg13g2_fill_1 FILLER_3_544 ();
 sg13g2_fill_2 FILLER_3_620 ();
 sg13g2_fill_2 FILLER_3_626 ();
 sg13g2_fill_1 FILLER_3_632 ();
 sg13g2_fill_2 FILLER_3_637 ();
 sg13g2_fill_1 FILLER_3_693 ();
 sg13g2_fill_2 FILLER_3_730 ();
 sg13g2_fill_1 FILLER_3_732 ();
 sg13g2_fill_1 FILLER_3_737 ();
 sg13g2_fill_1 FILLER_3_747 ();
 sg13g2_decap_4 FILLER_3_774 ();
 sg13g2_fill_2 FILLER_3_778 ();
 sg13g2_fill_1 FILLER_3_824 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_fill_2 FILLER_3_836 ();
 sg13g2_fill_2 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_901 ();
 sg13g2_fill_2 FILLER_3_913 ();
 sg13g2_fill_2 FILLER_3_945 ();
 sg13g2_decap_4 FILLER_3_969 ();
 sg13g2_fill_1 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_978 ();
 sg13g2_decap_8 FILLER_3_985 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_4 FILLER_3_1008 ();
 sg13g2_fill_2 FILLER_3_1020 ();
 sg13g2_fill_1 FILLER_3_1061 ();
 sg13g2_decap_4 FILLER_3_1101 ();
 sg13g2_fill_1 FILLER_3_1171 ();
 sg13g2_fill_2 FILLER_3_1181 ();
 sg13g2_fill_1 FILLER_3_1188 ();
 sg13g2_fill_1 FILLER_3_1223 ();
 sg13g2_fill_2 FILLER_3_1243 ();
 sg13g2_fill_1 FILLER_3_1245 ();
 sg13g2_fill_2 FILLER_3_1282 ();
 sg13g2_decap_8 FILLER_3_1318 ();
 sg13g2_decap_8 FILLER_3_1325 ();
 sg13g2_decap_8 FILLER_3_1342 ();
 sg13g2_fill_1 FILLER_3_1349 ();
 sg13g2_decap_4 FILLER_3_1376 ();
 sg13g2_fill_2 FILLER_3_1390 ();
 sg13g2_decap_8 FILLER_3_1415 ();
 sg13g2_fill_2 FILLER_3_1468 ();
 sg13g2_fill_1 FILLER_3_1470 ();
 sg13g2_fill_2 FILLER_3_1536 ();
 sg13g2_fill_1 FILLER_3_1574 ();
 sg13g2_decap_4 FILLER_3_1593 ();
 sg13g2_fill_2 FILLER_3_1663 ();
 sg13g2_fill_1 FILLER_3_1665 ();
 sg13g2_fill_1 FILLER_3_1670 ();
 sg13g2_fill_2 FILLER_3_1675 ();
 sg13g2_fill_2 FILLER_3_1681 ();
 sg13g2_fill_2 FILLER_3_1709 ();
 sg13g2_fill_1 FILLER_3_1741 ();
 sg13g2_fill_1 FILLER_3_1771 ();
 sg13g2_fill_1 FILLER_3_1778 ();
 sg13g2_decap_4 FILLER_3_1799 ();
 sg13g2_fill_1 FILLER_3_1860 ();
 sg13g2_fill_1 FILLER_3_1891 ();
 sg13g2_decap_4 FILLER_3_1895 ();
 sg13g2_decap_4 FILLER_3_1928 ();
 sg13g2_fill_2 FILLER_3_1932 ();
 sg13g2_fill_2 FILLER_3_1944 ();
 sg13g2_fill_1 FILLER_3_1950 ();
 sg13g2_decap_4 FILLER_3_1972 ();
 sg13g2_fill_2 FILLER_3_1976 ();
 sg13g2_fill_2 FILLER_3_1988 ();
 sg13g2_fill_2 FILLER_3_2000 ();
 sg13g2_decap_4 FILLER_3_2033 ();
 sg13g2_fill_2 FILLER_3_2090 ();
 sg13g2_decap_4 FILLER_3_2128 ();
 sg13g2_fill_1 FILLER_3_2132 ();
 sg13g2_fill_2 FILLER_3_2176 ();
 sg13g2_fill_2 FILLER_3_2265 ();
 sg13g2_fill_2 FILLER_3_2271 ();
 sg13g2_fill_1 FILLER_3_2273 ();
 sg13g2_decap_8 FILLER_3_2308 ();
 sg13g2_decap_4 FILLER_3_2315 ();
 sg13g2_fill_1 FILLER_3_2319 ();
 sg13g2_decap_8 FILLER_3_2343 ();
 sg13g2_decap_8 FILLER_3_2350 ();
 sg13g2_decap_8 FILLER_3_2357 ();
 sg13g2_decap_8 FILLER_3_2364 ();
 sg13g2_fill_2 FILLER_3_2384 ();
 sg13g2_fill_2 FILLER_3_2420 ();
 sg13g2_fill_1 FILLER_3_2422 ();
 sg13g2_decap_4 FILLER_3_2447 ();
 sg13g2_fill_1 FILLER_3_2451 ();
 sg13g2_decap_8 FILLER_3_2456 ();
 sg13g2_decap_8 FILLER_3_2463 ();
 sg13g2_fill_1 FILLER_3_2480 ();
 sg13g2_fill_2 FILLER_3_2491 ();
 sg13g2_fill_2 FILLER_3_2503 ();
 sg13g2_fill_1 FILLER_3_2505 ();
 sg13g2_fill_2 FILLER_3_2568 ();
 sg13g2_fill_1 FILLER_3_2570 ();
 sg13g2_decap_8 FILLER_3_2597 ();
 sg13g2_decap_8 FILLER_3_2604 ();
 sg13g2_decap_8 FILLER_3_2611 ();
 sg13g2_decap_8 FILLER_3_2618 ();
 sg13g2_decap_8 FILLER_3_2625 ();
 sg13g2_decap_8 FILLER_3_2632 ();
 sg13g2_decap_8 FILLER_3_2639 ();
 sg13g2_decap_8 FILLER_3_2646 ();
 sg13g2_decap_8 FILLER_3_2653 ();
 sg13g2_decap_8 FILLER_3_2660 ();
 sg13g2_fill_2 FILLER_3_2667 ();
 sg13g2_fill_1 FILLER_3_2669 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_14 ();
 sg13g2_fill_1 FILLER_4_16 ();
 sg13g2_decap_8 FILLER_4_47 ();
 sg13g2_fill_1 FILLER_4_54 ();
 sg13g2_fill_2 FILLER_4_64 ();
 sg13g2_fill_2 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_4 FILLER_4_137 ();
 sg13g2_fill_1 FILLER_4_141 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_166 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_187 ();
 sg13g2_decap_4 FILLER_4_199 ();
 sg13g2_fill_2 FILLER_4_203 ();
 sg13g2_fill_2 FILLER_4_220 ();
 sg13g2_fill_2 FILLER_4_227 ();
 sg13g2_decap_4 FILLER_4_233 ();
 sg13g2_decap_4 FILLER_4_250 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_4 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_fill_2 FILLER_4_296 ();
 sg13g2_fill_2 FILLER_4_308 ();
 sg13g2_decap_4 FILLER_4_324 ();
 sg13g2_fill_2 FILLER_4_337 ();
 sg13g2_fill_1 FILLER_4_339 ();
 sg13g2_fill_2 FILLER_4_344 ();
 sg13g2_fill_1 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_383 ();
 sg13g2_fill_2 FILLER_4_389 ();
 sg13g2_fill_1 FILLER_4_391 ();
 sg13g2_fill_1 FILLER_4_410 ();
 sg13g2_decap_4 FILLER_4_416 ();
 sg13g2_fill_2 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_426 ();
 sg13g2_decap_4 FILLER_4_437 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_4 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_491 ();
 sg13g2_decap_8 FILLER_4_498 ();
 sg13g2_fill_1 FILLER_4_509 ();
 sg13g2_fill_1 FILLER_4_520 ();
 sg13g2_decap_8 FILLER_4_531 ();
 sg13g2_decap_4 FILLER_4_538 ();
 sg13g2_fill_1 FILLER_4_582 ();
 sg13g2_fill_2 FILLER_4_588 ();
 sg13g2_fill_2 FILLER_4_638 ();
 sg13g2_decap_4 FILLER_4_649 ();
 sg13g2_fill_1 FILLER_4_653 ();
 sg13g2_decap_4 FILLER_4_658 ();
 sg13g2_fill_1 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_667 ();
 sg13g2_decap_4 FILLER_4_674 ();
 sg13g2_fill_2 FILLER_4_678 ();
 sg13g2_fill_2 FILLER_4_695 ();
 sg13g2_fill_1 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_4 FILLER_4_732 ();
 sg13g2_fill_2 FILLER_4_760 ();
 sg13g2_fill_2 FILLER_4_768 ();
 sg13g2_fill_2 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_4 FILLER_4_830 ();
 sg13g2_decap_4 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_4 FILLER_4_923 ();
 sg13g2_fill_2 FILLER_4_927 ();
 sg13g2_decap_4 FILLER_4_933 ();
 sg13g2_fill_2 FILLER_4_937 ();
 sg13g2_fill_2 FILLER_4_970 ();
 sg13g2_fill_2 FILLER_4_976 ();
 sg13g2_fill_2 FILLER_4_1004 ();
 sg13g2_decap_4 FILLER_4_1011 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_decap_8 FILLER_4_1059 ();
 sg13g2_decap_4 FILLER_4_1066 ();
 sg13g2_fill_2 FILLER_4_1070 ();
 sg13g2_fill_2 FILLER_4_1081 ();
 sg13g2_fill_1 FILLER_4_1104 ();
 sg13g2_fill_2 FILLER_4_1110 ();
 sg13g2_fill_1 FILLER_4_1133 ();
 sg13g2_fill_1 FILLER_4_1139 ();
 sg13g2_fill_1 FILLER_4_1145 ();
 sg13g2_fill_1 FILLER_4_1189 ();
 sg13g2_fill_2 FILLER_4_1198 ();
 sg13g2_decap_8 FILLER_4_1221 ();
 sg13g2_decap_8 FILLER_4_1228 ();
 sg13g2_decap_8 FILLER_4_1235 ();
 sg13g2_decap_8 FILLER_4_1242 ();
 sg13g2_fill_1 FILLER_4_1249 ();
 sg13g2_fill_2 FILLER_4_1271 ();
 sg13g2_fill_1 FILLER_4_1273 ();
 sg13g2_decap_8 FILLER_4_1311 ();
 sg13g2_fill_2 FILLER_4_1318 ();
 sg13g2_fill_1 FILLER_4_1320 ();
 sg13g2_decap_8 FILLER_4_1347 ();
 sg13g2_decap_4 FILLER_4_1354 ();
 sg13g2_fill_1 FILLER_4_1358 ();
 sg13g2_decap_8 FILLER_4_1425 ();
 sg13g2_fill_1 FILLER_4_1432 ();
 sg13g2_fill_1 FILLER_4_1437 ();
 sg13g2_fill_2 FILLER_4_1442 ();
 sg13g2_decap_8 FILLER_4_1454 ();
 sg13g2_fill_2 FILLER_4_1461 ();
 sg13g2_fill_1 FILLER_4_1463 ();
 sg13g2_decap_8 FILLER_4_1490 ();
 sg13g2_fill_2 FILLER_4_1497 ();
 sg13g2_decap_4 FILLER_4_1513 ();
 sg13g2_decap_8 FILLER_4_1525 ();
 sg13g2_decap_8 FILLER_4_1532 ();
 sg13g2_decap_8 FILLER_4_1539 ();
 sg13g2_fill_2 FILLER_4_1546 ();
 sg13g2_fill_1 FILLER_4_1548 ();
 sg13g2_fill_2 FILLER_4_1563 ();
 sg13g2_fill_1 FILLER_4_1565 ();
 sg13g2_decap_4 FILLER_4_1592 ();
 sg13g2_fill_1 FILLER_4_1596 ();
 sg13g2_decap_8 FILLER_4_1614 ();
 sg13g2_decap_8 FILLER_4_1621 ();
 sg13g2_fill_2 FILLER_4_1628 ();
 sg13g2_decap_8 FILLER_4_1666 ();
 sg13g2_decap_8 FILLER_4_1673 ();
 sg13g2_decap_8 FILLER_4_1680 ();
 sg13g2_fill_2 FILLER_4_1687 ();
 sg13g2_decap_8 FILLER_4_1693 ();
 sg13g2_decap_8 FILLER_4_1700 ();
 sg13g2_decap_8 FILLER_4_1707 ();
 sg13g2_decap_8 FILLER_4_1714 ();
 sg13g2_fill_1 FILLER_4_1721 ();
 sg13g2_fill_2 FILLER_4_1746 ();
 sg13g2_fill_2 FILLER_4_1754 ();
 sg13g2_fill_1 FILLER_4_1766 ();
 sg13g2_fill_2 FILLER_4_1782 ();
 sg13g2_fill_2 FILLER_4_1788 ();
 sg13g2_decap_8 FILLER_4_1796 ();
 sg13g2_fill_2 FILLER_4_1803 ();
 sg13g2_fill_1 FILLER_4_1805 ();
 sg13g2_fill_1 FILLER_4_1837 ();
 sg13g2_fill_1 FILLER_4_1856 ();
 sg13g2_fill_2 FILLER_4_1895 ();
 sg13g2_fill_2 FILLER_4_1937 ();
 sg13g2_fill_1 FILLER_4_1939 ();
 sg13g2_decap_8 FILLER_4_1950 ();
 sg13g2_fill_2 FILLER_4_1974 ();
 sg13g2_fill_1 FILLER_4_1976 ();
 sg13g2_decap_8 FILLER_4_2003 ();
 sg13g2_decap_8 FILLER_4_2014 ();
 sg13g2_decap_8 FILLER_4_2021 ();
 sg13g2_decap_8 FILLER_4_2028 ();
 sg13g2_decap_8 FILLER_4_2035 ();
 sg13g2_decap_8 FILLER_4_2042 ();
 sg13g2_decap_4 FILLER_4_2049 ();
 sg13g2_decap_8 FILLER_4_2057 ();
 sg13g2_decap_4 FILLER_4_2064 ();
 sg13g2_fill_1 FILLER_4_2068 ();
 sg13g2_decap_4 FILLER_4_2081 ();
 sg13g2_fill_1 FILLER_4_2085 ();
 sg13g2_decap_8 FILLER_4_2096 ();
 sg13g2_fill_2 FILLER_4_2103 ();
 sg13g2_fill_2 FILLER_4_2113 ();
 sg13g2_fill_1 FILLER_4_2115 ();
 sg13g2_fill_2 FILLER_4_2159 ();
 sg13g2_fill_1 FILLER_4_2161 ();
 sg13g2_fill_1 FILLER_4_2172 ();
 sg13g2_fill_2 FILLER_4_2223 ();
 sg13g2_fill_1 FILLER_4_2225 ();
 sg13g2_decap_8 FILLER_4_2287 ();
 sg13g2_fill_2 FILLER_4_2294 ();
 sg13g2_fill_1 FILLER_4_2296 ();
 sg13g2_decap_8 FILLER_4_2389 ();
 sg13g2_fill_2 FILLER_4_2396 ();
 sg13g2_fill_1 FILLER_4_2398 ();
 sg13g2_decap_4 FILLER_4_2439 ();
 sg13g2_decap_4 FILLER_4_2479 ();
 sg13g2_decap_8 FILLER_4_2517 ();
 sg13g2_decap_4 FILLER_4_2524 ();
 sg13g2_fill_2 FILLER_4_2528 ();
 sg13g2_fill_2 FILLER_4_2570 ();
 sg13g2_decap_8 FILLER_4_2602 ();
 sg13g2_decap_8 FILLER_4_2609 ();
 sg13g2_decap_8 FILLER_4_2616 ();
 sg13g2_decap_8 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_4 FILLER_4_2665 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_33 ();
 sg13g2_fill_1 FILLER_5_40 ();
 sg13g2_decap_8 FILLER_5_45 ();
 sg13g2_decap_4 FILLER_5_52 ();
 sg13g2_decap_4 FILLER_5_61 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_2 FILLER_5_71 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_fill_2 FILLER_5_79 ();
 sg13g2_fill_1 FILLER_5_89 ();
 sg13g2_decap_8 FILLER_5_100 ();
 sg13g2_decap_4 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_111 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_decap_8 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_136 ();
 sg13g2_fill_1 FILLER_5_141 ();
 sg13g2_fill_2 FILLER_5_157 ();
 sg13g2_fill_1 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_174 ();
 sg13g2_fill_2 FILLER_5_181 ();
 sg13g2_fill_1 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_4 FILLER_5_210 ();
 sg13g2_fill_2 FILLER_5_214 ();
 sg13g2_fill_1 FILLER_5_225 ();
 sg13g2_fill_1 FILLER_5_232 ();
 sg13g2_fill_1 FILLER_5_244 ();
 sg13g2_decap_8 FILLER_5_261 ();
 sg13g2_fill_2 FILLER_5_268 ();
 sg13g2_fill_1 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_282 ();
 sg13g2_fill_1 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_4 FILLER_5_346 ();
 sg13g2_fill_2 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_4 FILLER_5_372 ();
 sg13g2_fill_1 FILLER_5_376 ();
 sg13g2_fill_1 FILLER_5_382 ();
 sg13g2_fill_1 FILLER_5_392 ();
 sg13g2_fill_1 FILLER_5_411 ();
 sg13g2_fill_1 FILLER_5_416 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_fill_2 FILLER_5_435 ();
 sg13g2_fill_1 FILLER_5_437 ();
 sg13g2_decap_8 FILLER_5_464 ();
 sg13g2_decap_4 FILLER_5_471 ();
 sg13g2_fill_1 FILLER_5_475 ();
 sg13g2_decap_4 FILLER_5_485 ();
 sg13g2_fill_1 FILLER_5_489 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_fill_2 FILLER_5_526 ();
 sg13g2_decap_8 FILLER_5_534 ();
 sg13g2_decap_8 FILLER_5_541 ();
 sg13g2_fill_2 FILLER_5_548 ();
 sg13g2_fill_2 FILLER_5_554 ();
 sg13g2_decap_4 FILLER_5_565 ();
 sg13g2_fill_1 FILLER_5_569 ();
 sg13g2_fill_2 FILLER_5_575 ();
 sg13g2_decap_4 FILLER_5_581 ();
 sg13g2_fill_2 FILLER_5_598 ();
 sg13g2_fill_1 FILLER_5_610 ();
 sg13g2_fill_2 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_fill_1 FILLER_5_648 ();
 sg13g2_fill_2 FILLER_5_659 ();
 sg13g2_fill_1 FILLER_5_661 ();
 sg13g2_decap_8 FILLER_5_671 ();
 sg13g2_decap_8 FILLER_5_678 ();
 sg13g2_fill_2 FILLER_5_685 ();
 sg13g2_decap_8 FILLER_5_695 ();
 sg13g2_decap_8 FILLER_5_702 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_fill_2 FILLER_5_723 ();
 sg13g2_fill_1 FILLER_5_725 ();
 sg13g2_fill_1 FILLER_5_744 ();
 sg13g2_fill_2 FILLER_5_759 ();
 sg13g2_fill_2 FILLER_5_766 ();
 sg13g2_fill_1 FILLER_5_774 ();
 sg13g2_fill_1 FILLER_5_786 ();
 sg13g2_fill_2 FILLER_5_797 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_4 FILLER_5_830 ();
 sg13g2_fill_1 FILLER_5_874 ();
 sg13g2_decap_8 FILLER_5_895 ();
 sg13g2_decap_8 FILLER_5_902 ();
 sg13g2_decap_8 FILLER_5_909 ();
 sg13g2_fill_1 FILLER_5_916 ();
 sg13g2_fill_1 FILLER_5_952 ();
 sg13g2_fill_1 FILLER_5_984 ();
 sg13g2_fill_2 FILLER_5_989 ();
 sg13g2_fill_1 FILLER_5_996 ();
 sg13g2_fill_2 FILLER_5_1001 ();
 sg13g2_decap_4 FILLER_5_1029 ();
 sg13g2_fill_2 FILLER_5_1033 ();
 sg13g2_decap_8 FILLER_5_1040 ();
 sg13g2_decap_8 FILLER_5_1047 ();
 sg13g2_decap_8 FILLER_5_1054 ();
 sg13g2_decap_8 FILLER_5_1061 ();
 sg13g2_decap_4 FILLER_5_1068 ();
 sg13g2_fill_2 FILLER_5_1072 ();
 sg13g2_decap_4 FILLER_5_1079 ();
 sg13g2_decap_8 FILLER_5_1087 ();
 sg13g2_decap_4 FILLER_5_1094 ();
 sg13g2_fill_2 FILLER_5_1098 ();
 sg13g2_fill_2 FILLER_5_1104 ();
 sg13g2_decap_8 FILLER_5_1132 ();
 sg13g2_fill_2 FILLER_5_1148 ();
 sg13g2_decap_8 FILLER_5_1207 ();
 sg13g2_decap_8 FILLER_5_1214 ();
 sg13g2_decap_8 FILLER_5_1221 ();
 sg13g2_decap_8 FILLER_5_1228 ();
 sg13g2_decap_4 FILLER_5_1235 ();
 sg13g2_fill_1 FILLER_5_1239 ();
 sg13g2_decap_4 FILLER_5_1266 ();
 sg13g2_fill_1 FILLER_5_1270 ();
 sg13g2_decap_8 FILLER_5_1285 ();
 sg13g2_decap_8 FILLER_5_1292 ();
 sg13g2_decap_8 FILLER_5_1299 ();
 sg13g2_decap_8 FILLER_5_1306 ();
 sg13g2_decap_8 FILLER_5_1313 ();
 sg13g2_decap_8 FILLER_5_1320 ();
 sg13g2_fill_2 FILLER_5_1327 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_4 FILLER_5_1340 ();
 sg13g2_fill_2 FILLER_5_1344 ();
 sg13g2_fill_1 FILLER_5_1382 ();
 sg13g2_fill_1 FILLER_5_1387 ();
 sg13g2_fill_2 FILLER_5_1406 ();
 sg13g2_decap_4 FILLER_5_1412 ();
 sg13g2_decap_8 FILLER_5_1446 ();
 sg13g2_decap_4 FILLER_5_1453 ();
 sg13g2_fill_2 FILLER_5_1457 ();
 sg13g2_fill_2 FILLER_5_1479 ();
 sg13g2_fill_1 FILLER_5_1481 ();
 sg13g2_fill_1 FILLER_5_1518 ();
 sg13g2_decap_8 FILLER_5_1555 ();
 sg13g2_decap_4 FILLER_5_1566 ();
 sg13g2_fill_2 FILLER_5_1570 ();
 sg13g2_decap_8 FILLER_5_1582 ();
 sg13g2_fill_2 FILLER_5_1589 ();
 sg13g2_fill_1 FILLER_5_1591 ();
 sg13g2_decap_8 FILLER_5_1622 ();
 sg13g2_decap_4 FILLER_5_1629 ();
 sg13g2_fill_1 FILLER_5_1633 ();
 sg13g2_decap_8 FILLER_5_1638 ();
 sg13g2_decap_8 FILLER_5_1645 ();
 sg13g2_fill_1 FILLER_5_1652 ();
 sg13g2_decap_8 FILLER_5_1657 ();
 sg13g2_decap_8 FILLER_5_1664 ();
 sg13g2_decap_4 FILLER_5_1707 ();
 sg13g2_fill_1 FILLER_5_1711 ();
 sg13g2_decap_8 FILLER_5_1716 ();
 sg13g2_decap_8 FILLER_5_1723 ();
 sg13g2_decap_8 FILLER_5_1730 ();
 sg13g2_fill_1 FILLER_5_1737 ();
 sg13g2_decap_4 FILLER_5_1770 ();
 sg13g2_decap_4 FILLER_5_1783 ();
 sg13g2_fill_2 FILLER_5_1787 ();
 sg13g2_fill_2 FILLER_5_1794 ();
 sg13g2_decap_8 FILLER_5_1804 ();
 sg13g2_fill_2 FILLER_5_1811 ();
 sg13g2_fill_2 FILLER_5_1818 ();
 sg13g2_fill_2 FILLER_5_1860 ();
 sg13g2_fill_1 FILLER_5_1883 ();
 sg13g2_fill_2 FILLER_5_1887 ();
 sg13g2_decap_8 FILLER_5_1907 ();
 sg13g2_decap_8 FILLER_5_1914 ();
 sg13g2_decap_8 FILLER_5_1921 ();
 sg13g2_decap_4 FILLER_5_1928 ();
 sg13g2_fill_2 FILLER_5_1932 ();
 sg13g2_decap_8 FILLER_5_1964 ();
 sg13g2_decap_8 FILLER_5_1971 ();
 sg13g2_decap_4 FILLER_5_1978 ();
 sg13g2_fill_1 FILLER_5_1982 ();
 sg13g2_decap_4 FILLER_5_1987 ();
 sg13g2_fill_2 FILLER_5_1991 ();
 sg13g2_decap_8 FILLER_5_2003 ();
 sg13g2_decap_8 FILLER_5_2010 ();
 sg13g2_decap_8 FILLER_5_2017 ();
 sg13g2_fill_2 FILLER_5_2024 ();
 sg13g2_fill_1 FILLER_5_2040 ();
 sg13g2_fill_2 FILLER_5_2059 ();
 sg13g2_fill_1 FILLER_5_2061 ();
 sg13g2_decap_8 FILLER_5_2066 ();
 sg13g2_decap_8 FILLER_5_2073 ();
 sg13g2_fill_2 FILLER_5_2080 ();
 sg13g2_fill_1 FILLER_5_2082 ();
 sg13g2_fill_2 FILLER_5_2093 ();
 sg13g2_fill_2 FILLER_5_2129 ();
 sg13g2_fill_1 FILLER_5_2131 ();
 sg13g2_decap_8 FILLER_5_2158 ();
 sg13g2_fill_2 FILLER_5_2165 ();
 sg13g2_fill_1 FILLER_5_2188 ();
 sg13g2_decap_8 FILLER_5_2193 ();
 sg13g2_decap_8 FILLER_5_2200 ();
 sg13g2_decap_8 FILLER_5_2207 ();
 sg13g2_fill_2 FILLER_5_2214 ();
 sg13g2_fill_1 FILLER_5_2216 ();
 sg13g2_decap_8 FILLER_5_2247 ();
 sg13g2_fill_2 FILLER_5_2254 ();
 sg13g2_fill_2 FILLER_5_2260 ();
 sg13g2_fill_1 FILLER_5_2262 ();
 sg13g2_decap_8 FILLER_5_2286 ();
 sg13g2_decap_8 FILLER_5_2293 ();
 sg13g2_decap_4 FILLER_5_2300 ();
 sg13g2_fill_1 FILLER_5_2304 ();
 sg13g2_fill_1 FILLER_5_2351 ();
 sg13g2_decap_4 FILLER_5_2360 ();
 sg13g2_fill_1 FILLER_5_2364 ();
 sg13g2_decap_4 FILLER_5_2370 ();
 sg13g2_fill_2 FILLER_5_2400 ();
 sg13g2_fill_1 FILLER_5_2419 ();
 sg13g2_decap_8 FILLER_5_2446 ();
 sg13g2_decap_8 FILLER_5_2453 ();
 sg13g2_decap_4 FILLER_5_2460 ();
 sg13g2_fill_1 FILLER_5_2464 ();
 sg13g2_fill_2 FILLER_5_2496 ();
 sg13g2_fill_1 FILLER_5_2498 ();
 sg13g2_decap_4 FILLER_5_2509 ();
 sg13g2_decap_8 FILLER_5_2523 ();
 sg13g2_fill_2 FILLER_5_2530 ();
 sg13g2_fill_1 FILLER_5_2532 ();
 sg13g2_decap_4 FILLER_5_2624 ();
 sg13g2_decap_8 FILLER_5_2632 ();
 sg13g2_decap_8 FILLER_5_2639 ();
 sg13g2_decap_8 FILLER_5_2646 ();
 sg13g2_decap_8 FILLER_5_2653 ();
 sg13g2_decap_8 FILLER_5_2660 ();
 sg13g2_fill_2 FILLER_5_2667 ();
 sg13g2_fill_1 FILLER_5_2669 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_8 ();
 sg13g2_decap_4 FILLER_6_39 ();
 sg13g2_fill_2 FILLER_6_43 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_4 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_decap_4 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_149 ();
 sg13g2_fill_2 FILLER_6_155 ();
 sg13g2_fill_1 FILLER_6_171 ();
 sg13g2_decap_8 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_208 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_fill_2 FILLER_6_291 ();
 sg13g2_decap_4 FILLER_6_350 ();
 sg13g2_fill_2 FILLER_6_384 ();
 sg13g2_fill_1 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_4 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_413 ();
 sg13g2_fill_1 FILLER_6_433 ();
 sg13g2_decap_8 FILLER_6_470 ();
 sg13g2_fill_2 FILLER_6_477 ();
 sg13g2_fill_1 FILLER_6_509 ();
 sg13g2_fill_2 FILLER_6_514 ();
 sg13g2_decap_4 FILLER_6_551 ();
 sg13g2_fill_1 FILLER_6_555 ();
 sg13g2_decap_4 FILLER_6_561 ();
 sg13g2_fill_1 FILLER_6_565 ();
 sg13g2_decap_8 FILLER_6_575 ();
 sg13g2_decap_8 FILLER_6_582 ();
 sg13g2_decap_8 FILLER_6_589 ();
 sg13g2_decap_8 FILLER_6_596 ();
 sg13g2_decap_8 FILLER_6_603 ();
 sg13g2_decap_8 FILLER_6_610 ();
 sg13g2_decap_4 FILLER_6_617 ();
 sg13g2_fill_1 FILLER_6_621 ();
 sg13g2_decap_4 FILLER_6_661 ();
 sg13g2_fill_1 FILLER_6_665 ();
 sg13g2_fill_1 FILLER_6_670 ();
 sg13g2_fill_1 FILLER_6_675 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_fill_2 FILLER_6_714 ();
 sg13g2_fill_1 FILLER_6_716 ();
 sg13g2_fill_1 FILLER_6_752 ();
 sg13g2_fill_1 FILLER_6_757 ();
 sg13g2_fill_1 FILLER_6_763 ();
 sg13g2_fill_1 FILLER_6_768 ();
 sg13g2_fill_1 FILLER_6_774 ();
 sg13g2_fill_2 FILLER_6_780 ();
 sg13g2_fill_2 FILLER_6_786 ();
 sg13g2_fill_1 FILLER_6_792 ();
 sg13g2_decap_8 FILLER_6_829 ();
 sg13g2_decap_8 FILLER_6_836 ();
 sg13g2_decap_8 FILLER_6_848 ();
 sg13g2_decap_4 FILLER_6_855 ();
 sg13g2_fill_2 FILLER_6_859 ();
 sg13g2_decap_8 FILLER_6_871 ();
 sg13g2_decap_8 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_909 ();
 sg13g2_fill_2 FILLER_6_916 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_4 FILLER_6_980 ();
 sg13g2_fill_2 FILLER_6_984 ();
 sg13g2_fill_1 FILLER_6_1037 ();
 sg13g2_decap_4 FILLER_6_1047 ();
 sg13g2_decap_8 FILLER_6_1077 ();
 sg13g2_decap_8 FILLER_6_1084 ();
 sg13g2_decap_8 FILLER_6_1091 ();
 sg13g2_decap_8 FILLER_6_1098 ();
 sg13g2_decap_8 FILLER_6_1105 ();
 sg13g2_fill_2 FILLER_6_1112 ();
 sg13g2_fill_1 FILLER_6_1114 ();
 sg13g2_fill_2 FILLER_6_1120 ();
 sg13g2_fill_1 FILLER_6_1122 ();
 sg13g2_decap_8 FILLER_6_1127 ();
 sg13g2_decap_8 FILLER_6_1134 ();
 sg13g2_fill_1 FILLER_6_1141 ();
 sg13g2_decap_4 FILLER_6_1150 ();
 sg13g2_fill_2 FILLER_6_1154 ();
 sg13g2_decap_8 FILLER_6_1160 ();
 sg13g2_decap_8 FILLER_6_1167 ();
 sg13g2_decap_4 FILLER_6_1174 ();
 sg13g2_fill_1 FILLER_6_1178 ();
 sg13g2_decap_4 FILLER_6_1183 ();
 sg13g2_fill_1 FILLER_6_1187 ();
 sg13g2_fill_2 FILLER_6_1219 ();
 sg13g2_fill_1 FILLER_6_1221 ();
 sg13g2_decap_8 FILLER_6_1232 ();
 sg13g2_fill_1 FILLER_6_1239 ();
 sg13g2_fill_1 FILLER_6_1271 ();
 sg13g2_fill_2 FILLER_6_1298 ();
 sg13g2_decap_8 FILLER_6_1304 ();
 sg13g2_decap_8 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1318 ();
 sg13g2_decap_4 FILLER_6_1325 ();
 sg13g2_fill_1 FILLER_6_1329 ();
 sg13g2_decap_8 FILLER_6_1438 ();
 sg13g2_decap_8 FILLER_6_1445 ();
 sg13g2_fill_2 FILLER_6_1452 ();
 sg13g2_decap_8 FILLER_6_1458 ();
 sg13g2_decap_8 FILLER_6_1479 ();
 sg13g2_fill_1 FILLER_6_1512 ();
 sg13g2_fill_1 FILLER_6_1523 ();
 sg13g2_fill_1 FILLER_6_1528 ();
 sg13g2_decap_4 FILLER_6_1581 ();
 sg13g2_fill_1 FILLER_6_1585 ();
 sg13g2_decap_8 FILLER_6_1622 ();
 sg13g2_decap_8 FILLER_6_1629 ();
 sg13g2_fill_1 FILLER_6_1672 ();
 sg13g2_decap_4 FILLER_6_1742 ();
 sg13g2_fill_2 FILLER_6_1746 ();
 sg13g2_fill_2 FILLER_6_1751 ();
 sg13g2_decap_8 FILLER_6_1756 ();
 sg13g2_decap_4 FILLER_6_1763 ();
 sg13g2_fill_2 FILLER_6_1767 ();
 sg13g2_fill_1 FILLER_6_1774 ();
 sg13g2_fill_2 FILLER_6_1780 ();
 sg13g2_fill_1 FILLER_6_1782 ();
 sg13g2_fill_1 FILLER_6_1792 ();
 sg13g2_decap_8 FILLER_6_1798 ();
 sg13g2_decap_4 FILLER_6_1810 ();
 sg13g2_fill_1 FILLER_6_1819 ();
 sg13g2_fill_1 FILLER_6_1837 ();
 sg13g2_decap_4 FILLER_6_1844 ();
 sg13g2_fill_1 FILLER_6_1848 ();
 sg13g2_fill_1 FILLER_6_1853 ();
 sg13g2_fill_2 FILLER_6_1860 ();
 sg13g2_decap_8 FILLER_6_1866 ();
 sg13g2_decap_4 FILLER_6_1873 ();
 sg13g2_fill_2 FILLER_6_1877 ();
 sg13g2_fill_2 FILLER_6_1887 ();
 sg13g2_fill_1 FILLER_6_1894 ();
 sg13g2_decap_8 FILLER_6_1925 ();
 sg13g2_decap_8 FILLER_6_1932 ();
 sg13g2_decap_8 FILLER_6_1939 ();
 sg13g2_decap_4 FILLER_6_1946 ();
 sg13g2_decap_8 FILLER_6_1960 ();
 sg13g2_decap_8 FILLER_6_1967 ();
 sg13g2_fill_1 FILLER_6_1974 ();
 sg13g2_decap_4 FILLER_6_2015 ();
 sg13g2_fill_1 FILLER_6_2019 ();
 sg13g2_decap_4 FILLER_6_2050 ();
 sg13g2_fill_2 FILLER_6_2054 ();
 sg13g2_fill_1 FILLER_6_2138 ();
 sg13g2_decap_8 FILLER_6_2194 ();
 sg13g2_decap_4 FILLER_6_2201 ();
 sg13g2_fill_1 FILLER_6_2205 ();
 sg13g2_fill_2 FILLER_6_2236 ();
 sg13g2_fill_1 FILLER_6_2238 ();
 sg13g2_decap_8 FILLER_6_2275 ();
 sg13g2_decap_8 FILLER_6_2282 ();
 sg13g2_decap_8 FILLER_6_2289 ();
 sg13g2_fill_2 FILLER_6_2296 ();
 sg13g2_fill_1 FILLER_6_2298 ();
 sg13g2_fill_1 FILLER_6_2346 ();
 sg13g2_fill_2 FILLER_6_2373 ();
 sg13g2_fill_1 FILLER_6_2375 ();
 sg13g2_fill_2 FILLER_6_2416 ();
 sg13g2_fill_1 FILLER_6_2418 ();
 sg13g2_fill_1 FILLER_6_2445 ();
 sg13g2_fill_1 FILLER_6_2472 ();
 sg13g2_decap_8 FILLER_6_2486 ();
 sg13g2_decap_8 FILLER_6_2509 ();
 sg13g2_decap_8 FILLER_6_2516 ();
 sg13g2_decap_8 FILLER_6_2523 ();
 sg13g2_decap_4 FILLER_6_2530 ();
 sg13g2_fill_2 FILLER_6_2601 ();
 sg13g2_decap_8 FILLER_6_2611 ();
 sg13g2_fill_2 FILLER_6_2618 ();
 sg13g2_decap_8 FILLER_6_2650 ();
 sg13g2_decap_8 FILLER_6_2657 ();
 sg13g2_decap_4 FILLER_6_2664 ();
 sg13g2_fill_2 FILLER_6_2668 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_fill_1 FILLER_7_19 ();
 sg13g2_fill_2 FILLER_7_24 ();
 sg13g2_fill_2 FILLER_7_30 ();
 sg13g2_fill_1 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_38 ();
 sg13g2_fill_1 FILLER_7_40 ();
 sg13g2_fill_2 FILLER_7_45 ();
 sg13g2_fill_1 FILLER_7_70 ();
 sg13g2_decap_4 FILLER_7_87 ();
 sg13g2_fill_2 FILLER_7_91 ();
 sg13g2_decap_4 FILLER_7_106 ();
 sg13g2_fill_2 FILLER_7_156 ();
 sg13g2_fill_2 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_194 ();
 sg13g2_fill_2 FILLER_7_200 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_235 ();
 sg13g2_fill_2 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_264 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_fill_2 FILLER_7_282 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_decap_4 FILLER_7_289 ();
 sg13g2_decap_4 FILLER_7_307 ();
 sg13g2_fill_1 FILLER_7_355 ();
 sg13g2_fill_2 FILLER_7_361 ();
 sg13g2_fill_1 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_395 ();
 sg13g2_fill_2 FILLER_7_402 ();
 sg13g2_fill_2 FILLER_7_414 ();
 sg13g2_fill_1 FILLER_7_416 ();
 sg13g2_fill_2 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_592 ();
 sg13g2_decap_4 FILLER_7_599 ();
 sg13g2_fill_2 FILLER_7_607 ();
 sg13g2_decap_4 FILLER_7_615 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_fill_2 FILLER_7_637 ();
 sg13g2_fill_1 FILLER_7_652 ();
 sg13g2_fill_2 FILLER_7_687 ();
 sg13g2_decap_8 FILLER_7_694 ();
 sg13g2_fill_2 FILLER_7_707 ();
 sg13g2_fill_1 FILLER_7_713 ();
 sg13g2_fill_2 FILLER_7_745 ();
 sg13g2_fill_1 FILLER_7_747 ();
 sg13g2_fill_2 FILLER_7_752 ();
 sg13g2_fill_1 FILLER_7_754 ();
 sg13g2_fill_1 FILLER_7_765 ();
 sg13g2_fill_1 FILLER_7_771 ();
 sg13g2_decap_4 FILLER_7_832 ();
 sg13g2_fill_2 FILLER_7_840 ();
 sg13g2_decap_4 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_898 ();
 sg13g2_decap_4 FILLER_7_905 ();
 sg13g2_decap_8 FILLER_7_965 ();
 sg13g2_decap_8 FILLER_7_972 ();
 sg13g2_decap_8 FILLER_7_979 ();
 sg13g2_decap_8 FILLER_7_986 ();
 sg13g2_decap_8 FILLER_7_993 ();
 sg13g2_fill_2 FILLER_7_1000 ();
 sg13g2_fill_1 FILLER_7_1002 ();
 sg13g2_decap_8 FILLER_7_1032 ();
 sg13g2_fill_2 FILLER_7_1095 ();
 sg13g2_fill_1 FILLER_7_1097 ();
 sg13g2_fill_2 FILLER_7_1102 ();
 sg13g2_fill_1 FILLER_7_1104 ();
 sg13g2_decap_8 FILLER_7_1110 ();
 sg13g2_decap_8 FILLER_7_1117 ();
 sg13g2_decap_4 FILLER_7_1124 ();
 sg13g2_fill_2 FILLER_7_1128 ();
 sg13g2_fill_2 FILLER_7_1156 ();
 sg13g2_fill_1 FILLER_7_1158 ();
 sg13g2_fill_1 FILLER_7_1167 ();
 sg13g2_decap_4 FILLER_7_1172 ();
 sg13g2_fill_1 FILLER_7_1176 ();
 sg13g2_fill_1 FILLER_7_1182 ();
 sg13g2_fill_1 FILLER_7_1187 ();
 sg13g2_fill_2 FILLER_7_1237 ();
 sg13g2_decap_4 FILLER_7_1265 ();
 sg13g2_fill_2 FILLER_7_1279 ();
 sg13g2_decap_4 FILLER_7_1307 ();
 sg13g2_decap_8 FILLER_7_1412 ();
 sg13g2_decap_4 FILLER_7_1419 ();
 sg13g2_fill_1 FILLER_7_1423 ();
 sg13g2_decap_4 FILLER_7_1428 ();
 sg13g2_fill_1 FILLER_7_1436 ();
 sg13g2_decap_8 FILLER_7_1503 ();
 sg13g2_decap_8 FILLER_7_1510 ();
 sg13g2_decap_8 FILLER_7_1517 ();
 sg13g2_decap_8 FILLER_7_1573 ();
 sg13g2_decap_8 FILLER_7_1580 ();
 sg13g2_decap_8 FILLER_7_1587 ();
 sg13g2_fill_2 FILLER_7_1594 ();
 sg13g2_decap_4 FILLER_7_1600 ();
 sg13g2_fill_1 FILLER_7_1604 ();
 sg13g2_fill_1 FILLER_7_1615 ();
 sg13g2_fill_1 FILLER_7_1665 ();
 sg13g2_decap_8 FILLER_7_1685 ();
 sg13g2_fill_1 FILLER_7_1692 ();
 sg13g2_decap_8 FILLER_7_1697 ();
 sg13g2_fill_1 FILLER_7_1704 ();
 sg13g2_decap_8 FILLER_7_1713 ();
 sg13g2_decap_8 FILLER_7_1720 ();
 sg13g2_decap_4 FILLER_7_1735 ();
 sg13g2_fill_2 FILLER_7_1749 ();
 sg13g2_fill_1 FILLER_7_1756 ();
 sg13g2_decap_4 FILLER_7_1762 ();
 sg13g2_fill_2 FILLER_7_1766 ();
 sg13g2_fill_1 FILLER_7_1781 ();
 sg13g2_decap_8 FILLER_7_1787 ();
 sg13g2_fill_2 FILLER_7_1794 ();
 sg13g2_fill_1 FILLER_7_1796 ();
 sg13g2_fill_2 FILLER_7_1802 ();
 sg13g2_decap_4 FILLER_7_1809 ();
 sg13g2_fill_1 FILLER_7_1813 ();
 sg13g2_fill_2 FILLER_7_1854 ();
 sg13g2_decap_8 FILLER_7_1873 ();
 sg13g2_decap_4 FILLER_7_1880 ();
 sg13g2_fill_2 FILLER_7_1889 ();
 sg13g2_fill_1 FILLER_7_1891 ();
 sg13g2_fill_1 FILLER_7_1896 ();
 sg13g2_decap_8 FILLER_7_1933 ();
 sg13g2_fill_2 FILLER_7_1940 ();
 sg13g2_fill_2 FILLER_7_1968 ();
 sg13g2_decap_4 FILLER_7_2026 ();
 sg13g2_fill_1 FILLER_7_2082 ();
 sg13g2_fill_2 FILLER_7_2122 ();
 sg13g2_fill_1 FILLER_7_2124 ();
 sg13g2_decap_8 FILLER_7_2203 ();
 sg13g2_decap_4 FILLER_7_2210 ();
 sg13g2_fill_2 FILLER_7_2214 ();
 sg13g2_fill_2 FILLER_7_2268 ();
 sg13g2_fill_1 FILLER_7_2334 ();
 sg13g2_decap_4 FILLER_7_2390 ();
 sg13g2_fill_2 FILLER_7_2429 ();
 sg13g2_fill_1 FILLER_7_2437 ();
 sg13g2_fill_1 FILLER_7_2478 ();
 sg13g2_fill_1 FILLER_7_2505 ();
 sg13g2_fill_1 FILLER_7_2532 ();
 sg13g2_decap_4 FILLER_7_2537 ();
 sg13g2_fill_1 FILLER_7_2541 ();
 sg13g2_decap_8 FILLER_7_2552 ();
 sg13g2_decap_8 FILLER_7_2559 ();
 sg13g2_decap_8 FILLER_7_2566 ();
 sg13g2_fill_2 FILLER_7_2573 ();
 sg13g2_fill_1 FILLER_7_2575 ();
 sg13g2_fill_2 FILLER_7_2586 ();
 sg13g2_fill_1 FILLER_7_2588 ();
 sg13g2_decap_4 FILLER_7_2615 ();
 sg13g2_decap_4 FILLER_7_2665 ();
 sg13g2_fill_1 FILLER_7_2669 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_1 FILLER_8_118 ();
 sg13g2_fill_2 FILLER_8_132 ();
 sg13g2_decap_4 FILLER_8_150 ();
 sg13g2_fill_2 FILLER_8_170 ();
 sg13g2_decap_8 FILLER_8_176 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_242 ();
 sg13g2_fill_1 FILLER_8_247 ();
 sg13g2_fill_1 FILLER_8_254 ();
 sg13g2_fill_2 FILLER_8_260 ();
 sg13g2_decap_4 FILLER_8_292 ();
 sg13g2_fill_1 FILLER_8_296 ();
 sg13g2_fill_1 FILLER_8_317 ();
 sg13g2_fill_1 FILLER_8_327 ();
 sg13g2_fill_1 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_fill_1 FILLER_8_354 ();
 sg13g2_fill_1 FILLER_8_364 ();
 sg13g2_fill_2 FILLER_8_370 ();
 sg13g2_fill_1 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_381 ();
 sg13g2_decap_4 FILLER_8_419 ();
 sg13g2_fill_1 FILLER_8_474 ();
 sg13g2_fill_2 FILLER_8_484 ();
 sg13g2_fill_2 FILLER_8_500 ();
 sg13g2_fill_1 FILLER_8_519 ();
 sg13g2_fill_2 FILLER_8_543 ();
 sg13g2_fill_1 FILLER_8_585 ();
 sg13g2_fill_1 FILLER_8_626 ();
 sg13g2_decap_8 FILLER_8_631 ();
 sg13g2_decap_8 FILLER_8_638 ();
 sg13g2_fill_2 FILLER_8_645 ();
 sg13g2_fill_1 FILLER_8_647 ();
 sg13g2_fill_1 FILLER_8_693 ();
 sg13g2_decap_4 FILLER_8_737 ();
 sg13g2_fill_2 FILLER_8_755 ();
 sg13g2_fill_2 FILLER_8_788 ();
 sg13g2_fill_2 FILLER_8_808 ();
 sg13g2_fill_1 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_836 ();
 sg13g2_fill_1 FILLER_8_863 ();
 sg13g2_fill_2 FILLER_8_945 ();
 sg13g2_decap_4 FILLER_8_973 ();
 sg13g2_decap_4 FILLER_8_1003 ();
 sg13g2_fill_2 FILLER_8_1012 ();
 sg13g2_fill_1 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1019 ();
 sg13g2_fill_1 FILLER_8_1057 ();
 sg13g2_fill_2 FILLER_8_1062 ();
 sg13g2_fill_1 FILLER_8_1064 ();
 sg13g2_fill_2 FILLER_8_1091 ();
 sg13g2_fill_2 FILLER_8_1250 ();
 sg13g2_fill_2 FILLER_8_1317 ();
 sg13g2_fill_2 FILLER_8_1323 ();
 sg13g2_decap_4 FILLER_8_1335 ();
 sg13g2_fill_2 FILLER_8_1349 ();
 sg13g2_fill_2 FILLER_8_1362 ();
 sg13g2_fill_1 FILLER_8_1374 ();
 sg13g2_fill_2 FILLER_8_1404 ();
 sg13g2_fill_1 FILLER_8_1410 ();
 sg13g2_fill_1 FILLER_8_1416 ();
 sg13g2_fill_2 FILLER_8_1446 ();
 sg13g2_fill_1 FILLER_8_1448 ();
 sg13g2_decap_8 FILLER_8_1497 ();
 sg13g2_decap_8 FILLER_8_1504 ();
 sg13g2_decap_8 FILLER_8_1511 ();
 sg13g2_decap_8 FILLER_8_1518 ();
 sg13g2_fill_1 FILLER_8_1552 ();
 sg13g2_fill_2 FILLER_8_1622 ();
 sg13g2_fill_1 FILLER_8_1624 ();
 sg13g2_fill_1 FILLER_8_1635 ();
 sg13g2_fill_2 FILLER_8_1640 ();
 sg13g2_fill_1 FILLER_8_1642 ();
 sg13g2_decap_4 FILLER_8_1673 ();
 sg13g2_decap_4 FILLER_8_1713 ();
 sg13g2_fill_2 FILLER_8_1717 ();
 sg13g2_decap_4 FILLER_8_1755 ();
 sg13g2_fill_2 FILLER_8_1759 ();
 sg13g2_fill_1 FILLER_8_1805 ();
 sg13g2_fill_2 FILLER_8_1837 ();
 sg13g2_fill_1 FILLER_8_1839 ();
 sg13g2_fill_2 FILLER_8_1845 ();
 sg13g2_fill_2 FILLER_8_1851 ();
 sg13g2_fill_1 FILLER_8_1853 ();
 sg13g2_decap_8 FILLER_8_1884 ();
 sg13g2_decap_4 FILLER_8_1896 ();
 sg13g2_fill_2 FILLER_8_1904 ();
 sg13g2_decap_4 FILLER_8_1924 ();
 sg13g2_decap_8 FILLER_8_1932 ();
 sg13g2_fill_1 FILLER_8_1939 ();
 sg13g2_fill_2 FILLER_8_1950 ();
 sg13g2_fill_1 FILLER_8_1952 ();
 sg13g2_fill_2 FILLER_8_1974 ();
 sg13g2_fill_1 FILLER_8_1976 ();
 sg13g2_decap_4 FILLER_8_1991 ();
 sg13g2_fill_1 FILLER_8_1995 ();
 sg13g2_fill_2 FILLER_8_2038 ();
 sg13g2_fill_1 FILLER_8_2040 ();
 sg13g2_fill_1 FILLER_8_2090 ();
 sg13g2_decap_4 FILLER_8_2106 ();
 sg13g2_fill_1 FILLER_8_2110 ();
 sg13g2_fill_2 FILLER_8_2116 ();
 sg13g2_fill_2 FILLER_8_2154 ();
 sg13g2_fill_1 FILLER_8_2218 ();
 sg13g2_fill_2 FILLER_8_2245 ();
 sg13g2_decap_8 FILLER_8_2251 ();
 sg13g2_decap_4 FILLER_8_2258 ();
 sg13g2_fill_1 FILLER_8_2262 ();
 sg13g2_decap_4 FILLER_8_2273 ();
 sg13g2_fill_1 FILLER_8_2277 ();
 sg13g2_decap_4 FILLER_8_2282 ();
 sg13g2_fill_2 FILLER_8_2286 ();
 sg13g2_decap_8 FILLER_8_2292 ();
 sg13g2_decap_4 FILLER_8_2299 ();
 sg13g2_fill_2 FILLER_8_2307 ();
 sg13g2_fill_2 FILLER_8_2319 ();
 sg13g2_fill_2 FILLER_8_2344 ();
 sg13g2_fill_2 FILLER_8_2378 ();
 sg13g2_fill_1 FILLER_8_2380 ();
 sg13g2_fill_1 FILLER_8_2406 ();
 sg13g2_decap_4 FILLER_8_2419 ();
 sg13g2_fill_1 FILLER_8_2423 ();
 sg13g2_fill_2 FILLER_8_2429 ();
 sg13g2_decap_4 FILLER_8_2436 ();
 sg13g2_fill_2 FILLER_8_2463 ();
 sg13g2_fill_2 FILLER_8_2475 ();
 sg13g2_decap_4 FILLER_8_2503 ();
 sg13g2_fill_2 FILLER_8_2507 ();
 sg13g2_fill_1 FILLER_8_2539 ();
 sg13g2_fill_2 FILLER_8_2551 ();
 sg13g2_fill_2 FILLER_8_2579 ();
 sg13g2_fill_1 FILLER_8_2607 ();
 sg13g2_fill_2 FILLER_8_2668 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_2 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_17 ();
 sg13g2_fill_2 FILLER_9_24 ();
 sg13g2_fill_2 FILLER_9_34 ();
 sg13g2_fill_1 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_45 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_decap_8 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_8 FILLER_9_103 ();
 sg13g2_decap_4 FILLER_9_110 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_148 ();
 sg13g2_fill_1 FILLER_9_150 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_decap_8 FILLER_9_164 ();
 sg13g2_decap_4 FILLER_9_171 ();
 sg13g2_fill_1 FILLER_9_175 ();
 sg13g2_fill_1 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_fill_2 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_4 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_281 ();
 sg13g2_decap_4 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_292 ();
 sg13g2_fill_2 FILLER_9_313 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_2 FILLER_9_367 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_410 ();
 sg13g2_fill_2 FILLER_9_417 ();
 sg13g2_decap_4 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_431 ();
 sg13g2_fill_2 FILLER_9_437 ();
 sg13g2_fill_2 FILLER_9_444 ();
 sg13g2_decap_8 FILLER_9_450 ();
 sg13g2_decap_8 FILLER_9_470 ();
 sg13g2_decap_8 FILLER_9_477 ();
 sg13g2_fill_1 FILLER_9_484 ();
 sg13g2_fill_2 FILLER_9_507 ();
 sg13g2_fill_2 FILLER_9_526 ();
 sg13g2_fill_1 FILLER_9_536 ();
 sg13g2_fill_1 FILLER_9_547 ();
 sg13g2_fill_1 FILLER_9_552 ();
 sg13g2_fill_1 FILLER_9_564 ();
 sg13g2_fill_2 FILLER_9_586 ();
 sg13g2_fill_2 FILLER_9_623 ();
 sg13g2_fill_1 FILLER_9_625 ();
 sg13g2_fill_1 FILLER_9_656 ();
 sg13g2_decap_4 FILLER_9_661 ();
 sg13g2_fill_2 FILLER_9_665 ();
 sg13g2_fill_1 FILLER_9_672 ();
 sg13g2_fill_1 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_683 ();
 sg13g2_fill_1 FILLER_9_714 ();
 sg13g2_decap_4 FILLER_9_719 ();
 sg13g2_decap_4 FILLER_9_727 ();
 sg13g2_decap_4 FILLER_9_741 ();
 sg13g2_fill_1 FILLER_9_804 ();
 sg13g2_decap_8 FILLER_9_836 ();
 sg13g2_fill_1 FILLER_9_843 ();
 sg13g2_decap_4 FILLER_9_848 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_fill_1 FILLER_9_917 ();
 sg13g2_fill_1 FILLER_9_935 ();
 sg13g2_fill_1 FILLER_9_957 ();
 sg13g2_decap_8 FILLER_9_962 ();
 sg13g2_fill_1 FILLER_9_969 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1055 ();
 sg13g2_decap_4 FILLER_9_1065 ();
 sg13g2_fill_2 FILLER_9_1077 ();
 sg13g2_fill_1 FILLER_9_1079 ();
 sg13g2_fill_2 FILLER_9_1093 ();
 sg13g2_decap_8 FILLER_9_1104 ();
 sg13g2_fill_1 FILLER_9_1111 ();
 sg13g2_fill_2 FILLER_9_1116 ();
 sg13g2_fill_1 FILLER_9_1118 ();
 sg13g2_fill_1 FILLER_9_1123 ();
 sg13g2_fill_1 FILLER_9_1128 ();
 sg13g2_fill_1 FILLER_9_1134 ();
 sg13g2_fill_1 FILLER_9_1139 ();
 sg13g2_fill_2 FILLER_9_1206 ();
 sg13g2_fill_1 FILLER_9_1221 ();
 sg13g2_fill_1 FILLER_9_1227 ();
 sg13g2_fill_2 FILLER_9_1233 ();
 sg13g2_fill_1 FILLER_9_1235 ();
 sg13g2_fill_2 FILLER_9_1269 ();
 sg13g2_decap_8 FILLER_9_1289 ();
 sg13g2_fill_2 FILLER_9_1296 ();
 sg13g2_decap_8 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1309 ();
 sg13g2_decap_8 FILLER_9_1316 ();
 sg13g2_decap_4 FILLER_9_1323 ();
 sg13g2_fill_1 FILLER_9_1327 ();
 sg13g2_fill_1 FILLER_9_1366 ();
 sg13g2_fill_1 FILLER_9_1370 ();
 sg13g2_fill_1 FILLER_9_1375 ();
 sg13g2_fill_2 FILLER_9_1389 ();
 sg13g2_fill_1 FILLER_9_1417 ();
 sg13g2_fill_2 FILLER_9_1423 ();
 sg13g2_fill_2 FILLER_9_1429 ();
 sg13g2_fill_2 FILLER_9_1457 ();
 sg13g2_fill_1 FILLER_9_1467 ();
 sg13g2_fill_1 FILLER_9_1504 ();
 sg13g2_decap_8 FILLER_9_1508 ();
 sg13g2_decap_8 FILLER_9_1515 ();
 sg13g2_fill_1 FILLER_9_1522 ();
 sg13g2_fill_2 FILLER_9_1580 ();
 sg13g2_fill_1 FILLER_9_1582 ();
 sg13g2_fill_2 FILLER_9_1593 ();
 sg13g2_fill_2 FILLER_9_1599 ();
 sg13g2_fill_1 FILLER_9_1601 ();
 sg13g2_decap_4 FILLER_9_1648 ();
 sg13g2_fill_2 FILLER_9_1656 ();
 sg13g2_decap_4 FILLER_9_1710 ();
 sg13g2_decap_8 FILLER_9_1750 ();
 sg13g2_fill_1 FILLER_9_1757 ();
 sg13g2_fill_1 FILLER_9_1767 ();
 sg13g2_fill_2 FILLER_9_1788 ();
 sg13g2_fill_1 FILLER_9_1790 ();
 sg13g2_fill_2 FILLER_9_1801 ();
 sg13g2_fill_2 FILLER_9_1808 ();
 sg13g2_fill_1 FILLER_9_1810 ();
 sg13g2_decap_8 FILLER_9_1880 ();
 sg13g2_decap_8 FILLER_9_1887 ();
 sg13g2_decap_8 FILLER_9_1894 ();
 sg13g2_fill_2 FILLER_9_1901 ();
 sg13g2_fill_1 FILLER_9_1903 ();
 sg13g2_fill_2 FILLER_9_1930 ();
 sg13g2_fill_1 FILLER_9_1932 ();
 sg13g2_fill_2 FILLER_9_1937 ();
 sg13g2_decap_8 FILLER_9_1975 ();
 sg13g2_decap_8 FILLER_9_1982 ();
 sg13g2_decap_8 FILLER_9_1989 ();
 sg13g2_decap_8 FILLER_9_1996 ();
 sg13g2_decap_8 FILLER_9_2003 ();
 sg13g2_decap_8 FILLER_9_2010 ();
 sg13g2_fill_2 FILLER_9_2017 ();
 sg13g2_fill_1 FILLER_9_2019 ();
 sg13g2_decap_4 FILLER_9_2034 ();
 sg13g2_decap_4 FILLER_9_2042 ();
 sg13g2_fill_2 FILLER_9_2046 ();
 sg13g2_decap_8 FILLER_9_2052 ();
 sg13g2_decap_8 FILLER_9_2059 ();
 sg13g2_decap_4 FILLER_9_2066 ();
 sg13g2_fill_2 FILLER_9_2070 ();
 sg13g2_decap_8 FILLER_9_2076 ();
 sg13g2_fill_2 FILLER_9_2092 ();
 sg13g2_fill_2 FILLER_9_2133 ();
 sg13g2_fill_1 FILLER_9_2135 ();
 sg13g2_fill_2 FILLER_9_2140 ();
 sg13g2_fill_2 FILLER_9_2181 ();
 sg13g2_decap_4 FILLER_9_2205 ();
 sg13g2_fill_1 FILLER_9_2209 ();
 sg13g2_fill_1 FILLER_9_2244 ();
 sg13g2_decap_4 FILLER_9_2276 ();
 sg13g2_fill_2 FILLER_9_2336 ();
 sg13g2_decap_8 FILLER_9_2365 ();
 sg13g2_decap_8 FILLER_9_2372 ();
 sg13g2_fill_1 FILLER_9_2379 ();
 sg13g2_decap_8 FILLER_9_2384 ();
 sg13g2_fill_2 FILLER_9_2391 ();
 sg13g2_fill_1 FILLER_9_2393 ();
 sg13g2_decap_4 FILLER_9_2409 ();
 sg13g2_fill_1 FILLER_9_2453 ();
 sg13g2_fill_1 FILLER_9_2523 ();
 sg13g2_fill_1 FILLER_9_2568 ();
 sg13g2_fill_1 FILLER_9_2579 ();
 sg13g2_fill_1 FILLER_9_2590 ();
 sg13g2_fill_1 FILLER_9_2595 ();
 sg13g2_fill_2 FILLER_9_2600 ();
 sg13g2_decap_8 FILLER_9_2661 ();
 sg13g2_fill_2 FILLER_9_2668 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_decap_8 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_94 ();
 sg13g2_decap_8 FILLER_10_104 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_125 ();
 sg13g2_fill_1 FILLER_10_127 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_decap_4 FILLER_10_152 ();
 sg13g2_fill_2 FILLER_10_156 ();
 sg13g2_fill_2 FILLER_10_162 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_2 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_253 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_344 ();
 sg13g2_decap_4 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_fill_2 FILLER_10_393 ();
 sg13g2_fill_1 FILLER_10_395 ();
 sg13g2_decap_4 FILLER_10_400 ();
 sg13g2_fill_1 FILLER_10_404 ();
 sg13g2_decap_4 FILLER_10_409 ();
 sg13g2_fill_1 FILLER_10_413 ();
 sg13g2_decap_4 FILLER_10_418 ();
 sg13g2_fill_1 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_fill_2 FILLER_10_452 ();
 sg13g2_fill_1 FILLER_10_480 ();
 sg13g2_fill_2 FILLER_10_491 ();
 sg13g2_fill_2 FILLER_10_528 ();
 sg13g2_fill_2 FILLER_10_538 ();
 sg13g2_decap_4 FILLER_10_595 ();
 sg13g2_fill_2 FILLER_10_599 ();
 sg13g2_fill_2 FILLER_10_605 ();
 sg13g2_fill_1 FILLER_10_607 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_4 FILLER_10_620 ();
 sg13g2_fill_2 FILLER_10_624 ();
 sg13g2_fill_2 FILLER_10_635 ();
 sg13g2_fill_1 FILLER_10_637 ();
 sg13g2_fill_1 FILLER_10_642 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_4 FILLER_10_700 ();
 sg13g2_fill_1 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_8 FILLER_10_737 ();
 sg13g2_decap_8 FILLER_10_744 ();
 sg13g2_fill_1 FILLER_10_751 ();
 sg13g2_fill_2 FILLER_10_760 ();
 sg13g2_fill_1 FILLER_10_771 ();
 sg13g2_fill_2 FILLER_10_776 ();
 sg13g2_fill_2 FILLER_10_788 ();
 sg13g2_fill_1 FILLER_10_796 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_fill_2 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_888 ();
 sg13g2_decap_8 FILLER_10_895 ();
 sg13g2_decap_8 FILLER_10_902 ();
 sg13g2_decap_8 FILLER_10_909 ();
 sg13g2_fill_1 FILLER_10_916 ();
 sg13g2_fill_2 FILLER_10_922 ();
 sg13g2_fill_2 FILLER_10_933 ();
 sg13g2_decap_8 FILLER_10_948 ();
 sg13g2_decap_4 FILLER_10_955 ();
 sg13g2_fill_2 FILLER_10_959 ();
 sg13g2_decap_4 FILLER_10_970 ();
 sg13g2_fill_2 FILLER_10_974 ();
 sg13g2_fill_1 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1011 ();
 sg13g2_decap_8 FILLER_10_1018 ();
 sg13g2_decap_4 FILLER_10_1025 ();
 sg13g2_fill_2 FILLER_10_1029 ();
 sg13g2_fill_1 FILLER_10_1057 ();
 sg13g2_fill_1 FILLER_10_1063 ();
 sg13g2_fill_1 FILLER_10_1068 ();
 sg13g2_fill_1 FILLER_10_1074 ();
 sg13g2_fill_1 FILLER_10_1079 ();
 sg13g2_fill_2 FILLER_10_1088 ();
 sg13g2_fill_1 FILLER_10_1095 ();
 sg13g2_fill_2 FILLER_10_1105 ();
 sg13g2_fill_2 FILLER_10_1168 ();
 sg13g2_fill_2 FILLER_10_1174 ();
 sg13g2_fill_1 FILLER_10_1181 ();
 sg13g2_fill_1 FILLER_10_1186 ();
 sg13g2_fill_1 FILLER_10_1208 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_decap_8 FILLER_10_1246 ();
 sg13g2_fill_2 FILLER_10_1253 ();
 sg13g2_decap_8 FILLER_10_1265 ();
 sg13g2_decap_8 FILLER_10_1272 ();
 sg13g2_decap_8 FILLER_10_1279 ();
 sg13g2_fill_1 FILLER_10_1286 ();
 sg13g2_decap_8 FILLER_10_1296 ();
 sg13g2_decap_8 FILLER_10_1303 ();
 sg13g2_decap_8 FILLER_10_1310 ();
 sg13g2_decap_8 FILLER_10_1317 ();
 sg13g2_decap_8 FILLER_10_1324 ();
 sg13g2_decap_8 FILLER_10_1331 ();
 sg13g2_decap_8 FILLER_10_1338 ();
 sg13g2_decap_8 FILLER_10_1345 ();
 sg13g2_fill_1 FILLER_10_1352 ();
 sg13g2_fill_1 FILLER_10_1397 ();
 sg13g2_decap_8 FILLER_10_1410 ();
 sg13g2_decap_8 FILLER_10_1417 ();
 sg13g2_decap_8 FILLER_10_1424 ();
 sg13g2_decap_4 FILLER_10_1474 ();
 sg13g2_fill_1 FILLER_10_1478 ();
 sg13g2_decap_8 FILLER_10_1483 ();
 sg13g2_decap_4 FILLER_10_1490 ();
 sg13g2_fill_2 FILLER_10_1494 ();
 sg13g2_fill_1 FILLER_10_1502 ();
 sg13g2_fill_2 FILLER_10_1506 ();
 sg13g2_fill_2 FILLER_10_1548 ();
 sg13g2_fill_2 FILLER_10_1559 ();
 sg13g2_decap_8 FILLER_10_1587 ();
 sg13g2_decap_8 FILLER_10_1594 ();
 sg13g2_decap_8 FILLER_10_1601 ();
 sg13g2_decap_8 FILLER_10_1608 ();
 sg13g2_decap_8 FILLER_10_1615 ();
 sg13g2_decap_8 FILLER_10_1622 ();
 sg13g2_decap_8 FILLER_10_1629 ();
 sg13g2_decap_4 FILLER_10_1636 ();
 sg13g2_decap_8 FILLER_10_1662 ();
 sg13g2_decap_4 FILLER_10_1669 ();
 sg13g2_fill_2 FILLER_10_1673 ();
 sg13g2_fill_2 FILLER_10_1711 ();
 sg13g2_fill_1 FILLER_10_1713 ();
 sg13g2_fill_2 FILLER_10_1740 ();
 sg13g2_fill_2 FILLER_10_1766 ();
 sg13g2_fill_1 FILLER_10_1812 ();
 sg13g2_fill_2 FILLER_10_1826 ();
 sg13g2_decap_4 FILLER_10_1833 ();
 sg13g2_fill_2 FILLER_10_1847 ();
 sg13g2_fill_1 FILLER_10_1849 ();
 sg13g2_fill_2 FILLER_10_1854 ();
 sg13g2_fill_2 FILLER_10_1882 ();
 sg13g2_fill_1 FILLER_10_1884 ();
 sg13g2_decap_8 FILLER_10_1970 ();
 sg13g2_decap_4 FILLER_10_1977 ();
 sg13g2_fill_2 FILLER_10_1981 ();
 sg13g2_decap_8 FILLER_10_2030 ();
 sg13g2_decap_8 FILLER_10_2037 ();
 sg13g2_fill_2 FILLER_10_2044 ();
 sg13g2_decap_4 FILLER_10_2077 ();
 sg13g2_fill_2 FILLER_10_2081 ();
 sg13g2_decap_8 FILLER_10_2114 ();
 sg13g2_decap_8 FILLER_10_2121 ();
 sg13g2_decap_8 FILLER_10_2128 ();
 sg13g2_fill_2 FILLER_10_2135 ();
 sg13g2_fill_1 FILLER_10_2137 ();
 sg13g2_decap_8 FILLER_10_2142 ();
 sg13g2_decap_8 FILLER_10_2149 ();
 sg13g2_decap_8 FILLER_10_2156 ();
 sg13g2_decap_8 FILLER_10_2163 ();
 sg13g2_decap_8 FILLER_10_2170 ();
 sg13g2_decap_8 FILLER_10_2177 ();
 sg13g2_decap_8 FILLER_10_2184 ();
 sg13g2_decap_8 FILLER_10_2191 ();
 sg13g2_decap_8 FILLER_10_2198 ();
 sg13g2_fill_2 FILLER_10_2205 ();
 sg13g2_fill_1 FILLER_10_2207 ();
 sg13g2_decap_8 FILLER_10_2242 ();
 sg13g2_decap_8 FILLER_10_2249 ();
 sg13g2_fill_1 FILLER_10_2256 ();
 sg13g2_decap_8 FILLER_10_2293 ();
 sg13g2_fill_1 FILLER_10_2300 ();
 sg13g2_fill_2 FILLER_10_2327 ();
 sg13g2_fill_2 FILLER_10_2344 ();
 sg13g2_fill_2 FILLER_10_2377 ();
 sg13g2_fill_1 FILLER_10_2379 ();
 sg13g2_fill_2 FILLER_10_2390 ();
 sg13g2_fill_1 FILLER_10_2396 ();
 sg13g2_decap_8 FILLER_10_2402 ();
 sg13g2_fill_2 FILLER_10_2409 ();
 sg13g2_fill_1 FILLER_10_2411 ();
 sg13g2_fill_2 FILLER_10_2448 ();
 sg13g2_fill_1 FILLER_10_2450 ();
 sg13g2_decap_8 FILLER_10_2461 ();
 sg13g2_decap_4 FILLER_10_2472 ();
 sg13g2_fill_1 FILLER_10_2476 ();
 sg13g2_decap_8 FILLER_10_2483 ();
 sg13g2_decap_8 FILLER_10_2490 ();
 sg13g2_fill_2 FILLER_10_2497 ();
 sg13g2_fill_1 FILLER_10_2499 ();
 sg13g2_fill_1 FILLER_10_2520 ();
 sg13g2_decap_8 FILLER_10_2536 ();
 sg13g2_decap_8 FILLER_10_2543 ();
 sg13g2_fill_1 FILLER_10_2550 ();
 sg13g2_fill_2 FILLER_10_2561 ();
 sg13g2_fill_1 FILLER_10_2567 ();
 sg13g2_decap_4 FILLER_10_2574 ();
 sg13g2_fill_2 FILLER_10_2578 ();
 sg13g2_decap_8 FILLER_10_2585 ();
 sg13g2_fill_2 FILLER_10_2592 ();
 sg13g2_fill_1 FILLER_10_2608 ();
 sg13g2_decap_4 FILLER_10_2616 ();
 sg13g2_fill_2 FILLER_10_2636 ();
 sg13g2_fill_1 FILLER_10_2641 ();
 sg13g2_fill_2 FILLER_10_2668 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_fill_1 FILLER_11_56 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_136 ();
 sg13g2_fill_1 FILLER_11_152 ();
 sg13g2_fill_1 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_267 ();
 sg13g2_fill_2 FILLER_11_319 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_fill_2 FILLER_11_385 ();
 sg13g2_fill_1 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_397 ();
 sg13g2_decap_8 FILLER_11_451 ();
 sg13g2_decap_4 FILLER_11_458 ();
 sg13g2_fill_2 FILLER_11_462 ();
 sg13g2_fill_1 FILLER_11_490 ();
 sg13g2_fill_2 FILLER_11_505 ();
 sg13g2_fill_2 FILLER_11_523 ();
 sg13g2_fill_1 FILLER_11_551 ();
 sg13g2_fill_1 FILLER_11_556 ();
 sg13g2_fill_1 FILLER_11_592 ();
 sg13g2_fill_1 FILLER_11_598 ();
 sg13g2_fill_2 FILLER_11_608 ();
 sg13g2_fill_2 FILLER_11_614 ();
 sg13g2_fill_1 FILLER_11_647 ();
 sg13g2_decap_8 FILLER_11_674 ();
 sg13g2_decap_4 FILLER_11_681 ();
 sg13g2_fill_2 FILLER_11_685 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_fill_2 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_737 ();
 sg13g2_decap_8 FILLER_11_744 ();
 sg13g2_decap_8 FILLER_11_751 ();
 sg13g2_decap_4 FILLER_11_758 ();
 sg13g2_fill_1 FILLER_11_777 ();
 sg13g2_fill_2 FILLER_11_783 ();
 sg13g2_fill_1 FILLER_11_789 ();
 sg13g2_fill_2 FILLER_11_843 ();
 sg13g2_fill_1 FILLER_11_845 ();
 sg13g2_fill_2 FILLER_11_874 ();
 sg13g2_fill_2 FILLER_11_908 ();
 sg13g2_fill_1 FILLER_11_910 ();
 sg13g2_fill_1 FILLER_11_924 ();
 sg13g2_fill_2 FILLER_11_951 ();
 sg13g2_fill_1 FILLER_11_953 ();
 sg13g2_decap_4 FILLER_11_1084 ();
 sg13g2_fill_2 FILLER_11_1088 ();
 sg13g2_fill_2 FILLER_11_1137 ();
 sg13g2_fill_1 FILLER_11_1139 ();
 sg13g2_fill_2 FILLER_11_1175 ();
 sg13g2_decap_4 FILLER_11_1181 ();
 sg13g2_fill_1 FILLER_11_1189 ();
 sg13g2_fill_1 FILLER_11_1197 ();
 sg13g2_fill_2 FILLER_11_1245 ();
 sg13g2_fill_2 FILLER_11_1309 ();
 sg13g2_fill_1 FILLER_11_1311 ();
 sg13g2_decap_4 FILLER_11_1338 ();
 sg13g2_fill_2 FILLER_11_1342 ();
 sg13g2_fill_1 FILLER_11_1374 ();
 sg13g2_fill_2 FILLER_11_1380 ();
 sg13g2_fill_2 FILLER_11_1399 ();
 sg13g2_fill_1 FILLER_11_1401 ();
 sg13g2_fill_2 FILLER_11_1409 ();
 sg13g2_decap_8 FILLER_11_1419 ();
 sg13g2_decap_8 FILLER_11_1426 ();
 sg13g2_fill_2 FILLER_11_1453 ();
 sg13g2_decap_8 FILLER_11_1477 ();
 sg13g2_decap_4 FILLER_11_1484 ();
 sg13g2_fill_2 FILLER_11_1525 ();
 sg13g2_decap_8 FILLER_11_1530 ();
 sg13g2_decap_8 FILLER_11_1537 ();
 sg13g2_decap_4 FILLER_11_1544 ();
 sg13g2_fill_2 FILLER_11_1548 ();
 sg13g2_decap_8 FILLER_11_1566 ();
 sg13g2_decap_4 FILLER_11_1573 ();
 sg13g2_decap_8 FILLER_11_1582 ();
 sg13g2_fill_2 FILLER_11_1589 ();
 sg13g2_decap_8 FILLER_11_1601 ();
 sg13g2_decap_8 FILLER_11_1608 ();
 sg13g2_decap_4 FILLER_11_1615 ();
 sg13g2_fill_1 FILLER_11_1619 ();
 sg13g2_fill_1 FILLER_11_1639 ();
 sg13g2_fill_2 FILLER_11_1645 ();
 sg13g2_fill_1 FILLER_11_1659 ();
 sg13g2_decap_4 FILLER_11_1686 ();
 sg13g2_fill_1 FILLER_11_1690 ();
 sg13g2_fill_1 FILLER_11_1695 ();
 sg13g2_fill_2 FILLER_11_1700 ();
 sg13g2_decap_8 FILLER_11_1706 ();
 sg13g2_decap_8 FILLER_11_1713 ();
 sg13g2_fill_2 FILLER_11_1780 ();
 sg13g2_decap_4 FILLER_11_1813 ();
 sg13g2_fill_1 FILLER_11_1817 ();
 sg13g2_fill_1 FILLER_11_1839 ();
 sg13g2_fill_2 FILLER_11_1846 ();
 sg13g2_decap_8 FILLER_11_1852 ();
 sg13g2_decap_8 FILLER_11_1859 ();
 sg13g2_decap_4 FILLER_11_1887 ();
 sg13g2_fill_1 FILLER_11_1891 ();
 sg13g2_fill_1 FILLER_11_1899 ();
 sg13g2_fill_1 FILLER_11_1947 ();
 sg13g2_fill_2 FILLER_11_1974 ();
 sg13g2_fill_2 FILLER_11_2002 ();
 sg13g2_fill_1 FILLER_11_2030 ();
 sg13g2_decap_4 FILLER_11_2067 ();
 sg13g2_fill_2 FILLER_11_2092 ();
 sg13g2_fill_1 FILLER_11_2094 ();
 sg13g2_decap_4 FILLER_11_2121 ();
 sg13g2_fill_2 FILLER_11_2125 ();
 sg13g2_fill_2 FILLER_11_2137 ();
 sg13g2_fill_1 FILLER_11_2139 ();
 sg13g2_decap_4 FILLER_11_2161 ();
 sg13g2_fill_2 FILLER_11_2165 ();
 sg13g2_decap_8 FILLER_11_2201 ();
 sg13g2_decap_8 FILLER_11_2208 ();
 sg13g2_decap_8 FILLER_11_2215 ();
 sg13g2_decap_8 FILLER_11_2222 ();
 sg13g2_fill_2 FILLER_11_2229 ();
 sg13g2_fill_1 FILLER_11_2239 ();
 sg13g2_decap_8 FILLER_11_2289 ();
 sg13g2_decap_4 FILLER_11_2296 ();
 sg13g2_fill_1 FILLER_11_2300 ();
 sg13g2_fill_1 FILLER_11_2337 ();
 sg13g2_decap_8 FILLER_11_2341 ();
 sg13g2_decap_8 FILLER_11_2348 ();
 sg13g2_decap_4 FILLER_11_2355 ();
 sg13g2_fill_2 FILLER_11_2359 ();
 sg13g2_decap_4 FILLER_11_2371 ();
 sg13g2_fill_1 FILLER_11_2375 ();
 sg13g2_fill_1 FILLER_11_2412 ();
 sg13g2_decap_8 FILLER_11_2417 ();
 sg13g2_decap_4 FILLER_11_2424 ();
 sg13g2_fill_1 FILLER_11_2428 ();
 sg13g2_decap_8 FILLER_11_2446 ();
 sg13g2_decap_8 FILLER_11_2502 ();
 sg13g2_fill_2 FILLER_11_2509 ();
 sg13g2_fill_1 FILLER_11_2511 ();
 sg13g2_decap_8 FILLER_11_2542 ();
 sg13g2_decap_8 FILLER_11_2549 ();
 sg13g2_decap_8 FILLER_11_2556 ();
 sg13g2_decap_4 FILLER_11_2563 ();
 sg13g2_fill_2 FILLER_11_2567 ();
 sg13g2_fill_2 FILLER_11_2582 ();
 sg13g2_fill_1 FILLER_11_2584 ();
 sg13g2_fill_1 FILLER_11_2620 ();
 sg13g2_decap_8 FILLER_11_2661 ();
 sg13g2_fill_2 FILLER_11_2668 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_41 ();
 sg13g2_fill_2 FILLER_12_48 ();
 sg13g2_fill_1 FILLER_12_50 ();
 sg13g2_fill_2 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_145 ();
 sg13g2_fill_2 FILLER_12_173 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_decap_8 FILLER_12_279 ();
 sg13g2_decap_4 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_fill_2 FILLER_12_340 ();
 sg13g2_fill_1 FILLER_12_430 ();
 sg13g2_fill_2 FILLER_12_457 ();
 sg13g2_fill_1 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_464 ();
 sg13g2_decap_8 FILLER_12_471 ();
 sg13g2_fill_2 FILLER_12_521 ();
 sg13g2_fill_1 FILLER_12_583 ();
 sg13g2_fill_2 FILLER_12_614 ();
 sg13g2_fill_1 FILLER_12_629 ();
 sg13g2_fill_1 FILLER_12_649 ();
 sg13g2_fill_1 FILLER_12_668 ();
 sg13g2_fill_2 FILLER_12_675 ();
 sg13g2_fill_2 FILLER_12_694 ();
 sg13g2_fill_2 FILLER_12_700 ();
 sg13g2_fill_1 FILLER_12_707 ();
 sg13g2_fill_2 FILLER_12_713 ();
 sg13g2_fill_2 FILLER_12_801 ();
 sg13g2_fill_2 FILLER_12_806 ();
 sg13g2_fill_2 FILLER_12_814 ();
 sg13g2_fill_1 FILLER_12_829 ();
 sg13g2_decap_4 FILLER_12_867 ();
 sg13g2_fill_2 FILLER_12_871 ();
 sg13g2_decap_4 FILLER_12_915 ();
 sg13g2_fill_1 FILLER_12_919 ();
 sg13g2_decap_8 FILLER_12_971 ();
 sg13g2_fill_1 FILLER_12_978 ();
 sg13g2_decap_8 FILLER_12_1000 ();
 sg13g2_decap_8 FILLER_12_1007 ();
 sg13g2_decap_8 FILLER_12_1018 ();
 sg13g2_decap_8 FILLER_12_1025 ();
 sg13g2_decap_4 FILLER_12_1032 ();
 sg13g2_fill_1 FILLER_12_1044 ();
 sg13g2_fill_2 FILLER_12_1054 ();
 sg13g2_fill_1 FILLER_12_1056 ();
 sg13g2_fill_2 FILLER_12_1087 ();
 sg13g2_fill_1 FILLER_12_1089 ();
 sg13g2_decap_8 FILLER_12_1125 ();
 sg13g2_decap_8 FILLER_12_1132 ();
 sg13g2_decap_8 FILLER_12_1139 ();
 sg13g2_decap_4 FILLER_12_1146 ();
 sg13g2_fill_1 FILLER_12_1167 ();
 sg13g2_decap_8 FILLER_12_1180 ();
 sg13g2_fill_1 FILLER_12_1187 ();
 sg13g2_fill_2 FILLER_12_1196 ();
 sg13g2_fill_1 FILLER_12_1198 ();
 sg13g2_fill_1 FILLER_12_1208 ();
 sg13g2_decap_4 FILLER_12_1227 ();
 sg13g2_fill_1 FILLER_12_1231 ();
 sg13g2_decap_8 FILLER_12_1284 ();
 sg13g2_decap_8 FILLER_12_1291 ();
 sg13g2_decap_8 FILLER_12_1298 ();
 sg13g2_fill_2 FILLER_12_1305 ();
 sg13g2_fill_1 FILLER_12_1321 ();
 sg13g2_fill_1 FILLER_12_1348 ();
 sg13g2_fill_1 FILLER_12_1354 ();
 sg13g2_decap_8 FILLER_12_1359 ();
 sg13g2_decap_4 FILLER_12_1366 ();
 sg13g2_fill_2 FILLER_12_1373 ();
 sg13g2_fill_2 FILLER_12_1380 ();
 sg13g2_fill_1 FILLER_12_1386 ();
 sg13g2_fill_2 FILLER_12_1402 ();
 sg13g2_fill_2 FILLER_12_1409 ();
 sg13g2_fill_1 FILLER_12_1411 ();
 sg13g2_fill_2 FILLER_12_1417 ();
 sg13g2_fill_2 FILLER_12_1426 ();
 sg13g2_fill_1 FILLER_12_1428 ();
 sg13g2_fill_1 FILLER_12_1434 ();
 sg13g2_fill_1 FILLER_12_1495 ();
 sg13g2_fill_2 FILLER_12_1501 ();
 sg13g2_fill_2 FILLER_12_1605 ();
 sg13g2_decap_4 FILLER_12_1622 ();
 sg13g2_fill_2 FILLER_12_1626 ();
 sg13g2_fill_1 FILLER_12_1650 ();
 sg13g2_decap_8 FILLER_12_1656 ();
 sg13g2_decap_4 FILLER_12_1663 ();
 sg13g2_fill_2 FILLER_12_1667 ();
 sg13g2_decap_8 FILLER_12_1683 ();
 sg13g2_decap_8 FILLER_12_1690 ();
 sg13g2_decap_8 FILLER_12_1697 ();
 sg13g2_decap_8 FILLER_12_1704 ();
 sg13g2_decap_8 FILLER_12_1711 ();
 sg13g2_fill_2 FILLER_12_1718 ();
 sg13g2_fill_2 FILLER_12_1724 ();
 sg13g2_fill_2 FILLER_12_1730 ();
 sg13g2_fill_1 FILLER_12_1732 ();
 sg13g2_fill_2 FILLER_12_1737 ();
 sg13g2_fill_1 FILLER_12_1739 ();
 sg13g2_fill_2 FILLER_12_1745 ();
 sg13g2_fill_1 FILLER_12_1747 ();
 sg13g2_fill_2 FILLER_12_1758 ();
 sg13g2_fill_1 FILLER_12_1760 ();
 sg13g2_fill_2 FILLER_12_1779 ();
 sg13g2_fill_1 FILLER_12_1781 ();
 sg13g2_decap_4 FILLER_12_1786 ();
 sg13g2_fill_1 FILLER_12_1805 ();
 sg13g2_fill_2 FILLER_12_1811 ();
 sg13g2_fill_1 FILLER_12_1836 ();
 sg13g2_decap_8 FILLER_12_1889 ();
 sg13g2_fill_2 FILLER_12_1896 ();
 sg13g2_fill_1 FILLER_12_1921 ();
 sg13g2_fill_2 FILLER_12_1934 ();
 sg13g2_fill_1 FILLER_12_1936 ();
 sg13g2_fill_2 FILLER_12_1945 ();
 sg13g2_fill_2 FILLER_12_1997 ();
 sg13g2_fill_1 FILLER_12_2087 ();
 sg13g2_fill_2 FILLER_12_2118 ();
 sg13g2_fill_1 FILLER_12_2120 ();
 sg13g2_fill_2 FILLER_12_2161 ();
 sg13g2_fill_2 FILLER_12_2199 ();
 sg13g2_fill_1 FILLER_12_2201 ();
 sg13g2_decap_8 FILLER_12_2254 ();
 sg13g2_fill_2 FILLER_12_2261 ();
 sg13g2_fill_1 FILLER_12_2276 ();
 sg13g2_decap_4 FILLER_12_2303 ();
 sg13g2_fill_2 FILLER_12_2307 ();
 sg13g2_decap_4 FILLER_12_2313 ();
 sg13g2_decap_8 FILLER_12_2321 ();
 sg13g2_decap_8 FILLER_12_2328 ();
 sg13g2_decap_4 FILLER_12_2335 ();
 sg13g2_fill_2 FILLER_12_2339 ();
 sg13g2_fill_2 FILLER_12_2346 ();
 sg13g2_fill_2 FILLER_12_2456 ();
 sg13g2_decap_8 FILLER_12_2467 ();
 sg13g2_decap_4 FILLER_12_2474 ();
 sg13g2_decap_4 FILLER_12_2514 ();
 sg13g2_fill_1 FILLER_12_2518 ();
 sg13g2_fill_2 FILLER_12_2529 ();
 sg13g2_decap_8 FILLER_12_2535 ();
 sg13g2_decap_4 FILLER_12_2542 ();
 sg13g2_fill_1 FILLER_12_2546 ();
 sg13g2_fill_2 FILLER_12_2573 ();
 sg13g2_fill_1 FILLER_12_2575 ();
 sg13g2_fill_1 FILLER_12_2641 ();
 sg13g2_fill_2 FILLER_12_2668 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_12 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_66 ();
 sg13g2_fill_2 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_102 ();
 sg13g2_decap_4 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_decap_8 FILLER_13_166 ();
 sg13g2_decap_4 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_177 ();
 sg13g2_fill_1 FILLER_13_190 ();
 sg13g2_fill_2 FILLER_13_230 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_298 ();
 sg13g2_decap_4 FILLER_13_322 ();
 sg13g2_fill_1 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_382 ();
 sg13g2_fill_1 FILLER_13_388 ();
 sg13g2_decap_4 FILLER_13_394 ();
 sg13g2_fill_2 FILLER_13_398 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_fill_1 FILLER_13_417 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_decap_4 FILLER_13_434 ();
 sg13g2_fill_1 FILLER_13_477 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_fill_1 FILLER_13_538 ();
 sg13g2_fill_1 FILLER_13_573 ();
 sg13g2_fill_1 FILLER_13_587 ();
 sg13g2_fill_1 FILLER_13_627 ();
 sg13g2_decap_4 FILLER_13_637 ();
 sg13g2_fill_2 FILLER_13_650 ();
 sg13g2_fill_1 FILLER_13_687 ();
 sg13g2_fill_2 FILLER_13_700 ();
 sg13g2_decap_4 FILLER_13_713 ();
 sg13g2_fill_2 FILLER_13_717 ();
 sg13g2_fill_1 FILLER_13_723 ();
 sg13g2_fill_1 FILLER_13_729 ();
 sg13g2_decap_4 FILLER_13_739 ();
 sg13g2_fill_1 FILLER_13_743 ();
 sg13g2_fill_1 FILLER_13_754 ();
 sg13g2_fill_2 FILLER_13_768 ();
 sg13g2_fill_1 FILLER_13_819 ();
 sg13g2_fill_2 FILLER_13_827 ();
 sg13g2_fill_1 FILLER_13_837 ();
 sg13g2_decap_4 FILLER_13_841 ();
 sg13g2_fill_2 FILLER_13_845 ();
 sg13g2_fill_2 FILLER_13_873 ();
 sg13g2_decap_8 FILLER_13_947 ();
 sg13g2_decap_8 FILLER_13_954 ();
 sg13g2_fill_2 FILLER_13_987 ();
 sg13g2_fill_1 FILLER_13_989 ();
 sg13g2_decap_8 FILLER_13_1024 ();
 sg13g2_decap_8 FILLER_13_1031 ();
 sg13g2_decap_4 FILLER_13_1038 ();
 sg13g2_decap_4 FILLER_13_1046 ();
 sg13g2_fill_1 FILLER_13_1050 ();
 sg13g2_fill_2 FILLER_13_1060 ();
 sg13g2_fill_1 FILLER_13_1062 ();
 sg13g2_decap_8 FILLER_13_1084 ();
 sg13g2_decap_4 FILLER_13_1091 ();
 sg13g2_fill_2 FILLER_13_1095 ();
 sg13g2_decap_8 FILLER_13_1105 ();
 sg13g2_decap_4 FILLER_13_1112 ();
 sg13g2_fill_1 FILLER_13_1116 ();
 sg13g2_decap_4 FILLER_13_1122 ();
 sg13g2_decap_8 FILLER_13_1131 ();
 sg13g2_fill_2 FILLER_13_1142 ();
 sg13g2_fill_1 FILLER_13_1144 ();
 sg13g2_decap_4 FILLER_13_1166 ();
 sg13g2_fill_2 FILLER_13_1170 ();
 sg13g2_fill_2 FILLER_13_1213 ();
 sg13g2_decap_4 FILLER_13_1270 ();
 sg13g2_fill_1 FILLER_13_1274 ();
 sg13g2_decap_4 FILLER_13_1314 ();
 sg13g2_fill_1 FILLER_13_1318 ();
 sg13g2_decap_8 FILLER_13_1337 ();
 sg13g2_fill_1 FILLER_13_1344 ();
 sg13g2_decap_8 FILLER_13_1379 ();
 sg13g2_fill_2 FILLER_13_1415 ();
 sg13g2_decap_4 FILLER_13_1442 ();
 sg13g2_fill_2 FILLER_13_1446 ();
 sg13g2_fill_1 FILLER_13_1452 ();
 sg13g2_fill_1 FILLER_13_1458 ();
 sg13g2_fill_1 FILLER_13_1535 ();
 sg13g2_decap_4 FILLER_13_1546 ();
 sg13g2_fill_2 FILLER_13_1554 ();
 sg13g2_fill_2 FILLER_13_1562 ();
 sg13g2_fill_1 FILLER_13_1585 ();
 sg13g2_fill_2 FILLER_13_1596 ();
 sg13g2_fill_1 FILLER_13_1614 ();
 sg13g2_fill_2 FILLER_13_1637 ();
 sg13g2_fill_2 FILLER_13_1666 ();
 sg13g2_fill_1 FILLER_13_1668 ();
 sg13g2_decap_8 FILLER_13_1675 ();
 sg13g2_decap_8 FILLER_13_1682 ();
 sg13g2_fill_1 FILLER_13_1689 ();
 sg13g2_fill_1 FILLER_13_1699 ();
 sg13g2_fill_1 FILLER_13_1710 ();
 sg13g2_fill_2 FILLER_13_1715 ();
 sg13g2_fill_1 FILLER_13_1717 ();
 sg13g2_fill_1 FILLER_13_1723 ();
 sg13g2_decap_4 FILLER_13_1728 ();
 sg13g2_fill_2 FILLER_13_1732 ();
 sg13g2_decap_4 FILLER_13_1752 ();
 sg13g2_fill_1 FILLER_13_1756 ();
 sg13g2_fill_2 FILLER_13_1777 ();
 sg13g2_decap_8 FILLER_13_1810 ();
 sg13g2_decap_4 FILLER_13_1817 ();
 sg13g2_fill_2 FILLER_13_1821 ();
 sg13g2_decap_8 FILLER_13_1853 ();
 sg13g2_decap_8 FILLER_13_1860 ();
 sg13g2_fill_1 FILLER_13_1867 ();
 sg13g2_fill_1 FILLER_13_1881 ();
 sg13g2_decap_8 FILLER_13_1888 ();
 sg13g2_fill_2 FILLER_13_1895 ();
 sg13g2_fill_1 FILLER_13_1897 ();
 sg13g2_fill_1 FILLER_13_1913 ();
 sg13g2_decap_8 FILLER_13_1963 ();
 sg13g2_decap_8 FILLER_13_1970 ();
 sg13g2_decap_8 FILLER_13_1977 ();
 sg13g2_decap_4 FILLER_13_1984 ();
 sg13g2_fill_2 FILLER_13_1988 ();
 sg13g2_decap_4 FILLER_13_1994 ();
 sg13g2_fill_2 FILLER_13_1998 ();
 sg13g2_fill_2 FILLER_13_2010 ();
 sg13g2_decap_4 FILLER_13_2020 ();
 sg13g2_fill_1 FILLER_13_2029 ();
 sg13g2_fill_1 FILLER_13_2048 ();
 sg13g2_decap_4 FILLER_13_2085 ();
 sg13g2_fill_2 FILLER_13_2089 ();
 sg13g2_fill_2 FILLER_13_2101 ();
 sg13g2_fill_2 FILLER_13_2107 ();
 sg13g2_fill_1 FILLER_13_2146 ();
 sg13g2_fill_1 FILLER_13_2215 ();
 sg13g2_decap_8 FILLER_13_2298 ();
 sg13g2_decap_8 FILLER_13_2305 ();
 sg13g2_fill_1 FILLER_13_2343 ();
 sg13g2_fill_1 FILLER_13_2370 ();
 sg13g2_decap_4 FILLER_13_2381 ();
 sg13g2_fill_1 FILLER_13_2385 ();
 sg13g2_decap_8 FILLER_13_2410 ();
 sg13g2_fill_1 FILLER_13_2417 ();
 sg13g2_decap_8 FILLER_13_2428 ();
 sg13g2_fill_1 FILLER_13_2435 ();
 sg13g2_decap_4 FILLER_13_2440 ();
 sg13g2_fill_1 FILLER_13_2444 ();
 sg13g2_decap_8 FILLER_13_2481 ();
 sg13g2_decap_8 FILLER_13_2488 ();
 sg13g2_fill_2 FILLER_13_2495 ();
 sg13g2_decap_8 FILLER_13_2523 ();
 sg13g2_decap_8 FILLER_13_2530 ();
 sg13g2_fill_2 FILLER_13_2537 ();
 sg13g2_decap_4 FILLER_13_2549 ();
 sg13g2_fill_1 FILLER_13_2553 ();
 sg13g2_decap_8 FILLER_13_2558 ();
 sg13g2_decap_4 FILLER_13_2565 ();
 sg13g2_fill_1 FILLER_13_2569 ();
 sg13g2_fill_2 FILLER_13_2580 ();
 sg13g2_fill_2 FILLER_13_2624 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_13 ();
 sg13g2_fill_1 FILLER_14_17 ();
 sg13g2_fill_2 FILLER_14_23 ();
 sg13g2_fill_2 FILLER_14_29 ();
 sg13g2_fill_1 FILLER_14_31 ();
 sg13g2_fill_2 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_38 ();
 sg13g2_fill_1 FILLER_14_47 ();
 sg13g2_fill_1 FILLER_14_53 ();
 sg13g2_fill_2 FILLER_14_77 ();
 sg13g2_decap_4 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_1 FILLER_14_114 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_148 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_decap_8 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_174 ();
 sg13g2_fill_1 FILLER_14_176 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_260 ();
 sg13g2_fill_2 FILLER_14_271 ();
 sg13g2_fill_1 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_282 ();
 sg13g2_decap_8 FILLER_14_289 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_1 FILLER_14_333 ();
 sg13g2_fill_2 FILLER_14_355 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_fill_2 FILLER_14_367 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_380 ();
 sg13g2_fill_1 FILLER_14_387 ();
 sg13g2_decap_4 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_410 ();
 sg13g2_decap_4 FILLER_14_417 ();
 sg13g2_fill_1 FILLER_14_421 ();
 sg13g2_decap_8 FILLER_14_426 ();
 sg13g2_fill_1 FILLER_14_433 ();
 sg13g2_fill_2 FILLER_14_448 ();
 sg13g2_fill_1 FILLER_14_450 ();
 sg13g2_fill_1 FILLER_14_456 ();
 sg13g2_fill_2 FILLER_14_463 ();
 sg13g2_fill_1 FILLER_14_465 ();
 sg13g2_fill_2 FILLER_14_475 ();
 sg13g2_fill_1 FILLER_14_477 ();
 sg13g2_decap_4 FILLER_14_492 ();
 sg13g2_fill_1 FILLER_14_496 ();
 sg13g2_fill_2 FILLER_14_502 ();
 sg13g2_fill_1 FILLER_14_504 ();
 sg13g2_fill_1 FILLER_14_509 ();
 sg13g2_fill_2 FILLER_14_521 ();
 sg13g2_fill_2 FILLER_14_536 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_fill_1 FILLER_14_598 ();
 sg13g2_fill_1 FILLER_14_604 ();
 sg13g2_fill_1 FILLER_14_613 ();
 sg13g2_fill_1 FILLER_14_619 ();
 sg13g2_fill_2 FILLER_14_655 ();
 sg13g2_fill_2 FILLER_14_687 ();
 sg13g2_fill_1 FILLER_14_700 ();
 sg13g2_fill_1 FILLER_14_706 ();
 sg13g2_fill_2 FILLER_14_721 ();
 sg13g2_fill_2 FILLER_14_748 ();
 sg13g2_fill_2 FILLER_14_790 ();
 sg13g2_fill_2 FILLER_14_801 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_1 FILLER_14_811 ();
 sg13g2_decap_8 FILLER_14_817 ();
 sg13g2_decap_4 FILLER_14_834 ();
 sg13g2_fill_1 FILLER_14_838 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_decap_4 FILLER_14_919 ();
 sg13g2_fill_2 FILLER_14_923 ();
 sg13g2_fill_2 FILLER_14_935 ();
 sg13g2_fill_1 FILLER_14_937 ();
 sg13g2_fill_2 FILLER_14_942 ();
 sg13g2_fill_1 FILLER_14_944 ();
 sg13g2_decap_8 FILLER_14_949 ();
 sg13g2_decap_8 FILLER_14_956 ();
 sg13g2_fill_1 FILLER_14_963 ();
 sg13g2_fill_1 FILLER_14_968 ();
 sg13g2_decap_4 FILLER_14_1055 ();
 sg13g2_fill_2 FILLER_14_1067 ();
 sg13g2_fill_1 FILLER_14_1074 ();
 sg13g2_decap_8 FILLER_14_1079 ();
 sg13g2_decap_8 FILLER_14_1086 ();
 sg13g2_fill_2 FILLER_14_1097 ();
 sg13g2_fill_1 FILLER_14_1099 ();
 sg13g2_decap_8 FILLER_14_1197 ();
 sg13g2_decap_8 FILLER_14_1204 ();
 sg13g2_decap_8 FILLER_14_1211 ();
 sg13g2_fill_2 FILLER_14_1218 ();
 sg13g2_fill_2 FILLER_14_1228 ();
 sg13g2_fill_1 FILLER_14_1230 ();
 sg13g2_fill_2 FILLER_14_1241 ();
 sg13g2_decap_8 FILLER_14_1274 ();
 sg13g2_fill_2 FILLER_14_1320 ();
 sg13g2_fill_2 FILLER_14_1351 ();
 sg13g2_decap_8 FILLER_14_1357 ();
 sg13g2_fill_2 FILLER_14_1364 ();
 sg13g2_decap_4 FILLER_14_1370 ();
 sg13g2_decap_4 FILLER_14_1399 ();
 sg13g2_fill_1 FILLER_14_1419 ();
 sg13g2_decap_4 FILLER_14_1424 ();
 sg13g2_decap_8 FILLER_14_1434 ();
 sg13g2_decap_8 FILLER_14_1441 ();
 sg13g2_decap_4 FILLER_14_1448 ();
 sg13g2_fill_2 FILLER_14_1452 ();
 sg13g2_decap_4 FILLER_14_1504 ();
 sg13g2_decap_4 FILLER_14_1518 ();
 sg13g2_fill_2 FILLER_14_1527 ();
 sg13g2_fill_1 FILLER_14_1546 ();
 sg13g2_fill_1 FILLER_14_1555 ();
 sg13g2_fill_1 FILLER_14_1570 ();
 sg13g2_fill_1 FILLER_14_1590 ();
 sg13g2_fill_1 FILLER_14_1623 ();
 sg13g2_decap_4 FILLER_14_1632 ();
 sg13g2_decap_8 FILLER_14_1650 ();
 sg13g2_decap_8 FILLER_14_1657 ();
 sg13g2_decap_8 FILLER_14_1664 ();
 sg13g2_decap_8 FILLER_14_1671 ();
 sg13g2_fill_2 FILLER_14_1678 ();
 sg13g2_fill_1 FILLER_14_1718 ();
 sg13g2_fill_1 FILLER_14_1733 ();
 sg13g2_decap_4 FILLER_14_1744 ();
 sg13g2_fill_1 FILLER_14_1748 ();
 sg13g2_fill_2 FILLER_14_1754 ();
 sg13g2_fill_1 FILLER_14_1756 ();
 sg13g2_fill_2 FILLER_14_1761 ();
 sg13g2_fill_1 FILLER_14_1763 ();
 sg13g2_decap_4 FILLER_14_1768 ();
 sg13g2_fill_2 FILLER_14_1772 ();
 sg13g2_fill_2 FILLER_14_1809 ();
 sg13g2_fill_2 FILLER_14_1816 ();
 sg13g2_fill_2 FILLER_14_1875 ();
 sg13g2_fill_2 FILLER_14_1883 ();
 sg13g2_fill_1 FILLER_14_1885 ();
 sg13g2_fill_2 FILLER_14_1891 ();
 sg13g2_fill_1 FILLER_14_1893 ();
 sg13g2_fill_1 FILLER_14_1904 ();
 sg13g2_fill_1 FILLER_14_1909 ();
 sg13g2_fill_1 FILLER_14_1919 ();
 sg13g2_decap_8 FILLER_14_1957 ();
 sg13g2_decap_8 FILLER_14_1964 ();
 sg13g2_decap_8 FILLER_14_1971 ();
 sg13g2_decap_8 FILLER_14_1978 ();
 sg13g2_decap_4 FILLER_14_1990 ();
 sg13g2_fill_2 FILLER_14_1994 ();
 sg13g2_decap_8 FILLER_14_2010 ();
 sg13g2_fill_2 FILLER_14_2017 ();
 sg13g2_fill_2 FILLER_14_2023 ();
 sg13g2_fill_1 FILLER_14_2038 ();
 sg13g2_fill_1 FILLER_14_2042 ();
 sg13g2_decap_8 FILLER_14_2083 ();
 sg13g2_decap_4 FILLER_14_2090 ();
 sg13g2_fill_1 FILLER_14_2094 ();
 sg13g2_fill_1 FILLER_14_2106 ();
 sg13g2_decap_4 FILLER_14_2133 ();
 sg13g2_fill_1 FILLER_14_2163 ();
 sg13g2_fill_2 FILLER_14_2168 ();
 sg13g2_decap_8 FILLER_14_2194 ();
 sg13g2_fill_2 FILLER_14_2237 ();
 sg13g2_decap_4 FILLER_14_2260 ();
 sg13g2_decap_8 FILLER_14_2290 ();
 sg13g2_decap_8 FILLER_14_2297 ();
 sg13g2_decap_4 FILLER_14_2304 ();
 sg13g2_fill_2 FILLER_14_2308 ();
 sg13g2_fill_2 FILLER_14_2346 ();
 sg13g2_fill_1 FILLER_14_2362 ();
 sg13g2_decap_8 FILLER_14_2367 ();
 sg13g2_decap_4 FILLER_14_2374 ();
 sg13g2_fill_1 FILLER_14_2378 ();
 sg13g2_fill_2 FILLER_14_2402 ();
 sg13g2_fill_1 FILLER_14_2404 ();
 sg13g2_fill_2 FILLER_14_2411 ();
 sg13g2_fill_2 FILLER_14_2423 ();
 sg13g2_fill_2 FILLER_14_2451 ();
 sg13g2_decap_4 FILLER_14_2513 ();
 sg13g2_decap_8 FILLER_14_2557 ();
 sg13g2_decap_8 FILLER_14_2564 ();
 sg13g2_decap_4 FILLER_14_2571 ();
 sg13g2_fill_2 FILLER_14_2575 ();
 sg13g2_fill_2 FILLER_14_2601 ();
 sg13g2_decap_4 FILLER_14_2607 ();
 sg13g2_fill_2 FILLER_14_2611 ();
 sg13g2_decap_8 FILLER_14_2660 ();
 sg13g2_fill_2 FILLER_14_2667 ();
 sg13g2_fill_1 FILLER_14_2669 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_decap_4 FILLER_15_38 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_112 ();
 sg13g2_fill_2 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_fill_1 FILLER_15_224 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_250 ();
 sg13g2_decap_8 FILLER_15_257 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_271 ();
 sg13g2_decap_8 FILLER_15_278 ();
 sg13g2_decap_4 FILLER_15_285 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_decap_4 FILLER_15_386 ();
 sg13g2_fill_2 FILLER_15_390 ();
 sg13g2_decap_4 FILLER_15_418 ();
 sg13g2_fill_1 FILLER_15_422 ();
 sg13g2_decap_8 FILLER_15_432 ();
 sg13g2_fill_2 FILLER_15_439 ();
 sg13g2_fill_1 FILLER_15_441 ();
 sg13g2_decap_4 FILLER_15_446 ();
 sg13g2_fill_1 FILLER_15_450 ();
 sg13g2_decap_4 FILLER_15_456 ();
 sg13g2_fill_2 FILLER_15_477 ();
 sg13g2_fill_1 FILLER_15_479 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_fill_2 FILLER_15_494 ();
 sg13g2_fill_1 FILLER_15_511 ();
 sg13g2_fill_2 FILLER_15_522 ();
 sg13g2_fill_1 FILLER_15_524 ();
 sg13g2_decap_8 FILLER_15_528 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_decap_4 FILLER_15_542 ();
 sg13g2_fill_2 FILLER_15_546 ();
 sg13g2_fill_2 FILLER_15_590 ();
 sg13g2_fill_2 FILLER_15_596 ();
 sg13g2_fill_1 FILLER_15_598 ();
 sg13g2_decap_8 FILLER_15_608 ();
 sg13g2_decap_8 FILLER_15_615 ();
 sg13g2_decap_8 FILLER_15_622 ();
 sg13g2_decap_4 FILLER_15_629 ();
 sg13g2_fill_2 FILLER_15_633 ();
 sg13g2_fill_1 FILLER_15_660 ();
 sg13g2_fill_1 FILLER_15_680 ();
 sg13g2_fill_2 FILLER_15_695 ();
 sg13g2_fill_2 FILLER_15_761 ();
 sg13g2_fill_1 FILLER_15_763 ();
 sg13g2_fill_1 FILLER_15_773 ();
 sg13g2_decap_4 FILLER_15_783 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_fill_1 FILLER_15_799 ();
 sg13g2_fill_1 FILLER_15_835 ();
 sg13g2_fill_1 FILLER_15_862 ();
 sg13g2_fill_1 FILLER_15_873 ();
 sg13g2_fill_2 FILLER_15_916 ();
 sg13g2_fill_1 FILLER_15_979 ();
 sg13g2_fill_1 FILLER_15_984 ();
 sg13g2_fill_1 FILLER_15_1000 ();
 sg13g2_fill_1 FILLER_15_1005 ();
 sg13g2_fill_2 FILLER_15_1010 ();
 sg13g2_fill_2 FILLER_15_1038 ();
 sg13g2_fill_1 FILLER_15_1113 ();
 sg13g2_decap_4 FILLER_15_1118 ();
 sg13g2_fill_1 FILLER_15_1157 ();
 sg13g2_fill_1 FILLER_15_1183 ();
 sg13g2_fill_2 FILLER_15_1188 ();
 sg13g2_fill_1 FILLER_15_1190 ();
 sg13g2_fill_1 FILLER_15_1196 ();
 sg13g2_decap_8 FILLER_15_1202 ();
 sg13g2_decap_8 FILLER_15_1209 ();
 sg13g2_decap_8 FILLER_15_1220 ();
 sg13g2_decap_4 FILLER_15_1227 ();
 sg13g2_decap_4 FILLER_15_1236 ();
 sg13g2_fill_1 FILLER_15_1240 ();
 sg13g2_decap_8 FILLER_15_1272 ();
 sg13g2_decap_4 FILLER_15_1279 ();
 sg13g2_fill_2 FILLER_15_1313 ();
 sg13g2_fill_1 FILLER_15_1315 ();
 sg13g2_fill_2 FILLER_15_1320 ();
 sg13g2_fill_1 FILLER_15_1322 ();
 sg13g2_fill_2 FILLER_15_1328 ();
 sg13g2_fill_1 FILLER_15_1330 ();
 sg13g2_fill_2 FILLER_15_1339 ();
 sg13g2_fill_2 FILLER_15_1345 ();
 sg13g2_decap_8 FILLER_15_1357 ();
 sg13g2_decap_8 FILLER_15_1364 ();
 sg13g2_decap_4 FILLER_15_1371 ();
 sg13g2_fill_2 FILLER_15_1389 ();
 sg13g2_fill_1 FILLER_15_1391 ();
 sg13g2_decap_4 FILLER_15_1397 ();
 sg13g2_fill_2 FILLER_15_1436 ();
 sg13g2_fill_1 FILLER_15_1438 ();
 sg13g2_fill_1 FILLER_15_1488 ();
 sg13g2_decap_4 FILLER_15_1493 ();
 sg13g2_fill_1 FILLER_15_1509 ();
 sg13g2_fill_2 FILLER_15_1515 ();
 sg13g2_fill_2 FILLER_15_1522 ();
 sg13g2_fill_1 FILLER_15_1533 ();
 sg13g2_fill_1 FILLER_15_1539 ();
 sg13g2_fill_1 FILLER_15_1545 ();
 sg13g2_fill_1 FILLER_15_1596 ();
 sg13g2_fill_1 FILLER_15_1604 ();
 sg13g2_decap_4 FILLER_15_1617 ();
 sg13g2_fill_1 FILLER_15_1621 ();
 sg13g2_fill_2 FILLER_15_1632 ();
 sg13g2_fill_2 FILLER_15_1697 ();
 sg13g2_fill_1 FILLER_15_1699 ();
 sg13g2_fill_1 FILLER_15_1713 ();
 sg13g2_fill_1 FILLER_15_1736 ();
 sg13g2_fill_1 FILLER_15_1744 ();
 sg13g2_fill_1 FILLER_15_1750 ();
 sg13g2_fill_2 FILLER_15_1756 ();
 sg13g2_decap_8 FILLER_15_1767 ();
 sg13g2_fill_1 FILLER_15_1774 ();
 sg13g2_decap_8 FILLER_15_1794 ();
 sg13g2_decap_8 FILLER_15_1801 ();
 sg13g2_fill_1 FILLER_15_1808 ();
 sg13g2_fill_1 FILLER_15_1835 ();
 sg13g2_decap_8 FILLER_15_1840 ();
 sg13g2_decap_8 FILLER_15_1847 ();
 sg13g2_decap_8 FILLER_15_1854 ();
 sg13g2_decap_8 FILLER_15_1861 ();
 sg13g2_decap_4 FILLER_15_1868 ();
 sg13g2_fill_2 FILLER_15_1875 ();
 sg13g2_fill_2 FILLER_15_1881 ();
 sg13g2_fill_2 FILLER_15_1891 ();
 sg13g2_fill_1 FILLER_15_1893 ();
 sg13g2_fill_1 FILLER_15_1935 ();
 sg13g2_fill_2 FILLER_15_1962 ();
 sg13g2_fill_2 FILLER_15_1974 ();
 sg13g2_fill_2 FILLER_15_2002 ();
 sg13g2_fill_1 FILLER_15_2004 ();
 sg13g2_decap_8 FILLER_15_2015 ();
 sg13g2_decap_8 FILLER_15_2022 ();
 sg13g2_fill_2 FILLER_15_2029 ();
 sg13g2_fill_1 FILLER_15_2031 ();
 sg13g2_decap_8 FILLER_15_2075 ();
 sg13g2_decap_8 FILLER_15_2082 ();
 sg13g2_decap_8 FILLER_15_2089 ();
 sg13g2_fill_1 FILLER_15_2102 ();
 sg13g2_fill_2 FILLER_15_2113 ();
 sg13g2_fill_2 FILLER_15_2147 ();
 sg13g2_decap_8 FILLER_15_2153 ();
 sg13g2_decap_8 FILLER_15_2160 ();
 sg13g2_decap_8 FILLER_15_2199 ();
 sg13g2_fill_2 FILLER_15_2206 ();
 sg13g2_fill_1 FILLER_15_2208 ();
 sg13g2_decap_8 FILLER_15_2213 ();
 sg13g2_fill_2 FILLER_15_2220 ();
 sg13g2_fill_1 FILLER_15_2222 ();
 sg13g2_fill_2 FILLER_15_2253 ();
 sg13g2_decap_4 FILLER_15_2291 ();
 sg13g2_fill_1 FILLER_15_2295 ();
 sg13g2_decap_8 FILLER_15_2326 ();
 sg13g2_fill_1 FILLER_15_2333 ();
 sg13g2_decap_4 FILLER_15_2344 ();
 sg13g2_fill_2 FILLER_15_2348 ();
 sg13g2_decap_8 FILLER_15_2376 ();
 sg13g2_fill_1 FILLER_15_2414 ();
 sg13g2_decap_8 FILLER_15_2445 ();
 sg13g2_decap_4 FILLER_15_2452 ();
 sg13g2_fill_1 FILLER_15_2456 ();
 sg13g2_fill_1 FILLER_15_2477 ();
 sg13g2_decap_4 FILLER_15_2488 ();
 sg13g2_fill_2 FILLER_15_2496 ();
 sg13g2_decap_8 FILLER_15_2518 ();
 sg13g2_fill_2 FILLER_15_2561 ();
 sg13g2_fill_1 FILLER_15_2563 ();
 sg13g2_decap_8 FILLER_15_2616 ();
 sg13g2_fill_1 FILLER_15_2623 ();
 sg13g2_fill_1 FILLER_15_2628 ();
 sg13g2_fill_1 FILLER_15_2641 ();
 sg13g2_fill_2 FILLER_15_2668 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_13 ();
 sg13g2_fill_2 FILLER_16_20 ();
 sg13g2_fill_1 FILLER_16_22 ();
 sg13g2_decap_4 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_36 ();
 sg13g2_fill_2 FILLER_16_41 ();
 sg13g2_fill_1 FILLER_16_43 ();
 sg13g2_fill_2 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_fill_1 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_277 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_decap_4 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_fill_2 FILLER_16_409 ();
 sg13g2_fill_2 FILLER_16_477 ();
 sg13g2_fill_2 FILLER_16_510 ();
 sg13g2_fill_1 FILLER_16_512 ();
 sg13g2_decap_4 FILLER_16_519 ();
 sg13g2_decap_4 FILLER_16_529 ();
 sg13g2_fill_1 FILLER_16_533 ();
 sg13g2_fill_2 FILLER_16_569 ();
 sg13g2_decap_4 FILLER_16_575 ();
 sg13g2_fill_2 FILLER_16_579 ();
 sg13g2_fill_2 FILLER_16_618 ();
 sg13g2_fill_1 FILLER_16_620 ();
 sg13g2_fill_2 FILLER_16_625 ();
 sg13g2_fill_1 FILLER_16_627 ();
 sg13g2_fill_2 FILLER_16_675 ();
 sg13g2_fill_2 FILLER_16_685 ();
 sg13g2_fill_2 FILLER_16_690 ();
 sg13g2_fill_2 FILLER_16_698 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_fill_1 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_824 ();
 sg13g2_decap_8 FILLER_16_831 ();
 sg13g2_decap_8 FILLER_16_838 ();
 sg13g2_decap_4 FILLER_16_845 ();
 sg13g2_decap_4 FILLER_16_867 ();
 sg13g2_fill_2 FILLER_16_871 ();
 sg13g2_decap_4 FILLER_16_883 ();
 sg13g2_fill_1 FILLER_16_887 ();
 sg13g2_decap_8 FILLER_16_898 ();
 sg13g2_decap_4 FILLER_16_905 ();
 sg13g2_decap_4 FILLER_16_935 ();
 sg13g2_fill_1 FILLER_16_939 ();
 sg13g2_fill_1 FILLER_16_965 ();
 sg13g2_fill_2 FILLER_16_971 ();
 sg13g2_decap_8 FILLER_16_981 ();
 sg13g2_decap_8 FILLER_16_988 ();
 sg13g2_decap_4 FILLER_16_1000 ();
 sg13g2_fill_2 FILLER_16_1017 ();
 sg13g2_fill_1 FILLER_16_1019 ();
 sg13g2_fill_1 FILLER_16_1041 ();
 sg13g2_fill_1 FILLER_16_1093 ();
 sg13g2_fill_2 FILLER_16_1112 ();
 sg13g2_decap_4 FILLER_16_1119 ();
 sg13g2_fill_1 FILLER_16_1123 ();
 sg13g2_fill_2 FILLER_16_1159 ();
 sg13g2_fill_1 FILLER_16_1161 ();
 sg13g2_decap_4 FILLER_16_1166 ();
 sg13g2_fill_1 FILLER_16_1170 ();
 sg13g2_decap_8 FILLER_16_1179 ();
 sg13g2_fill_2 FILLER_16_1186 ();
 sg13g2_fill_1 FILLER_16_1188 ();
 sg13g2_fill_1 FILLER_16_1194 ();
 sg13g2_decap_8 FILLER_16_1261 ();
 sg13g2_fill_2 FILLER_16_1268 ();
 sg13g2_fill_1 FILLER_16_1270 ();
 sg13g2_fill_1 FILLER_16_1286 ();
 sg13g2_fill_2 FILLER_16_1325 ();
 sg13g2_fill_1 FILLER_16_1327 ();
 sg13g2_decap_8 FILLER_16_1359 ();
 sg13g2_decap_4 FILLER_16_1366 ();
 sg13g2_fill_1 FILLER_16_1370 ();
 sg13g2_fill_1 FILLER_16_1375 ();
 sg13g2_fill_1 FILLER_16_1402 ();
 sg13g2_fill_1 FILLER_16_1408 ();
 sg13g2_fill_1 FILLER_16_1414 ();
 sg13g2_fill_1 FILLER_16_1420 ();
 sg13g2_fill_1 FILLER_16_1436 ();
 sg13g2_fill_2 FILLER_16_1447 ();
 sg13g2_fill_1 FILLER_16_1449 ();
 sg13g2_decap_8 FILLER_16_1454 ();
 sg13g2_fill_2 FILLER_16_1461 ();
 sg13g2_fill_1 FILLER_16_1473 ();
 sg13g2_fill_1 FILLER_16_1483 ();
 sg13g2_decap_8 FILLER_16_1489 ();
 sg13g2_fill_1 FILLER_16_1506 ();
 sg13g2_fill_2 FILLER_16_1513 ();
 sg13g2_fill_1 FILLER_16_1515 ();
 sg13g2_fill_1 FILLER_16_1531 ();
 sg13g2_fill_2 FILLER_16_1540 ();
 sg13g2_decap_8 FILLER_16_1554 ();
 sg13g2_decap_4 FILLER_16_1561 ();
 sg13g2_fill_1 FILLER_16_1565 ();
 sg13g2_fill_2 FILLER_16_1574 ();
 sg13g2_fill_2 FILLER_16_1586 ();
 sg13g2_fill_1 FILLER_16_1588 ();
 sg13g2_fill_1 FILLER_16_1606 ();
 sg13g2_fill_1 FILLER_16_1632 ();
 sg13g2_decap_8 FILLER_16_1639 ();
 sg13g2_decap_4 FILLER_16_1646 ();
 sg13g2_decap_4 FILLER_16_1686 ();
 sg13g2_fill_1 FILLER_16_1690 ();
 sg13g2_fill_1 FILLER_16_1711 ();
 sg13g2_fill_1 FILLER_16_1745 ();
 sg13g2_decap_4 FILLER_16_1755 ();
 sg13g2_fill_2 FILLER_16_1759 ();
 sg13g2_fill_2 FILLER_16_1766 ();
 sg13g2_fill_1 FILLER_16_1785 ();
 sg13g2_fill_1 FILLER_16_1790 ();
 sg13g2_decap_4 FILLER_16_1795 ();
 sg13g2_fill_2 FILLER_16_1811 ();
 sg13g2_fill_1 FILLER_16_1816 ();
 sg13g2_fill_2 FILLER_16_1827 ();
 sg13g2_decap_4 FILLER_16_1834 ();
 sg13g2_decap_8 FILLER_16_1846 ();
 sg13g2_decap_8 FILLER_16_1853 ();
 sg13g2_decap_8 FILLER_16_1860 ();
 sg13g2_decap_8 FILLER_16_1867 ();
 sg13g2_fill_2 FILLER_16_1874 ();
 sg13g2_fill_1 FILLER_16_1876 ();
 sg13g2_fill_2 FILLER_16_1886 ();
 sg13g2_decap_4 FILLER_16_1898 ();
 sg13g2_fill_2 FILLER_16_1907 ();
 sg13g2_fill_1 FILLER_16_1909 ();
 sg13g2_fill_1 FILLER_16_1914 ();
 sg13g2_fill_1 FILLER_16_1920 ();
 sg13g2_decap_4 FILLER_16_1929 ();
 sg13g2_fill_1 FILLER_16_1933 ();
 sg13g2_fill_1 FILLER_16_1938 ();
 sg13g2_decap_8 FILLER_16_1953 ();
 sg13g2_fill_2 FILLER_16_1986 ();
 sg13g2_fill_1 FILLER_16_2038 ();
 sg13g2_fill_1 FILLER_16_2092 ();
 sg13g2_fill_2 FILLER_16_2100 ();
 sg13g2_fill_1 FILLER_16_2102 ();
 sg13g2_decap_4 FILLER_16_2106 ();
 sg13g2_fill_2 FILLER_16_2110 ();
 sg13g2_fill_1 FILLER_16_2136 ();
 sg13g2_decap_8 FILLER_16_2145 ();
 sg13g2_fill_1 FILLER_16_2152 ();
 sg13g2_decap_4 FILLER_16_2209 ();
 sg13g2_decap_4 FILLER_16_2217 ();
 sg13g2_decap_8 FILLER_16_2247 ();
 sg13g2_decap_8 FILLER_16_2264 ();
 sg13g2_fill_1 FILLER_16_2275 ();
 sg13g2_decap_8 FILLER_16_2280 ();
 sg13g2_decap_8 FILLER_16_2287 ();
 sg13g2_decap_8 FILLER_16_2294 ();
 sg13g2_fill_1 FILLER_16_2301 ();
 sg13g2_decap_4 FILLER_16_2306 ();
 sg13g2_fill_1 FILLER_16_2310 ();
 sg13g2_decap_8 FILLER_16_2335 ();
 sg13g2_decap_8 FILLER_16_2342 ();
 sg13g2_decap_8 FILLER_16_2349 ();
 sg13g2_fill_1 FILLER_16_2356 ();
 sg13g2_fill_2 FILLER_16_2408 ();
 sg13g2_fill_1 FILLER_16_2410 ();
 sg13g2_fill_2 FILLER_16_2421 ();
 sg13g2_fill_1 FILLER_16_2423 ();
 sg13g2_decap_8 FILLER_16_2450 ();
 sg13g2_fill_2 FILLER_16_2457 ();
 sg13g2_fill_2 FILLER_16_2485 ();
 sg13g2_fill_2 FILLER_16_2491 ();
 sg13g2_decap_8 FILLER_16_2519 ();
 sg13g2_decap_4 FILLER_16_2526 ();
 sg13g2_fill_2 FILLER_16_2530 ();
 sg13g2_decap_4 FILLER_16_2580 ();
 sg13g2_decap_8 FILLER_16_2601 ();
 sg13g2_decap_8 FILLER_16_2608 ();
 sg13g2_decap_8 FILLER_16_2615 ();
 sg13g2_decap_4 FILLER_16_2622 ();
 sg13g2_decap_8 FILLER_16_2645 ();
 sg13g2_decap_8 FILLER_16_2652 ();
 sg13g2_decap_8 FILLER_16_2659 ();
 sg13g2_decap_4 FILLER_16_2666 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_34 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_fill_2 FILLER_17_154 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_decap_4 FILLER_17_177 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_226 ();
 sg13g2_fill_1 FILLER_17_231 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_fill_2 FILLER_17_269 ();
 sg13g2_fill_2 FILLER_17_336 ();
 sg13g2_fill_2 FILLER_17_348 ();
 sg13g2_fill_1 FILLER_17_355 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_decap_4 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_402 ();
 sg13g2_fill_1 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_478 ();
 sg13g2_fill_1 FILLER_17_480 ();
 sg13g2_fill_1 FILLER_17_526 ();
 sg13g2_decap_8 FILLER_17_531 ();
 sg13g2_decap_8 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_545 ();
 sg13g2_fill_1 FILLER_17_565 ();
 sg13g2_fill_1 FILLER_17_575 ();
 sg13g2_decap_4 FILLER_17_581 ();
 sg13g2_fill_1 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_593 ();
 sg13g2_decap_8 FILLER_17_600 ();
 sg13g2_fill_1 FILLER_17_662 ();
 sg13g2_decap_4 FILLER_17_693 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_decap_4 FILLER_17_712 ();
 sg13g2_fill_1 FILLER_17_716 ();
 sg13g2_fill_1 FILLER_17_722 ();
 sg13g2_fill_2 FILLER_17_749 ();
 sg13g2_fill_1 FILLER_17_751 ();
 sg13g2_fill_1 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_769 ();
 sg13g2_fill_2 FILLER_17_781 ();
 sg13g2_fill_1 FILLER_17_783 ();
 sg13g2_fill_2 FILLER_17_788 ();
 sg13g2_fill_1 FILLER_17_790 ();
 sg13g2_fill_2 FILLER_17_795 ();
 sg13g2_fill_1 FILLER_17_797 ();
 sg13g2_fill_1 FILLER_17_808 ();
 sg13g2_decap_8 FILLER_17_813 ();
 sg13g2_decap_8 FILLER_17_820 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_fill_1 FILLER_17_841 ();
 sg13g2_decap_8 FILLER_17_894 ();
 sg13g2_fill_1 FILLER_17_901 ();
 sg13g2_fill_1 FILLER_17_948 ();
 sg13g2_fill_1 FILLER_17_954 ();
 sg13g2_fill_2 FILLER_17_963 ();
 sg13g2_fill_1 FILLER_17_965 ();
 sg13g2_decap_8 FILLER_17_992 ();
 sg13g2_decap_4 FILLER_17_999 ();
 sg13g2_fill_1 FILLER_17_1003 ();
 sg13g2_decap_4 FILLER_17_1017 ();
 sg13g2_fill_2 FILLER_17_1021 ();
 sg13g2_fill_2 FILLER_17_1032 ();
 sg13g2_fill_1 FILLER_17_1052 ();
 sg13g2_fill_2 FILLER_17_1114 ();
 sg13g2_decap_4 FILLER_17_1125 ();
 sg13g2_fill_1 FILLER_17_1129 ();
 sg13g2_decap_8 FILLER_17_1143 ();
 sg13g2_decap_4 FILLER_17_1150 ();
 sg13g2_fill_2 FILLER_17_1154 ();
 sg13g2_decap_4 FILLER_17_1197 ();
 sg13g2_fill_1 FILLER_17_1201 ();
 sg13g2_decap_8 FILLER_17_1238 ();
 sg13g2_fill_2 FILLER_17_1245 ();
 sg13g2_decap_8 FILLER_17_1273 ();
 sg13g2_decap_8 FILLER_17_1280 ();
 sg13g2_fill_2 FILLER_17_1305 ();
 sg13g2_decap_4 FILLER_17_1311 ();
 sg13g2_decap_8 FILLER_17_1319 ();
 sg13g2_fill_2 FILLER_17_1326 ();
 sg13g2_fill_1 FILLER_17_1328 ();
 sg13g2_fill_2 FILLER_17_1350 ();
 sg13g2_fill_2 FILLER_17_1388 ();
 sg13g2_fill_1 FILLER_17_1410 ();
 sg13g2_fill_1 FILLER_17_1416 ();
 sg13g2_fill_1 FILLER_17_1421 ();
 sg13g2_fill_1 FILLER_17_1431 ();
 sg13g2_decap_8 FILLER_17_1441 ();
 sg13g2_decap_4 FILLER_17_1448 ();
 sg13g2_fill_1 FILLER_17_1452 ();
 sg13g2_decap_8 FILLER_17_1462 ();
 sg13g2_decap_8 FILLER_17_1469 ();
 sg13g2_fill_1 FILLER_17_1533 ();
 sg13g2_fill_2 FILLER_17_1546 ();
 sg13g2_fill_2 FILLER_17_1573 ();
 sg13g2_fill_1 FILLER_17_1575 ();
 sg13g2_fill_1 FILLER_17_1586 ();
 sg13g2_decap_8 FILLER_17_1592 ();
 sg13g2_fill_2 FILLER_17_1599 ();
 sg13g2_fill_2 FILLER_17_1606 ();
 sg13g2_fill_1 FILLER_17_1622 ();
 sg13g2_fill_1 FILLER_17_1641 ();
 sg13g2_decap_8 FILLER_17_1646 ();
 sg13g2_decap_8 FILLER_17_1653 ();
 sg13g2_decap_8 FILLER_17_1660 ();
 sg13g2_decap_8 FILLER_17_1675 ();
 sg13g2_decap_8 FILLER_17_1682 ();
 sg13g2_decap_8 FILLER_17_1689 ();
 sg13g2_fill_2 FILLER_17_1696 ();
 sg13g2_fill_1 FILLER_17_1698 ();
 sg13g2_fill_1 FILLER_17_1733 ();
 sg13g2_fill_1 FILLER_17_1738 ();
 sg13g2_fill_2 FILLER_17_1753 ();
 sg13g2_fill_1 FILLER_17_1769 ();
 sg13g2_fill_2 FILLER_17_1780 ();
 sg13g2_fill_1 FILLER_17_1782 ();
 sg13g2_fill_2 FILLER_17_1789 ();
 sg13g2_fill_2 FILLER_17_1796 ();
 sg13g2_fill_1 FILLER_17_1812 ();
 sg13g2_fill_1 FILLER_17_1823 ();
 sg13g2_fill_2 FILLER_17_1834 ();
 sg13g2_fill_1 FILLER_17_1836 ();
 sg13g2_decap_8 FILLER_17_1899 ();
 sg13g2_fill_1 FILLER_17_1906 ();
 sg13g2_decap_8 FILLER_17_1911 ();
 sg13g2_decap_8 FILLER_17_1918 ();
 sg13g2_fill_2 FILLER_17_1925 ();
 sg13g2_fill_1 FILLER_17_1927 ();
 sg13g2_fill_2 FILLER_17_1938 ();
 sg13g2_fill_1 FILLER_17_1940 ();
 sg13g2_decap_8 FILLER_17_1971 ();
 sg13g2_fill_2 FILLER_17_1978 ();
 sg13g2_fill_1 FILLER_17_2020 ();
 sg13g2_fill_1 FILLER_17_2025 ();
 sg13g2_fill_2 FILLER_17_2052 ();
 sg13g2_decap_8 FILLER_17_2085 ();
 sg13g2_decap_4 FILLER_17_2092 ();
 sg13g2_fill_1 FILLER_17_2125 ();
 sg13g2_fill_2 FILLER_17_2230 ();
 sg13g2_fill_1 FILLER_17_2232 ();
 sg13g2_decap_8 FILLER_17_2243 ();
 sg13g2_decap_8 FILLER_17_2250 ();
 sg13g2_decap_8 FILLER_17_2257 ();
 sg13g2_decap_4 FILLER_17_2264 ();
 sg13g2_fill_1 FILLER_17_2268 ();
 sg13g2_decap_8 FILLER_17_2273 ();
 sg13g2_decap_8 FILLER_17_2280 ();
 sg13g2_decap_8 FILLER_17_2287 ();
 sg13g2_fill_2 FILLER_17_2294 ();
 sg13g2_decap_4 FILLER_17_2332 ();
 sg13g2_decap_4 FILLER_17_2342 ();
 sg13g2_fill_1 FILLER_17_2378 ();
 sg13g2_fill_1 FILLER_17_2389 ();
 sg13g2_fill_1 FILLER_17_2400 ();
 sg13g2_fill_1 FILLER_17_2407 ();
 sg13g2_fill_1 FILLER_17_2414 ();
 sg13g2_fill_1 FILLER_17_2441 ();
 sg13g2_decap_8 FILLER_17_2446 ();
 sg13g2_fill_2 FILLER_17_2453 ();
 sg13g2_decap_8 FILLER_17_2471 ();
 sg13g2_fill_2 FILLER_17_2478 ();
 sg13g2_fill_1 FILLER_17_2480 ();
 sg13g2_decap_4 FILLER_17_2507 ();
 sg13g2_fill_2 FILLER_17_2511 ();
 sg13g2_decap_8 FILLER_17_2519 ();
 sg13g2_fill_2 FILLER_17_2526 ();
 sg13g2_decap_4 FILLER_17_2534 ();
 sg13g2_fill_1 FILLER_17_2538 ();
 sg13g2_fill_2 FILLER_17_2549 ();
 sg13g2_decap_4 FILLER_17_2561 ();
 sg13g2_fill_1 FILLER_17_2565 ();
 sg13g2_fill_2 FILLER_17_2570 ();
 sg13g2_fill_1 FILLER_17_2572 ();
 sg13g2_fill_2 FILLER_17_2609 ();
 sg13g2_fill_1 FILLER_17_2611 ();
 sg13g2_fill_2 FILLER_17_2616 ();
 sg13g2_fill_1 FILLER_17_2618 ();
 sg13g2_fill_1 FILLER_17_2629 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_2 FILLER_18_44 ();
 sg13g2_fill_2 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_109 ();
 sg13g2_fill_1 FILLER_18_128 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_177 ();
 sg13g2_fill_2 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_193 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_decap_4 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_4 FILLER_18_301 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_312 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_fill_2 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_18_378 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_fill_2 FILLER_18_393 ();
 sg13g2_fill_1 FILLER_18_395 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_fill_2 FILLER_18_447 ();
 sg13g2_fill_2 FILLER_18_455 ();
 sg13g2_decap_4 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_474 ();
 sg13g2_fill_2 FILLER_18_480 ();
 sg13g2_fill_1 FILLER_18_495 ();
 sg13g2_fill_1 FILLER_18_505 ();
 sg13g2_fill_1 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_538 ();
 sg13g2_decap_8 FILLER_18_545 ();
 sg13g2_fill_1 FILLER_18_552 ();
 sg13g2_fill_2 FILLER_18_593 ();
 sg13g2_fill_2 FILLER_18_621 ();
 sg13g2_fill_1 FILLER_18_623 ();
 sg13g2_fill_1 FILLER_18_652 ();
 sg13g2_decap_8 FILLER_18_699 ();
 sg13g2_decap_4 FILLER_18_706 ();
 sg13g2_decap_4 FILLER_18_715 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_fill_2 FILLER_18_735 ();
 sg13g2_fill_2 FILLER_18_763 ();
 sg13g2_fill_1 FILLER_18_765 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_fill_1 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_782 ();
 sg13g2_decap_8 FILLER_18_789 ();
 sg13g2_fill_2 FILLER_18_796 ();
 sg13g2_fill_1 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_decap_8 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_829 ();
 sg13g2_decap_8 FILLER_18_836 ();
 sg13g2_fill_2 FILLER_18_879 ();
 sg13g2_fill_1 FILLER_18_881 ();
 sg13g2_fill_2 FILLER_18_908 ();
 sg13g2_fill_1 FILLER_18_954 ();
 sg13g2_decap_4 FILLER_18_1001 ();
 sg13g2_fill_2 FILLER_18_1005 ();
 sg13g2_fill_2 FILLER_18_1042 ();
 sg13g2_fill_2 FILLER_18_1062 ();
 sg13g2_fill_1 FILLER_18_1064 ();
 sg13g2_fill_1 FILLER_18_1070 ();
 sg13g2_decap_8 FILLER_18_1120 ();
 sg13g2_fill_2 FILLER_18_1127 ();
 sg13g2_decap_8 FILLER_18_1134 ();
 sg13g2_decap_4 FILLER_18_1141 ();
 sg13g2_fill_1 FILLER_18_1145 ();
 sg13g2_decap_8 FILLER_18_1151 ();
 sg13g2_decap_4 FILLER_18_1158 ();
 sg13g2_fill_1 FILLER_18_1162 ();
 sg13g2_fill_2 FILLER_18_1189 ();
 sg13g2_fill_1 FILLER_18_1191 ();
 sg13g2_fill_1 FILLER_18_1213 ();
 sg13g2_fill_2 FILLER_18_1254 ();
 sg13g2_fill_1 FILLER_18_1256 ();
 sg13g2_decap_8 FILLER_18_1266 ();
 sg13g2_decap_8 FILLER_18_1273 ();
 sg13g2_decap_4 FILLER_18_1323 ();
 sg13g2_fill_2 FILLER_18_1327 ();
 sg13g2_fill_2 FILLER_18_1339 ();
 sg13g2_fill_1 FILLER_18_1341 ();
 sg13g2_decap_4 FILLER_18_1355 ();
 sg13g2_fill_1 FILLER_18_1371 ();
 sg13g2_fill_1 FILLER_18_1419 ();
 sg13g2_fill_2 FILLER_18_1430 ();
 sg13g2_fill_1 FILLER_18_1439 ();
 sg13g2_decap_4 FILLER_18_1445 ();
 sg13g2_fill_2 FILLER_18_1449 ();
 sg13g2_fill_1 FILLER_18_1457 ();
 sg13g2_decap_8 FILLER_18_1469 ();
 sg13g2_fill_2 FILLER_18_1476 ();
 sg13g2_fill_2 FILLER_18_1491 ();
 sg13g2_fill_1 FILLER_18_1493 ();
 sg13g2_fill_1 FILLER_18_1553 ();
 sg13g2_fill_2 FILLER_18_1573 ();
 sg13g2_fill_1 FILLER_18_1575 ();
 sg13g2_decap_4 FILLER_18_1583 ();
 sg13g2_fill_2 FILLER_18_1587 ();
 sg13g2_decap_4 FILLER_18_1595 ();
 sg13g2_fill_2 FILLER_18_1599 ();
 sg13g2_fill_2 FILLER_18_1606 ();
 sg13g2_fill_1 FILLER_18_1608 ();
 sg13g2_fill_2 FILLER_18_1642 ();
 sg13g2_fill_2 FILLER_18_1719 ();
 sg13g2_decap_8 FILLER_18_1726 ();
 sg13g2_fill_2 FILLER_18_1733 ();
 sg13g2_fill_1 FILLER_18_1735 ();
 sg13g2_decap_4 FILLER_18_1758 ();
 sg13g2_fill_1 FILLER_18_1762 ();
 sg13g2_fill_2 FILLER_18_1789 ();
 sg13g2_fill_2 FILLER_18_1801 ();
 sg13g2_fill_1 FILLER_18_1890 ();
 sg13g2_decap_8 FILLER_18_1962 ();
 sg13g2_decap_8 FILLER_18_1969 ();
 sg13g2_decap_8 FILLER_18_1976 ();
 sg13g2_decap_8 FILLER_18_1993 ();
 sg13g2_fill_1 FILLER_18_2000 ();
 sg13g2_fill_1 FILLER_18_2005 ();
 sg13g2_fill_2 FILLER_18_2032 ();
 sg13g2_decap_4 FILLER_18_2081 ();
 sg13g2_fill_2 FILLER_18_2085 ();
 sg13g2_fill_2 FILLER_18_2134 ();
 sg13g2_fill_1 FILLER_18_2136 ();
 sg13g2_fill_2 FILLER_18_2183 ();
 sg13g2_fill_1 FILLER_18_2211 ();
 sg13g2_decap_8 FILLER_18_2221 ();
 sg13g2_fill_1 FILLER_18_2228 ();
 sg13g2_decap_4 FILLER_18_2233 ();
 sg13g2_fill_1 FILLER_18_2237 ();
 sg13g2_fill_1 FILLER_18_2252 ();
 sg13g2_decap_8 FILLER_18_2289 ();
 sg13g2_fill_1 FILLER_18_2296 ();
 sg13g2_fill_1 FILLER_18_2301 ();
 sg13g2_fill_2 FILLER_18_2310 ();
 sg13g2_fill_1 FILLER_18_2312 ();
 sg13g2_decap_8 FILLER_18_2339 ();
 sg13g2_fill_2 FILLER_18_2352 ();
 sg13g2_decap_8 FILLER_18_2358 ();
 sg13g2_fill_2 FILLER_18_2365 ();
 sg13g2_fill_1 FILLER_18_2367 ();
 sg13g2_decap_4 FILLER_18_2384 ();
 sg13g2_fill_1 FILLER_18_2388 ();
 sg13g2_fill_2 FILLER_18_2418 ();
 sg13g2_decap_8 FILLER_18_2432 ();
 sg13g2_decap_4 FILLER_18_2439 ();
 sg13g2_fill_2 FILLER_18_2443 ();
 sg13g2_fill_2 FILLER_18_2451 ();
 sg13g2_fill_1 FILLER_18_2453 ();
 sg13g2_decap_8 FILLER_18_2462 ();
 sg13g2_fill_2 FILLER_18_2469 ();
 sg13g2_decap_8 FILLER_18_2481 ();
 sg13g2_fill_1 FILLER_18_2488 ();
 sg13g2_fill_1 FILLER_18_2524 ();
 sg13g2_decap_8 FILLER_18_2551 ();
 sg13g2_decap_8 FILLER_18_2558 ();
 sg13g2_fill_2 FILLER_18_2565 ();
 sg13g2_decap_4 FILLER_18_2664 ();
 sg13g2_fill_2 FILLER_18_2668 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_7 ();
 sg13g2_fill_1 FILLER_19_13 ();
 sg13g2_fill_1 FILLER_19_18 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_116 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_184 ();
 sg13g2_fill_1 FILLER_19_212 ();
 sg13g2_fill_1 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_234 ();
 sg13g2_fill_1 FILLER_19_244 ();
 sg13g2_fill_1 FILLER_19_255 ();
 sg13g2_fill_1 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_decap_4 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_fill_2 FILLER_19_282 ();
 sg13g2_fill_2 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_346 ();
 sg13g2_fill_1 FILLER_19_416 ();
 sg13g2_decap_4 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_4 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_decap_8 FILLER_19_542 ();
 sg13g2_decap_4 FILLER_19_549 ();
 sg13g2_fill_1 FILLER_19_553 ();
 sg13g2_fill_2 FILLER_19_577 ();
 sg13g2_fill_1 FILLER_19_601 ();
 sg13g2_fill_1 FILLER_19_606 ();
 sg13g2_fill_1 FILLER_19_616 ();
 sg13g2_fill_1 FILLER_19_642 ();
 sg13g2_decap_8 FILLER_19_647 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_fill_2 FILLER_19_704 ();
 sg13g2_fill_1 FILLER_19_706 ();
 sg13g2_fill_2 FILLER_19_735 ();
 sg13g2_fill_1 FILLER_19_737 ();
 sg13g2_decap_8 FILLER_19_750 ();
 sg13g2_decap_4 FILLER_19_757 ();
 sg13g2_decap_8 FILLER_19_766 ();
 sg13g2_decap_4 FILLER_19_773 ();
 sg13g2_decap_8 FILLER_19_834 ();
 sg13g2_decap_4 FILLER_19_841 ();
 sg13g2_fill_1 FILLER_19_845 ();
 sg13g2_fill_2 FILLER_19_891 ();
 sg13g2_fill_1 FILLER_19_893 ();
 sg13g2_fill_2 FILLER_19_898 ();
 sg13g2_fill_1 FILLER_19_900 ();
 sg13g2_decap_8 FILLER_19_922 ();
 sg13g2_decap_8 FILLER_19_929 ();
 sg13g2_decap_8 FILLER_19_936 ();
 sg13g2_decap_4 FILLER_19_943 ();
 sg13g2_fill_1 FILLER_19_968 ();
 sg13g2_decap_4 FILLER_19_1004 ();
 sg13g2_fill_1 FILLER_19_1008 ();
 sg13g2_decap_4 FILLER_19_1035 ();
 sg13g2_fill_1 FILLER_19_1039 ();
 sg13g2_fill_1 FILLER_19_1074 ();
 sg13g2_fill_2 FILLER_19_1078 ();
 sg13g2_fill_1 FILLER_19_1080 ();
 sg13g2_fill_1 FILLER_19_1114 ();
 sg13g2_fill_1 FILLER_19_1124 ();
 sg13g2_fill_2 FILLER_19_1156 ();
 sg13g2_fill_1 FILLER_19_1158 ();
 sg13g2_decap_8 FILLER_19_1215 ();
 sg13g2_decap_8 FILLER_19_1222 ();
 sg13g2_decap_8 FILLER_19_1229 ();
 sg13g2_decap_4 FILLER_19_1236 ();
 sg13g2_fill_2 FILLER_19_1240 ();
 sg13g2_decap_8 FILLER_19_1246 ();
 sg13g2_decap_8 FILLER_19_1253 ();
 sg13g2_fill_2 FILLER_19_1260 ();
 sg13g2_fill_2 FILLER_19_1327 ();
 sg13g2_fill_1 FILLER_19_1355 ();
 sg13g2_decap_8 FILLER_19_1363 ();
 sg13g2_decap_4 FILLER_19_1370 ();
 sg13g2_fill_1 FILLER_19_1402 ();
 sg13g2_fill_1 FILLER_19_1416 ();
 sg13g2_fill_2 FILLER_19_1430 ();
 sg13g2_decap_8 FILLER_19_1438 ();
 sg13g2_fill_1 FILLER_19_1445 ();
 sg13g2_fill_1 FILLER_19_1471 ();
 sg13g2_fill_1 FILLER_19_1513 ();
 sg13g2_fill_2 FILLER_19_1540 ();
 sg13g2_fill_2 FILLER_19_1551 ();
 sg13g2_fill_1 FILLER_19_1553 ();
 sg13g2_decap_4 FILLER_19_1558 ();
 sg13g2_fill_1 FILLER_19_1562 ();
 sg13g2_decap_8 FILLER_19_1581 ();
 sg13g2_fill_2 FILLER_19_1588 ();
 sg13g2_fill_1 FILLER_19_1590 ();
 sg13g2_fill_2 FILLER_19_1601 ();
 sg13g2_fill_1 FILLER_19_1603 ();
 sg13g2_fill_1 FILLER_19_1614 ();
 sg13g2_fill_1 FILLER_19_1625 ();
 sg13g2_fill_1 FILLER_19_1631 ();
 sg13g2_fill_2 FILLER_19_1651 ();
 sg13g2_decap_8 FILLER_19_1679 ();
 sg13g2_fill_2 FILLER_19_1686 ();
 sg13g2_fill_1 FILLER_19_1688 ();
 sg13g2_fill_2 FILLER_19_1722 ();
 sg13g2_fill_1 FILLER_19_1752 ();
 sg13g2_fill_2 FILLER_19_1757 ();
 sg13g2_fill_1 FILLER_19_1759 ();
 sg13g2_fill_2 FILLER_19_1764 ();
 sg13g2_fill_1 FILLER_19_1775 ();
 sg13g2_fill_1 FILLER_19_1780 ();
 sg13g2_fill_2 FILLER_19_1786 ();
 sg13g2_fill_1 FILLER_19_1788 ();
 sg13g2_fill_1 FILLER_19_1816 ();
 sg13g2_decap_4 FILLER_19_1873 ();
 sg13g2_fill_1 FILLER_19_1877 ();
 sg13g2_fill_2 FILLER_19_1882 ();
 sg13g2_fill_1 FILLER_19_1884 ();
 sg13g2_decap_4 FILLER_19_1890 ();
 sg13g2_fill_1 FILLER_19_1936 ();
 sg13g2_decap_8 FILLER_19_1958 ();
 sg13g2_fill_2 FILLER_19_1965 ();
 sg13g2_fill_1 FILLER_19_1967 ();
 sg13g2_fill_2 FILLER_19_2020 ();
 sg13g2_fill_1 FILLER_19_2034 ();
 sg13g2_fill_1 FILLER_19_2065 ();
 sg13g2_decap_8 FILLER_19_2074 ();
 sg13g2_decap_8 FILLER_19_2081 ();
 sg13g2_fill_1 FILLER_19_2110 ();
 sg13g2_fill_2 FILLER_19_2137 ();
 sg13g2_fill_2 FILLER_19_2153 ();
 sg13g2_fill_2 FILLER_19_2180 ();
 sg13g2_fill_1 FILLER_19_2182 ();
 sg13g2_decap_4 FILLER_19_2196 ();
 sg13g2_decap_8 FILLER_19_2236 ();
 sg13g2_fill_2 FILLER_19_2243 ();
 sg13g2_fill_1 FILLER_19_2245 ();
 sg13g2_decap_8 FILLER_19_2282 ();
 sg13g2_fill_1 FILLER_19_2289 ();
 sg13g2_fill_2 FILLER_19_2303 ();
 sg13g2_fill_1 FILLER_19_2305 ();
 sg13g2_decap_8 FILLER_19_2348 ();
 sg13g2_fill_2 FILLER_19_2355 ();
 sg13g2_decap_4 FILLER_19_2361 ();
 sg13g2_decap_8 FILLER_19_2375 ();
 sg13g2_fill_1 FILLER_19_2404 ();
 sg13g2_fill_2 FILLER_19_2417 ();
 sg13g2_fill_1 FILLER_19_2419 ();
 sg13g2_decap_8 FILLER_19_2478 ();
 sg13g2_fill_1 FILLER_19_2508 ();
 sg13g2_fill_1 FILLER_19_2521 ();
 sg13g2_fill_2 FILLER_19_2564 ();
 sg13g2_fill_2 FILLER_19_2574 ();
 sg13g2_fill_2 FILLER_19_2588 ();
 sg13g2_decap_4 FILLER_19_2626 ();
 sg13g2_fill_2 FILLER_19_2630 ();
 sg13g2_fill_1 FILLER_19_2646 ();
 sg13g2_decap_8 FILLER_19_2655 ();
 sg13g2_decap_8 FILLER_19_2662 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_fill_2 FILLER_20_75 ();
 sg13g2_fill_1 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_94 ();
 sg13g2_fill_2 FILLER_20_150 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_188 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_fill_2 FILLER_20_206 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_fill_2 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_decap_4 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_decap_4 FILLER_20_347 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_378 ();
 sg13g2_fill_1 FILLER_20_393 ();
 sg13g2_fill_2 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_409 ();
 sg13g2_decap_4 FILLER_20_415 ();
 sg13g2_fill_1 FILLER_20_419 ();
 sg13g2_fill_2 FILLER_20_429 ();
 sg13g2_fill_1 FILLER_20_431 ();
 sg13g2_fill_1 FILLER_20_463 ();
 sg13g2_decap_4 FILLER_20_491 ();
 sg13g2_fill_1 FILLER_20_495 ();
 sg13g2_fill_2 FILLER_20_528 ();
 sg13g2_fill_2 FILLER_20_535 ();
 sg13g2_fill_2 FILLER_20_543 ();
 sg13g2_fill_1 FILLER_20_575 ();
 sg13g2_fill_1 FILLER_20_589 ();
 sg13g2_fill_2 FILLER_20_593 ();
 sg13g2_fill_1 FILLER_20_595 ();
 sg13g2_fill_2 FILLER_20_601 ();
 sg13g2_decap_8 FILLER_20_612 ();
 sg13g2_decap_8 FILLER_20_628 ();
 sg13g2_fill_1 FILLER_20_635 ();
 sg13g2_fill_1 FILLER_20_650 ();
 sg13g2_decap_4 FILLER_20_661 ();
 sg13g2_fill_1 FILLER_20_665 ();
 sg13g2_fill_2 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_689 ();
 sg13g2_decap_8 FILLER_20_696 ();
 sg13g2_fill_2 FILLER_20_703 ();
 sg13g2_fill_1 FILLER_20_714 ();
 sg13g2_decap_4 FILLER_20_719 ();
 sg13g2_fill_1 FILLER_20_723 ();
 sg13g2_decap_4 FILLER_20_733 ();
 sg13g2_fill_1 FILLER_20_737 ();
 sg13g2_fill_2 FILLER_20_742 ();
 sg13g2_fill_1 FILLER_20_744 ();
 sg13g2_decap_8 FILLER_20_750 ();
 sg13g2_fill_1 FILLER_20_757 ();
 sg13g2_fill_2 FILLER_20_798 ();
 sg13g2_fill_2 FILLER_20_804 ();
 sg13g2_decap_4 FILLER_20_811 ();
 sg13g2_decap_4 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_849 ();
 sg13g2_fill_2 FILLER_20_856 ();
 sg13g2_decap_4 FILLER_20_884 ();
 sg13g2_fill_2 FILLER_20_888 ();
 sg13g2_decap_8 FILLER_20_895 ();
 sg13g2_decap_4 FILLER_20_902 ();
 sg13g2_fill_2 FILLER_20_912 ();
 sg13g2_decap_4 FILLER_20_954 ();
 sg13g2_fill_2 FILLER_20_958 ();
 sg13g2_decap_8 FILLER_20_994 ();
 sg13g2_decap_4 FILLER_20_1001 ();
 sg13g2_fill_1 FILLER_20_1005 ();
 sg13g2_fill_2 FILLER_20_1058 ();
 sg13g2_decap_4 FILLER_20_1068 ();
 sg13g2_fill_1 FILLER_20_1072 ();
 sg13g2_fill_2 FILLER_20_1082 ();
 sg13g2_decap_8 FILLER_20_1101 ();
 sg13g2_fill_2 FILLER_20_1108 ();
 sg13g2_fill_1 FILLER_20_1110 ();
 sg13g2_fill_2 FILLER_20_1132 ();
 sg13g2_decap_8 FILLER_20_1138 ();
 sg13g2_decap_4 FILLER_20_1145 ();
 sg13g2_fill_1 FILLER_20_1149 ();
 sg13g2_fill_1 FILLER_20_1185 ();
 sg13g2_decap_8 FILLER_20_1190 ();
 sg13g2_decap_4 FILLER_20_1197 ();
 sg13g2_fill_2 FILLER_20_1201 ();
 sg13g2_fill_2 FILLER_20_1229 ();
 sg13g2_fill_1 FILLER_20_1258 ();
 sg13g2_fill_2 FILLER_20_1292 ();
 sg13g2_fill_2 FILLER_20_1304 ();
 sg13g2_fill_1 FILLER_20_1306 ();
 sg13g2_fill_1 FILLER_20_1333 ();
 sg13g2_decap_8 FILLER_20_1342 ();
 sg13g2_fill_2 FILLER_20_1349 ();
 sg13g2_fill_1 FILLER_20_1351 ();
 sg13g2_fill_2 FILLER_20_1356 ();
 sg13g2_fill_1 FILLER_20_1358 ();
 sg13g2_decap_8 FILLER_20_1362 ();
 sg13g2_decap_8 FILLER_20_1369 ();
 sg13g2_fill_1 FILLER_20_1379 ();
 sg13g2_fill_1 FILLER_20_1390 ();
 sg13g2_fill_1 FILLER_20_1401 ();
 sg13g2_fill_2 FILLER_20_1421 ();
 sg13g2_decap_4 FILLER_20_1428 ();
 sg13g2_fill_1 FILLER_20_1432 ();
 sg13g2_fill_1 FILLER_20_1454 ();
 sg13g2_decap_4 FILLER_20_1462 ();
 sg13g2_fill_1 FILLER_20_1471 ();
 sg13g2_fill_1 FILLER_20_1476 ();
 sg13g2_fill_2 FILLER_20_1482 ();
 sg13g2_fill_2 FILLER_20_1491 ();
 sg13g2_fill_1 FILLER_20_1493 ();
 sg13g2_fill_2 FILLER_20_1514 ();
 sg13g2_fill_1 FILLER_20_1516 ();
 sg13g2_decap_4 FILLER_20_1530 ();
 sg13g2_fill_1 FILLER_20_1539 ();
 sg13g2_fill_1 FILLER_20_1545 ();
 sg13g2_fill_1 FILLER_20_1550 ();
 sg13g2_fill_1 FILLER_20_1560 ();
 sg13g2_fill_2 FILLER_20_1566 ();
 sg13g2_fill_1 FILLER_20_1568 ();
 sg13g2_decap_4 FILLER_20_1574 ();
 sg13g2_fill_2 FILLER_20_1639 ();
 sg13g2_fill_1 FILLER_20_1641 ();
 sg13g2_fill_1 FILLER_20_1678 ();
 sg13g2_fill_1 FILLER_20_1691 ();
 sg13g2_fill_1 FILLER_20_1699 ();
 sg13g2_fill_1 FILLER_20_1770 ();
 sg13g2_fill_2 FILLER_20_1776 ();
 sg13g2_fill_2 FILLER_20_1791 ();
 sg13g2_fill_2 FILLER_20_1798 ();
 sg13g2_fill_1 FILLER_20_1804 ();
 sg13g2_fill_1 FILLER_20_1808 ();
 sg13g2_fill_1 FILLER_20_1812 ();
 sg13g2_fill_1 FILLER_20_1845 ();
 sg13g2_fill_1 FILLER_20_1850 ();
 sg13g2_fill_1 FILLER_20_1855 ();
 sg13g2_fill_2 FILLER_20_1877 ();
 sg13g2_fill_1 FILLER_20_1918 ();
 sg13g2_decap_8 FILLER_20_1955 ();
 sg13g2_decap_8 FILLER_20_1962 ();
 sg13g2_fill_1 FILLER_20_1995 ();
 sg13g2_decap_8 FILLER_20_2062 ();
 sg13g2_decap_8 FILLER_20_2069 ();
 sg13g2_fill_1 FILLER_20_2076 ();
 sg13g2_fill_2 FILLER_20_2085 ();
 sg13g2_fill_1 FILLER_20_2087 ();
 sg13g2_decap_8 FILLER_20_2123 ();
 sg13g2_fill_1 FILLER_20_2130 ();
 sg13g2_fill_2 FILLER_20_2163 ();
 sg13g2_decap_8 FILLER_20_2172 ();
 sg13g2_fill_2 FILLER_20_2179 ();
 sg13g2_fill_1 FILLER_20_2181 ();
 sg13g2_fill_2 FILLER_20_2262 ();
 sg13g2_fill_2 FILLER_20_2316 ();
 sg13g2_fill_2 FILLER_20_2332 ();
 sg13g2_fill_1 FILLER_20_2334 ();
 sg13g2_fill_1 FILLER_20_2339 ();
 sg13g2_fill_2 FILLER_20_2344 ();
 sg13g2_decap_4 FILLER_20_2376 ();
 sg13g2_fill_1 FILLER_20_2380 ();
 sg13g2_fill_1 FILLER_20_2390 ();
 sg13g2_fill_1 FILLER_20_2417 ();
 sg13g2_fill_2 FILLER_20_2474 ();
 sg13g2_decap_8 FILLER_20_2518 ();
 sg13g2_fill_2 FILLER_20_2529 ();
 sg13g2_fill_1 FILLER_20_2531 ();
 sg13g2_fill_1 FILLER_20_2592 ();
 sg13g2_decap_4 FILLER_20_2599 ();
 sg13g2_fill_2 FILLER_20_2609 ();
 sg13g2_fill_2 FILLER_20_2628 ();
 sg13g2_fill_1 FILLER_20_2630 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_4 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_44 ();
 sg13g2_fill_1 FILLER_21_55 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_134 ();
 sg13g2_decap_8 FILLER_21_171 ();
 sg13g2_fill_2 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_186 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_195 ();
 sg13g2_decap_4 FILLER_21_201 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_211 ();
 sg13g2_decap_8 FILLER_21_218 ();
 sg13g2_decap_8 FILLER_21_225 ();
 sg13g2_decap_4 FILLER_21_232 ();
 sg13g2_decap_4 FILLER_21_241 ();
 sg13g2_fill_1 FILLER_21_245 ();
 sg13g2_fill_1 FILLER_21_258 ();
 sg13g2_decap_4 FILLER_21_269 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_342 ();
 sg13g2_decap_4 FILLER_21_349 ();
 sg13g2_fill_1 FILLER_21_353 ();
 sg13g2_fill_2 FILLER_21_359 ();
 sg13g2_fill_2 FILLER_21_365 ();
 sg13g2_fill_1 FILLER_21_367 ();
 sg13g2_decap_4 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_4 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_fill_1 FILLER_21_412 ();
 sg13g2_fill_2 FILLER_21_423 ();
 sg13g2_fill_1 FILLER_21_474 ();
 sg13g2_fill_1 FILLER_21_510 ();
 sg13g2_decap_8 FILLER_21_543 ();
 sg13g2_fill_2 FILLER_21_550 ();
 sg13g2_fill_1 FILLER_21_552 ();
 sg13g2_decap_4 FILLER_21_557 ();
 sg13g2_fill_1 FILLER_21_565 ();
 sg13g2_fill_2 FILLER_21_571 ();
 sg13g2_fill_1 FILLER_21_573 ();
 sg13g2_fill_1 FILLER_21_590 ();
 sg13g2_fill_2 FILLER_21_596 ();
 sg13g2_fill_1 FILLER_21_602 ();
 sg13g2_fill_1 FILLER_21_608 ();
 sg13g2_fill_1 FILLER_21_620 ();
 sg13g2_decap_4 FILLER_21_662 ();
 sg13g2_fill_2 FILLER_21_666 ();
 sg13g2_decap_4 FILLER_21_673 ();
 sg13g2_fill_1 FILLER_21_677 ();
 sg13g2_fill_1 FILLER_21_683 ();
 sg13g2_fill_2 FILLER_21_692 ();
 sg13g2_fill_1 FILLER_21_694 ();
 sg13g2_decap_4 FILLER_21_700 ();
 sg13g2_fill_1 FILLER_21_704 ();
 sg13g2_fill_2 FILLER_21_719 ();
 sg13g2_fill_1 FILLER_21_721 ();
 sg13g2_fill_1 FILLER_21_728 ();
 sg13g2_fill_2 FILLER_21_734 ();
 sg13g2_fill_1 FILLER_21_741 ();
 sg13g2_fill_2 FILLER_21_747 ();
 sg13g2_decap_8 FILLER_21_753 ();
 sg13g2_fill_2 FILLER_21_760 ();
 sg13g2_fill_1 FILLER_21_762 ();
 sg13g2_fill_1 FILLER_21_768 ();
 sg13g2_fill_2 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_4 FILLER_21_803 ();
 sg13g2_fill_2 FILLER_21_812 ();
 sg13g2_fill_1 FILLER_21_814 ();
 sg13g2_fill_1 FILLER_21_820 ();
 sg13g2_decap_4 FILLER_21_827 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_842 ();
 sg13g2_decap_8 FILLER_21_849 ();
 sg13g2_fill_2 FILLER_21_856 ();
 sg13g2_fill_1 FILLER_21_858 ();
 sg13g2_fill_1 FILLER_21_875 ();
 sg13g2_fill_1 FILLER_21_916 ();
 sg13g2_fill_2 FILLER_21_927 ();
 sg13g2_decap_8 FILLER_21_959 ();
 sg13g2_decap_8 FILLER_21_966 ();
 sg13g2_fill_1 FILLER_21_973 ();
 sg13g2_decap_8 FILLER_21_995 ();
 sg13g2_decap_4 FILLER_21_1002 ();
 sg13g2_fill_2 FILLER_21_1006 ();
 sg13g2_fill_2 FILLER_21_1012 ();
 sg13g2_fill_1 FILLER_21_1014 ();
 sg13g2_decap_8 FILLER_21_1027 ();
 sg13g2_decap_8 FILLER_21_1034 ();
 sg13g2_decap_8 FILLER_21_1041 ();
 sg13g2_decap_8 FILLER_21_1052 ();
 sg13g2_fill_2 FILLER_21_1059 ();
 sg13g2_fill_2 FILLER_21_1070 ();
 sg13g2_fill_1 FILLER_21_1072 ();
 sg13g2_fill_1 FILLER_21_1109 ();
 sg13g2_decap_8 FILLER_21_1149 ();
 sg13g2_decap_8 FILLER_21_1156 ();
 sg13g2_fill_1 FILLER_21_1163 ();
 sg13g2_fill_2 FILLER_21_1168 ();
 sg13g2_fill_1 FILLER_21_1249 ();
 sg13g2_fill_2 FILLER_21_1260 ();
 sg13g2_fill_1 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1276 ();
 sg13g2_fill_2 FILLER_21_1283 ();
 sg13g2_fill_1 FILLER_21_1285 ();
 sg13g2_fill_1 FILLER_21_1315 ();
 sg13g2_fill_2 FILLER_21_1320 ();
 sg13g2_decap_8 FILLER_21_1326 ();
 sg13g2_fill_1 FILLER_21_1369 ();
 sg13g2_fill_2 FILLER_21_1379 ();
 sg13g2_fill_1 FILLER_21_1396 ();
 sg13g2_fill_1 FILLER_21_1408 ();
 sg13g2_decap_8 FILLER_21_1424 ();
 sg13g2_fill_1 FILLER_21_1460 ();
 sg13g2_fill_2 FILLER_21_1470 ();
 sg13g2_fill_2 FILLER_21_1477 ();
 sg13g2_fill_1 FILLER_21_1479 ();
 sg13g2_fill_2 FILLER_21_1485 ();
 sg13g2_fill_2 FILLER_21_1492 ();
 sg13g2_fill_1 FILLER_21_1515 ();
 sg13g2_decap_4 FILLER_21_1522 ();
 sg13g2_fill_1 FILLER_21_1526 ();
 sg13g2_decap_4 FILLER_21_1532 ();
 sg13g2_fill_2 FILLER_21_1536 ();
 sg13g2_decap_8 FILLER_21_1568 ();
 sg13g2_fill_1 FILLER_21_1575 ();
 sg13g2_fill_2 FILLER_21_1582 ();
 sg13g2_decap_4 FILLER_21_1588 ();
 sg13g2_fill_2 FILLER_21_1603 ();
 sg13g2_fill_1 FILLER_21_1618 ();
 sg13g2_decap_8 FILLER_21_1641 ();
 sg13g2_decap_4 FILLER_21_1648 ();
 sg13g2_fill_2 FILLER_21_1652 ();
 sg13g2_fill_1 FILLER_21_1658 ();
 sg13g2_fill_1 FILLER_21_1695 ();
 sg13g2_fill_2 FILLER_21_1708 ();
 sg13g2_fill_2 FILLER_21_1753 ();
 sg13g2_decap_8 FILLER_21_1772 ();
 sg13g2_fill_2 FILLER_21_1790 ();
 sg13g2_fill_2 FILLER_21_1800 ();
 sg13g2_fill_2 FILLER_21_1812 ();
 sg13g2_decap_8 FILLER_21_1833 ();
 sg13g2_fill_2 FILLER_21_1840 ();
 sg13g2_decap_8 FILLER_21_1848 ();
 sg13g2_decap_8 FILLER_21_1855 ();
 sg13g2_decap_8 FILLER_21_1862 ();
 sg13g2_fill_2 FILLER_21_1869 ();
 sg13g2_fill_1 FILLER_21_1871 ();
 sg13g2_fill_1 FILLER_21_1876 ();
 sg13g2_fill_1 FILLER_21_1882 ();
 sg13g2_fill_1 FILLER_21_1888 ();
 sg13g2_fill_1 FILLER_21_1894 ();
 sg13g2_fill_2 FILLER_21_1899 ();
 sg13g2_fill_2 FILLER_21_1911 ();
 sg13g2_fill_1 FILLER_21_1936 ();
 sg13g2_fill_2 FILLER_21_1963 ();
 sg13g2_fill_1 FILLER_21_1965 ();
 sg13g2_fill_2 FILLER_21_1976 ();
 sg13g2_fill_1 FILLER_21_1978 ();
 sg13g2_fill_2 FILLER_21_2005 ();
 sg13g2_fill_2 FILLER_21_2050 ();
 sg13g2_fill_2 FILLER_21_2062 ();
 sg13g2_fill_2 FILLER_21_2108 ();
 sg13g2_fill_2 FILLER_21_2120 ();
 sg13g2_fill_1 FILLER_21_2122 ();
 sg13g2_decap_4 FILLER_21_2185 ();
 sg13g2_fill_2 FILLER_21_2189 ();
 sg13g2_decap_4 FILLER_21_2201 ();
 sg13g2_fill_2 FILLER_21_2205 ();
 sg13g2_fill_1 FILLER_21_2211 ();
 sg13g2_decap_8 FILLER_21_2246 ();
 sg13g2_decap_4 FILLER_21_2253 ();
 sg13g2_fill_1 FILLER_21_2257 ();
 sg13g2_decap_8 FILLER_21_2279 ();
 sg13g2_decap_8 FILLER_21_2286 ();
 sg13g2_decap_8 FILLER_21_2293 ();
 sg13g2_decap_4 FILLER_21_2300 ();
 sg13g2_fill_1 FILLER_21_2304 ();
 sg13g2_fill_1 FILLER_21_2334 ();
 sg13g2_fill_1 FILLER_21_2339 ();
 sg13g2_fill_1 FILLER_21_2346 ();
 sg13g2_fill_1 FILLER_21_2351 ();
 sg13g2_decap_8 FILLER_21_2356 ();
 sg13g2_fill_2 FILLER_21_2369 ();
 sg13g2_fill_2 FILLER_21_2402 ();
 sg13g2_fill_1 FILLER_21_2404 ();
 sg13g2_fill_1 FILLER_21_2415 ();
 sg13g2_fill_2 FILLER_21_2430 ();
 sg13g2_fill_1 FILLER_21_2432 ();
 sg13g2_decap_4 FILLER_21_2437 ();
 sg13g2_fill_2 FILLER_21_2455 ();
 sg13g2_fill_1 FILLER_21_2457 ();
 sg13g2_fill_2 FILLER_21_2468 ();
 sg13g2_fill_1 FILLER_21_2470 ();
 sg13g2_decap_8 FILLER_21_2505 ();
 sg13g2_decap_8 FILLER_21_2512 ();
 sg13g2_fill_2 FILLER_21_2519 ();
 sg13g2_decap_8 FILLER_21_2551 ();
 sg13g2_decap_8 FILLER_21_2558 ();
 sg13g2_decap_8 FILLER_21_2565 ();
 sg13g2_fill_2 FILLER_21_2582 ();
 sg13g2_fill_2 FILLER_21_2594 ();
 sg13g2_fill_1 FILLER_21_2596 ();
 sg13g2_decap_4 FILLER_21_2638 ();
 sg13g2_fill_2 FILLER_21_2668 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_7 ();
 sg13g2_decap_4 FILLER_22_16 ();
 sg13g2_fill_2 FILLER_22_20 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_162 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_2 FILLER_22_296 ();
 sg13g2_fill_1 FILLER_22_302 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_fill_2 FILLER_22_393 ();
 sg13g2_fill_1 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_decap_4 FILLER_22_429 ();
 sg13g2_fill_2 FILLER_22_433 ();
 sg13g2_fill_2 FILLER_22_466 ();
 sg13g2_fill_1 FILLER_22_468 ();
 sg13g2_fill_1 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_509 ();
 sg13g2_decap_8 FILLER_22_516 ();
 sg13g2_fill_2 FILLER_22_523 ();
 sg13g2_fill_1 FILLER_22_525 ();
 sg13g2_fill_2 FILLER_22_535 ();
 sg13g2_fill_1 FILLER_22_537 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_fill_1 FILLER_22_566 ();
 sg13g2_fill_2 FILLER_22_593 ();
 sg13g2_fill_1 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_631 ();
 sg13g2_fill_2 FILLER_22_695 ();
 sg13g2_fill_1 FILLER_22_697 ();
 sg13g2_fill_2 FILLER_22_703 ();
 sg13g2_fill_2 FILLER_22_757 ();
 sg13g2_fill_1 FILLER_22_764 ();
 sg13g2_fill_1 FILLER_22_769 ();
 sg13g2_fill_2 FILLER_22_801 ();
 sg13g2_decap_4 FILLER_22_816 ();
 sg13g2_fill_1 FILLER_22_820 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_decap_4 FILLER_22_840 ();
 sg13g2_fill_2 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_fill_1 FILLER_22_914 ();
 sg13g2_fill_2 FILLER_22_946 ();
 sg13g2_decap_8 FILLER_22_973 ();
 sg13g2_decap_8 FILLER_22_980 ();
 sg13g2_decap_8 FILLER_22_987 ();
 sg13g2_decap_8 FILLER_22_994 ();
 sg13g2_decap_8 FILLER_22_1001 ();
 sg13g2_decap_8 FILLER_22_1008 ();
 sg13g2_decap_8 FILLER_22_1015 ();
 sg13g2_decap_8 FILLER_22_1022 ();
 sg13g2_decap_4 FILLER_22_1029 ();
 sg13g2_fill_2 FILLER_22_1033 ();
 sg13g2_decap_8 FILLER_22_1039 ();
 sg13g2_decap_8 FILLER_22_1046 ();
 sg13g2_fill_2 FILLER_22_1053 ();
 sg13g2_fill_1 FILLER_22_1055 ();
 sg13g2_decap_8 FILLER_22_1147 ();
 sg13g2_decap_8 FILLER_22_1154 ();
 sg13g2_decap_8 FILLER_22_1161 ();
 sg13g2_fill_1 FILLER_22_1168 ();
 sg13g2_fill_1 FILLER_22_1240 ();
 sg13g2_fill_2 FILLER_22_1244 ();
 sg13g2_fill_1 FILLER_22_1249 ();
 sg13g2_decap_8 FILLER_22_1279 ();
 sg13g2_fill_2 FILLER_22_1286 ();
 sg13g2_fill_1 FILLER_22_1288 ();
 sg13g2_decap_8 FILLER_22_1292 ();
 sg13g2_decap_8 FILLER_22_1299 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_decap_4 FILLER_22_1313 ();
 sg13g2_decap_8 FILLER_22_1351 ();
 sg13g2_decap_8 FILLER_22_1358 ();
 sg13g2_decap_8 FILLER_22_1365 ();
 sg13g2_decap_8 FILLER_22_1372 ();
 sg13g2_decap_4 FILLER_22_1379 ();
 sg13g2_fill_1 FILLER_22_1383 ();
 sg13g2_fill_2 FILLER_22_1394 ();
 sg13g2_fill_1 FILLER_22_1401 ();
 sg13g2_decap_4 FILLER_22_1407 ();
 sg13g2_fill_1 FILLER_22_1418 ();
 sg13g2_fill_2 FILLER_22_1424 ();
 sg13g2_decap_4 FILLER_22_1432 ();
 sg13g2_fill_2 FILLER_22_1436 ();
 sg13g2_decap_4 FILLER_22_1467 ();
 sg13g2_fill_2 FILLER_22_1471 ();
 sg13g2_fill_1 FILLER_22_1478 ();
 sg13g2_fill_2 FILLER_22_1484 ();
 sg13g2_decap_4 FILLER_22_1503 ();
 sg13g2_fill_2 FILLER_22_1517 ();
 sg13g2_fill_1 FILLER_22_1519 ();
 sg13g2_decap_4 FILLER_22_1532 ();
 sg13g2_fill_2 FILLER_22_1536 ();
 sg13g2_decap_4 FILLER_22_1553 ();
 sg13g2_decap_4 FILLER_22_1574 ();
 sg13g2_fill_2 FILLER_22_1582 ();
 sg13g2_fill_1 FILLER_22_1584 ();
 sg13g2_fill_2 FILLER_22_1593 ();
 sg13g2_fill_1 FILLER_22_1595 ();
 sg13g2_decap_8 FILLER_22_1636 ();
 sg13g2_decap_8 FILLER_22_1643 ();
 sg13g2_decap_4 FILLER_22_1650 ();
 sg13g2_fill_1 FILLER_22_1654 ();
 sg13g2_fill_2 FILLER_22_1674 ();
 sg13g2_fill_1 FILLER_22_1705 ();
 sg13g2_fill_1 FILLER_22_1718 ();
 sg13g2_fill_1 FILLER_22_1726 ();
 sg13g2_fill_2 FILLER_22_1754 ();
 sg13g2_fill_1 FILLER_22_1772 ();
 sg13g2_fill_1 FILLER_22_1807 ();
 sg13g2_decap_8 FILLER_22_1859 ();
 sg13g2_decap_8 FILLER_22_1866 ();
 sg13g2_decap_4 FILLER_22_1873 ();
 sg13g2_fill_1 FILLER_22_1895 ();
 sg13g2_decap_8 FILLER_22_1900 ();
 sg13g2_decap_4 FILLER_22_1907 ();
 sg13g2_fill_1 FILLER_22_1911 ();
 sg13g2_decap_4 FILLER_22_1916 ();
 sg13g2_fill_2 FILLER_22_1934 ();
 sg13g2_fill_1 FILLER_22_1946 ();
 sg13g2_decap_8 FILLER_22_1951 ();
 sg13g2_decap_8 FILLER_22_1958 ();
 sg13g2_fill_1 FILLER_22_1965 ();
 sg13g2_fill_2 FILLER_22_2007 ();
 sg13g2_fill_2 FILLER_22_2076 ();
 sg13g2_fill_1 FILLER_22_2078 ();
 sg13g2_decap_4 FILLER_22_2093 ();
 sg13g2_fill_1 FILLER_22_2123 ();
 sg13g2_decap_4 FILLER_22_2170 ();
 sg13g2_fill_1 FILLER_22_2174 ();
 sg13g2_fill_2 FILLER_22_2188 ();
 sg13g2_decap_4 FILLER_22_2194 ();
 sg13g2_fill_1 FILLER_22_2228 ();
 sg13g2_decap_8 FILLER_22_2239 ();
 sg13g2_decap_8 FILLER_22_2246 ();
 sg13g2_fill_2 FILLER_22_2253 ();
 sg13g2_fill_1 FILLER_22_2255 ();
 sg13g2_fill_1 FILLER_22_2266 ();
 sg13g2_decap_8 FILLER_22_2293 ();
 sg13g2_fill_2 FILLER_22_2300 ();
 sg13g2_fill_2 FILLER_22_2328 ();
 sg13g2_fill_1 FILLER_22_2330 ();
 sg13g2_fill_2 FILLER_22_2341 ();
 sg13g2_decap_8 FILLER_22_2348 ();
 sg13g2_decap_8 FILLER_22_2355 ();
 sg13g2_decap_4 FILLER_22_2362 ();
 sg13g2_fill_1 FILLER_22_2366 ();
 sg13g2_decap_8 FILLER_22_2391 ();
 sg13g2_decap_8 FILLER_22_2398 ();
 sg13g2_fill_2 FILLER_22_2405 ();
 sg13g2_fill_1 FILLER_22_2407 ();
 sg13g2_decap_8 FILLER_22_2414 ();
 sg13g2_decap_8 FILLER_22_2421 ();
 sg13g2_decap_8 FILLER_22_2428 ();
 sg13g2_decap_8 FILLER_22_2435 ();
 sg13g2_decap_8 FILLER_22_2442 ();
 sg13g2_decap_8 FILLER_22_2449 ();
 sg13g2_fill_1 FILLER_22_2456 ();
 sg13g2_fill_2 FILLER_22_2468 ();
 sg13g2_fill_1 FILLER_22_2470 ();
 sg13g2_fill_1 FILLER_22_2476 ();
 sg13g2_fill_2 FILLER_22_2491 ();
 sg13g2_decap_8 FILLER_22_2503 ();
 sg13g2_decap_8 FILLER_22_2510 ();
 sg13g2_fill_2 FILLER_22_2517 ();
 sg13g2_fill_1 FILLER_22_2519 ();
 sg13g2_fill_2 FILLER_22_2530 ();
 sg13g2_fill_1 FILLER_22_2532 ();
 sg13g2_decap_4 FILLER_22_2539 ();
 sg13g2_fill_1 FILLER_22_2543 ();
 sg13g2_decap_4 FILLER_22_2549 ();
 sg13g2_fill_1 FILLER_22_2553 ();
 sg13g2_decap_4 FILLER_22_2558 ();
 sg13g2_decap_8 FILLER_22_2566 ();
 sg13g2_decap_8 FILLER_22_2573 ();
 sg13g2_decap_8 FILLER_22_2585 ();
 sg13g2_decap_8 FILLER_22_2592 ();
 sg13g2_decap_4 FILLER_22_2599 ();
 sg13g2_fill_2 FILLER_22_2603 ();
 sg13g2_decap_8 FILLER_22_2609 ();
 sg13g2_decap_8 FILLER_22_2616 ();
 sg13g2_decap_8 FILLER_22_2623 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_32 ();
 sg13g2_fill_1 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_fill_1 FILLER_23_123 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_214 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_decap_4 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_318 ();
 sg13g2_decap_4 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_2 FILLER_23_339 ();
 sg13g2_fill_1 FILLER_23_341 ();
 sg13g2_decap_4 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_fill_2 FILLER_23_403 ();
 sg13g2_fill_1 FILLER_23_405 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_419 ();
 sg13g2_fill_1 FILLER_23_426 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_fill_1 FILLER_23_488 ();
 sg13g2_fill_1 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_fill_2 FILLER_23_525 ();
 sg13g2_fill_1 FILLER_23_527 ();
 sg13g2_decap_4 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_542 ();
 sg13g2_fill_1 FILLER_23_548 ();
 sg13g2_decap_8 FILLER_23_584 ();
 sg13g2_decap_8 FILLER_23_591 ();
 sg13g2_fill_1 FILLER_23_598 ();
 sg13g2_decap_8 FILLER_23_625 ();
 sg13g2_decap_8 FILLER_23_632 ();
 sg13g2_decap_4 FILLER_23_639 ();
 sg13g2_fill_2 FILLER_23_643 ();
 sg13g2_decap_8 FILLER_23_649 ();
 sg13g2_fill_2 FILLER_23_656 ();
 sg13g2_fill_1 FILLER_23_658 ();
 sg13g2_fill_1 FILLER_23_675 ();
 sg13g2_decap_8 FILLER_23_680 ();
 sg13g2_fill_1 FILLER_23_687 ();
 sg13g2_fill_2 FILLER_23_721 ();
 sg13g2_fill_2 FILLER_23_728 ();
 sg13g2_fill_1 FILLER_23_730 ();
 sg13g2_decap_4 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_739 ();
 sg13g2_fill_1 FILLER_23_774 ();
 sg13g2_fill_2 FILLER_23_798 ();
 sg13g2_decap_4 FILLER_23_840 ();
 sg13g2_fill_1 FILLER_23_879 ();
 sg13g2_fill_2 FILLER_23_890 ();
 sg13g2_fill_1 FILLER_23_935 ();
 sg13g2_fill_2 FILLER_23_941 ();
 sg13g2_decap_8 FILLER_23_974 ();
 sg13g2_fill_1 FILLER_23_981 ();
 sg13g2_decap_8 FILLER_23_995 ();
 sg13g2_fill_2 FILLER_23_1002 ();
 sg13g2_fill_2 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1036 ();
 sg13g2_decap_4 FILLER_23_1043 ();
 sg13g2_fill_1 FILLER_23_1081 ();
 sg13g2_fill_1 FILLER_23_1107 ();
 sg13g2_fill_1 FILLER_23_1113 ();
 sg13g2_fill_1 FILLER_23_1127 ();
 sg13g2_fill_2 FILLER_23_1133 ();
 sg13g2_fill_2 FILLER_23_1160 ();
 sg13g2_fill_1 FILLER_23_1192 ();
 sg13g2_fill_2 FILLER_23_1202 ();
 sg13g2_decap_8 FILLER_23_1257 ();
 sg13g2_decap_8 FILLER_23_1264 ();
 sg13g2_decap_8 FILLER_23_1271 ();
 sg13g2_fill_2 FILLER_23_1282 ();
 sg13g2_decap_8 FILLER_23_1310 ();
 sg13g2_fill_2 FILLER_23_1317 ();
 sg13g2_fill_1 FILLER_23_1319 ();
 sg13g2_decap_8 FILLER_23_1340 ();
 sg13g2_decap_8 FILLER_23_1347 ();
 sg13g2_decap_8 FILLER_23_1354 ();
 sg13g2_decap_8 FILLER_23_1361 ();
 sg13g2_decap_8 FILLER_23_1404 ();
 sg13g2_fill_2 FILLER_23_1416 ();
 sg13g2_fill_1 FILLER_23_1418 ();
 sg13g2_decap_8 FILLER_23_1423 ();
 sg13g2_decap_8 FILLER_23_1430 ();
 sg13g2_decap_8 FILLER_23_1437 ();
 sg13g2_decap_4 FILLER_23_1444 ();
 sg13g2_decap_4 FILLER_23_1468 ();
 sg13g2_fill_2 FILLER_23_1472 ();
 sg13g2_decap_8 FILLER_23_1478 ();
 sg13g2_decap_4 FILLER_23_1494 ();
 sg13g2_fill_1 FILLER_23_1503 ();
 sg13g2_fill_2 FILLER_23_1531 ();
 sg13g2_fill_2 FILLER_23_1542 ();
 sg13g2_decap_8 FILLER_23_1549 ();
 sg13g2_decap_4 FILLER_23_1556 ();
 sg13g2_fill_1 FILLER_23_1560 ();
 sg13g2_decap_8 FILLER_23_1582 ();
 sg13g2_decap_4 FILLER_23_1589 ();
 sg13g2_fill_1 FILLER_23_1593 ();
 sg13g2_decap_4 FILLER_23_1607 ();
 sg13g2_decap_8 FILLER_23_1651 ();
 sg13g2_fill_2 FILLER_23_1658 ();
 sg13g2_fill_1 FILLER_23_1660 ();
 sg13g2_decap_4 FILLER_23_1664 ();
 sg13g2_fill_1 FILLER_23_1668 ();
 sg13g2_fill_2 FILLER_23_1676 ();
 sg13g2_fill_1 FILLER_23_1700 ();
 sg13g2_fill_2 FILLER_23_1722 ();
 sg13g2_fill_2 FILLER_23_1732 ();
 sg13g2_fill_2 FILLER_23_1798 ();
 sg13g2_fill_1 FILLER_23_1919 ();
 sg13g2_fill_2 FILLER_23_1924 ();
 sg13g2_fill_1 FILLER_23_1926 ();
 sg13g2_decap_8 FILLER_23_1945 ();
 sg13g2_decap_4 FILLER_23_1952 ();
 sg13g2_fill_2 FILLER_23_1956 ();
 sg13g2_fill_2 FILLER_23_1967 ();
 sg13g2_fill_1 FILLER_23_1969 ();
 sg13g2_fill_1 FILLER_23_1977 ();
 sg13g2_fill_1 FILLER_23_1983 ();
 sg13g2_fill_2 FILLER_23_2015 ();
 sg13g2_fill_2 FILLER_23_2027 ();
 sg13g2_fill_2 FILLER_23_2066 ();
 sg13g2_fill_1 FILLER_23_2068 ();
 sg13g2_fill_2 FILLER_23_2084 ();
 sg13g2_fill_1 FILLER_23_2112 ();
 sg13g2_fill_1 FILLER_23_2134 ();
 sg13g2_decap_4 FILLER_23_2165 ();
 sg13g2_fill_2 FILLER_23_2169 ();
 sg13g2_fill_2 FILLER_23_2192 ();
 sg13g2_fill_1 FILLER_23_2194 ();
 sg13g2_decap_8 FILLER_23_2199 ();
 sg13g2_fill_2 FILLER_23_2206 ();
 sg13g2_decap_8 FILLER_23_2218 ();
 sg13g2_decap_4 FILLER_23_2225 ();
 sg13g2_decap_8 FILLER_23_2289 ();
 sg13g2_decap_8 FILLER_23_2296 ();
 sg13g2_decap_4 FILLER_23_2303 ();
 sg13g2_fill_2 FILLER_23_2307 ();
 sg13g2_decap_8 FILLER_23_2313 ();
 sg13g2_decap_8 FILLER_23_2320 ();
 sg13g2_decap_8 FILLER_23_2327 ();
 sg13g2_fill_1 FILLER_23_2334 ();
 sg13g2_fill_2 FILLER_23_2348 ();
 sg13g2_fill_2 FILLER_23_2391 ();
 sg13g2_fill_2 FILLER_23_2399 ();
 sg13g2_fill_1 FILLER_23_2411 ();
 sg13g2_decap_8 FILLER_23_2417 ();
 sg13g2_decap_8 FILLER_23_2424 ();
 sg13g2_decap_8 FILLER_23_2431 ();
 sg13g2_fill_1 FILLER_23_2438 ();
 sg13g2_fill_2 FILLER_23_2449 ();
 sg13g2_fill_1 FILLER_23_2451 ();
 sg13g2_decap_4 FILLER_23_2536 ();
 sg13g2_fill_2 FILLER_23_2590 ();
 sg13g2_fill_1 FILLER_23_2602 ();
 sg13g2_fill_1 FILLER_23_2629 ();
 sg13g2_fill_1 FILLER_23_2656 ();
 sg13g2_decap_8 FILLER_23_2661 ();
 sg13g2_fill_2 FILLER_23_2668 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_51 ();
 sg13g2_fill_2 FILLER_24_71 ();
 sg13g2_fill_1 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_157 ();
 sg13g2_fill_1 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_248 ();
 sg13g2_fill_2 FILLER_24_259 ();
 sg13g2_fill_2 FILLER_24_274 ();
 sg13g2_decap_8 FILLER_24_281 ();
 sg13g2_decap_8 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_fill_1 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_426 ();
 sg13g2_fill_1 FILLER_24_428 ();
 sg13g2_fill_1 FILLER_24_439 ();
 sg13g2_decap_4 FILLER_24_449 ();
 sg13g2_decap_8 FILLER_24_463 ();
 sg13g2_decap_8 FILLER_24_470 ();
 sg13g2_decap_8 FILLER_24_477 ();
 sg13g2_fill_2 FILLER_24_484 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_4 FILLER_24_504 ();
 sg13g2_fill_1 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_545 ();
 sg13g2_fill_2 FILLER_24_552 ();
 sg13g2_fill_1 FILLER_24_554 ();
 sg13g2_decap_4 FILLER_24_559 ();
 sg13g2_fill_1 FILLER_24_563 ();
 sg13g2_fill_1 FILLER_24_569 ();
 sg13g2_fill_1 FILLER_24_586 ();
 sg13g2_fill_1 FILLER_24_590 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_fill_1 FILLER_24_620 ();
 sg13g2_fill_2 FILLER_24_634 ();
 sg13g2_fill_1 FILLER_24_636 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_fill_2 FILLER_24_674 ();
 sg13g2_fill_2 FILLER_24_706 ();
 sg13g2_fill_1 FILLER_24_708 ();
 sg13g2_decap_4 FILLER_24_713 ();
 sg13g2_fill_1 FILLER_24_717 ();
 sg13g2_decap_4 FILLER_24_722 ();
 sg13g2_fill_1 FILLER_24_726 ();
 sg13g2_fill_1 FILLER_24_842 ();
 sg13g2_fill_2 FILLER_24_892 ();
 sg13g2_decap_8 FILLER_24_915 ();
 sg13g2_fill_1 FILLER_24_941 ();
 sg13g2_decap_8 FILLER_24_959 ();
 sg13g2_decap_4 FILLER_24_966 ();
 sg13g2_fill_2 FILLER_24_1001 ();
 sg13g2_fill_1 FILLER_24_1003 ();
 sg13g2_decap_4 FILLER_24_1029 ();
 sg13g2_fill_2 FILLER_24_1033 ();
 sg13g2_decap_8 FILLER_24_1039 ();
 sg13g2_fill_2 FILLER_24_1046 ();
 sg13g2_fill_1 FILLER_24_1048 ();
 sg13g2_decap_8 FILLER_24_1062 ();
 sg13g2_decap_8 FILLER_24_1069 ();
 sg13g2_fill_1 FILLER_24_1085 ();
 sg13g2_fill_2 FILLER_24_1108 ();
 sg13g2_fill_1 FILLER_24_1110 ();
 sg13g2_decap_4 FILLER_24_1116 ();
 sg13g2_fill_2 FILLER_24_1159 ();
 sg13g2_fill_2 FILLER_24_1169 ();
 sg13g2_fill_1 FILLER_24_1171 ();
 sg13g2_fill_2 FILLER_24_1177 ();
 sg13g2_fill_1 FILLER_24_1179 ();
 sg13g2_fill_2 FILLER_24_1184 ();
 sg13g2_fill_1 FILLER_24_1186 ();
 sg13g2_fill_2 FILLER_24_1217 ();
 sg13g2_fill_1 FILLER_24_1219 ();
 sg13g2_fill_2 FILLER_24_1225 ();
 sg13g2_fill_2 FILLER_24_1234 ();
 sg13g2_decap_8 FILLER_24_1267 ();
 sg13g2_decap_8 FILLER_24_1274 ();
 sg13g2_decap_4 FILLER_24_1281 ();
 sg13g2_fill_1 FILLER_24_1299 ();
 sg13g2_decap_4 FILLER_24_1326 ();
 sg13g2_fill_2 FILLER_24_1340 ();
 sg13g2_fill_1 FILLER_24_1342 ();
 sg13g2_decap_4 FILLER_24_1369 ();
 sg13g2_fill_2 FILLER_24_1373 ();
 sg13g2_fill_2 FILLER_24_1387 ();
 sg13g2_fill_2 FILLER_24_1393 ();
 sg13g2_fill_2 FILLER_24_1400 ();
 sg13g2_fill_1 FILLER_24_1402 ();
 sg13g2_fill_2 FILLER_24_1485 ();
 sg13g2_fill_2 FILLER_24_1497 ();
 sg13g2_fill_1 FILLER_24_1499 ();
 sg13g2_fill_1 FILLER_24_1538 ();
 sg13g2_fill_1 FILLER_24_1543 ();
 sg13g2_decap_4 FILLER_24_1551 ();
 sg13g2_decap_4 FILLER_24_1559 ();
 sg13g2_fill_2 FILLER_24_1563 ();
 sg13g2_fill_1 FILLER_24_1575 ();
 sg13g2_fill_1 FILLER_24_1580 ();
 sg13g2_fill_2 FILLER_24_1593 ();
 sg13g2_fill_1 FILLER_24_1595 ();
 sg13g2_decap_8 FILLER_24_1614 ();
 sg13g2_fill_2 FILLER_24_1621 ();
 sg13g2_fill_1 FILLER_24_1623 ();
 sg13g2_decap_8 FILLER_24_1660 ();
 sg13g2_fill_2 FILLER_24_1667 ();
 sg13g2_fill_1 FILLER_24_1685 ();
 sg13g2_fill_1 FILLER_24_1694 ();
 sg13g2_fill_1 FILLER_24_1721 ();
 sg13g2_fill_1 FILLER_24_1732 ();
 sg13g2_fill_1 FILLER_24_1738 ();
 sg13g2_fill_1 FILLER_24_1744 ();
 sg13g2_fill_1 FILLER_24_1759 ();
 sg13g2_fill_2 FILLER_24_1793 ();
 sg13g2_fill_2 FILLER_24_1818 ();
 sg13g2_fill_1 FILLER_24_1820 ();
 sg13g2_fill_2 FILLER_24_1824 ();
 sg13g2_fill_2 FILLER_24_1841 ();
 sg13g2_fill_1 FILLER_24_1843 ();
 sg13g2_decap_8 FILLER_24_1864 ();
 sg13g2_decap_4 FILLER_24_1871 ();
 sg13g2_fill_1 FILLER_24_1895 ();
 sg13g2_fill_2 FILLER_24_1901 ();
 sg13g2_fill_1 FILLER_24_1903 ();
 sg13g2_fill_1 FILLER_24_1908 ();
 sg13g2_fill_2 FILLER_24_1981 ();
 sg13g2_fill_2 FILLER_24_2015 ();
 sg13g2_fill_2 FILLER_24_2053 ();
 sg13g2_decap_4 FILLER_24_2059 ();
 sg13g2_fill_1 FILLER_24_2127 ();
 sg13g2_decap_8 FILLER_24_2132 ();
 sg13g2_fill_2 FILLER_24_2139 ();
 sg13g2_fill_1 FILLER_24_2141 ();
 sg13g2_fill_2 FILLER_24_2152 ();
 sg13g2_fill_1 FILLER_24_2154 ();
 sg13g2_decap_8 FILLER_24_2192 ();
 sg13g2_fill_2 FILLER_24_2199 ();
 sg13g2_fill_1 FILLER_24_2201 ();
 sg13g2_fill_1 FILLER_24_2225 ();
 sg13g2_fill_2 FILLER_24_2256 ();
 sg13g2_fill_1 FILLER_24_2258 ();
 sg13g2_fill_1 FILLER_24_2273 ();
 sg13g2_fill_2 FILLER_24_2300 ();
 sg13g2_fill_2 FILLER_24_2335 ();
 sg13g2_fill_1 FILLER_24_2337 ();
 sg13g2_decap_8 FILLER_24_2346 ();
 sg13g2_fill_1 FILLER_24_2390 ();
 sg13g2_decap_4 FILLER_24_2423 ();
 sg13g2_fill_2 FILLER_24_2518 ();
 sg13g2_fill_1 FILLER_24_2520 ();
 sg13g2_decap_4 FILLER_24_2573 ();
 sg13g2_fill_2 FILLER_24_2577 ();
 sg13g2_fill_1 FILLER_24_2584 ();
 sg13g2_decap_8 FILLER_24_2661 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_12 ();
 sg13g2_fill_2 FILLER_25_19 ();
 sg13g2_fill_2 FILLER_25_40 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_76 ();
 sg13g2_fill_1 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_1 FILLER_25_195 ();
 sg13g2_decap_4 FILLER_25_244 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_fill_2 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_275 ();
 sg13g2_decap_8 FILLER_25_282 ();
 sg13g2_decap_8 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_310 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_359 ();
 sg13g2_decap_4 FILLER_25_365 ();
 sg13g2_fill_1 FILLER_25_369 ();
 sg13g2_decap_4 FILLER_25_375 ();
 sg13g2_fill_1 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_398 ();
 sg13g2_fill_1 FILLER_25_400 ();
 sg13g2_fill_1 FILLER_25_450 ();
 sg13g2_decap_8 FILLER_25_461 ();
 sg13g2_decap_8 FILLER_25_468 ();
 sg13g2_decap_8 FILLER_25_475 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_fill_1 FILLER_25_493 ();
 sg13g2_fill_2 FILLER_25_510 ();
 sg13g2_decap_8 FILLER_25_548 ();
 sg13g2_decap_4 FILLER_25_555 ();
 sg13g2_fill_1 FILLER_25_559 ();
 sg13g2_fill_1 FILLER_25_579 ();
 sg13g2_decap_8 FILLER_25_614 ();
 sg13g2_decap_4 FILLER_25_621 ();
 sg13g2_fill_1 FILLER_25_625 ();
 sg13g2_fill_2 FILLER_25_630 ();
 sg13g2_fill_2 FILLER_25_637 ();
 sg13g2_fill_1 FILLER_25_644 ();
 sg13g2_fill_1 FILLER_25_655 ();
 sg13g2_fill_1 FILLER_25_661 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_4 FILLER_25_674 ();
 sg13g2_decap_4 FILLER_25_682 ();
 sg13g2_fill_1 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_698 ();
 sg13g2_fill_2 FILLER_25_705 ();
 sg13g2_decap_8 FILLER_25_712 ();
 sg13g2_fill_1 FILLER_25_729 ();
 sg13g2_fill_2 FILLER_25_735 ();
 sg13g2_fill_1 FILLER_25_742 ();
 sg13g2_fill_2 FILLER_25_748 ();
 sg13g2_fill_2 FILLER_25_754 ();
 sg13g2_decap_4 FILLER_25_766 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_4 FILLER_25_812 ();
 sg13g2_fill_1 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_827 ();
 sg13g2_decap_8 FILLER_25_834 ();
 sg13g2_decap_8 FILLER_25_841 ();
 sg13g2_decap_4 FILLER_25_848 ();
 sg13g2_fill_1 FILLER_25_876 ();
 sg13g2_fill_1 FILLER_25_891 ();
 sg13g2_decap_4 FILLER_25_932 ();
 sg13g2_fill_1 FILLER_25_940 ();
 sg13g2_fill_1 FILLER_25_966 ();
 sg13g2_fill_1 FILLER_25_971 ();
 sg13g2_fill_1 FILLER_25_998 ();
 sg13g2_fill_2 FILLER_25_1004 ();
 sg13g2_fill_1 FILLER_25_1024 ();
 sg13g2_fill_2 FILLER_25_1039 ();
 sg13g2_fill_1 FILLER_25_1046 ();
 sg13g2_decap_4 FILLER_25_1096 ();
 sg13g2_decap_4 FILLER_25_1105 ();
 sg13g2_fill_2 FILLER_25_1109 ();
 sg13g2_fill_2 FILLER_25_1146 ();
 sg13g2_fill_1 FILLER_25_1148 ();
 sg13g2_decap_8 FILLER_25_1210 ();
 sg13g2_decap_4 FILLER_25_1217 ();
 sg13g2_fill_2 FILLER_25_1225 ();
 sg13g2_fill_1 FILLER_25_1240 ();
 sg13g2_fill_1 FILLER_25_1250 ();
 sg13g2_fill_1 FILLER_25_1314 ();
 sg13g2_decap_8 FILLER_25_1359 ();
 sg13g2_fill_2 FILLER_25_1366 ();
 sg13g2_decap_4 FILLER_25_1388 ();
 sg13g2_fill_2 FILLER_25_1414 ();
 sg13g2_decap_4 FILLER_25_1420 ();
 sg13g2_decap_4 FILLER_25_1429 ();
 sg13g2_fill_2 FILLER_25_1433 ();
 sg13g2_decap_8 FILLER_25_1447 ();
 sg13g2_decap_8 FILLER_25_1454 ();
 sg13g2_fill_1 FILLER_25_1466 ();
 sg13g2_fill_1 FILLER_25_1472 ();
 sg13g2_decap_8 FILLER_25_1491 ();
 sg13g2_fill_1 FILLER_25_1498 ();
 sg13g2_fill_2 FILLER_25_1503 ();
 sg13g2_fill_1 FILLER_25_1505 ();
 sg13g2_fill_2 FILLER_25_1515 ();
 sg13g2_decap_4 FILLER_25_1547 ();
 sg13g2_decap_8 FILLER_25_1608 ();
 sg13g2_decap_8 FILLER_25_1615 ();
 sg13g2_fill_2 FILLER_25_1622 ();
 sg13g2_decap_4 FILLER_25_1636 ();
 sg13g2_fill_1 FILLER_25_1640 ();
 sg13g2_decap_8 FILLER_25_1645 ();
 sg13g2_decap_8 FILLER_25_1652 ();
 sg13g2_decap_8 FILLER_25_1659 ();
 sg13g2_decap_8 FILLER_25_1666 ();
 sg13g2_fill_2 FILLER_25_1673 ();
 sg13g2_fill_1 FILLER_25_1675 ();
 sg13g2_fill_1 FILLER_25_1701 ();
 sg13g2_decap_4 FILLER_25_1738 ();
 sg13g2_fill_2 FILLER_25_1742 ();
 sg13g2_fill_2 FILLER_25_1749 ();
 sg13g2_fill_1 FILLER_25_1761 ();
 sg13g2_fill_2 FILLER_25_1766 ();
 sg13g2_fill_1 FILLER_25_1768 ();
 sg13g2_fill_1 FILLER_25_1773 ();
 sg13g2_fill_2 FILLER_25_1792 ();
 sg13g2_fill_1 FILLER_25_1794 ();
 sg13g2_fill_2 FILLER_25_1801 ();
 sg13g2_fill_1 FILLER_25_1803 ();
 sg13g2_fill_2 FILLER_25_1808 ();
 sg13g2_decap_8 FILLER_25_1815 ();
 sg13g2_fill_2 FILLER_25_1822 ();
 sg13g2_fill_1 FILLER_25_1842 ();
 sg13g2_fill_1 FILLER_25_1848 ();
 sg13g2_fill_1 FILLER_25_1875 ();
 sg13g2_decap_8 FILLER_25_1886 ();
 sg13g2_decap_8 FILLER_25_1893 ();
 sg13g2_decap_4 FILLER_25_1900 ();
 sg13g2_fill_2 FILLER_25_1904 ();
 sg13g2_fill_1 FILLER_25_1910 ();
 sg13g2_fill_2 FILLER_25_1937 ();
 sg13g2_fill_1 FILLER_25_1965 ();
 sg13g2_fill_2 FILLER_25_2044 ();
 sg13g2_fill_1 FILLER_25_2075 ();
 sg13g2_decap_8 FILLER_25_2097 ();
 sg13g2_decap_4 FILLER_25_2104 ();
 sg13g2_fill_2 FILLER_25_2126 ();
 sg13g2_fill_2 FILLER_25_2194 ();
 sg13g2_fill_1 FILLER_25_2196 ();
 sg13g2_fill_2 FILLER_25_2249 ();
 sg13g2_fill_1 FILLER_25_2251 ();
 sg13g2_decap_4 FILLER_25_2265 ();
 sg13g2_decap_8 FILLER_25_2299 ();
 sg13g2_fill_2 FILLER_25_2306 ();
 sg13g2_fill_1 FILLER_25_2308 ();
 sg13g2_decap_8 FILLER_25_2345 ();
 sg13g2_decap_4 FILLER_25_2352 ();
 sg13g2_fill_1 FILLER_25_2356 ();
 sg13g2_fill_1 FILLER_25_2361 ();
 sg13g2_fill_1 FILLER_25_2372 ();
 sg13g2_fill_2 FILLER_25_2387 ();
 sg13g2_fill_2 FILLER_25_2429 ();
 sg13g2_fill_1 FILLER_25_2431 ();
 sg13g2_fill_2 FILLER_25_2461 ();
 sg13g2_fill_1 FILLER_25_2505 ();
 sg13g2_fill_2 FILLER_25_2512 ();
 sg13g2_fill_2 FILLER_25_2523 ();
 sg13g2_fill_1 FILLER_25_2525 ();
 sg13g2_decap_4 FILLER_25_2537 ();
 sg13g2_fill_1 FILLER_25_2541 ();
 sg13g2_fill_2 FILLER_25_2557 ();
 sg13g2_fill_1 FILLER_25_2559 ();
 sg13g2_fill_1 FILLER_25_2568 ();
 sg13g2_fill_2 FILLER_25_2595 ();
 sg13g2_fill_2 FILLER_25_2601 ();
 sg13g2_fill_2 FILLER_25_2607 ();
 sg13g2_fill_1 FILLER_25_2631 ();
 sg13g2_decap_4 FILLER_25_2654 ();
 sg13g2_fill_2 FILLER_25_2658 ();
 sg13g2_decap_8 FILLER_25_2663 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_16 ();
 sg13g2_fill_2 FILLER_26_40 ();
 sg13g2_fill_1 FILLER_26_42 ();
 sg13g2_fill_1 FILLER_26_51 ();
 sg13g2_fill_1 FILLER_26_60 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_126 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_decap_4 FILLER_26_176 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_202 ();
 sg13g2_fill_2 FILLER_26_225 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_4 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_4 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_406 ();
 sg13g2_fill_2 FILLER_26_468 ();
 sg13g2_decap_4 FILLER_26_475 ();
 sg13g2_fill_1 FILLER_26_479 ();
 sg13g2_fill_1 FILLER_26_494 ();
 sg13g2_fill_1 FILLER_26_530 ();
 sg13g2_fill_1 FILLER_26_571 ();
 sg13g2_fill_2 FILLER_26_592 ();
 sg13g2_fill_1 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_608 ();
 sg13g2_fill_1 FILLER_26_615 ();
 sg13g2_decap_8 FILLER_26_661 ();
 sg13g2_fill_1 FILLER_26_668 ();
 sg13g2_decap_4 FILLER_26_698 ();
 sg13g2_fill_2 FILLER_26_702 ();
 sg13g2_fill_1 FILLER_26_780 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_fill_2 FILLER_26_852 ();
 sg13g2_fill_1 FILLER_26_854 ();
 sg13g2_fill_1 FILLER_26_914 ();
 sg13g2_fill_1 FILLER_26_941 ();
 sg13g2_fill_1 FILLER_26_946 ();
 sg13g2_fill_2 FILLER_26_977 ();
 sg13g2_fill_1 FILLER_26_979 ();
 sg13g2_fill_1 FILLER_26_1054 ();
 sg13g2_decap_8 FILLER_26_1059 ();
 sg13g2_fill_2 FILLER_26_1066 ();
 sg13g2_fill_2 FILLER_26_1094 ();
 sg13g2_decap_4 FILLER_26_1135 ();
 sg13g2_fill_2 FILLER_26_1149 ();
 sg13g2_fill_1 FILLER_26_1151 ();
 sg13g2_fill_1 FILLER_26_1193 ();
 sg13g2_fill_1 FILLER_26_1207 ();
 sg13g2_fill_1 FILLER_26_1218 ();
 sg13g2_fill_2 FILLER_26_1245 ();
 sg13g2_fill_1 FILLER_26_1250 ();
 sg13g2_decap_4 FILLER_26_1275 ();
 sg13g2_fill_2 FILLER_26_1279 ();
 sg13g2_fill_2 FILLER_26_1311 ();
 sg13g2_fill_1 FILLER_26_1313 ();
 sg13g2_fill_2 FILLER_26_1334 ();
 sg13g2_decap_8 FILLER_26_1362 ();
 sg13g2_decap_8 FILLER_26_1369 ();
 sg13g2_decap_4 FILLER_26_1398 ();
 sg13g2_fill_1 FILLER_26_1402 ();
 sg13g2_fill_1 FILLER_26_1431 ();
 sg13g2_fill_2 FILLER_26_1447 ();
 sg13g2_fill_2 FILLER_26_1466 ();
 sg13g2_fill_1 FILLER_26_1468 ();
 sg13g2_decap_8 FILLER_26_1495 ();
 sg13g2_fill_2 FILLER_26_1502 ();
 sg13g2_fill_1 FILLER_26_1504 ();
 sg13g2_fill_2 FILLER_26_1509 ();
 sg13g2_fill_1 FILLER_26_1511 ();
 sg13g2_decap_4 FILLER_26_1517 ();
 sg13g2_fill_2 FILLER_26_1521 ();
 sg13g2_decap_4 FILLER_26_1527 ();
 sg13g2_fill_1 FILLER_26_1566 ();
 sg13g2_decap_4 FILLER_26_1589 ();
 sg13g2_decap_4 FILLER_26_1614 ();
 sg13g2_fill_1 FILLER_26_1618 ();
 sg13g2_fill_2 FILLER_26_1669 ();
 sg13g2_decap_4 FILLER_26_1680 ();
 sg13g2_decap_4 FILLER_26_1694 ();
 sg13g2_fill_1 FILLER_26_1698 ();
 sg13g2_decap_8 FILLER_26_1716 ();
 sg13g2_fill_2 FILLER_26_1723 ();
 sg13g2_fill_2 FILLER_26_1733 ();
 sg13g2_fill_1 FILLER_26_1735 ();
 sg13g2_fill_1 FILLER_26_1740 ();
 sg13g2_decap_8 FILLER_26_1747 ();
 sg13g2_decap_8 FILLER_26_1754 ();
 sg13g2_decap_4 FILLER_26_1761 ();
 sg13g2_fill_2 FILLER_26_1778 ();
 sg13g2_fill_1 FILLER_26_1780 ();
 sg13g2_fill_2 FILLER_26_1787 ();
 sg13g2_fill_1 FILLER_26_1789 ();
 sg13g2_fill_2 FILLER_26_1800 ();
 sg13g2_decap_8 FILLER_26_1806 ();
 sg13g2_decap_8 FILLER_26_1813 ();
 sg13g2_fill_1 FILLER_26_1845 ();
 sg13g2_decap_4 FILLER_26_1872 ();
 sg13g2_fill_1 FILLER_26_1876 ();
 sg13g2_decap_4 FILLER_26_1887 ();
 sg13g2_fill_1 FILLER_26_1891 ();
 sg13g2_decap_4 FILLER_26_1902 ();
 sg13g2_fill_2 FILLER_26_1906 ();
 sg13g2_decap_8 FILLER_26_1914 ();
 sg13g2_fill_2 FILLER_26_1921 ();
 sg13g2_fill_2 FILLER_26_1935 ();
 sg13g2_fill_2 FILLER_26_1962 ();
 sg13g2_fill_2 FILLER_26_2049 ();
 sg13g2_fill_2 FILLER_26_2079 ();
 sg13g2_fill_1 FILLER_26_2081 ();
 sg13g2_decap_8 FILLER_26_2086 ();
 sg13g2_fill_2 FILLER_26_2093 ();
 sg13g2_fill_1 FILLER_26_2095 ();
 sg13g2_decap_8 FILLER_26_2122 ();
 sg13g2_decap_4 FILLER_26_2129 ();
 sg13g2_fill_2 FILLER_26_2133 ();
 sg13g2_decap_4 FILLER_26_2181 ();
 sg13g2_fill_2 FILLER_26_2215 ();
 sg13g2_decap_4 FILLER_26_2227 ();
 sg13g2_decap_8 FILLER_26_2235 ();
 sg13g2_decap_8 FILLER_26_2242 ();
 sg13g2_decap_8 FILLER_26_2253 ();
 sg13g2_decap_4 FILLER_26_2260 ();
 sg13g2_fill_2 FILLER_26_2264 ();
 sg13g2_decap_8 FILLER_26_2290 ();
 sg13g2_decap_8 FILLER_26_2297 ();
 sg13g2_decap_8 FILLER_26_2304 ();
 sg13g2_fill_2 FILLER_26_2311 ();
 sg13g2_fill_2 FILLER_26_2337 ();
 sg13g2_fill_1 FILLER_26_2339 ();
 sg13g2_decap_4 FILLER_26_2350 ();
 sg13g2_fill_2 FILLER_26_2354 ();
 sg13g2_decap_4 FILLER_26_2361 ();
 sg13g2_fill_1 FILLER_26_2365 ();
 sg13g2_decap_4 FILLER_26_2378 ();
 sg13g2_fill_1 FILLER_26_2382 ();
 sg13g2_fill_1 FILLER_26_2388 ();
 sg13g2_fill_2 FILLER_26_2406 ();
 sg13g2_fill_1 FILLER_26_2417 ();
 sg13g2_fill_1 FILLER_26_2428 ();
 sg13g2_decap_8 FILLER_26_2435 ();
 sg13g2_fill_1 FILLER_26_2442 ();
 sg13g2_fill_2 FILLER_26_2452 ();
 sg13g2_fill_2 FILLER_26_2480 ();
 sg13g2_fill_1 FILLER_26_2482 ();
 sg13g2_fill_2 FILLER_26_2509 ();
 sg13g2_decap_4 FILLER_26_2516 ();
 sg13g2_decap_8 FILLER_26_2530 ();
 sg13g2_decap_8 FILLER_26_2537 ();
 sg13g2_decap_4 FILLER_26_2584 ();
 sg13g2_fill_2 FILLER_26_2588 ();
 sg13g2_fill_1 FILLER_26_2626 ();
 sg13g2_fill_1 FILLER_26_2641 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_57 ();
 sg13g2_decap_8 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_91 ();
 sg13g2_fill_1 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_fill_2 FILLER_27_109 ();
 sg13g2_decap_4 FILLER_27_115 ();
 sg13g2_fill_1 FILLER_27_122 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_2 FILLER_27_142 ();
 sg13g2_fill_1 FILLER_27_144 ();
 sg13g2_decap_4 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_fill_2 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_4 FILLER_27_209 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_223 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_240 ();
 sg13g2_fill_2 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_decap_4 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_342 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_2 FILLER_27_416 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_fill_1 FILLER_27_447 ();
 sg13g2_decap_8 FILLER_27_479 ();
 sg13g2_decap_4 FILLER_27_486 ();
 sg13g2_fill_2 FILLER_27_533 ();
 sg13g2_fill_2 FILLER_27_557 ();
 sg13g2_fill_1 FILLER_27_572 ();
 sg13g2_fill_2 FILLER_27_577 ();
 sg13g2_fill_2 FILLER_27_587 ();
 sg13g2_fill_1 FILLER_27_615 ();
 sg13g2_fill_1 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_fill_2 FILLER_27_699 ();
 sg13g2_fill_1 FILLER_27_701 ();
 sg13g2_fill_2 FILLER_27_716 ();
 sg13g2_fill_1 FILLER_27_718 ();
 sg13g2_fill_2 FILLER_27_745 ();
 sg13g2_fill_1 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_771 ();
 sg13g2_decap_8 FILLER_27_778 ();
 sg13g2_fill_2 FILLER_27_785 ();
 sg13g2_fill_2 FILLER_27_796 ();
 sg13g2_fill_1 FILLER_27_798 ();
 sg13g2_fill_2 FILLER_27_809 ();
 sg13g2_fill_2 FILLER_27_821 ();
 sg13g2_fill_1 FILLER_27_823 ();
 sg13g2_decap_8 FILLER_27_850 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_fill_2 FILLER_27_895 ();
 sg13g2_fill_2 FILLER_27_946 ();
 sg13g2_decap_8 FILLER_27_969 ();
 sg13g2_decap_8 FILLER_27_976 ();
 sg13g2_decap_8 FILLER_27_983 ();
 sg13g2_decap_8 FILLER_27_990 ();
 sg13g2_decap_8 FILLER_27_997 ();
 sg13g2_decap_4 FILLER_27_1004 ();
 sg13g2_fill_2 FILLER_27_1008 ();
 sg13g2_fill_2 FILLER_27_1081 ();
 sg13g2_fill_1 FILLER_27_1083 ();
 sg13g2_decap_4 FILLER_27_1140 ();
 sg13g2_decap_8 FILLER_27_1165 ();
 sg13g2_fill_1 FILLER_27_1212 ();
 sg13g2_fill_1 FILLER_27_1249 ();
 sg13g2_fill_2 FILLER_27_1295 ();
 sg13g2_fill_1 FILLER_27_1297 ();
 sg13g2_decap_8 FILLER_27_1324 ();
 sg13g2_fill_2 FILLER_27_1331 ();
 sg13g2_decap_8 FILLER_27_1336 ();
 sg13g2_fill_1 FILLER_27_1343 ();
 sg13g2_fill_1 FILLER_27_1406 ();
 sg13g2_fill_2 FILLER_27_1423 ();
 sg13g2_decap_8 FILLER_27_1430 ();
 sg13g2_fill_2 FILLER_27_1442 ();
 sg13g2_decap_8 FILLER_27_1448 ();
 sg13g2_fill_2 FILLER_27_1455 ();
 sg13g2_fill_1 FILLER_27_1470 ();
 sg13g2_decap_4 FILLER_27_1488 ();
 sg13g2_fill_2 FILLER_27_1492 ();
 sg13g2_fill_1 FILLER_27_1513 ();
 sg13g2_fill_2 FILLER_27_1528 ();
 sg13g2_fill_1 FILLER_27_1535 ();
 sg13g2_fill_2 FILLER_27_1542 ();
 sg13g2_fill_2 FILLER_27_1549 ();
 sg13g2_fill_1 FILLER_27_1556 ();
 sg13g2_fill_2 FILLER_27_1569 ();
 sg13g2_fill_1 FILLER_27_1576 ();
 sg13g2_fill_1 FILLER_27_1584 ();
 sg13g2_fill_2 FILLER_27_1589 ();
 sg13g2_fill_1 FILLER_27_1591 ();
 sg13g2_decap_4 FILLER_27_1596 ();
 sg13g2_fill_1 FILLER_27_1692 ();
 sg13g2_decap_8 FILLER_27_1703 ();
 sg13g2_decap_8 FILLER_27_1710 ();
 sg13g2_fill_1 FILLER_27_1717 ();
 sg13g2_decap_4 FILLER_27_1744 ();
 sg13g2_fill_1 FILLER_27_1748 ();
 sg13g2_decap_4 FILLER_27_1760 ();
 sg13g2_decap_4 FILLER_27_1846 ();
 sg13g2_fill_2 FILLER_27_1855 ();
 sg13g2_decap_8 FILLER_27_1861 ();
 sg13g2_decap_8 FILLER_27_1868 ();
 sg13g2_decap_4 FILLER_27_1875 ();
 sg13g2_decap_4 FILLER_27_1884 ();
 sg13g2_fill_1 FILLER_27_1888 ();
 sg13g2_fill_1 FILLER_27_1904 ();
 sg13g2_fill_2 FILLER_27_1925 ();
 sg13g2_fill_1 FILLER_27_1927 ();
 sg13g2_fill_2 FILLER_27_1933 ();
 sg13g2_fill_2 FILLER_27_1961 ();
 sg13g2_fill_1 FILLER_27_1963 ();
 sg13g2_fill_1 FILLER_27_1969 ();
 sg13g2_decap_8 FILLER_27_1988 ();
 sg13g2_decap_4 FILLER_27_1995 ();
 sg13g2_fill_1 FILLER_27_1999 ();
 sg13g2_decap_8 FILLER_27_2004 ();
 sg13g2_decap_4 FILLER_27_2011 ();
 sg13g2_fill_2 FILLER_27_2015 ();
 sg13g2_fill_1 FILLER_27_2025 ();
 sg13g2_decap_8 FILLER_27_2043 ();
 sg13g2_fill_2 FILLER_27_2076 ();
 sg13g2_decap_4 FILLER_27_2104 ();
 sg13g2_decap_4 FILLER_27_2118 ();
 sg13g2_fill_1 FILLER_27_2122 ();
 sg13g2_fill_1 FILLER_27_2166 ();
 sg13g2_decap_8 FILLER_27_2175 ();
 sg13g2_fill_1 FILLER_27_2182 ();
 sg13g2_decap_8 FILLER_27_2223 ();
 sg13g2_decap_4 FILLER_27_2235 ();
 sg13g2_fill_2 FILLER_27_2239 ();
 sg13g2_fill_2 FILLER_27_2262 ();
 sg13g2_decap_8 FILLER_27_2285 ();
 sg13g2_decap_8 FILLER_27_2292 ();
 sg13g2_decap_4 FILLER_27_2299 ();
 sg13g2_fill_1 FILLER_27_2303 ();
 sg13g2_fill_2 FILLER_27_2330 ();
 sg13g2_fill_1 FILLER_27_2336 ();
 sg13g2_fill_1 FILLER_27_2343 ();
 sg13g2_fill_1 FILLER_27_2376 ();
 sg13g2_fill_2 FILLER_27_2383 ();
 sg13g2_decap_8 FILLER_27_2404 ();
 sg13g2_fill_2 FILLER_27_2411 ();
 sg13g2_decap_4 FILLER_27_2422 ();
 sg13g2_fill_2 FILLER_27_2426 ();
 sg13g2_decap_8 FILLER_27_2434 ();
 sg13g2_fill_1 FILLER_27_2451 ();
 sg13g2_fill_1 FILLER_27_2456 ();
 sg13g2_fill_1 FILLER_27_2465 ();
 sg13g2_fill_2 FILLER_27_2500 ();
 sg13g2_fill_1 FILLER_27_2502 ();
 sg13g2_decap_8 FILLER_27_2535 ();
 sg13g2_decap_4 FILLER_27_2542 ();
 sg13g2_fill_2 FILLER_27_2555 ();
 sg13g2_fill_2 FILLER_27_2571 ();
 sg13g2_fill_1 FILLER_27_2573 ();
 sg13g2_decap_8 FILLER_27_2580 ();
 sg13g2_fill_2 FILLER_27_2587 ();
 sg13g2_fill_1 FILLER_27_2601 ();
 sg13g2_fill_2 FILLER_27_2608 ();
 sg13g2_fill_1 FILLER_27_2610 ();
 sg13g2_fill_1 FILLER_27_2669 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_decap_4 FILLER_28_75 ();
 sg13g2_decap_4 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_113 ();
 sg13g2_fill_1 FILLER_28_117 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_decap_4 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_fill_1 FILLER_28_216 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_fill_2 FILLER_28_274 ();
 sg13g2_decap_8 FILLER_28_295 ();
 sg13g2_fill_2 FILLER_28_302 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_326 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_4 FILLER_28_352 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_decap_4 FILLER_28_361 ();
 sg13g2_fill_2 FILLER_28_365 ();
 sg13g2_decap_4 FILLER_28_403 ();
 sg13g2_decap_8 FILLER_28_416 ();
 sg13g2_decap_4 FILLER_28_423 ();
 sg13g2_fill_2 FILLER_28_427 ();
 sg13g2_fill_1 FILLER_28_473 ();
 sg13g2_fill_1 FILLER_28_484 ();
 sg13g2_fill_2 FILLER_28_504 ();
 sg13g2_fill_1 FILLER_28_506 ();
 sg13g2_fill_2 FILLER_28_515 ();
 sg13g2_fill_1 FILLER_28_517 ();
 sg13g2_fill_2 FILLER_28_523 ();
 sg13g2_fill_2 FILLER_28_544 ();
 sg13g2_decap_4 FILLER_28_554 ();
 sg13g2_fill_2 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_579 ();
 sg13g2_fill_2 FILLER_28_586 ();
 sg13g2_fill_1 FILLER_28_588 ();
 sg13g2_fill_1 FILLER_28_594 ();
 sg13g2_fill_2 FILLER_28_600 ();
 sg13g2_fill_2 FILLER_28_612 ();
 sg13g2_fill_1 FILLER_28_614 ();
 sg13g2_fill_1 FILLER_28_641 ();
 sg13g2_fill_1 FILLER_28_647 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_fill_2 FILLER_28_679 ();
 sg13g2_fill_1 FILLER_28_706 ();
 sg13g2_fill_2 FILLER_28_736 ();
 sg13g2_fill_1 FILLER_28_738 ();
 sg13g2_fill_2 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_774 ();
 sg13g2_decap_8 FILLER_28_781 ();
 sg13g2_decap_8 FILLER_28_788 ();
 sg13g2_decap_4 FILLER_28_795 ();
 sg13g2_fill_1 FILLER_28_829 ();
 sg13g2_decap_8 FILLER_28_837 ();
 sg13g2_decap_4 FILLER_28_844 ();
 sg13g2_fill_2 FILLER_28_848 ();
 sg13g2_fill_1 FILLER_28_905 ();
 sg13g2_fill_1 FILLER_28_919 ();
 sg13g2_decap_4 FILLER_28_960 ();
 sg13g2_fill_1 FILLER_28_964 ();
 sg13g2_fill_2 FILLER_28_969 ();
 sg13g2_decap_4 FILLER_28_997 ();
 sg13g2_decap_4 FILLER_28_1006 ();
 sg13g2_fill_1 FILLER_28_1010 ();
 sg13g2_decap_8 FILLER_28_1111 ();
 sg13g2_decap_4 FILLER_28_1118 ();
 sg13g2_decap_8 FILLER_28_1156 ();
 sg13g2_decap_8 FILLER_28_1163 ();
 sg13g2_fill_2 FILLER_28_1170 ();
 sg13g2_fill_1 FILLER_28_1172 ();
 sg13g2_fill_2 FILLER_28_1191 ();
 sg13g2_fill_1 FILLER_28_1193 ();
 sg13g2_fill_2 FILLER_28_1203 ();
 sg13g2_fill_1 FILLER_28_1205 ();
 sg13g2_decap_4 FILLER_28_1236 ();
 sg13g2_fill_2 FILLER_28_1240 ();
 sg13g2_decap_8 FILLER_28_1278 ();
 sg13g2_decap_4 FILLER_28_1285 ();
 sg13g2_fill_1 FILLER_28_1289 ();
 sg13g2_decap_8 FILLER_28_1294 ();
 sg13g2_decap_4 FILLER_28_1301 ();
 sg13g2_fill_2 FILLER_28_1305 ();
 sg13g2_decap_8 FILLER_28_1311 ();
 sg13g2_decap_8 FILLER_28_1318 ();
 sg13g2_decap_4 FILLER_28_1325 ();
 sg13g2_fill_1 FILLER_28_1329 ();
 sg13g2_fill_2 FILLER_28_1343 ();
 sg13g2_fill_1 FILLER_28_1345 ();
 sg13g2_decap_8 FILLER_28_1389 ();
 sg13g2_fill_2 FILLER_28_1417 ();
 sg13g2_decap_4 FILLER_28_1432 ();
 sg13g2_fill_2 FILLER_28_1436 ();
 sg13g2_decap_8 FILLER_28_1443 ();
 sg13g2_fill_2 FILLER_28_1468 ();
 sg13g2_fill_1 FILLER_28_1470 ();
 sg13g2_decap_8 FILLER_28_1476 ();
 sg13g2_fill_2 FILLER_28_1483 ();
 sg13g2_fill_1 FILLER_28_1489 ();
 sg13g2_fill_1 FILLER_28_1494 ();
 sg13g2_decap_8 FILLER_28_1507 ();
 sg13g2_decap_8 FILLER_28_1514 ();
 sg13g2_decap_4 FILLER_28_1521 ();
 sg13g2_fill_2 FILLER_28_1530 ();
 sg13g2_fill_1 FILLER_28_1594 ();
 sg13g2_fill_1 FILLER_28_1626 ();
 sg13g2_fill_2 FILLER_28_1637 ();
 sg13g2_fill_1 FILLER_28_1639 ();
 sg13g2_decap_8 FILLER_28_1692 ();
 sg13g2_decap_8 FILLER_28_1699 ();
 sg13g2_decap_8 FILLER_28_1706 ();
 sg13g2_fill_2 FILLER_28_1713 ();
 sg13g2_fill_1 FILLER_28_1715 ();
 sg13g2_fill_1 FILLER_28_1742 ();
 sg13g2_fill_2 FILLER_28_1757 ();
 sg13g2_fill_1 FILLER_28_1775 ();
 sg13g2_fill_2 FILLER_28_1780 ();
 sg13g2_fill_1 FILLER_28_1782 ();
 sg13g2_fill_1 FILLER_28_1813 ();
 sg13g2_fill_2 FILLER_28_1818 ();
 sg13g2_fill_1 FILLER_28_1820 ();
 sg13g2_fill_2 FILLER_28_1825 ();
 sg13g2_fill_1 FILLER_28_1902 ();
 sg13g2_fill_2 FILLER_28_1907 ();
 sg13g2_fill_1 FILLER_28_1909 ();
 sg13g2_decap_8 FILLER_28_1977 ();
 sg13g2_decap_8 FILLER_28_1984 ();
 sg13g2_decap_8 FILLER_28_1991 ();
 sg13g2_fill_2 FILLER_28_1998 ();
 sg13g2_decap_8 FILLER_28_2052 ();
 sg13g2_fill_2 FILLER_28_2059 ();
 sg13g2_fill_1 FILLER_28_2061 ();
 sg13g2_fill_2 FILLER_28_2066 ();
 sg13g2_fill_1 FILLER_28_2068 ();
 sg13g2_decap_4 FILLER_28_2126 ();
 sg13g2_fill_2 FILLER_28_2130 ();
 sg13g2_fill_1 FILLER_28_2136 ();
 sg13g2_fill_1 FILLER_28_2160 ();
 sg13g2_fill_1 FILLER_28_2187 ();
 sg13g2_decap_8 FILLER_28_2268 ();
 sg13g2_decap_8 FILLER_28_2275 ();
 sg13g2_decap_8 FILLER_28_2282 ();
 sg13g2_decap_8 FILLER_28_2289 ();
 sg13g2_decap_8 FILLER_28_2296 ();
 sg13g2_decap_8 FILLER_28_2303 ();
 sg13g2_fill_2 FILLER_28_2310 ();
 sg13g2_fill_1 FILLER_28_2342 ();
 sg13g2_fill_1 FILLER_28_2428 ();
 sg13g2_fill_1 FILLER_28_2491 ();
 sg13g2_fill_1 FILLER_28_2515 ();
 sg13g2_fill_2 FILLER_28_2526 ();
 sg13g2_fill_1 FILLER_28_2528 ();
 sg13g2_decap_4 FILLER_28_2535 ();
 sg13g2_fill_2 FILLER_28_2539 ();
 sg13g2_fill_2 FILLER_28_2581 ();
 sg13g2_decap_8 FILLER_28_2588 ();
 sg13g2_decap_8 FILLER_28_2595 ();
 sg13g2_decap_4 FILLER_28_2602 ();
 sg13g2_fill_1 FILLER_28_2606 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_4 FILLER_29_46 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_decap_8 FILLER_29_69 ();
 sg13g2_decap_8 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_decap_4 FILLER_29_101 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_110 ();
 sg13g2_decap_4 FILLER_29_115 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_decap_4 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_fill_1 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_fill_2 FILLER_29_374 ();
 sg13g2_decap_8 FILLER_29_451 ();
 sg13g2_decap_4 FILLER_29_458 ();
 sg13g2_fill_2 FILLER_29_495 ();
 sg13g2_fill_1 FILLER_29_497 ();
 sg13g2_fill_1 FILLER_29_518 ();
 sg13g2_fill_1 FILLER_29_523 ();
 sg13g2_decap_4 FILLER_29_550 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_fill_2 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_fill_2 FILLER_29_665 ();
 sg13g2_fill_1 FILLER_29_667 ();
 sg13g2_fill_1 FILLER_29_694 ();
 sg13g2_decap_4 FILLER_29_709 ();
 sg13g2_fill_1 FILLER_29_713 ();
 sg13g2_fill_1 FILLER_29_723 ();
 sg13g2_fill_2 FILLER_29_728 ();
 sg13g2_fill_2 FILLER_29_779 ();
 sg13g2_fill_1 FILLER_29_781 ();
 sg13g2_fill_1 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_843 ();
 sg13g2_fill_2 FILLER_29_850 ();
 sg13g2_fill_2 FILLER_29_862 ();
 sg13g2_fill_1 FILLER_29_932 ();
 sg13g2_fill_2 FILLER_29_940 ();
 sg13g2_fill_1 FILLER_29_942 ();
 sg13g2_fill_2 FILLER_29_947 ();
 sg13g2_fill_1 FILLER_29_949 ();
 sg13g2_fill_2 FILLER_29_976 ();
 sg13g2_decap_4 FILLER_29_982 ();
 sg13g2_fill_2 FILLER_29_986 ();
 sg13g2_decap_4 FILLER_29_1018 ();
 sg13g2_fill_1 FILLER_29_1022 ();
 sg13g2_decap_8 FILLER_29_1027 ();
 sg13g2_decap_4 FILLER_29_1034 ();
 sg13g2_fill_2 FILLER_29_1038 ();
 sg13g2_decap_8 FILLER_29_1074 ();
 sg13g2_fill_2 FILLER_29_1085 ();
 sg13g2_fill_1 FILLER_29_1087 ();
 sg13g2_decap_4 FILLER_29_1092 ();
 sg13g2_fill_2 FILLER_29_1096 ();
 sg13g2_fill_1 FILLER_29_1102 ();
 sg13g2_decap_8 FILLER_29_1107 ();
 sg13g2_decap_8 FILLER_29_1114 ();
 sg13g2_fill_1 FILLER_29_1121 ();
 sg13g2_fill_1 FILLER_29_1156 ();
 sg13g2_fill_1 FILLER_29_1165 ();
 sg13g2_fill_2 FILLER_29_1170 ();
 sg13g2_fill_2 FILLER_29_1177 ();
 sg13g2_fill_2 FILLER_29_1184 ();
 sg13g2_fill_1 FILLER_29_1186 ();
 sg13g2_fill_1 FILLER_29_1192 ();
 sg13g2_fill_2 FILLER_29_1198 ();
 sg13g2_fill_1 FILLER_29_1200 ();
 sg13g2_fill_1 FILLER_29_1205 ();
 sg13g2_decap_4 FILLER_29_1211 ();
 sg13g2_fill_1 FILLER_29_1215 ();
 sg13g2_fill_2 FILLER_29_1226 ();
 sg13g2_fill_1 FILLER_29_1228 ();
 sg13g2_fill_2 FILLER_29_1233 ();
 sg13g2_fill_1 FILLER_29_1235 ();
 sg13g2_fill_2 FILLER_29_1254 ();
 sg13g2_fill_1 FILLER_29_1256 ();
 sg13g2_decap_8 FILLER_29_1261 ();
 sg13g2_fill_1 FILLER_29_1268 ();
 sg13g2_fill_2 FILLER_29_1331 ();
 sg13g2_fill_1 FILLER_29_1333 ();
 sg13g2_fill_2 FILLER_29_1337 ();
 sg13g2_fill_1 FILLER_29_1339 ();
 sg13g2_decap_4 FILLER_29_1373 ();
 sg13g2_fill_2 FILLER_29_1403 ();
 sg13g2_fill_1 FILLER_29_1405 ();
 sg13g2_fill_1 FILLER_29_1421 ();
 sg13g2_fill_1 FILLER_29_1447 ();
 sg13g2_decap_4 FILLER_29_1452 ();
 sg13g2_fill_2 FILLER_29_1461 ();
 sg13g2_decap_4 FILLER_29_1477 ();
 sg13g2_fill_2 FILLER_29_1481 ();
 sg13g2_decap_4 FILLER_29_1488 ();
 sg13g2_fill_1 FILLER_29_1497 ();
 sg13g2_decap_4 FILLER_29_1517 ();
 sg13g2_fill_2 FILLER_29_1521 ();
 sg13g2_fill_2 FILLER_29_1527 ();
 sg13g2_fill_1 FILLER_29_1529 ();
 sg13g2_decap_4 FILLER_29_1539 ();
 sg13g2_fill_2 FILLER_29_1553 ();
 sg13g2_decap_4 FILLER_29_1565 ();
 sg13g2_decap_8 FILLER_29_1602 ();
 sg13g2_fill_2 FILLER_29_1622 ();
 sg13g2_fill_1 FILLER_29_1624 ();
 sg13g2_fill_1 FILLER_29_1655 ();
 sg13g2_decap_4 FILLER_29_1666 ();
 sg13g2_fill_1 FILLER_29_1670 ();
 sg13g2_decap_8 FILLER_29_1705 ();
 sg13g2_fill_1 FILLER_29_1712 ();
 sg13g2_fill_1 FILLER_29_1743 ();
 sg13g2_fill_1 FILLER_29_1780 ();
 sg13g2_fill_2 FILLER_29_1795 ();
 sg13g2_fill_1 FILLER_29_1797 ();
 sg13g2_fill_2 FILLER_29_1820 ();
 sg13g2_fill_1 FILLER_29_1822 ();
 sg13g2_fill_1 FILLER_29_1831 ();
 sg13g2_fill_1 FILLER_29_1873 ();
 sg13g2_decap_8 FILLER_29_1878 ();
 sg13g2_decap_8 FILLER_29_1885 ();
 sg13g2_fill_2 FILLER_29_1928 ();
 sg13g2_decap_8 FILLER_29_1966 ();
 sg13g2_fill_1 FILLER_29_1973 ();
 sg13g2_fill_1 FILLER_29_2093 ();
 sg13g2_decap_4 FILLER_29_2106 ();
 sg13g2_fill_2 FILLER_29_2115 ();
 sg13g2_decap_8 FILLER_29_2153 ();
 sg13g2_decap_8 FILLER_29_2160 ();
 sg13g2_fill_2 FILLER_29_2167 ();
 sg13g2_decap_8 FILLER_29_2173 ();
 sg13g2_decap_8 FILLER_29_2180 ();
 sg13g2_decap_4 FILLER_29_2187 ();
 sg13g2_decap_4 FILLER_29_2231 ();
 sg13g2_fill_1 FILLER_29_2235 ();
 sg13g2_fill_2 FILLER_29_2266 ();
 sg13g2_decap_4 FILLER_29_2304 ();
 sg13g2_decap_8 FILLER_29_2312 ();
 sg13g2_decap_4 FILLER_29_2329 ();
 sg13g2_fill_1 FILLER_29_2333 ();
 sg13g2_decap_4 FILLER_29_2349 ();
 sg13g2_fill_1 FILLER_29_2353 ();
 sg13g2_decap_4 FILLER_29_2414 ();
 sg13g2_fill_1 FILLER_29_2418 ();
 sg13g2_fill_2 FILLER_29_2429 ();
 sg13g2_fill_1 FILLER_29_2431 ();
 sg13g2_decap_4 FILLER_29_2445 ();
 sg13g2_fill_1 FILLER_29_2449 ();
 sg13g2_fill_2 FILLER_29_2460 ();
 sg13g2_fill_2 FILLER_29_2472 ();
 sg13g2_decap_8 FILLER_29_2478 ();
 sg13g2_fill_2 FILLER_29_2485 ();
 sg13g2_fill_1 FILLER_29_2596 ();
 sg13g2_fill_1 FILLER_29_2641 ();
 sg13g2_fill_2 FILLER_29_2668 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_decap_4 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_4 FILLER_30_147 ();
 sg13g2_fill_2 FILLER_30_151 ();
 sg13g2_fill_1 FILLER_30_174 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_268 ();
 sg13g2_decap_4 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_fill_2 FILLER_30_399 ();
 sg13g2_fill_1 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_decap_4 FILLER_30_411 ();
 sg13g2_decap_4 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_432 ();
 sg13g2_decap_4 FILLER_30_439 ();
 sg13g2_decap_8 FILLER_30_451 ();
 sg13g2_decap_8 FILLER_30_475 ();
 sg13g2_decap_8 FILLER_30_482 ();
 sg13g2_fill_2 FILLER_30_493 ();
 sg13g2_fill_1 FILLER_30_495 ();
 sg13g2_fill_2 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_fill_1 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_565 ();
 sg13g2_decap_8 FILLER_30_572 ();
 sg13g2_decap_8 FILLER_30_579 ();
 sg13g2_decap_4 FILLER_30_586 ();
 sg13g2_fill_2 FILLER_30_595 ();
 sg13g2_fill_1 FILLER_30_597 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_4 FILLER_30_616 ();
 sg13g2_fill_1 FILLER_30_624 ();
 sg13g2_decap_8 FILLER_30_659 ();
 sg13g2_decap_8 FILLER_30_666 ();
 sg13g2_fill_2 FILLER_30_673 ();
 sg13g2_fill_1 FILLER_30_675 ();
 sg13g2_fill_2 FILLER_30_685 ();
 sg13g2_fill_1 FILLER_30_687 ();
 sg13g2_fill_2 FILLER_30_692 ();
 sg13g2_fill_1 FILLER_30_694 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_fill_2 FILLER_30_716 ();
 sg13g2_decap_4 FILLER_30_740 ();
 sg13g2_fill_2 FILLER_30_744 ();
 sg13g2_fill_1 FILLER_30_750 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_4 FILLER_30_763 ();
 sg13g2_fill_1 FILLER_30_767 ();
 sg13g2_fill_2 FILLER_30_779 ();
 sg13g2_fill_1 FILLER_30_807 ();
 sg13g2_decap_4 FILLER_30_818 ();
 sg13g2_fill_2 FILLER_30_822 ();
 sg13g2_decap_8 FILLER_30_834 ();
 sg13g2_decap_4 FILLER_30_841 ();
 sg13g2_fill_1 FILLER_30_845 ();
 sg13g2_fill_1 FILLER_30_891 ();
 sg13g2_decap_8 FILLER_30_930 ();
 sg13g2_decap_4 FILLER_30_937 ();
 sg13g2_fill_1 FILLER_30_941 ();
 sg13g2_decap_4 FILLER_30_947 ();
 sg13g2_fill_1 FILLER_30_951 ();
 sg13g2_decap_4 FILLER_30_1003 ();
 sg13g2_decap_4 FILLER_30_1012 ();
 sg13g2_fill_2 FILLER_30_1042 ();
 sg13g2_fill_1 FILLER_30_1044 ();
 sg13g2_fill_2 FILLER_30_1076 ();
 sg13g2_fill_1 FILLER_30_1078 ();
 sg13g2_fill_1 FILLER_30_1089 ();
 sg13g2_fill_2 FILLER_30_1112 ();
 sg13g2_fill_1 FILLER_30_1114 ();
 sg13g2_decap_4 FILLER_30_1120 ();
 sg13g2_fill_1 FILLER_30_1124 ();
 sg13g2_fill_1 FILLER_30_1138 ();
 sg13g2_fill_2 FILLER_30_1188 ();
 sg13g2_fill_1 FILLER_30_1190 ();
 sg13g2_decap_4 FILLER_30_1195 ();
 sg13g2_decap_8 FILLER_30_1203 ();
 sg13g2_decap_4 FILLER_30_1210 ();
 sg13g2_fill_1 FILLER_30_1214 ();
 sg13g2_fill_2 FILLER_30_1246 ();
 sg13g2_fill_1 FILLER_30_1248 ();
 sg13g2_decap_8 FILLER_30_1279 ();
 sg13g2_fill_2 FILLER_30_1286 ();
 sg13g2_fill_1 FILLER_30_1288 ();
 sg13g2_fill_2 FILLER_30_1299 ();
 sg13g2_fill_1 FILLER_30_1301 ();
 sg13g2_decap_4 FILLER_30_1311 ();
 sg13g2_fill_2 FILLER_30_1315 ();
 sg13g2_fill_2 FILLER_30_1344 ();
 sg13g2_fill_1 FILLER_30_1346 ();
 sg13g2_decap_8 FILLER_30_1351 ();
 sg13g2_decap_8 FILLER_30_1358 ();
 sg13g2_fill_2 FILLER_30_1365 ();
 sg13g2_decap_4 FILLER_30_1380 ();
 sg13g2_fill_2 FILLER_30_1394 ();
 sg13g2_fill_1 FILLER_30_1400 ();
 sg13g2_fill_2 FILLER_30_1447 ();
 sg13g2_decap_8 FILLER_30_1459 ();
 sg13g2_decap_4 FILLER_30_1466 ();
 sg13g2_fill_2 FILLER_30_1470 ();
 sg13g2_decap_4 FILLER_30_1489 ();
 sg13g2_fill_2 FILLER_30_1493 ();
 sg13g2_decap_8 FILLER_30_1504 ();
 sg13g2_fill_2 FILLER_30_1511 ();
 sg13g2_fill_1 FILLER_30_1517 ();
 sg13g2_fill_2 FILLER_30_1542 ();
 sg13g2_fill_1 FILLER_30_1544 ();
 sg13g2_fill_2 FILLER_30_1550 ();
 sg13g2_fill_1 FILLER_30_1552 ();
 sg13g2_decap_4 FILLER_30_1572 ();
 sg13g2_fill_2 FILLER_30_1584 ();
 sg13g2_decap_8 FILLER_30_1591 ();
 sg13g2_fill_2 FILLER_30_1607 ();
 sg13g2_fill_1 FILLER_30_1609 ();
 sg13g2_fill_2 FILLER_30_1615 ();
 sg13g2_fill_1 FILLER_30_1617 ();
 sg13g2_decap_8 FILLER_30_1622 ();
 sg13g2_fill_2 FILLER_30_1629 ();
 sg13g2_fill_1 FILLER_30_1631 ();
 sg13g2_fill_2 FILLER_30_1650 ();
 sg13g2_decap_8 FILLER_30_1662 ();
 sg13g2_decap_8 FILLER_30_1669 ();
 sg13g2_decap_8 FILLER_30_1676 ();
 sg13g2_decap_8 FILLER_30_1683 ();
 sg13g2_decap_8 FILLER_30_1690 ();
 sg13g2_decap_8 FILLER_30_1697 ();
 sg13g2_decap_8 FILLER_30_1704 ();
 sg13g2_decap_8 FILLER_30_1711 ();
 sg13g2_decap_4 FILLER_30_1718 ();
 sg13g2_fill_2 FILLER_30_1722 ();
 sg13g2_decap_4 FILLER_30_1728 ();
 sg13g2_fill_1 FILLER_30_1732 ();
 sg13g2_fill_1 FILLER_30_1747 ();
 sg13g2_fill_1 FILLER_30_1786 ();
 sg13g2_fill_2 FILLER_30_1797 ();
 sg13g2_decap_8 FILLER_30_1814 ();
 sg13g2_fill_2 FILLER_30_1821 ();
 sg13g2_fill_1 FILLER_30_1823 ();
 sg13g2_decap_8 FILLER_30_1832 ();
 sg13g2_fill_2 FILLER_30_1839 ();
 sg13g2_fill_1 FILLER_30_1852 ();
 sg13g2_fill_2 FILLER_30_1857 ();
 sg13g2_fill_2 FILLER_30_1880 ();
 sg13g2_decap_8 FILLER_30_1887 ();
 sg13g2_fill_2 FILLER_30_1894 ();
 sg13g2_fill_1 FILLER_30_1896 ();
 sg13g2_decap_8 FILLER_30_1901 ();
 sg13g2_decap_4 FILLER_30_1908 ();
 sg13g2_fill_2 FILLER_30_1912 ();
 sg13g2_decap_8 FILLER_30_1946 ();
 sg13g2_fill_2 FILLER_30_1953 ();
 sg13g2_fill_1 FILLER_30_1955 ();
 sg13g2_fill_1 FILLER_30_1960 ();
 sg13g2_decap_8 FILLER_30_1997 ();
 sg13g2_fill_1 FILLER_30_2004 ();
 sg13g2_decap_4 FILLER_30_2009 ();
 sg13g2_fill_2 FILLER_30_2022 ();
 sg13g2_fill_1 FILLER_30_2024 ();
 sg13g2_decap_8 FILLER_30_2029 ();
 sg13g2_fill_1 FILLER_30_2036 ();
 sg13g2_fill_2 FILLER_30_2047 ();
 sg13g2_decap_8 FILLER_30_2070 ();
 sg13g2_decap_4 FILLER_30_2077 ();
 sg13g2_fill_1 FILLER_30_2091 ();
 sg13g2_fill_1 FILLER_30_2100 ();
 sg13g2_decap_8 FILLER_30_2111 ();
 sg13g2_decap_8 FILLER_30_2118 ();
 sg13g2_decap_8 FILLER_30_2125 ();
 sg13g2_fill_2 FILLER_30_2132 ();
 sg13g2_fill_1 FILLER_30_2134 ();
 sg13g2_decap_8 FILLER_30_2171 ();
 sg13g2_decap_4 FILLER_30_2178 ();
 sg13g2_fill_1 FILLER_30_2182 ();
 sg13g2_fill_1 FILLER_30_2193 ();
 sg13g2_fill_2 FILLER_30_2260 ();
 sg13g2_decap_8 FILLER_30_2283 ();
 sg13g2_decap_8 FILLER_30_2290 ();
 sg13g2_decap_4 FILLER_30_2297 ();
 sg13g2_fill_1 FILLER_30_2301 ();
 sg13g2_fill_1 FILLER_30_2332 ();
 sg13g2_fill_2 FILLER_30_2337 ();
 sg13g2_decap_8 FILLER_30_2344 ();
 sg13g2_fill_1 FILLER_30_2351 ();
 sg13g2_decap_4 FILLER_30_2362 ();
 sg13g2_fill_1 FILLER_30_2366 ();
 sg13g2_decap_4 FILLER_30_2371 ();
 sg13g2_fill_1 FILLER_30_2375 ();
 sg13g2_decap_8 FILLER_30_2386 ();
 sg13g2_decap_8 FILLER_30_2407 ();
 sg13g2_decap_8 FILLER_30_2450 ();
 sg13g2_decap_8 FILLER_30_2457 ();
 sg13g2_fill_2 FILLER_30_2464 ();
 sg13g2_fill_2 FILLER_30_2491 ();
 sg13g2_decap_8 FILLER_30_2497 ();
 sg13g2_fill_2 FILLER_30_2504 ();
 sg13g2_fill_1 FILLER_30_2506 ();
 sg13g2_decap_8 FILLER_30_2515 ();
 sg13g2_fill_2 FILLER_30_2522 ();
 sg13g2_fill_1 FILLER_30_2524 ();
 sg13g2_decap_8 FILLER_30_2529 ();
 sg13g2_fill_2 FILLER_30_2536 ();
 sg13g2_fill_1 FILLER_30_2538 ();
 sg13g2_fill_1 FILLER_30_2553 ();
 sg13g2_fill_2 FILLER_30_2558 ();
 sg13g2_fill_1 FILLER_30_2560 ();
 sg13g2_decap_4 FILLER_30_2581 ();
 sg13g2_fill_1 FILLER_30_2595 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_15 ();
 sg13g2_decap_4 FILLER_31_22 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_fill_2 FILLER_31_33 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_86 ();
 sg13g2_decap_8 FILLER_31_117 ();
 sg13g2_decap_4 FILLER_31_124 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_fill_1 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_237 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_276 ();
 sg13g2_decap_4 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_293 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_decap_4 FILLER_31_331 ();
 sg13g2_decap_4 FILLER_31_398 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_fill_2 FILLER_31_426 ();
 sg13g2_fill_1 FILLER_31_428 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_fill_1 FILLER_31_441 ();
 sg13g2_fill_1 FILLER_31_503 ();
 sg13g2_fill_2 FILLER_31_555 ();
 sg13g2_fill_1 FILLER_31_557 ();
 sg13g2_fill_1 FILLER_31_571 ();
 sg13g2_fill_2 FILLER_31_582 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_fill_2 FILLER_31_609 ();
 sg13g2_fill_1 FILLER_31_611 ();
 sg13g2_decap_4 FILLER_31_621 ();
 sg13g2_fill_1 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_630 ();
 sg13g2_fill_2 FILLER_31_645 ();
 sg13g2_decap_8 FILLER_31_664 ();
 sg13g2_decap_8 FILLER_31_671 ();
 sg13g2_decap_8 FILLER_31_678 ();
 sg13g2_decap_8 FILLER_31_685 ();
 sg13g2_decap_8 FILLER_31_692 ();
 sg13g2_decap_4 FILLER_31_699 ();
 sg13g2_fill_2 FILLER_31_703 ();
 sg13g2_fill_1 FILLER_31_737 ();
 sg13g2_fill_2 FILLER_31_757 ();
 sg13g2_fill_1 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_fill_2 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_839 ();
 sg13g2_fill_1 FILLER_31_846 ();
 sg13g2_fill_2 FILLER_31_900 ();
 sg13g2_decap_8 FILLER_31_929 ();
 sg13g2_decap_8 FILLER_31_936 ();
 sg13g2_fill_2 FILLER_31_943 ();
 sg13g2_fill_1 FILLER_31_945 ();
 sg13g2_fill_2 FILLER_31_959 ();
 sg13g2_fill_1 FILLER_31_965 ();
 sg13g2_fill_2 FILLER_31_971 ();
 sg13g2_fill_2 FILLER_31_977 ();
 sg13g2_fill_1 FILLER_31_979 ();
 sg13g2_decap_4 FILLER_31_985 ();
 sg13g2_decap_8 FILLER_31_998 ();
 sg13g2_fill_2 FILLER_31_1005 ();
 sg13g2_decap_4 FILLER_31_1012 ();
 sg13g2_fill_1 FILLER_31_1046 ();
 sg13g2_fill_1 FILLER_31_1051 ();
 sg13g2_fill_1 FILLER_31_1056 ();
 sg13g2_fill_2 FILLER_31_1083 ();
 sg13g2_fill_1 FILLER_31_1085 ();
 sg13g2_fill_2 FILLER_31_1112 ();
 sg13g2_fill_1 FILLER_31_1114 ();
 sg13g2_decap_8 FILLER_31_1119 ();
 sg13g2_fill_2 FILLER_31_1126 ();
 sg13g2_fill_2 FILLER_31_1164 ();
 sg13g2_fill_2 FILLER_31_1170 ();
 sg13g2_fill_1 FILLER_31_1193 ();
 sg13g2_decap_4 FILLER_31_1198 ();
 sg13g2_fill_2 FILLER_31_1202 ();
 sg13g2_decap_4 FILLER_31_1243 ();
 sg13g2_fill_2 FILLER_31_1251 ();
 sg13g2_fill_1 FILLER_31_1253 ();
 sg13g2_decap_8 FILLER_31_1280 ();
 sg13g2_fill_2 FILLER_31_1287 ();
 sg13g2_decap_8 FILLER_31_1293 ();
 sg13g2_fill_2 FILLER_31_1300 ();
 sg13g2_fill_1 FILLER_31_1302 ();
 sg13g2_decap_8 FILLER_31_1337 ();
 sg13g2_fill_1 FILLER_31_1344 ();
 sg13g2_fill_2 FILLER_31_1349 ();
 sg13g2_fill_1 FILLER_31_1377 ();
 sg13g2_fill_2 FILLER_31_1412 ();
 sg13g2_fill_1 FILLER_31_1451 ();
 sg13g2_fill_1 FILLER_31_1492 ();
 sg13g2_fill_2 FILLER_31_1511 ();
 sg13g2_fill_1 FILLER_31_1546 ();
 sg13g2_fill_1 FILLER_31_1558 ();
 sg13g2_fill_1 FILLER_31_1565 ();
 sg13g2_decap_8 FILLER_31_1570 ();
 sg13g2_decap_8 FILLER_31_1577 ();
 sg13g2_decap_8 FILLER_31_1584 ();
 sg13g2_decap_8 FILLER_31_1591 ();
 sg13g2_decap_8 FILLER_31_1598 ();
 sg13g2_fill_1 FILLER_31_1605 ();
 sg13g2_fill_2 FILLER_31_1611 ();
 sg13g2_fill_2 FILLER_31_1618 ();
 sg13g2_fill_2 FILLER_31_1625 ();
 sg13g2_fill_1 FILLER_31_1627 ();
 sg13g2_decap_4 FILLER_31_1654 ();
 sg13g2_fill_2 FILLER_31_1658 ();
 sg13g2_fill_2 FILLER_31_1670 ();
 sg13g2_decap_8 FILLER_31_1686 ();
 sg13g2_fill_2 FILLER_31_1693 ();
 sg13g2_fill_1 FILLER_31_1695 ();
 sg13g2_decap_4 FILLER_31_1699 ();
 sg13g2_fill_1 FILLER_31_1703 ();
 sg13g2_decap_8 FILLER_31_1712 ();
 sg13g2_decap_8 FILLER_31_1719 ();
 sg13g2_fill_2 FILLER_31_1726 ();
 sg13g2_fill_1 FILLER_31_1728 ();
 sg13g2_fill_2 FILLER_31_1752 ();
 sg13g2_decap_4 FILLER_31_1764 ();
 sg13g2_decap_4 FILLER_31_1778 ();
 sg13g2_fill_1 FILLER_31_1782 ();
 sg13g2_fill_2 FILLER_31_1787 ();
 sg13g2_fill_2 FILLER_31_1795 ();
 sg13g2_fill_2 FILLER_31_1803 ();
 sg13g2_fill_2 FILLER_31_1831 ();
 sg13g2_decap_4 FILLER_31_1837 ();
 sg13g2_fill_1 FILLER_31_1875 ();
 sg13g2_decap_4 FILLER_31_1889 ();
 sg13g2_fill_1 FILLER_31_1893 ();
 sg13g2_fill_2 FILLER_31_1903 ();
 sg13g2_fill_1 FILLER_31_1924 ();
 sg13g2_fill_2 FILLER_31_1935 ();
 sg13g2_fill_2 FILLER_31_1941 ();
 sg13g2_fill_2 FILLER_31_1974 ();
 sg13g2_fill_1 FILLER_31_1976 ();
 sg13g2_decap_8 FILLER_31_1985 ();
 sg13g2_decap_8 FILLER_31_1992 ();
 sg13g2_decap_8 FILLER_31_1999 ();
 sg13g2_decap_8 FILLER_31_2006 ();
 sg13g2_decap_8 FILLER_31_2018 ();
 sg13g2_fill_2 FILLER_31_2025 ();
 sg13g2_fill_1 FILLER_31_2027 ();
 sg13g2_fill_2 FILLER_31_2048 ();
 sg13g2_fill_2 FILLER_31_2123 ();
 sg13g2_fill_1 FILLER_31_2125 ();
 sg13g2_fill_1 FILLER_31_2160 ();
 sg13g2_decap_8 FILLER_31_2182 ();
 sg13g2_fill_2 FILLER_31_2189 ();
 sg13g2_fill_1 FILLER_31_2191 ();
 sg13g2_fill_2 FILLER_31_2196 ();
 sg13g2_fill_1 FILLER_31_2198 ();
 sg13g2_decap_8 FILLER_31_2220 ();
 sg13g2_decap_4 FILLER_31_2227 ();
 sg13g2_fill_1 FILLER_31_2231 ();
 sg13g2_decap_8 FILLER_31_2246 ();
 sg13g2_fill_2 FILLER_31_2253 ();
 sg13g2_decap_4 FILLER_31_2260 ();
 sg13g2_fill_2 FILLER_31_2264 ();
 sg13g2_decap_8 FILLER_31_2310 ();
 sg13g2_decap_8 FILLER_31_2317 ();
 sg13g2_decap_8 FILLER_31_2324 ();
 sg13g2_decap_4 FILLER_31_2331 ();
 sg13g2_decap_4 FILLER_31_2338 ();
 sg13g2_fill_1 FILLER_31_2342 ();
 sg13g2_decap_4 FILLER_31_2346 ();
 sg13g2_fill_2 FILLER_31_2350 ();
 sg13g2_decap_8 FILLER_31_2356 ();
 sg13g2_decap_8 FILLER_31_2363 ();
 sg13g2_decap_8 FILLER_31_2370 ();
 sg13g2_decap_4 FILLER_31_2377 ();
 sg13g2_fill_2 FILLER_31_2385 ();
 sg13g2_fill_1 FILLER_31_2387 ();
 sg13g2_decap_4 FILLER_31_2392 ();
 sg13g2_fill_1 FILLER_31_2422 ();
 sg13g2_fill_1 FILLER_31_2448 ();
 sg13g2_decap_8 FILLER_31_2454 ();
 sg13g2_decap_4 FILLER_31_2461 ();
 sg13g2_fill_2 FILLER_31_2469 ();
 sg13g2_decap_4 FILLER_31_2497 ();
 sg13g2_fill_1 FILLER_31_2505 ();
 sg13g2_fill_1 FILLER_31_2511 ();
 sg13g2_decap_8 FILLER_31_2516 ();
 sg13g2_decap_8 FILLER_31_2523 ();
 sg13g2_decap_8 FILLER_31_2530 ();
 sg13g2_decap_8 FILLER_31_2537 ();
 sg13g2_decap_8 FILLER_31_2544 ();
 sg13g2_decap_8 FILLER_31_2551 ();
 sg13g2_decap_8 FILLER_31_2558 ();
 sg13g2_decap_4 FILLER_31_2565 ();
 sg13g2_fill_1 FILLER_31_2569 ();
 sg13g2_fill_1 FILLER_31_2575 ();
 sg13g2_fill_1 FILLER_31_2642 ();
 sg13g2_decap_4 FILLER_31_2657 ();
 sg13g2_fill_2 FILLER_31_2661 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_2 FILLER_32_61 ();
 sg13g2_fill_2 FILLER_32_71 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_4 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_fill_2 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_4 FILLER_32_322 ();
 sg13g2_fill_1 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_fill_2 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_367 ();
 sg13g2_decap_4 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_397 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_fill_1 FILLER_32_414 ();
 sg13g2_fill_2 FILLER_32_462 ();
 sg13g2_fill_1 FILLER_32_464 ();
 sg13g2_fill_1 FILLER_32_474 ();
 sg13g2_fill_2 FILLER_32_520 ();
 sg13g2_fill_1 FILLER_32_525 ();
 sg13g2_fill_1 FILLER_32_542 ();
 sg13g2_fill_1 FILLER_32_579 ();
 sg13g2_fill_1 FILLER_32_585 ();
 sg13g2_fill_1 FILLER_32_631 ();
 sg13g2_fill_2 FILLER_32_636 ();
 sg13g2_fill_2 FILLER_32_648 ();
 sg13g2_decap_8 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_683 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_696 ();
 sg13g2_fill_1 FILLER_32_703 ();
 sg13g2_decap_4 FILLER_32_718 ();
 sg13g2_fill_2 FILLER_32_722 ();
 sg13g2_fill_2 FILLER_32_734 ();
 sg13g2_fill_1 FILLER_32_736 ();
 sg13g2_fill_1 FILLER_32_742 ();
 sg13g2_fill_2 FILLER_32_751 ();
 sg13g2_decap_8 FILLER_32_779 ();
 sg13g2_decap_4 FILLER_32_786 ();
 sg13g2_fill_1 FILLER_32_790 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_4 FILLER_32_812 ();
 sg13g2_fill_2 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_825 ();
 sg13g2_decap_8 FILLER_32_832 ();
 sg13g2_decap_8 FILLER_32_839 ();
 sg13g2_decap_8 FILLER_32_846 ();
 sg13g2_decap_4 FILLER_32_853 ();
 sg13g2_decap_4 FILLER_32_861 ();
 sg13g2_fill_2 FILLER_32_901 ();
 sg13g2_fill_1 FILLER_32_929 ();
 sg13g2_fill_1 FILLER_32_956 ();
 sg13g2_fill_1 FILLER_32_983 ();
 sg13g2_decap_4 FILLER_32_988 ();
 sg13g2_fill_2 FILLER_32_992 ();
 sg13g2_decap_4 FILLER_32_1024 ();
 sg13g2_decap_8 FILLER_32_1032 ();
 sg13g2_decap_4 FILLER_32_1039 ();
 sg13g2_fill_1 FILLER_32_1043 ();
 sg13g2_decap_4 FILLER_32_1053 ();
 sg13g2_decap_8 FILLER_32_1061 ();
 sg13g2_fill_1 FILLER_32_1068 ();
 sg13g2_fill_1 FILLER_32_1074 ();
 sg13g2_decap_4 FILLER_32_1118 ();
 sg13g2_fill_1 FILLER_32_1122 ();
 sg13g2_decap_4 FILLER_32_1163 ();
 sg13g2_decap_4 FILLER_32_1203 ();
 sg13g2_decap_8 FILLER_32_1238 ();
 sg13g2_decap_4 FILLER_32_1245 ();
 sg13g2_fill_2 FILLER_32_1259 ();
 sg13g2_fill_1 FILLER_32_1265 ();
 sg13g2_fill_2 FILLER_32_1270 ();
 sg13g2_fill_2 FILLER_32_1298 ();
 sg13g2_fill_1 FILLER_32_1300 ();
 sg13g2_fill_2 FILLER_32_1327 ();
 sg13g2_fill_1 FILLER_32_1329 ();
 sg13g2_decap_4 FILLER_32_1356 ();
 sg13g2_decap_8 FILLER_32_1364 ();
 sg13g2_fill_1 FILLER_32_1371 ();
 sg13g2_decap_4 FILLER_32_1417 ();
 sg13g2_fill_1 FILLER_32_1421 ();
 sg13g2_fill_1 FILLER_32_1432 ();
 sg13g2_decap_8 FILLER_32_1438 ();
 sg13g2_decap_4 FILLER_32_1445 ();
 sg13g2_fill_2 FILLER_32_1449 ();
 sg13g2_decap_4 FILLER_32_1462 ();
 sg13g2_fill_2 FILLER_32_1493 ();
 sg13g2_fill_1 FILLER_32_1495 ();
 sg13g2_fill_2 FILLER_32_1518 ();
 sg13g2_fill_1 FILLER_32_1520 ();
 sg13g2_fill_1 FILLER_32_1526 ();
 sg13g2_fill_1 FILLER_32_1535 ();
 sg13g2_fill_1 FILLER_32_1542 ();
 sg13g2_decap_8 FILLER_32_1567 ();
 sg13g2_decap_4 FILLER_32_1574 ();
 sg13g2_fill_2 FILLER_32_1578 ();
 sg13g2_decap_4 FILLER_32_1584 ();
 sg13g2_decap_4 FILLER_32_1596 ();
 sg13g2_fill_1 FILLER_32_1708 ();
 sg13g2_decap_8 FILLER_32_1722 ();
 sg13g2_decap_8 FILLER_32_1729 ();
 sg13g2_decap_4 FILLER_32_1736 ();
 sg13g2_fill_2 FILLER_32_1766 ();
 sg13g2_fill_1 FILLER_32_1768 ();
 sg13g2_fill_1 FILLER_32_1795 ();
 sg13g2_fill_1 FILLER_32_1806 ();
 sg13g2_fill_1 FILLER_32_1833 ();
 sg13g2_decap_8 FILLER_32_1865 ();
 sg13g2_decap_8 FILLER_32_1872 ();
 sg13g2_decap_8 FILLER_32_1879 ();
 sg13g2_decap_8 FILLER_32_1886 ();
 sg13g2_decap_8 FILLER_32_1893 ();
 sg13g2_decap_8 FILLER_32_1900 ();
 sg13g2_decap_8 FILLER_32_1907 ();
 sg13g2_decap_8 FILLER_32_1914 ();
 sg13g2_fill_2 FILLER_32_1931 ();
 sg13g2_fill_1 FILLER_32_1933 ();
 sg13g2_decap_4 FILLER_32_1944 ();
 sg13g2_decap_8 FILLER_32_1952 ();
 sg13g2_decap_8 FILLER_32_1959 ();
 sg13g2_decap_8 FILLER_32_1966 ();
 sg13g2_decap_8 FILLER_32_1973 ();
 sg13g2_decap_4 FILLER_32_1980 ();
 sg13g2_fill_2 FILLER_32_1984 ();
 sg13g2_decap_4 FILLER_32_2006 ();
 sg13g2_fill_1 FILLER_32_2030 ();
 sg13g2_fill_2 FILLER_32_2035 ();
 sg13g2_decap_8 FILLER_32_2049 ();
 sg13g2_decap_8 FILLER_32_2056 ();
 sg13g2_fill_2 FILLER_32_2063 ();
 sg13g2_decap_4 FILLER_32_2078 ();
 sg13g2_fill_1 FILLER_32_2082 ();
 sg13g2_fill_1 FILLER_32_2095 ();
 sg13g2_fill_2 FILLER_32_2178 ();
 sg13g2_fill_2 FILLER_32_2206 ();
 sg13g2_fill_1 FILLER_32_2208 ();
 sg13g2_decap_8 FILLER_32_2235 ();
 sg13g2_decap_8 FILLER_32_2242 ();
 sg13g2_fill_1 FILLER_32_2249 ();
 sg13g2_decap_4 FILLER_32_2286 ();
 sg13g2_decap_8 FILLER_32_2294 ();
 sg13g2_decap_4 FILLER_32_2301 ();
 sg13g2_fill_2 FILLER_32_2305 ();
 sg13g2_fill_1 FILLER_32_2380 ();
 sg13g2_fill_1 FILLER_32_2385 ();
 sg13g2_fill_2 FILLER_32_2400 ();
 sg13g2_fill_1 FILLER_32_2410 ();
 sg13g2_fill_2 FILLER_32_2430 ();
 sg13g2_fill_1 FILLER_32_2432 ();
 sg13g2_fill_2 FILLER_32_2438 ();
 sg13g2_fill_1 FILLER_32_2440 ();
 sg13g2_fill_1 FILLER_32_2447 ();
 sg13g2_fill_2 FILLER_32_2452 ();
 sg13g2_fill_1 FILLER_32_2454 ();
 sg13g2_fill_2 FILLER_32_2497 ();
 sg13g2_decap_8 FILLER_32_2547 ();
 sg13g2_decap_4 FILLER_32_2554 ();
 sg13g2_fill_1 FILLER_32_2562 ();
 sg13g2_fill_2 FILLER_32_2583 ();
 sg13g2_fill_1 FILLER_32_2595 ();
 sg13g2_fill_2 FILLER_32_2606 ();
 sg13g2_fill_2 FILLER_32_2621 ();
 sg13g2_decap_8 FILLER_32_2653 ();
 sg13g2_decap_8 FILLER_32_2660 ();
 sg13g2_fill_2 FILLER_32_2667 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_decap_4 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_2 FILLER_33_63 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_decap_4 FILLER_33_196 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_205 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_223 ();
 sg13g2_decap_8 FILLER_33_228 ();
 sg13g2_decap_8 FILLER_33_239 ();
 sg13g2_decap_4 FILLER_33_246 ();
 sg13g2_fill_2 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_297 ();
 sg13g2_decap_4 FILLER_33_303 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_decap_4 FILLER_33_390 ();
 sg13g2_decap_4 FILLER_33_420 ();
 sg13g2_fill_1 FILLER_33_438 ();
 sg13g2_fill_2 FILLER_33_443 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_fill_2 FILLER_33_462 ();
 sg13g2_fill_1 FILLER_33_464 ();
 sg13g2_fill_2 FILLER_33_474 ();
 sg13g2_fill_2 FILLER_33_502 ();
 sg13g2_fill_1 FILLER_33_513 ();
 sg13g2_fill_2 FILLER_33_548 ();
 sg13g2_fill_1 FILLER_33_615 ();
 sg13g2_fill_1 FILLER_33_650 ();
 sg13g2_fill_1 FILLER_33_660 ();
 sg13g2_decap_4 FILLER_33_666 ();
 sg13g2_fill_1 FILLER_33_670 ();
 sg13g2_fill_1 FILLER_33_731 ();
 sg13g2_fill_1 FILLER_33_737 ();
 sg13g2_fill_1 FILLER_33_747 ();
 sg13g2_fill_1 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_788 ();
 sg13g2_decap_8 FILLER_33_795 ();
 sg13g2_decap_8 FILLER_33_802 ();
 sg13g2_decap_8 FILLER_33_809 ();
 sg13g2_decap_8 FILLER_33_816 ();
 sg13g2_decap_8 FILLER_33_823 ();
 sg13g2_decap_8 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_837 ();
 sg13g2_decap_4 FILLER_33_844 ();
 sg13g2_fill_1 FILLER_33_848 ();
 sg13g2_fill_1 FILLER_33_885 ();
 sg13g2_fill_2 FILLER_33_912 ();
 sg13g2_fill_1 FILLER_33_918 ();
 sg13g2_fill_1 FILLER_33_924 ();
 sg13g2_fill_2 FILLER_33_951 ();
 sg13g2_fill_2 FILLER_33_958 ();
 sg13g2_fill_1 FILLER_33_965 ();
 sg13g2_fill_2 FILLER_33_970 ();
 sg13g2_fill_2 FILLER_33_998 ();
 sg13g2_fill_2 FILLER_33_1004 ();
 sg13g2_fill_1 FILLER_33_1006 ();
 sg13g2_decap_4 FILLER_33_1012 ();
 sg13g2_decap_8 FILLER_33_1020 ();
 sg13g2_decap_8 FILLER_33_1027 ();
 sg13g2_decap_8 FILLER_33_1034 ();
 sg13g2_decap_8 FILLER_33_1041 ();
 sg13g2_decap_8 FILLER_33_1048 ();
 sg13g2_fill_2 FILLER_33_1055 ();
 sg13g2_fill_1 FILLER_33_1057 ();
 sg13g2_decap_4 FILLER_33_1084 ();
 sg13g2_fill_2 FILLER_33_1088 ();
 sg13g2_fill_1 FILLER_33_1116 ();
 sg13g2_fill_2 FILLER_33_1121 ();
 sg13g2_decap_4 FILLER_33_1152 ();
 sg13g2_fill_2 FILLER_33_1156 ();
 sg13g2_fill_2 FILLER_33_1168 ();
 sg13g2_fill_2 FILLER_33_1174 ();
 sg13g2_decap_4 FILLER_33_1180 ();
 sg13g2_fill_2 FILLER_33_1184 ();
 sg13g2_decap_4 FILLER_33_1190 ();
 sg13g2_decap_4 FILLER_33_1211 ();
 sg13g2_fill_2 FILLER_33_1215 ();
 sg13g2_decap_4 FILLER_33_1227 ();
 sg13g2_decap_4 FILLER_33_1262 ();
 sg13g2_fill_2 FILLER_33_1270 ();
 sg13g2_fill_1 FILLER_33_1286 ();
 sg13g2_fill_2 FILLER_33_1297 ();
 sg13g2_fill_2 FILLER_33_1309 ();
 sg13g2_fill_1 FILLER_33_1311 ();
 sg13g2_fill_1 FILLER_33_1322 ();
 sg13g2_fill_2 FILLER_33_1333 ();
 sg13g2_fill_1 FILLER_33_1335 ();
 sg13g2_decap_8 FILLER_33_1340 ();
 sg13g2_decap_8 FILLER_33_1347 ();
 sg13g2_decap_4 FILLER_33_1373 ();
 sg13g2_fill_2 FILLER_33_1396 ();
 sg13g2_fill_1 FILLER_33_1410 ();
 sg13g2_decap_4 FILLER_33_1424 ();
 sg13g2_decap_8 FILLER_33_1439 ();
 sg13g2_decap_8 FILLER_33_1446 ();
 sg13g2_decap_4 FILLER_33_1453 ();
 sg13g2_fill_2 FILLER_33_1457 ();
 sg13g2_decap_4 FILLER_33_1464 ();
 sg13g2_fill_1 FILLER_33_1468 ();
 sg13g2_fill_2 FILLER_33_1494 ();
 sg13g2_fill_1 FILLER_33_1496 ();
 sg13g2_decap_8 FILLER_33_1506 ();
 sg13g2_fill_1 FILLER_33_1528 ();
 sg13g2_fill_2 FILLER_33_1534 ();
 sg13g2_decap_4 FILLER_33_1562 ();
 sg13g2_fill_1 FILLER_33_1566 ();
 sg13g2_fill_1 FILLER_33_1606 ();
 sg13g2_fill_2 FILLER_33_1612 ();
 sg13g2_decap_8 FILLER_33_1624 ();
 sg13g2_fill_1 FILLER_33_1631 ();
 sg13g2_decap_8 FILLER_33_1668 ();
 sg13g2_fill_1 FILLER_33_1675 ();
 sg13g2_fill_2 FILLER_33_1680 ();
 sg13g2_fill_1 FILLER_33_1682 ();
 sg13g2_decap_4 FILLER_33_1687 ();
 sg13g2_decap_8 FILLER_33_1716 ();
 sg13g2_decap_8 FILLER_33_1723 ();
 sg13g2_fill_2 FILLER_33_1767 ();
 sg13g2_fill_1 FILLER_33_1775 ();
 sg13g2_fill_1 FILLER_33_1802 ();
 sg13g2_fill_1 FILLER_33_1806 ();
 sg13g2_decap_8 FILLER_33_1852 ();
 sg13g2_decap_4 FILLER_33_1859 ();
 sg13g2_fill_1 FILLER_33_1863 ();
 sg13g2_decap_8 FILLER_33_1882 ();
 sg13g2_decap_8 FILLER_33_1889 ();
 sg13g2_decap_8 FILLER_33_1896 ();
 sg13g2_decap_8 FILLER_33_1903 ();
 sg13g2_decap_8 FILLER_33_1910 ();
 sg13g2_decap_8 FILLER_33_1917 ();
 sg13g2_fill_2 FILLER_33_1924 ();
 sg13g2_fill_1 FILLER_33_1926 ();
 sg13g2_decap_8 FILLER_33_1936 ();
 sg13g2_decap_8 FILLER_33_1943 ();
 sg13g2_fill_1 FILLER_33_1950 ();
 sg13g2_fill_2 FILLER_33_1955 ();
 sg13g2_fill_1 FILLER_33_1957 ();
 sg13g2_decap_8 FILLER_33_1962 ();
 sg13g2_decap_8 FILLER_33_1969 ();
 sg13g2_fill_2 FILLER_33_1976 ();
 sg13g2_fill_1 FILLER_33_2043 ();
 sg13g2_decap_8 FILLER_33_2070 ();
 sg13g2_decap_4 FILLER_33_2077 ();
 sg13g2_fill_2 FILLER_33_2127 ();
 sg13g2_fill_1 FILLER_33_2129 ();
 sg13g2_decap_8 FILLER_33_2154 ();
 sg13g2_fill_1 FILLER_33_2171 ();
 sg13g2_fill_2 FILLER_33_2186 ();
 sg13g2_fill_1 FILLER_33_2188 ();
 sg13g2_fill_1 FILLER_33_2193 ();
 sg13g2_fill_1 FILLER_33_2199 ();
 sg13g2_fill_1 FILLER_33_2210 ();
 sg13g2_decap_8 FILLER_33_2241 ();
 sg13g2_decap_8 FILLER_33_2248 ();
 sg13g2_decap_8 FILLER_33_2255 ();
 sg13g2_fill_2 FILLER_33_2272 ();
 sg13g2_fill_1 FILLER_33_2274 ();
 sg13g2_decap_8 FILLER_33_2301 ();
 sg13g2_decap_4 FILLER_33_2317 ();
 sg13g2_fill_1 FILLER_33_2321 ();
 sg13g2_fill_2 FILLER_33_2329 ();
 sg13g2_fill_1 FILLER_33_2338 ();
 sg13g2_fill_2 FILLER_33_2354 ();
 sg13g2_fill_2 FILLER_33_2387 ();
 sg13g2_fill_1 FILLER_33_2389 ();
 sg13g2_fill_2 FILLER_33_2416 ();
 sg13g2_fill_2 FILLER_33_2426 ();
 sg13g2_fill_2 FILLER_33_2432 ();
 sg13g2_fill_1 FILLER_33_2434 ();
 sg13g2_decap_8 FILLER_33_2488 ();
 sg13g2_fill_1 FILLER_33_2495 ();
 sg13g2_fill_2 FILLER_33_2543 ();
 sg13g2_fill_1 FILLER_33_2545 ();
 sg13g2_decap_8 FILLER_33_2635 ();
 sg13g2_fill_2 FILLER_33_2668 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_9 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_22 ();
 sg13g2_decap_4 FILLER_34_28 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_fill_2 FILLER_34_45 ();
 sg13g2_fill_1 FILLER_34_47 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_81 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_2 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_90 ();
 sg13g2_decap_8 FILLER_34_99 ();
 sg13g2_decap_8 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_141 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_218 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_2 FILLER_34_337 ();
 sg13g2_fill_1 FILLER_34_339 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_365 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_394 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_decap_8 FILLER_34_445 ();
 sg13g2_decap_4 FILLER_34_452 ();
 sg13g2_fill_2 FILLER_34_456 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_482 ();
 sg13g2_decap_8 FILLER_34_489 ();
 sg13g2_fill_1 FILLER_34_509 ();
 sg13g2_fill_2 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_549 ();
 sg13g2_fill_1 FILLER_34_556 ();
 sg13g2_fill_1 FILLER_34_561 ();
 sg13g2_fill_1 FILLER_34_582 ();
 sg13g2_fill_2 FILLER_34_592 ();
 sg13g2_fill_1 FILLER_34_602 ();
 sg13g2_fill_1 FILLER_34_608 ();
 sg13g2_fill_2 FILLER_34_667 ();
 sg13g2_decap_4 FILLER_34_677 ();
 sg13g2_fill_1 FILLER_34_681 ();
 sg13g2_fill_1 FILLER_34_691 ();
 sg13g2_fill_1 FILLER_34_701 ();
 sg13g2_fill_1 FILLER_34_720 ();
 sg13g2_fill_2 FILLER_34_727 ();
 sg13g2_fill_2 FILLER_34_755 ();
 sg13g2_fill_1 FILLER_34_789 ();
 sg13g2_fill_1 FILLER_34_794 ();
 sg13g2_fill_2 FILLER_34_810 ();
 sg13g2_decap_4 FILLER_34_842 ();
 sg13g2_fill_2 FILLER_34_880 ();
 sg13g2_fill_1 FILLER_34_882 ();
 sg13g2_fill_1 FILLER_34_897 ();
 sg13g2_fill_2 FILLER_34_919 ();
 sg13g2_fill_2 FILLER_34_1037 ();
 sg13g2_decap_8 FILLER_34_1073 ();
 sg13g2_decap_8 FILLER_34_1080 ();
 sg13g2_fill_1 FILLER_34_1087 ();
 sg13g2_decap_8 FILLER_34_1143 ();
 sg13g2_fill_2 FILLER_34_1150 ();
 sg13g2_decap_4 FILLER_34_1157 ();
 sg13g2_fill_2 FILLER_34_1161 ();
 sg13g2_fill_1 FILLER_34_1193 ();
 sg13g2_decap_4 FILLER_34_1208 ();
 sg13g2_fill_2 FILLER_34_1212 ();
 sg13g2_decap_8 FILLER_34_1218 ();
 sg13g2_decap_4 FILLER_34_1225 ();
 sg13g2_fill_1 FILLER_34_1229 ();
 sg13g2_decap_4 FILLER_34_1240 ();
 sg13g2_fill_2 FILLER_34_1244 ();
 sg13g2_fill_1 FILLER_34_1250 ();
 sg13g2_fill_2 FILLER_34_1277 ();
 sg13g2_fill_2 FILLER_34_1305 ();
 sg13g2_fill_2 FILLER_34_1333 ();
 sg13g2_fill_1 FILLER_34_1335 ();
 sg13g2_fill_1 FILLER_34_1340 ();
 sg13g2_fill_2 FILLER_34_1367 ();
 sg13g2_fill_1 FILLER_34_1376 ();
 sg13g2_fill_2 FILLER_34_1387 ();
 sg13g2_fill_2 FILLER_34_1415 ();
 sg13g2_decap_8 FILLER_34_1454 ();
 sg13g2_decap_8 FILLER_34_1461 ();
 sg13g2_fill_2 FILLER_34_1468 ();
 sg13g2_fill_1 FILLER_34_1470 ();
 sg13g2_fill_2 FILLER_34_1486 ();
 sg13g2_decap_4 FILLER_34_1516 ();
 sg13g2_decap_8 FILLER_34_1546 ();
 sg13g2_decap_8 FILLER_34_1553 ();
 sg13g2_fill_2 FILLER_34_1560 ();
 sg13g2_fill_2 FILLER_34_1572 ();
 sg13g2_fill_1 FILLER_34_1597 ();
 sg13g2_fill_2 FILLER_34_1611 ();
 sg13g2_fill_1 FILLER_34_1613 ();
 sg13g2_fill_2 FILLER_34_1618 ();
 sg13g2_decap_8 FILLER_34_1640 ();
 sg13g2_fill_1 FILLER_34_1647 ();
 sg13g2_decap_8 FILLER_34_1652 ();
 sg13g2_fill_1 FILLER_34_1659 ();
 sg13g2_fill_2 FILLER_34_1664 ();
 sg13g2_fill_1 FILLER_34_1666 ();
 sg13g2_decap_8 FILLER_34_1693 ();
 sg13g2_decap_4 FILLER_34_1700 ();
 sg13g2_fill_1 FILLER_34_1704 ();
 sg13g2_fill_2 FILLER_34_1711 ();
 sg13g2_fill_1 FILLER_34_1713 ();
 sg13g2_fill_2 FILLER_34_1744 ();
 sg13g2_fill_2 FILLER_34_1759 ();
 sg13g2_fill_1 FILLER_34_1787 ();
 sg13g2_fill_2 FILLER_34_1792 ();
 sg13g2_fill_2 FILLER_34_1797 ();
 sg13g2_fill_1 FILLER_34_1811 ();
 sg13g2_decap_8 FILLER_34_1835 ();
 sg13g2_decap_8 FILLER_34_1842 ();
 sg13g2_decap_8 FILLER_34_1849 ();
 sg13g2_decap_8 FILLER_34_1856 ();
 sg13g2_decap_8 FILLER_34_1863 ();
 sg13g2_decap_4 FILLER_34_1905 ();
 sg13g2_fill_1 FILLER_34_1923 ();
 sg13g2_fill_2 FILLER_34_1963 ();
 sg13g2_fill_1 FILLER_34_1965 ();
 sg13g2_fill_1 FILLER_34_1970 ();
 sg13g2_fill_1 FILLER_34_1979 ();
 sg13g2_fill_1 FILLER_34_1993 ();
 sg13g2_fill_1 FILLER_34_2020 ();
 sg13g2_fill_1 FILLER_34_2042 ();
 sg13g2_fill_1 FILLER_34_2055 ();
 sg13g2_decap_8 FILLER_34_2060 ();
 sg13g2_decap_8 FILLER_34_2067 ();
 sg13g2_decap_8 FILLER_34_2074 ();
 sg13g2_fill_2 FILLER_34_2081 ();
 sg13g2_fill_1 FILLER_34_2083 ();
 sg13g2_decap_8 FILLER_34_2122 ();
 sg13g2_decap_8 FILLER_34_2129 ();
 sg13g2_decap_8 FILLER_34_2136 ();
 sg13g2_decap_8 FILLER_34_2143 ();
 sg13g2_fill_2 FILLER_34_2150 ();
 sg13g2_fill_1 FILLER_34_2152 ();
 sg13g2_decap_4 FILLER_34_2173 ();
 sg13g2_decap_8 FILLER_34_2182 ();
 sg13g2_decap_8 FILLER_34_2189 ();
 sg13g2_fill_2 FILLER_34_2196 ();
 sg13g2_decap_8 FILLER_34_2230 ();
 sg13g2_fill_2 FILLER_34_2237 ();
 sg13g2_decap_8 FILLER_34_2249 ();
 sg13g2_fill_1 FILLER_34_2256 ();
 sg13g2_decap_8 FILLER_34_2302 ();
 sg13g2_decap_8 FILLER_34_2309 ();
 sg13g2_fill_1 FILLER_34_2316 ();
 sg13g2_fill_2 FILLER_34_2340 ();
 sg13g2_fill_2 FILLER_34_2347 ();
 sg13g2_fill_1 FILLER_34_2361 ();
 sg13g2_fill_1 FILLER_34_2377 ();
 sg13g2_decap_4 FILLER_34_2394 ();
 sg13g2_fill_1 FILLER_34_2398 ();
 sg13g2_fill_2 FILLER_34_2403 ();
 sg13g2_fill_2 FILLER_34_2409 ();
 sg13g2_fill_2 FILLER_34_2415 ();
 sg13g2_decap_4 FILLER_34_2422 ();
 sg13g2_fill_2 FILLER_34_2431 ();
 sg13g2_decap_8 FILLER_34_2437 ();
 sg13g2_decap_8 FILLER_34_2444 ();
 sg13g2_decap_8 FILLER_34_2451 ();
 sg13g2_decap_4 FILLER_34_2458 ();
 sg13g2_fill_2 FILLER_34_2462 ();
 sg13g2_decap_4 FILLER_34_2479 ();
 sg13g2_decap_4 FILLER_34_2493 ();
 sg13g2_fill_2 FILLER_34_2513 ();
 sg13g2_fill_1 FILLER_34_2515 ();
 sg13g2_fill_1 FILLER_34_2530 ();
 sg13g2_fill_1 FILLER_34_2583 ();
 sg13g2_fill_1 FILLER_34_2594 ();
 sg13g2_fill_2 FILLER_34_2601 ();
 sg13g2_decap_8 FILLER_34_2651 ();
 sg13g2_decap_8 FILLER_34_2658 ();
 sg13g2_decap_4 FILLER_34_2665 ();
 sg13g2_fill_1 FILLER_34_2669 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_5 ();
 sg13g2_fill_1 FILLER_35_9 ();
 sg13g2_fill_1 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_103 ();
 sg13g2_decap_4 FILLER_35_117 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_fill_2 FILLER_35_130 ();
 sg13g2_fill_1 FILLER_35_132 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_fill_2 FILLER_35_195 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_215 ();
 sg13g2_decap_8 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_229 ();
 sg13g2_fill_2 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_242 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_281 ();
 sg13g2_fill_1 FILLER_35_299 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_decap_4 FILLER_35_393 ();
 sg13g2_fill_2 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_430 ();
 sg13g2_decap_8 FILLER_35_544 ();
 sg13g2_decap_8 FILLER_35_551 ();
 sg13g2_decap_4 FILLER_35_558 ();
 sg13g2_fill_1 FILLER_35_562 ();
 sg13g2_fill_2 FILLER_35_567 ();
 sg13g2_fill_2 FILLER_35_630 ();
 sg13g2_fill_2 FILLER_35_675 ();
 sg13g2_fill_1 FILLER_35_685 ();
 sg13g2_fill_2 FILLER_35_696 ();
 sg13g2_fill_2 FILLER_35_713 ();
 sg13g2_fill_2 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_808 ();
 sg13g2_fill_2 FILLER_35_836 ();
 sg13g2_decap_4 FILLER_35_843 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_858 ();
 sg13g2_fill_1 FILLER_35_865 ();
 sg13g2_decap_8 FILLER_35_876 ();
 sg13g2_fill_2 FILLER_35_883 ();
 sg13g2_fill_2 FILLER_35_893 ();
 sg13g2_fill_1 FILLER_35_895 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_fill_1 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_940 ();
 sg13g2_decap_8 FILLER_35_947 ();
 sg13g2_decap_4 FILLER_35_954 ();
 sg13g2_fill_1 FILLER_35_962 ();
 sg13g2_decap_8 FILLER_35_976 ();
 sg13g2_decap_8 FILLER_35_983 ();
 sg13g2_decap_4 FILLER_35_990 ();
 sg13g2_fill_1 FILLER_35_994 ();
 sg13g2_fill_2 FILLER_35_1000 ();
 sg13g2_fill_1 FILLER_35_1002 ();
 sg13g2_decap_4 FILLER_35_1029 ();
 sg13g2_fill_2 FILLER_35_1033 ();
 sg13g2_fill_1 FILLER_35_1040 ();
 sg13g2_fill_1 FILLER_35_1045 ();
 sg13g2_fill_2 FILLER_35_1089 ();
 sg13g2_fill_1 FILLER_35_1091 ();
 sg13g2_fill_2 FILLER_35_1110 ();
 sg13g2_fill_2 FILLER_35_1151 ();
 sg13g2_fill_2 FILLER_35_1204 ();
 sg13g2_fill_1 FILLER_35_1232 ();
 sg13g2_fill_1 FILLER_35_1263 ();
 sg13g2_fill_2 FILLER_35_1277 ();
 sg13g2_fill_1 FILLER_35_1279 ();
 sg13g2_fill_2 FILLER_35_1285 ();
 sg13g2_decap_8 FILLER_35_1295 ();
 sg13g2_decap_8 FILLER_35_1302 ();
 sg13g2_decap_4 FILLER_35_1309 ();
 sg13g2_decap_8 FILLER_35_1317 ();
 sg13g2_fill_2 FILLER_35_1324 ();
 sg13g2_decap_8 FILLER_35_1361 ();
 sg13g2_decap_8 FILLER_35_1368 ();
 sg13g2_fill_1 FILLER_35_1375 ();
 sg13g2_fill_2 FILLER_35_1388 ();
 sg13g2_fill_1 FILLER_35_1390 ();
 sg13g2_decap_4 FILLER_35_1430 ();
 sg13g2_fill_2 FILLER_35_1434 ();
 sg13g2_decap_8 FILLER_35_1441 ();
 sg13g2_decap_4 FILLER_35_1448 ();
 sg13g2_fill_1 FILLER_35_1456 ();
 sg13g2_fill_1 FILLER_35_1462 ();
 sg13g2_fill_1 FILLER_35_1472 ();
 sg13g2_decap_8 FILLER_35_1507 ();
 sg13g2_decap_8 FILLER_35_1514 ();
 sg13g2_fill_2 FILLER_35_1521 ();
 sg13g2_decap_8 FILLER_35_1531 ();
 sg13g2_fill_2 FILLER_35_1538 ();
 sg13g2_fill_1 FILLER_35_1540 ();
 sg13g2_fill_1 FILLER_35_1610 ();
 sg13g2_decap_8 FILLER_35_1630 ();
 sg13g2_decap_8 FILLER_35_1637 ();
 sg13g2_decap_4 FILLER_35_1644 ();
 sg13g2_decap_8 FILLER_35_1658 ();
 sg13g2_decap_8 FILLER_35_1669 ();
 sg13g2_decap_8 FILLER_35_1702 ();
 sg13g2_decap_8 FILLER_35_1714 ();
 sg13g2_decap_4 FILLER_35_1721 ();
 sg13g2_fill_2 FILLER_35_1725 ();
 sg13g2_fill_1 FILLER_35_1741 ();
 sg13g2_decap_8 FILLER_35_1778 ();
 sg13g2_decap_8 FILLER_35_1785 ();
 sg13g2_fill_1 FILLER_35_1812 ();
 sg13g2_fill_1 FILLER_35_1817 ();
 sg13g2_decap_8 FILLER_35_1826 ();
 sg13g2_decap_8 FILLER_35_1833 ();
 sg13g2_decap_8 FILLER_35_1840 ();
 sg13g2_decap_8 FILLER_35_1847 ();
 sg13g2_decap_4 FILLER_35_1854 ();
 sg13g2_fill_2 FILLER_35_1858 ();
 sg13g2_decap_4 FILLER_35_1865 ();
 sg13g2_decap_4 FILLER_35_1896 ();
 sg13g2_fill_1 FILLER_35_1905 ();
 sg13g2_fill_1 FILLER_35_1944 ();
 sg13g2_fill_2 FILLER_35_1968 ();
 sg13g2_fill_1 FILLER_35_1975 ();
 sg13g2_decap_8 FILLER_35_1980 ();
 sg13g2_fill_1 FILLER_35_1987 ();
 sg13g2_decap_8 FILLER_35_1992 ();
 sg13g2_fill_1 FILLER_35_1999 ();
 sg13g2_decap_8 FILLER_35_2004 ();
 sg13g2_fill_2 FILLER_35_2011 ();
 sg13g2_fill_1 FILLER_35_2013 ();
 sg13g2_decap_4 FILLER_35_2040 ();
 sg13g2_fill_1 FILLER_35_2044 ();
 sg13g2_decap_4 FILLER_35_2069 ();
 sg13g2_decap_8 FILLER_35_2085 ();
 sg13g2_decap_4 FILLER_35_2092 ();
 sg13g2_fill_1 FILLER_35_2096 ();
 sg13g2_decap_8 FILLER_35_2107 ();
 sg13g2_fill_1 FILLER_35_2114 ();
 sg13g2_decap_8 FILLER_35_2125 ();
 sg13g2_decap_8 FILLER_35_2158 ();
 sg13g2_fill_1 FILLER_35_2186 ();
 sg13g2_fill_1 FILLER_35_2210 ();
 sg13g2_decap_8 FILLER_35_2296 ();
 sg13g2_decap_4 FILLER_35_2303 ();
 sg13g2_fill_1 FILLER_35_2307 ();
 sg13g2_fill_1 FILLER_35_2315 ();
 sg13g2_fill_1 FILLER_35_2359 ();
 sg13g2_fill_1 FILLER_35_2364 ();
 sg13g2_fill_1 FILLER_35_2392 ();
 sg13g2_decap_8 FILLER_35_2397 ();
 sg13g2_fill_2 FILLER_35_2404 ();
 sg13g2_fill_1 FILLER_35_2436 ();
 sg13g2_fill_1 FILLER_35_2441 ();
 sg13g2_fill_2 FILLER_35_2452 ();
 sg13g2_fill_1 FILLER_35_2458 ();
 sg13g2_fill_1 FILLER_35_2464 ();
 sg13g2_fill_1 FILLER_35_2475 ();
 sg13g2_fill_1 FILLER_35_2484 ();
 sg13g2_fill_1 FILLER_35_2525 ();
 sg13g2_decap_8 FILLER_35_2552 ();
 sg13g2_fill_2 FILLER_35_2559 ();
 sg13g2_fill_1 FILLER_35_2561 ();
 sg13g2_fill_2 FILLER_35_2571 ();
 sg13g2_decap_8 FILLER_35_2612 ();
 sg13g2_decap_8 FILLER_35_2619 ();
 sg13g2_fill_2 FILLER_35_2626 ();
 sg13g2_fill_1 FILLER_35_2628 ();
 sg13g2_fill_2 FILLER_35_2668 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_57 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_decap_4 FILLER_36_71 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_decap_4 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_4 FILLER_36_158 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_2 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_236 ();
 sg13g2_decap_4 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_247 ();
 sg13g2_fill_1 FILLER_36_271 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_379 ();
 sg13g2_fill_1 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_fill_2 FILLER_36_410 ();
 sg13g2_fill_2 FILLER_36_416 ();
 sg13g2_fill_2 FILLER_36_502 ();
 sg13g2_fill_1 FILLER_36_510 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_decap_4 FILLER_36_549 ();
 sg13g2_fill_2 FILLER_36_553 ();
 sg13g2_decap_4 FILLER_36_559 ();
 sg13g2_fill_2 FILLER_36_563 ();
 sg13g2_fill_1 FILLER_36_586 ();
 sg13g2_decap_4 FILLER_36_598 ();
 sg13g2_fill_2 FILLER_36_602 ();
 sg13g2_decap_4 FILLER_36_608 ();
 sg13g2_fill_1 FILLER_36_612 ();
 sg13g2_decap_4 FILLER_36_618 ();
 sg13g2_fill_2 FILLER_36_622 ();
 sg13g2_decap_4 FILLER_36_634 ();
 sg13g2_decap_4 FILLER_36_647 ();
 sg13g2_fill_2 FILLER_36_655 ();
 sg13g2_fill_2 FILLER_36_661 ();
 sg13g2_fill_2 FILLER_36_668 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_decap_4 FILLER_36_697 ();
 sg13g2_fill_2 FILLER_36_733 ();
 sg13g2_decap_4 FILLER_36_766 ();
 sg13g2_fill_1 FILLER_36_770 ();
 sg13g2_fill_2 FILLER_36_810 ();
 sg13g2_decap_4 FILLER_36_825 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_4 FILLER_36_847 ();
 sg13g2_fill_1 FILLER_36_851 ();
 sg13g2_decap_4 FILLER_36_878 ();
 sg13g2_fill_1 FILLER_36_882 ();
 sg13g2_decap_4 FILLER_36_909 ();
 sg13g2_fill_2 FILLER_36_913 ();
 sg13g2_fill_2 FILLER_36_955 ();
 sg13g2_fill_1 FILLER_36_957 ();
 sg13g2_decap_4 FILLER_36_987 ();
 sg13g2_fill_2 FILLER_36_991 ();
 sg13g2_fill_1 FILLER_36_1002 ();
 sg13g2_fill_2 FILLER_36_1007 ();
 sg13g2_fill_2 FILLER_36_1013 ();
 sg13g2_decap_8 FILLER_36_1019 ();
 sg13g2_decap_4 FILLER_36_1026 ();
 sg13g2_fill_1 FILLER_36_1030 ();
 sg13g2_decap_8 FILLER_36_1083 ();
 sg13g2_decap_4 FILLER_36_1120 ();
 sg13g2_fill_1 FILLER_36_1124 ();
 sg13g2_decap_4 FILLER_36_1154 ();
 sg13g2_decap_4 FILLER_36_1162 ();
 sg13g2_fill_2 FILLER_36_1166 ();
 sg13g2_fill_2 FILLER_36_1198 ();
 sg13g2_fill_1 FILLER_36_1200 ();
 sg13g2_decap_4 FILLER_36_1206 ();
 sg13g2_fill_1 FILLER_36_1210 ();
 sg13g2_decap_4 FILLER_36_1221 ();
 sg13g2_fill_1 FILLER_36_1225 ();
 sg13g2_fill_2 FILLER_36_1251 ();
 sg13g2_fill_1 FILLER_36_1253 ();
 sg13g2_decap_8 FILLER_36_1259 ();
 sg13g2_decap_8 FILLER_36_1296 ();
 sg13g2_decap_8 FILLER_36_1303 ();
 sg13g2_fill_1 FILLER_36_1310 ();
 sg13g2_decap_8 FILLER_36_1316 ();
 sg13g2_fill_1 FILLER_36_1323 ();
 sg13g2_fill_1 FILLER_36_1360 ();
 sg13g2_fill_2 FILLER_36_1371 ();
 sg13g2_fill_1 FILLER_36_1394 ();
 sg13g2_fill_1 FILLER_36_1411 ();
 sg13g2_fill_2 FILLER_36_1423 ();
 sg13g2_fill_2 FILLER_36_1456 ();
 sg13g2_decap_4 FILLER_36_1479 ();
 sg13g2_fill_1 FILLER_36_1498 ();
 sg13g2_decap_4 FILLER_36_1525 ();
 sg13g2_decap_8 FILLER_36_1533 ();
 sg13g2_decap_4 FILLER_36_1540 ();
 sg13g2_fill_1 FILLER_36_1554 ();
 sg13g2_decap_8 FILLER_36_1558 ();
 sg13g2_fill_2 FILLER_36_1565 ();
 sg13g2_decap_4 FILLER_36_1571 ();
 sg13g2_fill_1 FILLER_36_1575 ();
 sg13g2_decap_8 FILLER_36_1580 ();
 sg13g2_decap_4 FILLER_36_1591 ();
 sg13g2_fill_2 FILLER_36_1600 ();
 sg13g2_fill_1 FILLER_36_1602 ();
 sg13g2_decap_4 FILLER_36_1612 ();
 sg13g2_fill_2 FILLER_36_1616 ();
 sg13g2_fill_2 FILLER_36_1683 ();
 sg13g2_decap_8 FILLER_36_1734 ();
 sg13g2_decap_8 FILLER_36_1767 ();
 sg13g2_decap_8 FILLER_36_1774 ();
 sg13g2_decap_4 FILLER_36_1781 ();
 sg13g2_fill_2 FILLER_36_1810 ();
 sg13g2_decap_8 FILLER_36_1846 ();
 sg13g2_decap_4 FILLER_36_1858 ();
 sg13g2_fill_1 FILLER_36_1862 ();
 sg13g2_fill_2 FILLER_36_1884 ();
 sg13g2_fill_2 FILLER_36_1889 ();
 sg13g2_fill_1 FILLER_36_1900 ();
 sg13g2_fill_1 FILLER_36_1932 ();
 sg13g2_fill_1 FILLER_36_1955 ();
 sg13g2_fill_1 FILLER_36_1971 ();
 sg13g2_fill_1 FILLER_36_1986 ();
 sg13g2_decap_4 FILLER_36_1991 ();
 sg13g2_fill_1 FILLER_36_1995 ();
 sg13g2_decap_4 FILLER_36_2010 ();
 sg13g2_fill_1 FILLER_36_2014 ();
 sg13g2_fill_2 FILLER_36_2030 ();
 sg13g2_fill_1 FILLER_36_2032 ();
 sg13g2_fill_2 FILLER_36_2082 ();
 sg13g2_fill_1 FILLER_36_2084 ();
 sg13g2_fill_2 FILLER_36_2147 ();
 sg13g2_fill_2 FILLER_36_2175 ();
 sg13g2_fill_1 FILLER_36_2177 ();
 sg13g2_decap_4 FILLER_36_2213 ();
 sg13g2_decap_8 FILLER_36_2221 ();
 sg13g2_decap_8 FILLER_36_2228 ();
 sg13g2_decap_4 FILLER_36_2235 ();
 sg13g2_fill_2 FILLER_36_2279 ();
 sg13g2_decap_4 FILLER_36_2307 ();
 sg13g2_fill_1 FILLER_36_2311 ();
 sg13g2_fill_1 FILLER_36_2346 ();
 sg13g2_decap_4 FILLER_36_2379 ();
 sg13g2_fill_2 FILLER_36_2383 ();
 sg13g2_fill_2 FILLER_36_2430 ();
 sg13g2_fill_2 FILLER_36_2458 ();
 sg13g2_fill_1 FILLER_36_2460 ();
 sg13g2_fill_2 FILLER_36_2497 ();
 sg13g2_fill_1 FILLER_36_2499 ();
 sg13g2_fill_1 FILLER_36_2536 ();
 sg13g2_fill_1 FILLER_36_2541 ();
 sg13g2_fill_1 FILLER_36_2545 ();
 sg13g2_fill_2 FILLER_36_2617 ();
 sg13g2_fill_1 FILLER_36_2619 ();
 sg13g2_decap_8 FILLER_36_2660 ();
 sg13g2_fill_2 FILLER_36_2667 ();
 sg13g2_fill_1 FILLER_36_2669 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_decap_4 FILLER_37_47 ();
 sg13g2_decap_4 FILLER_37_68 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_fill_1 FILLER_37_135 ();
 sg13g2_fill_1 FILLER_37_175 ();
 sg13g2_decap_4 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_decap_4 FILLER_37_201 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_4 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_decap_4 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_305 ();
 sg13g2_decap_4 FILLER_37_310 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_fill_1 FILLER_37_333 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_decap_4 FILLER_37_395 ();
 sg13g2_decap_8 FILLER_37_403 ();
 sg13g2_decap_8 FILLER_37_410 ();
 sg13g2_fill_2 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_37_465 ();
 sg13g2_fill_2 FILLER_37_510 ();
 sg13g2_fill_1 FILLER_37_536 ();
 sg13g2_fill_2 FILLER_37_560 ();
 sg13g2_fill_1 FILLER_37_567 ();
 sg13g2_fill_2 FILLER_37_573 ();
 sg13g2_fill_2 FILLER_37_609 ();
 sg13g2_fill_1 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_631 ();
 sg13g2_decap_8 FILLER_37_638 ();
 sg13g2_fill_1 FILLER_37_645 ();
 sg13g2_fill_2 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_662 ();
 sg13g2_decap_8 FILLER_37_669 ();
 sg13g2_fill_2 FILLER_37_676 ();
 sg13g2_fill_1 FILLER_37_683 ();
 sg13g2_fill_1 FILLER_37_689 ();
 sg13g2_fill_2 FILLER_37_695 ();
 sg13g2_fill_1 FILLER_37_697 ();
 sg13g2_fill_2 FILLER_37_743 ();
 sg13g2_fill_2 FILLER_37_771 ();
 sg13g2_fill_1 FILLER_37_773 ();
 sg13g2_fill_2 FILLER_37_783 ();
 sg13g2_fill_1 FILLER_37_814 ();
 sg13g2_fill_2 FILLER_37_841 ();
 sg13g2_fill_1 FILLER_37_857 ();
 sg13g2_decap_4 FILLER_37_918 ();
 sg13g2_fill_2 FILLER_37_922 ();
 sg13g2_fill_2 FILLER_37_950 ();
 sg13g2_fill_1 FILLER_37_952 ();
 sg13g2_decap_4 FILLER_37_963 ();
 sg13g2_fill_2 FILLER_37_967 ();
 sg13g2_fill_1 FILLER_37_1009 ();
 sg13g2_decap_8 FILLER_37_1014 ();
 sg13g2_decap_8 FILLER_37_1021 ();
 sg13g2_decap_8 FILLER_37_1028 ();
 sg13g2_decap_4 FILLER_37_1035 ();
 sg13g2_fill_2 FILLER_37_1043 ();
 sg13g2_fill_1 FILLER_37_1045 ();
 sg13g2_decap_4 FILLER_37_1051 ();
 sg13g2_fill_1 FILLER_37_1055 ();
 sg13g2_fill_2 FILLER_37_1060 ();
 sg13g2_decap_4 FILLER_37_1066 ();
 sg13g2_decap_4 FILLER_37_1105 ();
 sg13g2_fill_1 FILLER_37_1109 ();
 sg13g2_fill_1 FILLER_37_1114 ();
 sg13g2_decap_4 FILLER_37_1120 ();
 sg13g2_fill_2 FILLER_37_1124 ();
 sg13g2_decap_8 FILLER_37_1152 ();
 sg13g2_fill_1 FILLER_37_1159 ();
 sg13g2_fill_1 FILLER_37_1169 ();
 sg13g2_fill_2 FILLER_37_1179 ();
 sg13g2_fill_1 FILLER_37_1181 ();
 sg13g2_decap_8 FILLER_37_1186 ();
 sg13g2_fill_2 FILLER_37_1193 ();
 sg13g2_fill_1 FILLER_37_1195 ();
 sg13g2_decap_4 FILLER_37_1219 ();
 sg13g2_decap_8 FILLER_37_1244 ();
 sg13g2_decap_8 FILLER_37_1251 ();
 sg13g2_decap_4 FILLER_37_1258 ();
 sg13g2_fill_1 FILLER_37_1262 ();
 sg13g2_fill_2 FILLER_37_1271 ();
 sg13g2_fill_1 FILLER_37_1281 ();
 sg13g2_fill_1 FILLER_37_1287 ();
 sg13g2_decap_8 FILLER_37_1318 ();
 sg13g2_decap_8 FILLER_37_1325 ();
 sg13g2_fill_1 FILLER_37_1332 ();
 sg13g2_fill_1 FILLER_37_1337 ();
 sg13g2_decap_8 FILLER_37_1360 ();
 sg13g2_fill_1 FILLER_37_1367 ();
 sg13g2_decap_4 FILLER_37_1371 ();
 sg13g2_fill_2 FILLER_37_1375 ();
 sg13g2_decap_4 FILLER_37_1382 ();
 sg13g2_fill_1 FILLER_37_1397 ();
 sg13g2_fill_2 FILLER_37_1424 ();
 sg13g2_fill_1 FILLER_37_1431 ();
 sg13g2_fill_2 FILLER_37_1438 ();
 sg13g2_fill_1 FILLER_37_1444 ();
 sg13g2_fill_1 FILLER_37_1450 ();
 sg13g2_fill_1 FILLER_37_1489 ();
 sg13g2_fill_2 FILLER_37_1509 ();
 sg13g2_fill_1 FILLER_37_1521 ();
 sg13g2_fill_1 FILLER_37_1548 ();
 sg13g2_fill_1 FILLER_37_1553 ();
 sg13g2_fill_1 FILLER_37_1580 ();
 sg13g2_fill_1 FILLER_37_1594 ();
 sg13g2_decap_8 FILLER_37_1608 ();
 sg13g2_fill_1 FILLER_37_1615 ();
 sg13g2_decap_8 FILLER_37_1662 ();
 sg13g2_decap_8 FILLER_37_1669 ();
 sg13g2_decap_4 FILLER_37_1676 ();
 sg13g2_fill_1 FILLER_37_1680 ();
 sg13g2_fill_2 FILLER_37_1692 ();
 sg13g2_decap_4 FILLER_37_1700 ();
 sg13g2_decap_8 FILLER_37_1708 ();
 sg13g2_decap_8 FILLER_37_1715 ();
 sg13g2_decap_8 FILLER_37_1722 ();
 sg13g2_fill_1 FILLER_37_1729 ();
 sg13g2_decap_4 FILLER_37_1735 ();
 sg13g2_fill_2 FILLER_37_1739 ();
 sg13g2_decap_8 FILLER_37_1759 ();
 sg13g2_fill_1 FILLER_37_1766 ();
 sg13g2_decap_8 FILLER_37_1803 ();
 sg13g2_decap_8 FILLER_37_1810 ();
 sg13g2_fill_2 FILLER_37_1817 ();
 sg13g2_decap_8 FILLER_37_1829 ();
 sg13g2_fill_2 FILLER_37_1836 ();
 sg13g2_fill_1 FILLER_37_1838 ();
 sg13g2_fill_2 FILLER_37_1843 ();
 sg13g2_fill_1 FILLER_37_1850 ();
 sg13g2_fill_1 FILLER_37_1855 ();
 sg13g2_fill_2 FILLER_37_1886 ();
 sg13g2_fill_2 FILLER_37_1892 ();
 sg13g2_fill_1 FILLER_37_1894 ();
 sg13g2_fill_2 FILLER_37_1904 ();
 sg13g2_fill_1 FILLER_37_1915 ();
 sg13g2_fill_1 FILLER_37_1926 ();
 sg13g2_fill_1 FILLER_37_1936 ();
 sg13g2_fill_2 FILLER_37_1941 ();
 sg13g2_fill_1 FILLER_37_1948 ();
 sg13g2_decap_8 FILLER_37_1992 ();
 sg13g2_decap_8 FILLER_37_1999 ();
 sg13g2_decap_8 FILLER_37_2006 ();
 sg13g2_fill_2 FILLER_37_2013 ();
 sg13g2_fill_1 FILLER_37_2015 ();
 sg13g2_decap_8 FILLER_37_2029 ();
 sg13g2_fill_2 FILLER_37_2036 ();
 sg13g2_fill_2 FILLER_37_2082 ();
 sg13g2_fill_1 FILLER_37_2110 ();
 sg13g2_decap_4 FILLER_37_2136 ();
 sg13g2_fill_2 FILLER_37_2140 ();
 sg13g2_fill_2 FILLER_37_2146 ();
 sg13g2_fill_1 FILLER_37_2158 ();
 sg13g2_decap_8 FILLER_37_2223 ();
 sg13g2_fill_1 FILLER_37_2243 ();
 sg13g2_decap_4 FILLER_37_2248 ();
 sg13g2_decap_8 FILLER_37_2260 ();
 sg13g2_decap_8 FILLER_37_2293 ();
 sg13g2_decap_4 FILLER_37_2300 ();
 sg13g2_fill_1 FILLER_37_2304 ();
 sg13g2_fill_1 FILLER_37_2331 ();
 sg13g2_fill_1 FILLER_37_2346 ();
 sg13g2_fill_1 FILLER_37_2376 ();
 sg13g2_fill_1 FILLER_37_2408 ();
 sg13g2_fill_1 FILLER_37_2413 ();
 sg13g2_fill_1 FILLER_37_2418 ();
 sg13g2_fill_1 FILLER_37_2427 ();
 sg13g2_fill_2 FILLER_37_2434 ();
 sg13g2_decap_4 FILLER_37_2450 ();
 sg13g2_fill_1 FILLER_37_2459 ();
 sg13g2_decap_8 FILLER_37_2500 ();
 sg13g2_decap_8 FILLER_37_2507 ();
 sg13g2_fill_2 FILLER_37_2514 ();
 sg13g2_fill_2 FILLER_37_2519 ();
 sg13g2_fill_1 FILLER_37_2521 ();
 sg13g2_fill_2 FILLER_37_2525 ();
 sg13g2_fill_1 FILLER_37_2532 ();
 sg13g2_fill_2 FILLER_37_2540 ();
 sg13g2_fill_2 FILLER_37_2563 ();
 sg13g2_decap_4 FILLER_37_2633 ();
 sg13g2_decap_8 FILLER_37_2641 ();
 sg13g2_fill_1 FILLER_37_2648 ();
 sg13g2_decap_8 FILLER_37_2653 ();
 sg13g2_decap_8 FILLER_37_2660 ();
 sg13g2_fill_2 FILLER_37_2667 ();
 sg13g2_fill_1 FILLER_37_2669 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_12 ();
 sg13g2_fill_2 FILLER_38_17 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_57 ();
 sg13g2_fill_2 FILLER_38_64 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_4 FILLER_38_165 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_fill_2 FILLER_38_174 ();
 sg13g2_fill_1 FILLER_38_176 ();
 sg13g2_decap_8 FILLER_38_181 ();
 sg13g2_decap_4 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_192 ();
 sg13g2_fill_2 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_222 ();
 sg13g2_fill_1 FILLER_38_224 ();
 sg13g2_decap_4 FILLER_38_282 ();
 sg13g2_decap_8 FILLER_38_290 ();
 sg13g2_decap_8 FILLER_38_297 ();
 sg13g2_decap_8 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_fill_1 FILLER_38_318 ();
 sg13g2_fill_2 FILLER_38_345 ();
 sg13g2_fill_1 FILLER_38_366 ();
 sg13g2_decap_4 FILLER_38_376 ();
 sg13g2_fill_1 FILLER_38_380 ();
 sg13g2_fill_2 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_413 ();
 sg13g2_fill_1 FILLER_38_422 ();
 sg13g2_fill_2 FILLER_38_432 ();
 sg13g2_fill_2 FILLER_38_468 ();
 sg13g2_fill_1 FILLER_38_515 ();
 sg13g2_fill_2 FILLER_38_533 ();
 sg13g2_fill_2 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_593 ();
 sg13g2_decap_4 FILLER_38_654 ();
 sg13g2_fill_1 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_667 ();
 sg13g2_decap_4 FILLER_38_674 ();
 sg13g2_fill_1 FILLER_38_678 ();
 sg13g2_fill_2 FILLER_38_684 ();
 sg13g2_fill_1 FILLER_38_686 ();
 sg13g2_fill_1 FILLER_38_692 ();
 sg13g2_fill_2 FILLER_38_724 ();
 sg13g2_fill_1 FILLER_38_726 ();
 sg13g2_fill_1 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_758 ();
 sg13g2_decap_8 FILLER_38_764 ();
 sg13g2_decap_4 FILLER_38_771 ();
 sg13g2_fill_1 FILLER_38_775 ();
 sg13g2_fill_2 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_790 ();
 sg13g2_decap_4 FILLER_38_797 ();
 sg13g2_fill_2 FILLER_38_801 ();
 sg13g2_fill_1 FILLER_38_813 ();
 sg13g2_decap_8 FILLER_38_850 ();
 sg13g2_decap_4 FILLER_38_857 ();
 sg13g2_fill_2 FILLER_38_861 ();
 sg13g2_decap_4 FILLER_38_921 ();
 sg13g2_decap_4 FILLER_38_976 ();
 sg13g2_fill_2 FILLER_38_980 ();
 sg13g2_decap_4 FILLER_38_986 ();
 sg13g2_fill_2 FILLER_38_990 ();
 sg13g2_fill_2 FILLER_38_1002 ();
 sg13g2_fill_1 FILLER_38_1060 ();
 sg13g2_decap_8 FILLER_38_1090 ();
 sg13g2_decap_8 FILLER_38_1097 ();
 sg13g2_decap_8 FILLER_38_1104 ();
 sg13g2_decap_4 FILLER_38_1119 ();
 sg13g2_fill_1 FILLER_38_1123 ();
 sg13g2_fill_1 FILLER_38_1154 ();
 sg13g2_fill_2 FILLER_38_1168 ();
 sg13g2_fill_1 FILLER_38_1174 ();
 sg13g2_fill_1 FILLER_38_1179 ();
 sg13g2_fill_1 FILLER_38_1184 ();
 sg13g2_decap_4 FILLER_38_1189 ();
 sg13g2_decap_4 FILLER_38_1197 ();
 sg13g2_fill_2 FILLER_38_1201 ();
 sg13g2_decap_4 FILLER_38_1285 ();
 sg13g2_fill_1 FILLER_38_1289 ();
 sg13g2_fill_2 FILLER_38_1299 ();
 sg13g2_fill_1 FILLER_38_1301 ();
 sg13g2_decap_4 FILLER_38_1384 ();
 sg13g2_fill_1 FILLER_38_1427 ();
 sg13g2_fill_2 FILLER_38_1433 ();
 sg13g2_fill_1 FILLER_38_1476 ();
 sg13g2_decap_8 FILLER_38_1491 ();
 sg13g2_decap_8 FILLER_38_1498 ();
 sg13g2_decap_4 FILLER_38_1505 ();
 sg13g2_fill_2 FILLER_38_1509 ();
 sg13g2_fill_2 FILLER_38_1516 ();
 sg13g2_fill_1 FILLER_38_1545 ();
 sg13g2_fill_1 FILLER_38_1577 ();
 sg13g2_decap_8 FILLER_38_1609 ();
 sg13g2_decap_8 FILLER_38_1616 ();
 sg13g2_decap_4 FILLER_38_1623 ();
 sg13g2_fill_2 FILLER_38_1636 ();
 sg13g2_decap_4 FILLER_38_1642 ();
 sg13g2_decap_4 FILLER_38_1651 ();
 sg13g2_fill_2 FILLER_38_1681 ();
 sg13g2_fill_1 FILLER_38_1683 ();
 sg13g2_decap_4 FILLER_38_1689 ();
 sg13g2_fill_1 FILLER_38_1693 ();
 sg13g2_decap_8 FILLER_38_1698 ();
 sg13g2_decap_8 FILLER_38_1705 ();
 sg13g2_decap_8 FILLER_38_1712 ();
 sg13g2_decap_8 FILLER_38_1719 ();
 sg13g2_decap_8 FILLER_38_1726 ();
 sg13g2_decap_8 FILLER_38_1733 ();
 sg13g2_fill_2 FILLER_38_1748 ();
 sg13g2_decap_8 FILLER_38_1760 ();
 sg13g2_decap_4 FILLER_38_1767 ();
 sg13g2_fill_1 FILLER_38_1771 ();
 sg13g2_decap_8 FILLER_38_1776 ();
 sg13g2_fill_2 FILLER_38_1783 ();
 sg13g2_fill_1 FILLER_38_1785 ();
 sg13g2_decap_8 FILLER_38_1820 ();
 sg13g2_decap_8 FILLER_38_1827 ();
 sg13g2_fill_2 FILLER_38_1834 ();
 sg13g2_fill_1 FILLER_38_1857 ();
 sg13g2_fill_2 FILLER_38_1878 ();
 sg13g2_fill_1 FILLER_38_1889 ();
 sg13g2_decap_4 FILLER_38_1895 ();
 sg13g2_fill_1 FILLER_38_1903 ();
 sg13g2_fill_1 FILLER_38_1909 ();
 sg13g2_decap_4 FILLER_38_1943 ();
 sg13g2_decap_4 FILLER_38_1987 ();
 sg13g2_fill_2 FILLER_38_1991 ();
 sg13g2_decap_8 FILLER_38_1996 ();
 sg13g2_decap_4 FILLER_38_2003 ();
 sg13g2_fill_1 FILLER_38_2007 ();
 sg13g2_fill_2 FILLER_38_2013 ();
 sg13g2_fill_1 FILLER_38_2022 ();
 sg13g2_fill_2 FILLER_38_2085 ();
 sg13g2_fill_2 FILLER_38_2128 ();
 sg13g2_fill_1 FILLER_38_2130 ();
 sg13g2_fill_1 FILLER_38_2141 ();
 sg13g2_fill_2 FILLER_38_2155 ();
 sg13g2_decap_8 FILLER_38_2175 ();
 sg13g2_fill_2 FILLER_38_2182 ();
 sg13g2_fill_2 FILLER_38_2218 ();
 sg13g2_fill_2 FILLER_38_2230 ();
 sg13g2_fill_2 FILLER_38_2258 ();
 sg13g2_fill_1 FILLER_38_2260 ();
 sg13g2_decap_8 FILLER_38_2297 ();
 sg13g2_decap_4 FILLER_38_2304 ();
 sg13g2_fill_1 FILLER_38_2308 ();
 sg13g2_decap_8 FILLER_38_2313 ();
 sg13g2_decap_8 FILLER_38_2320 ();
 sg13g2_decap_4 FILLER_38_2327 ();
 sg13g2_fill_1 FILLER_38_2331 ();
 sg13g2_decap_4 FILLER_38_2342 ();
 sg13g2_fill_1 FILLER_38_2346 ();
 sg13g2_fill_2 FILLER_38_2355 ();
 sg13g2_fill_1 FILLER_38_2357 ();
 sg13g2_decap_4 FILLER_38_2362 ();
 sg13g2_fill_2 FILLER_38_2366 ();
 sg13g2_fill_2 FILLER_38_2398 ();
 sg13g2_decap_4 FILLER_38_2404 ();
 sg13g2_fill_1 FILLER_38_2408 ();
 sg13g2_fill_1 FILLER_38_2413 ();
 sg13g2_fill_1 FILLER_38_2417 ();
 sg13g2_fill_1 FILLER_38_2423 ();
 sg13g2_fill_1 FILLER_38_2431 ();
 sg13g2_fill_1 FILLER_38_2437 ();
 sg13g2_fill_1 FILLER_38_2464 ();
 sg13g2_decap_8 FILLER_38_2479 ();
 sg13g2_decap_8 FILLER_38_2486 ();
 sg13g2_decap_8 FILLER_38_2493 ();
 sg13g2_decap_8 FILLER_38_2500 ();
 sg13g2_fill_1 FILLER_38_2521 ();
 sg13g2_fill_1 FILLER_38_2526 ();
 sg13g2_fill_1 FILLER_38_2532 ();
 sg13g2_fill_1 FILLER_38_2538 ();
 sg13g2_fill_2 FILLER_38_2562 ();
 sg13g2_fill_1 FILLER_38_2597 ();
 sg13g2_fill_2 FILLER_38_2602 ();
 sg13g2_decap_4 FILLER_38_2610 ();
 sg13g2_decap_8 FILLER_38_2618 ();
 sg13g2_fill_2 FILLER_38_2625 ();
 sg13g2_decap_8 FILLER_38_2656 ();
 sg13g2_decap_8 FILLER_38_2663 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_decap_4 FILLER_39_93 ();
 sg13g2_fill_1 FILLER_39_101 ();
 sg13g2_fill_1 FILLER_39_115 ();
 sg13g2_fill_1 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_fill_2 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_228 ();
 sg13g2_fill_2 FILLER_39_243 ();
 sg13g2_fill_1 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_289 ();
 sg13g2_decap_8 FILLER_39_300 ();
 sg13g2_decap_4 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_311 ();
 sg13g2_decap_4 FILLER_39_317 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_fill_2 FILLER_39_348 ();
 sg13g2_fill_1 FILLER_39_387 ();
 sg13g2_decap_4 FILLER_39_425 ();
 sg13g2_fill_2 FILLER_39_434 ();
 sg13g2_fill_2 FILLER_39_500 ();
 sg13g2_fill_2 FILLER_39_525 ();
 sg13g2_fill_2 FILLER_39_571 ();
 sg13g2_fill_1 FILLER_39_573 ();
 sg13g2_fill_2 FILLER_39_600 ();
 sg13g2_decap_8 FILLER_39_612 ();
 sg13g2_fill_1 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_628 ();
 sg13g2_decap_8 FILLER_39_635 ();
 sg13g2_decap_4 FILLER_39_642 ();
 sg13g2_fill_1 FILLER_39_646 ();
 sg13g2_fill_1 FILLER_39_661 ();
 sg13g2_fill_2 FILLER_39_693 ();
 sg13g2_fill_2 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_738 ();
 sg13g2_fill_1 FILLER_39_740 ();
 sg13g2_fill_2 FILLER_39_749 ();
 sg13g2_fill_1 FILLER_39_751 ();
 sg13g2_decap_8 FILLER_39_769 ();
 sg13g2_fill_1 FILLER_39_776 ();
 sg13g2_fill_1 FILLER_39_785 ();
 sg13g2_fill_1 FILLER_39_794 ();
 sg13g2_fill_2 FILLER_39_835 ();
 sg13g2_fill_1 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_848 ();
 sg13g2_fill_2 FILLER_39_855 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_4 FILLER_39_875 ();
 sg13g2_decap_4 FILLER_39_883 ();
 sg13g2_fill_1 FILLER_39_887 ();
 sg13g2_decap_4 FILLER_39_919 ();
 sg13g2_fill_1 FILLER_39_923 ();
 sg13g2_decap_4 FILLER_39_941 ();
 sg13g2_fill_1 FILLER_39_945 ();
 sg13g2_fill_2 FILLER_39_972 ();
 sg13g2_decap_4 FILLER_39_1004 ();
 sg13g2_fill_2 FILLER_39_1013 ();
 sg13g2_fill_1 FILLER_39_1015 ();
 sg13g2_decap_8 FILLER_39_1020 ();
 sg13g2_decap_4 FILLER_39_1027 ();
 sg13g2_fill_2 FILLER_39_1031 ();
 sg13g2_decap_8 FILLER_39_1080 ();
 sg13g2_decap_8 FILLER_39_1087 ();
 sg13g2_decap_8 FILLER_39_1094 ();
 sg13g2_fill_2 FILLER_39_1101 ();
 sg13g2_fill_1 FILLER_39_1103 ();
 sg13g2_fill_1 FILLER_39_1125 ();
 sg13g2_fill_2 FILLER_39_1140 ();
 sg13g2_fill_1 FILLER_39_1142 ();
 sg13g2_fill_2 FILLER_39_1147 ();
 sg13g2_fill_1 FILLER_39_1187 ();
 sg13g2_decap_8 FILLER_39_1197 ();
 sg13g2_decap_4 FILLER_39_1204 ();
 sg13g2_fill_1 FILLER_39_1208 ();
 sg13g2_decap_8 FILLER_39_1213 ();
 sg13g2_decap_4 FILLER_39_1220 ();
 sg13g2_decap_8 FILLER_39_1238 ();
 sg13g2_decap_8 FILLER_39_1245 ();
 sg13g2_fill_2 FILLER_39_1252 ();
 sg13g2_decap_8 FILLER_39_1298 ();
 sg13g2_fill_1 FILLER_39_1331 ();
 sg13g2_fill_1 FILLER_39_1345 ();
 sg13g2_fill_1 FILLER_39_1363 ();
 sg13g2_fill_1 FILLER_39_1377 ();
 sg13g2_fill_2 FILLER_39_1437 ();
 sg13g2_fill_1 FILLER_39_1480 ();
 sg13g2_decap_4 FILLER_39_1485 ();
 sg13g2_fill_1 FILLER_39_1489 ();
 sg13g2_decap_8 FILLER_39_1494 ();
 sg13g2_decap_8 FILLER_39_1501 ();
 sg13g2_decap_8 FILLER_39_1508 ();
 sg13g2_fill_2 FILLER_39_1515 ();
 sg13g2_fill_1 FILLER_39_1537 ();
 sg13g2_fill_2 FILLER_39_1546 ();
 sg13g2_decap_4 FILLER_39_1553 ();
 sg13g2_fill_2 FILLER_39_1561 ();
 sg13g2_decap_4 FILLER_39_1567 ();
 sg13g2_decap_4 FILLER_39_1576 ();
 sg13g2_fill_1 FILLER_39_1580 ();
 sg13g2_fill_1 FILLER_39_1594 ();
 sg13g2_decap_8 FILLER_39_1599 ();
 sg13g2_fill_1 FILLER_39_1606 ();
 sg13g2_fill_1 FILLER_39_1629 ();
 sg13g2_fill_2 FILLER_39_1635 ();
 sg13g2_decap_4 FILLER_39_1688 ();
 sg13g2_fill_1 FILLER_39_1692 ();
 sg13g2_decap_8 FILLER_39_1707 ();
 sg13g2_decap_4 FILLER_39_1714 ();
 sg13g2_decap_8 FILLER_39_1732 ();
 sg13g2_decap_8 FILLER_39_1765 ();
 sg13g2_fill_2 FILLER_39_1772 ();
 sg13g2_fill_1 FILLER_39_1774 ();
 sg13g2_decap_8 FILLER_39_1810 ();
 sg13g2_decap_8 FILLER_39_1817 ();
 sg13g2_fill_2 FILLER_39_1824 ();
 sg13g2_fill_1 FILLER_39_1826 ();
 sg13g2_fill_1 FILLER_39_1847 ();
 sg13g2_fill_2 FILLER_39_1867 ();
 sg13g2_fill_1 FILLER_39_1884 ();
 sg13g2_fill_2 FILLER_39_1890 ();
 sg13g2_fill_1 FILLER_39_1901 ();
 sg13g2_fill_1 FILLER_39_1907 ();
 sg13g2_fill_1 FILLER_39_1914 ();
 sg13g2_fill_1 FILLER_39_1938 ();
 sg13g2_fill_2 FILLER_39_1949 ();
 sg13g2_fill_2 FILLER_39_1964 ();
 sg13g2_fill_1 FILLER_39_1986 ();
 sg13g2_fill_1 FILLER_39_1999 ();
 sg13g2_fill_2 FILLER_39_2037 ();
 sg13g2_fill_1 FILLER_39_2100 ();
 sg13g2_fill_1 FILLER_39_2108 ();
 sg13g2_fill_2 FILLER_39_2143 ();
 sg13g2_decap_8 FILLER_39_2153 ();
 sg13g2_decap_8 FILLER_39_2160 ();
 sg13g2_fill_2 FILLER_39_2167 ();
 sg13g2_fill_2 FILLER_39_2211 ();
 sg13g2_fill_2 FILLER_39_2237 ();
 sg13g2_fill_2 FILLER_39_2266 ();
 sg13g2_fill_1 FILLER_39_2268 ();
 sg13g2_decap_8 FILLER_39_2321 ();
 sg13g2_decap_8 FILLER_39_2328 ();
 sg13g2_decap_8 FILLER_39_2345 ();
 sg13g2_decap_8 FILLER_39_2352 ();
 sg13g2_decap_8 FILLER_39_2359 ();
 sg13g2_decap_8 FILLER_39_2366 ();
 sg13g2_fill_2 FILLER_39_2373 ();
 sg13g2_fill_1 FILLER_39_2375 ();
 sg13g2_decap_8 FILLER_39_2380 ();
 sg13g2_decap_8 FILLER_39_2402 ();
 sg13g2_fill_2 FILLER_39_2422 ();
 sg13g2_fill_2 FILLER_39_2441 ();
 sg13g2_fill_1 FILLER_39_2449 ();
 sg13g2_decap_8 FILLER_39_2454 ();
 sg13g2_decap_4 FILLER_39_2461 ();
 sg13g2_fill_1 FILLER_39_2465 ();
 sg13g2_decap_8 FILLER_39_2470 ();
 sg13g2_decap_8 FILLER_39_2477 ();
 sg13g2_decap_8 FILLER_39_2484 ();
 sg13g2_decap_8 FILLER_39_2491 ();
 sg13g2_decap_8 FILLER_39_2498 ();
 sg13g2_decap_8 FILLER_39_2505 ();
 sg13g2_decap_4 FILLER_39_2512 ();
 sg13g2_fill_2 FILLER_39_2516 ();
 sg13g2_fill_2 FILLER_39_2530 ();
 sg13g2_fill_1 FILLER_39_2532 ();
 sg13g2_fill_2 FILLER_39_2542 ();
 sg13g2_fill_2 FILLER_39_2549 ();
 sg13g2_decap_4 FILLER_39_2583 ();
 sg13g2_fill_1 FILLER_39_2601 ();
 sg13g2_decap_8 FILLER_39_2606 ();
 sg13g2_decap_8 FILLER_39_2613 ();
 sg13g2_decap_8 FILLER_39_2620 ();
 sg13g2_decap_4 FILLER_39_2627 ();
 sg13g2_fill_1 FILLER_39_2631 ();
 sg13g2_fill_2 FILLER_39_2668 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_7 ();
 sg13g2_fill_1 FILLER_40_9 ();
 sg13g2_fill_1 FILLER_40_14 ();
 sg13g2_fill_2 FILLER_40_41 ();
 sg13g2_fill_2 FILLER_40_69 ();
 sg13g2_fill_1 FILLER_40_71 ();
 sg13g2_fill_2 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_decap_8 FILLER_40_96 ();
 sg13g2_fill_2 FILLER_40_103 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_fill_2 FILLER_40_119 ();
 sg13g2_decap_4 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_192 ();
 sg13g2_decap_4 FILLER_40_198 ();
 sg13g2_fill_1 FILLER_40_202 ();
 sg13g2_decap_8 FILLER_40_239 ();
 sg13g2_fill_1 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_268 ();
 sg13g2_fill_1 FILLER_40_274 ();
 sg13g2_fill_2 FILLER_40_285 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_fill_1 FILLER_40_324 ();
 sg13g2_fill_1 FILLER_40_360 ();
 sg13g2_fill_1 FILLER_40_396 ();
 sg13g2_fill_2 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_403 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_fill_1 FILLER_40_499 ();
 sg13g2_decap_8 FILLER_40_537 ();
 sg13g2_decap_4 FILLER_40_544 ();
 sg13g2_fill_1 FILLER_40_548 ();
 sg13g2_decap_4 FILLER_40_554 ();
 sg13g2_decap_4 FILLER_40_563 ();
 sg13g2_fill_2 FILLER_40_567 ();
 sg13g2_fill_1 FILLER_40_573 ();
 sg13g2_fill_1 FILLER_40_592 ();
 sg13g2_fill_2 FILLER_40_615 ();
 sg13g2_fill_1 FILLER_40_621 ();
 sg13g2_decap_4 FILLER_40_625 ();
 sg13g2_fill_2 FILLER_40_629 ();
 sg13g2_decap_8 FILLER_40_642 ();
 sg13g2_fill_1 FILLER_40_649 ();
 sg13g2_fill_2 FILLER_40_654 ();
 sg13g2_fill_1 FILLER_40_661 ();
 sg13g2_fill_1 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_678 ();
 sg13g2_decap_4 FILLER_40_685 ();
 sg13g2_fill_1 FILLER_40_705 ();
 sg13g2_fill_1 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_731 ();
 sg13g2_decap_8 FILLER_40_738 ();
 sg13g2_decap_8 FILLER_40_745 ();
 sg13g2_fill_1 FILLER_40_752 ();
 sg13g2_fill_1 FILLER_40_791 ();
 sg13g2_decap_4 FILLER_40_828 ();
 sg13g2_fill_1 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_874 ();
 sg13g2_fill_2 FILLER_40_881 ();
 sg13g2_fill_1 FILLER_40_883 ();
 sg13g2_decap_8 FILLER_40_908 ();
 sg13g2_decap_8 FILLER_40_915 ();
 sg13g2_decap_8 FILLER_40_922 ();
 sg13g2_decap_4 FILLER_40_929 ();
 sg13g2_fill_1 FILLER_40_933 ();
 sg13g2_fill_2 FILLER_40_992 ();
 sg13g2_decap_4 FILLER_40_1094 ();
 sg13g2_fill_2 FILLER_40_1103 ();
 sg13g2_fill_1 FILLER_40_1105 ();
 sg13g2_fill_2 FILLER_40_1136 ();
 sg13g2_fill_1 FILLER_40_1138 ();
 sg13g2_decap_8 FILLER_40_1152 ();
 sg13g2_decap_4 FILLER_40_1159 ();
 sg13g2_fill_1 FILLER_40_1163 ();
 sg13g2_fill_1 FILLER_40_1168 ();
 sg13g2_fill_1 FILLER_40_1178 ();
 sg13g2_decap_8 FILLER_40_1183 ();
 sg13g2_decap_8 FILLER_40_1190 ();
 sg13g2_decap_4 FILLER_40_1197 ();
 sg13g2_fill_2 FILLER_40_1201 ();
 sg13g2_decap_4 FILLER_40_1215 ();
 sg13g2_fill_2 FILLER_40_1219 ();
 sg13g2_decap_8 FILLER_40_1247 ();
 sg13g2_decap_8 FILLER_40_1254 ();
 sg13g2_decap_4 FILLER_40_1261 ();
 sg13g2_fill_2 FILLER_40_1265 ();
 sg13g2_decap_8 FILLER_40_1271 ();
 sg13g2_fill_2 FILLER_40_1278 ();
 sg13g2_fill_2 FILLER_40_1284 ();
 sg13g2_decap_4 FILLER_40_1296 ();
 sg13g2_fill_1 FILLER_40_1300 ();
 sg13g2_decap_8 FILLER_40_1305 ();
 sg13g2_fill_1 FILLER_40_1312 ();
 sg13g2_fill_1 FILLER_40_1317 ();
 sg13g2_decap_8 FILLER_40_1384 ();
 sg13g2_fill_1 FILLER_40_1397 ();
 sg13g2_fill_2 FILLER_40_1434 ();
 sg13g2_fill_1 FILLER_40_1446 ();
 sg13g2_fill_1 FILLER_40_1464 ();
 sg13g2_decap_8 FILLER_40_1469 ();
 sg13g2_fill_1 FILLER_40_1485 ();
 sg13g2_fill_1 FILLER_40_1494 ();
 sg13g2_decap_8 FILLER_40_1500 ();
 sg13g2_fill_2 FILLER_40_1507 ();
 sg13g2_fill_1 FILLER_40_1509 ();
 sg13g2_fill_2 FILLER_40_1534 ();
 sg13g2_fill_1 FILLER_40_1536 ();
 sg13g2_decap_4 FILLER_40_1541 ();
 sg13g2_fill_2 FILLER_40_1545 ();
 sg13g2_decap_8 FILLER_40_1551 ();
 sg13g2_decap_8 FILLER_40_1558 ();
 sg13g2_decap_4 FILLER_40_1565 ();
 sg13g2_fill_1 FILLER_40_1569 ();
 sg13g2_fill_1 FILLER_40_1592 ();
 sg13g2_decap_8 FILLER_40_1598 ();
 sg13g2_decap_8 FILLER_40_1605 ();
 sg13g2_decap_8 FILLER_40_1612 ();
 sg13g2_decap_8 FILLER_40_1619 ();
 sg13g2_decap_4 FILLER_40_1626 ();
 sg13g2_fill_2 FILLER_40_1652 ();
 sg13g2_decap_4 FILLER_40_1658 ();
 sg13g2_fill_2 FILLER_40_1666 ();
 sg13g2_decap_8 FILLER_40_1672 ();
 sg13g2_fill_2 FILLER_40_1679 ();
 sg13g2_fill_1 FILLER_40_1681 ();
 sg13g2_decap_4 FILLER_40_1686 ();
 sg13g2_decap_4 FILLER_40_1742 ();
 sg13g2_fill_1 FILLER_40_1746 ();
 sg13g2_decap_8 FILLER_40_1777 ();
 sg13g2_decap_4 FILLER_40_1784 ();
 sg13g2_fill_1 FILLER_40_1788 ();
 sg13g2_fill_2 FILLER_40_1793 ();
 sg13g2_fill_1 FILLER_40_1795 ();
 sg13g2_fill_1 FILLER_40_1808 ();
 sg13g2_decap_8 FILLER_40_1813 ();
 sg13g2_decap_8 FILLER_40_1820 ();
 sg13g2_decap_4 FILLER_40_1827 ();
 sg13g2_fill_2 FILLER_40_1831 ();
 sg13g2_fill_1 FILLER_40_1857 ();
 sg13g2_decap_4 FILLER_40_1863 ();
 sg13g2_fill_2 FILLER_40_1870 ();
 sg13g2_fill_2 FILLER_40_1897 ();
 sg13g2_fill_1 FILLER_40_1899 ();
 sg13g2_fill_1 FILLER_40_1910 ();
 sg13g2_fill_1 FILLER_40_1918 ();
 sg13g2_fill_1 FILLER_40_1933 ();
 sg13g2_fill_1 FILLER_40_1937 ();
 sg13g2_fill_1 FILLER_40_1973 ();
 sg13g2_fill_1 FILLER_40_1986 ();
 sg13g2_fill_2 FILLER_40_1995 ();
 sg13g2_decap_4 FILLER_40_2001 ();
 sg13g2_decap_4 FILLER_40_2009 ();
 sg13g2_fill_1 FILLER_40_2013 ();
 sg13g2_fill_2 FILLER_40_2026 ();
 sg13g2_fill_2 FILLER_40_2054 ();
 sg13g2_fill_1 FILLER_40_2062 ();
 sg13g2_fill_1 FILLER_40_2105 ();
 sg13g2_fill_1 FILLER_40_2145 ();
 sg13g2_decap_8 FILLER_40_2172 ();
 sg13g2_decap_8 FILLER_40_2179 ();
 sg13g2_decap_4 FILLER_40_2186 ();
 sg13g2_decap_4 FILLER_40_2204 ();
 sg13g2_decap_4 FILLER_40_2298 ();
 sg13g2_fill_1 FILLER_40_2302 ();
 sg13g2_decap_8 FILLER_40_2307 ();
 sg13g2_decap_4 FILLER_40_2314 ();
 sg13g2_decap_8 FILLER_40_2373 ();
 sg13g2_fill_2 FILLER_40_2380 ();
 sg13g2_fill_1 FILLER_40_2382 ();
 sg13g2_decap_4 FILLER_40_2387 ();
 sg13g2_fill_1 FILLER_40_2445 ();
 sg13g2_fill_2 FILLER_40_2492 ();
 sg13g2_decap_8 FILLER_40_2503 ();
 sg13g2_decap_8 FILLER_40_2510 ();
 sg13g2_fill_1 FILLER_40_2535 ();
 sg13g2_fill_1 FILLER_40_2584 ();
 sg13g2_decap_8 FILLER_40_2621 ();
 sg13g2_fill_2 FILLER_40_2628 ();
 sg13g2_fill_1 FILLER_40_2630 ();
 sg13g2_fill_2 FILLER_40_2667 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_43 ();
 sg13g2_fill_1 FILLER_41_60 ();
 sg13g2_decap_8 FILLER_41_107 ();
 sg13g2_decap_4 FILLER_41_114 ();
 sg13g2_decap_4 FILLER_41_131 ();
 sg13g2_decap_8 FILLER_41_143 ();
 sg13g2_fill_2 FILLER_41_150 ();
 sg13g2_fill_1 FILLER_41_156 ();
 sg13g2_fill_1 FILLER_41_183 ();
 sg13g2_decap_8 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_decap_8 FILLER_41_219 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_decap_8 FILLER_41_232 ();
 sg13g2_decap_8 FILLER_41_239 ();
 sg13g2_fill_2 FILLER_41_246 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_fill_1 FILLER_41_261 ();
 sg13g2_decap_4 FILLER_41_267 ();
 sg13g2_fill_2 FILLER_41_271 ();
 sg13g2_decap_4 FILLER_41_277 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_decap_4 FILLER_41_287 ();
 sg13g2_decap_4 FILLER_41_300 ();
 sg13g2_decap_4 FILLER_41_308 ();
 sg13g2_fill_1 FILLER_41_312 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_decap_4 FILLER_41_349 ();
 sg13g2_fill_1 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_41_393 ();
 sg13g2_decap_4 FILLER_41_400 ();
 sg13g2_fill_1 FILLER_41_404 ();
 sg13g2_decap_8 FILLER_41_409 ();
 sg13g2_decap_8 FILLER_41_416 ();
 sg13g2_decap_8 FILLER_41_423 ();
 sg13g2_fill_2 FILLER_41_430 ();
 sg13g2_fill_1 FILLER_41_441 ();
 sg13g2_fill_2 FILLER_41_494 ();
 sg13g2_fill_1 FILLER_41_496 ();
 sg13g2_fill_2 FILLER_41_533 ();
 sg13g2_decap_4 FILLER_41_554 ();
 sg13g2_decap_4 FILLER_41_563 ();
 sg13g2_fill_2 FILLER_41_567 ();
 sg13g2_fill_1 FILLER_41_579 ();
 sg13g2_decap_4 FILLER_41_586 ();
 sg13g2_fill_1 FILLER_41_599 ();
 sg13g2_fill_2 FILLER_41_608 ();
 sg13g2_fill_1 FILLER_41_610 ();
 sg13g2_decap_4 FILLER_41_635 ();
 sg13g2_fill_1 FILLER_41_650 ();
 sg13g2_fill_1 FILLER_41_657 ();
 sg13g2_fill_1 FILLER_41_662 ();
 sg13g2_decap_4 FILLER_41_668 ();
 sg13g2_fill_2 FILLER_41_676 ();
 sg13g2_decap_8 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_689 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_4 FILLER_41_700 ();
 sg13g2_decap_4 FILLER_41_708 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_decap_8 FILLER_41_717 ();
 sg13g2_decap_4 FILLER_41_724 ();
 sg13g2_fill_1 FILLER_41_728 ();
 sg13g2_fill_2 FILLER_41_733 ();
 sg13g2_fill_1 FILLER_41_735 ();
 sg13g2_fill_1 FILLER_41_762 ();
 sg13g2_fill_1 FILLER_41_784 ();
 sg13g2_fill_2 FILLER_41_815 ();
 sg13g2_decap_4 FILLER_41_825 ();
 sg13g2_fill_2 FILLER_41_829 ();
 sg13g2_fill_1 FILLER_41_848 ();
 sg13g2_fill_2 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_881 ();
 sg13g2_fill_1 FILLER_41_883 ();
 sg13g2_fill_2 FILLER_41_914 ();
 sg13g2_decap_8 FILLER_41_926 ();
 sg13g2_decap_8 FILLER_41_933 ();
 sg13g2_decap_8 FILLER_41_940 ();
 sg13g2_decap_8 FILLER_41_947 ();
 sg13g2_decap_8 FILLER_41_954 ();
 sg13g2_fill_2 FILLER_41_961 ();
 sg13g2_fill_1 FILLER_41_963 ();
 sg13g2_fill_1 FILLER_41_1016 ();
 sg13g2_decap_4 FILLER_41_1026 ();
 sg13g2_fill_2 FILLER_41_1030 ();
 sg13g2_fill_2 FILLER_41_1068 ();
 sg13g2_fill_1 FILLER_41_1070 ();
 sg13g2_fill_1 FILLER_41_1075 ();
 sg13g2_fill_1 FILLER_41_1102 ();
 sg13g2_fill_1 FILLER_41_1107 ();
 sg13g2_fill_1 FILLER_41_1113 ();
 sg13g2_fill_1 FILLER_41_1122 ();
 sg13g2_fill_2 FILLER_41_1128 ();
 sg13g2_fill_1 FILLER_41_1130 ();
 sg13g2_fill_1 FILLER_41_1136 ();
 sg13g2_decap_4 FILLER_41_1158 ();
 sg13g2_fill_1 FILLER_41_1167 ();
 sg13g2_decap_8 FILLER_41_1172 ();
 sg13g2_fill_2 FILLER_41_1179 ();
 sg13g2_fill_1 FILLER_41_1181 ();
 sg13g2_decap_8 FILLER_41_1187 ();
 sg13g2_fill_1 FILLER_41_1194 ();
 sg13g2_fill_2 FILLER_41_1208 ();
 sg13g2_fill_1 FILLER_41_1210 ();
 sg13g2_decap_4 FILLER_41_1221 ();
 sg13g2_fill_1 FILLER_41_1225 ();
 sg13g2_fill_2 FILLER_41_1266 ();
 sg13g2_decap_8 FILLER_41_1304 ();
 sg13g2_decap_4 FILLER_41_1311 ();
 sg13g2_fill_1 FILLER_41_1315 ();
 sg13g2_decap_4 FILLER_41_1326 ();
 sg13g2_fill_2 FILLER_41_1330 ();
 sg13g2_decap_4 FILLER_41_1343 ();
 sg13g2_fill_1 FILLER_41_1347 ();
 sg13g2_decap_8 FILLER_41_1398 ();
 sg13g2_decap_4 FILLER_41_1405 ();
 sg13g2_fill_1 FILLER_41_1409 ();
 sg13g2_fill_2 FILLER_41_1415 ();
 sg13g2_decap_8 FILLER_41_1423 ();
 sg13g2_fill_2 FILLER_41_1430 ();
 sg13g2_fill_2 FILLER_41_1437 ();
 sg13g2_fill_2 FILLER_41_1443 ();
 sg13g2_fill_1 FILLER_41_1445 ();
 sg13g2_fill_2 FILLER_41_1449 ();
 sg13g2_fill_1 FILLER_41_1462 ();
 sg13g2_decap_8 FILLER_41_1511 ();
 sg13g2_fill_2 FILLER_41_1518 ();
 sg13g2_fill_1 FILLER_41_1520 ();
 sg13g2_decap_4 FILLER_41_1533 ();
 sg13g2_fill_2 FILLER_41_1537 ();
 sg13g2_fill_1 FILLER_41_1543 ();
 sg13g2_decap_8 FILLER_41_1549 ();
 sg13g2_decap_8 FILLER_41_1556 ();
 sg13g2_decap_8 FILLER_41_1563 ();
 sg13g2_fill_2 FILLER_41_1580 ();
 sg13g2_fill_1 FILLER_41_1594 ();
 sg13g2_decap_8 FILLER_41_1598 ();
 sg13g2_decap_8 FILLER_41_1605 ();
 sg13g2_decap_8 FILLER_41_1612 ();
 sg13g2_decap_8 FILLER_41_1619 ();
 sg13g2_fill_2 FILLER_41_1626 ();
 sg13g2_decap_8 FILLER_41_1633 ();
 sg13g2_decap_8 FILLER_41_1640 ();
 sg13g2_decap_8 FILLER_41_1673 ();
 sg13g2_decap_4 FILLER_41_1680 ();
 sg13g2_fill_1 FILLER_41_1684 ();
 sg13g2_decap_4 FILLER_41_1691 ();
 sg13g2_fill_2 FILLER_41_1695 ();
 sg13g2_decap_8 FILLER_41_1701 ();
 sg13g2_decap_8 FILLER_41_1708 ();
 sg13g2_decap_4 FILLER_41_1715 ();
 sg13g2_decap_8 FILLER_41_1729 ();
 sg13g2_fill_2 FILLER_41_1736 ();
 sg13g2_decap_8 FILLER_41_1747 ();
 sg13g2_fill_1 FILLER_41_1754 ();
 sg13g2_decap_4 FILLER_41_1769 ();
 sg13g2_fill_1 FILLER_41_1773 ();
 sg13g2_decap_4 FILLER_41_1824 ();
 sg13g2_fill_1 FILLER_41_1834 ();
 sg13g2_fill_1 FILLER_41_1860 ();
 sg13g2_fill_2 FILLER_41_1868 ();
 sg13g2_fill_2 FILLER_41_1875 ();
 sg13g2_fill_2 FILLER_41_1882 ();
 sg13g2_fill_1 FILLER_41_1884 ();
 sg13g2_fill_1 FILLER_41_1894 ();
 sg13g2_fill_1 FILLER_41_1906 ();
 sg13g2_fill_1 FILLER_41_1912 ();
 sg13g2_fill_1 FILLER_41_1933 ();
 sg13g2_fill_2 FILLER_41_1939 ();
 sg13g2_fill_1 FILLER_41_1946 ();
 sg13g2_fill_1 FILLER_41_1952 ();
 sg13g2_fill_2 FILLER_41_1961 ();
 sg13g2_fill_1 FILLER_41_1963 ();
 sg13g2_fill_1 FILLER_41_1968 ();
 sg13g2_fill_2 FILLER_41_1974 ();
 sg13g2_fill_2 FILLER_41_1981 ();
 sg13g2_fill_1 FILLER_41_1983 ();
 sg13g2_decap_8 FILLER_41_1996 ();
 sg13g2_decap_8 FILLER_41_2003 ();
 sg13g2_decap_4 FILLER_41_2010 ();
 sg13g2_fill_1 FILLER_41_2014 ();
 sg13g2_decap_8 FILLER_41_2028 ();
 sg13g2_decap_4 FILLER_41_2035 ();
 sg13g2_fill_2 FILLER_41_2039 ();
 sg13g2_decap_8 FILLER_41_2045 ();
 sg13g2_fill_1 FILLER_41_2052 ();
 sg13g2_fill_1 FILLER_41_2101 ();
 sg13g2_fill_1 FILLER_41_2164 ();
 sg13g2_fill_2 FILLER_41_2179 ();
 sg13g2_fill_1 FILLER_41_2181 ();
 sg13g2_fill_2 FILLER_41_2187 ();
 sg13g2_fill_1 FILLER_41_2189 ();
 sg13g2_decap_4 FILLER_41_2251 ();
 sg13g2_decap_8 FILLER_41_2301 ();
 sg13g2_fill_1 FILLER_41_2308 ();
 sg13g2_fill_2 FILLER_41_2335 ();
 sg13g2_decap_4 FILLER_41_2363 ();
 sg13g2_fill_2 FILLER_41_2393 ();
 sg13g2_decap_4 FILLER_41_2421 ();
 sg13g2_decap_8 FILLER_41_2429 ();
 sg13g2_decap_8 FILLER_41_2436 ();
 sg13g2_decap_4 FILLER_41_2443 ();
 sg13g2_fill_2 FILLER_41_2447 ();
 sg13g2_fill_2 FILLER_41_2464 ();
 sg13g2_decap_4 FILLER_41_2523 ();
 sg13g2_fill_1 FILLER_41_2535 ();
 sg13g2_fill_1 FILLER_41_2590 ();
 sg13g2_fill_2 FILLER_41_2667 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_fill_2 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_37 ();
 sg13g2_decap_4 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_72 ();
 sg13g2_decap_8 FILLER_42_83 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_fill_1 FILLER_42_92 ();
 sg13g2_fill_1 FILLER_42_103 ();
 sg13g2_decap_4 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_124 ();
 sg13g2_decap_4 FILLER_42_131 ();
 sg13g2_fill_2 FILLER_42_143 ();
 sg13g2_decap_8 FILLER_42_209 ();
 sg13g2_decap_4 FILLER_42_216 ();
 sg13g2_fill_1 FILLER_42_220 ();
 sg13g2_fill_2 FILLER_42_234 ();
 sg13g2_fill_1 FILLER_42_236 ();
 sg13g2_fill_1 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_295 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_8 FILLER_42_330 ();
 sg13g2_decap_8 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_351 ();
 sg13g2_decap_8 FILLER_42_358 ();
 sg13g2_fill_2 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_fill_1 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_388 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_1 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_424 ();
 sg13g2_fill_1 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_decap_8 FILLER_42_440 ();
 sg13g2_fill_1 FILLER_42_447 ();
 sg13g2_fill_2 FILLER_42_461 ();
 sg13g2_fill_1 FILLER_42_463 ();
 sg13g2_fill_1 FILLER_42_468 ();
 sg13g2_decap_8 FILLER_42_482 ();
 sg13g2_decap_4 FILLER_42_489 ();
 sg13g2_fill_1 FILLER_42_493 ();
 sg13g2_fill_2 FILLER_42_511 ();
 sg13g2_fill_1 FILLER_42_523 ();
 sg13g2_decap_8 FILLER_42_529 ();
 sg13g2_decap_4 FILLER_42_536 ();
 sg13g2_decap_8 FILLER_42_550 ();
 sg13g2_fill_2 FILLER_42_557 ();
 sg13g2_fill_1 FILLER_42_564 ();
 sg13g2_fill_2 FILLER_42_590 ();
 sg13g2_fill_2 FILLER_42_604 ();
 sg13g2_fill_1 FILLER_42_642 ();
 sg13g2_decap_4 FILLER_42_677 ();
 sg13g2_fill_2 FILLER_42_702 ();
 sg13g2_fill_2 FILLER_42_728 ();
 sg13g2_fill_1 FILLER_42_769 ();
 sg13g2_decap_4 FILLER_42_775 ();
 sg13g2_fill_2 FILLER_42_799 ();
 sg13g2_decap_8 FILLER_42_815 ();
 sg13g2_decap_4 FILLER_42_822 ();
 sg13g2_fill_1 FILLER_42_826 ();
 sg13g2_fill_2 FILLER_42_835 ();
 sg13g2_fill_2 FILLER_42_946 ();
 sg13g2_fill_1 FILLER_42_948 ();
 sg13g2_decap_8 FILLER_42_953 ();
 sg13g2_fill_2 FILLER_42_960 ();
 sg13g2_fill_1 FILLER_42_962 ();
 sg13g2_fill_1 FILLER_42_993 ();
 sg13g2_decap_8 FILLER_42_1004 ();
 sg13g2_decap_8 FILLER_42_1011 ();
 sg13g2_fill_2 FILLER_42_1018 ();
 sg13g2_fill_1 FILLER_42_1020 ();
 sg13g2_decap_8 FILLER_42_1030 ();
 sg13g2_fill_1 FILLER_42_1041 ();
 sg13g2_fill_2 FILLER_42_1084 ();
 sg13g2_fill_1 FILLER_42_1147 ();
 sg13g2_decap_8 FILLER_42_1152 ();
 sg13g2_fill_2 FILLER_42_1194 ();
 sg13g2_fill_1 FILLER_42_1200 ();
 sg13g2_fill_1 FILLER_42_1222 ();
 sg13g2_fill_2 FILLER_42_1233 ();
 sg13g2_decap_8 FILLER_42_1256 ();
 sg13g2_decap_8 FILLER_42_1263 ();
 sg13g2_fill_2 FILLER_42_1270 ();
 sg13g2_fill_1 FILLER_42_1272 ();
 sg13g2_fill_2 FILLER_42_1303 ();
 sg13g2_fill_1 FILLER_42_1305 ();
 sg13g2_decap_4 FILLER_42_1372 ();
 sg13g2_decap_8 FILLER_42_1402 ();
 sg13g2_decap_8 FILLER_42_1409 ();
 sg13g2_fill_1 FILLER_42_1416 ();
 sg13g2_decap_8 FILLER_42_1422 ();
 sg13g2_decap_4 FILLER_42_1429 ();
 sg13g2_fill_2 FILLER_42_1449 ();
 sg13g2_decap_8 FILLER_42_1461 ();
 sg13g2_fill_2 FILLER_42_1468 ();
 sg13g2_decap_4 FILLER_42_1485 ();
 sg13g2_fill_2 FILLER_42_1489 ();
 sg13g2_fill_2 FILLER_42_1496 ();
 sg13g2_fill_2 FILLER_42_1507 ();
 sg13g2_fill_1 FILLER_42_1509 ();
 sg13g2_fill_2 FILLER_42_1542 ();
 sg13g2_decap_4 FILLER_42_1631 ();
 sg13g2_fill_2 FILLER_42_1635 ();
 sg13g2_fill_2 FILLER_42_1677 ();
 sg13g2_fill_1 FILLER_42_1679 ();
 sg13g2_decap_8 FILLER_42_1683 ();
 sg13g2_decap_8 FILLER_42_1690 ();
 sg13g2_decap_8 FILLER_42_1763 ();
 sg13g2_decap_4 FILLER_42_1770 ();
 sg13g2_fill_2 FILLER_42_1774 ();
 sg13g2_fill_2 FILLER_42_1839 ();
 sg13g2_decap_4 FILLER_42_1846 ();
 sg13g2_fill_2 FILLER_42_1850 ();
 sg13g2_fill_2 FILLER_42_1861 ();
 sg13g2_fill_2 FILLER_42_1869 ();
 sg13g2_decap_8 FILLER_42_1878 ();
 sg13g2_decap_4 FILLER_42_1885 ();
 sg13g2_fill_1 FILLER_42_1889 ();
 sg13g2_fill_1 FILLER_42_1898 ();
 sg13g2_decap_4 FILLER_42_1903 ();
 sg13g2_fill_2 FILLER_42_1922 ();
 sg13g2_fill_2 FILLER_42_1930 ();
 sg13g2_fill_2 FILLER_42_1937 ();
 sg13g2_fill_2 FILLER_42_1944 ();
 sg13g2_fill_2 FILLER_42_1961 ();
 sg13g2_fill_1 FILLER_42_1963 ();
 sg13g2_fill_2 FILLER_42_1973 ();
 sg13g2_fill_1 FILLER_42_1975 ();
 sg13g2_decap_4 FILLER_42_1986 ();
 sg13g2_decap_8 FILLER_42_2007 ();
 sg13g2_decap_4 FILLER_42_2014 ();
 sg13g2_decap_4 FILLER_42_2071 ();
 sg13g2_fill_2 FILLER_42_2075 ();
 sg13g2_fill_2 FILLER_42_2138 ();
 sg13g2_fill_2 FILLER_42_2161 ();
 sg13g2_fill_1 FILLER_42_2163 ();
 sg13g2_fill_1 FILLER_42_2190 ();
 sg13g2_decap_4 FILLER_42_2195 ();
 sg13g2_fill_2 FILLER_42_2199 ();
 sg13g2_fill_1 FILLER_42_2227 ();
 sg13g2_decap_8 FILLER_42_2232 ();
 sg13g2_decap_4 FILLER_42_2239 ();
 sg13g2_fill_2 FILLER_42_2243 ();
 sg13g2_decap_8 FILLER_42_2249 ();
 sg13g2_decap_8 FILLER_42_2256 ();
 sg13g2_decap_8 FILLER_42_2263 ();
 sg13g2_decap_4 FILLER_42_2270 ();
 sg13g2_decap_8 FILLER_42_2278 ();
 sg13g2_fill_2 FILLER_42_2285 ();
 sg13g2_fill_1 FILLER_42_2287 ();
 sg13g2_decap_8 FILLER_42_2300 ();
 sg13g2_decap_8 FILLER_42_2307 ();
 sg13g2_fill_1 FILLER_42_2343 ();
 sg13g2_fill_1 FILLER_42_2362 ();
 sg13g2_decap_4 FILLER_42_2368 ();
 sg13g2_fill_1 FILLER_42_2386 ();
 sg13g2_fill_2 FILLER_42_2397 ();
 sg13g2_fill_1 FILLER_42_2399 ();
 sg13g2_decap_8 FILLER_42_2409 ();
 sg13g2_fill_2 FILLER_42_2416 ();
 sg13g2_fill_1 FILLER_42_2418 ();
 sg13g2_decap_4 FILLER_42_2434 ();
 sg13g2_decap_8 FILLER_42_2473 ();
 sg13g2_fill_2 FILLER_42_2480 ();
 sg13g2_fill_1 FILLER_42_2529 ();
 sg13g2_fill_2 FILLER_42_2535 ();
 sg13g2_fill_1 FILLER_42_2543 ();
 sg13g2_fill_2 FILLER_42_2566 ();
 sg13g2_fill_1 FILLER_42_2590 ();
 sg13g2_fill_2 FILLER_42_2604 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_7 ();
 sg13g2_fill_1 FILLER_43_9 ();
 sg13g2_decap_4 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_23 ();
 sg13g2_fill_2 FILLER_43_43 ();
 sg13g2_fill_1 FILLER_43_55 ();
 sg13g2_fill_1 FILLER_43_82 ();
 sg13g2_fill_1 FILLER_43_135 ();
 sg13g2_fill_2 FILLER_43_144 ();
 sg13g2_fill_1 FILLER_43_146 ();
 sg13g2_fill_2 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_271 ();
 sg13g2_decap_4 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_281 ();
 sg13g2_fill_2 FILLER_43_296 ();
 sg13g2_fill_1 FILLER_43_298 ();
 sg13g2_fill_1 FILLER_43_330 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_4 FILLER_43_369 ();
 sg13g2_fill_2 FILLER_43_373 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_4 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_394 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_2 FILLER_43_444 ();
 sg13g2_fill_1 FILLER_43_446 ();
 sg13g2_decap_8 FILLER_43_451 ();
 sg13g2_decap_8 FILLER_43_458 ();
 sg13g2_decap_8 FILLER_43_465 ();
 sg13g2_decap_8 FILLER_43_472 ();
 sg13g2_decap_8 FILLER_43_479 ();
 sg13g2_fill_1 FILLER_43_486 ();
 sg13g2_decap_4 FILLER_43_491 ();
 sg13g2_fill_2 FILLER_43_495 ();
 sg13g2_decap_8 FILLER_43_500 ();
 sg13g2_decap_4 FILLER_43_507 ();
 sg13g2_fill_1 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_516 ();
 sg13g2_decap_8 FILLER_43_523 ();
 sg13g2_fill_2 FILLER_43_530 ();
 sg13g2_fill_1 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_548 ();
 sg13g2_fill_1 FILLER_43_555 ();
 sg13g2_fill_1 FILLER_43_566 ();
 sg13g2_fill_2 FILLER_43_571 ();
 sg13g2_fill_1 FILLER_43_595 ();
 sg13g2_fill_1 FILLER_43_610 ();
 sg13g2_fill_1 FILLER_43_616 ();
 sg13g2_fill_1 FILLER_43_629 ();
 sg13g2_fill_1 FILLER_43_651 ();
 sg13g2_fill_2 FILLER_43_657 ();
 sg13g2_fill_2 FILLER_43_663 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_decap_4 FILLER_43_677 ();
 sg13g2_decap_4 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_694 ();
 sg13g2_decap_4 FILLER_43_732 ();
 sg13g2_fill_1 FILLER_43_742 ();
 sg13g2_fill_1 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_764 ();
 sg13g2_decap_8 FILLER_43_771 ();
 sg13g2_decap_8 FILLER_43_778 ();
 sg13g2_decap_4 FILLER_43_793 ();
 sg13g2_fill_1 FILLER_43_797 ();
 sg13g2_fill_1 FILLER_43_808 ();
 sg13g2_decap_4 FILLER_43_817 ();
 sg13g2_fill_2 FILLER_43_821 ();
 sg13g2_fill_1 FILLER_43_827 ();
 sg13g2_fill_2 FILLER_43_845 ();
 sg13g2_fill_2 FILLER_43_851 ();
 sg13g2_fill_1 FILLER_43_863 ();
 sg13g2_decap_4 FILLER_43_872 ();
 sg13g2_fill_2 FILLER_43_876 ();
 sg13g2_fill_1 FILLER_43_881 ();
 sg13g2_decap_4 FILLER_43_890 ();
 sg13g2_fill_2 FILLER_43_925 ();
 sg13g2_fill_2 FILLER_43_931 ();
 sg13g2_decap_4 FILLER_43_969 ();
 sg13g2_fill_1 FILLER_43_973 ();
 sg13g2_decap_4 FILLER_43_1000 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_fill_1 FILLER_43_1029 ();
 sg13g2_decap_8 FILLER_43_1060 ();
 sg13g2_fill_1 FILLER_43_1067 ();
 sg13g2_fill_2 FILLER_43_1077 ();
 sg13g2_decap_4 FILLER_43_1118 ();
 sg13g2_decap_4 FILLER_43_1130 ();
 sg13g2_fill_1 FILLER_43_1155 ();
 sg13g2_fill_2 FILLER_43_1238 ();
 sg13g2_decap_8 FILLER_43_1266 ();
 sg13g2_decap_8 FILLER_43_1273 ();
 sg13g2_decap_4 FILLER_43_1294 ();
 sg13g2_decap_4 FILLER_43_1354 ();
 sg13g2_decap_8 FILLER_43_1368 ();
 sg13g2_decap_8 FILLER_43_1375 ();
 sg13g2_fill_2 FILLER_43_1382 ();
 sg13g2_fill_1 FILLER_43_1384 ();
 sg13g2_fill_1 FILLER_43_1389 ();
 sg13g2_decap_8 FILLER_43_1406 ();
 sg13g2_fill_1 FILLER_43_1443 ();
 sg13g2_fill_2 FILLER_43_1514 ();
 sg13g2_fill_1 FILLER_43_1521 ();
 sg13g2_fill_1 FILLER_43_1527 ();
 sg13g2_fill_2 FILLER_43_1541 ();
 sg13g2_fill_1 FILLER_43_1580 ();
 sg13g2_fill_1 FILLER_43_1590 ();
 sg13g2_fill_1 FILLER_43_1627 ();
 sg13g2_decap_4 FILLER_43_1654 ();
 sg13g2_fill_2 FILLER_43_1658 ();
 sg13g2_decap_8 FILLER_43_1664 ();
 sg13g2_decap_8 FILLER_43_1671 ();
 sg13g2_decap_8 FILLER_43_1678 ();
 sg13g2_decap_8 FILLER_43_1685 ();
 sg13g2_fill_1 FILLER_43_1692 ();
 sg13g2_decap_8 FILLER_43_1698 ();
 sg13g2_fill_2 FILLER_43_1705 ();
 sg13g2_fill_1 FILLER_43_1707 ();
 sg13g2_fill_2 FILLER_43_1713 ();
 sg13g2_decap_8 FILLER_43_1724 ();
 sg13g2_fill_1 FILLER_43_1735 ();
 sg13g2_fill_1 FILLER_43_1766 ();
 sg13g2_fill_2 FILLER_43_1772 ();
 sg13g2_fill_1 FILLER_43_1784 ();
 sg13g2_fill_1 FILLER_43_1818 ();
 sg13g2_fill_2 FILLER_43_1829 ();
 sg13g2_decap_8 FILLER_43_1834 ();
 sg13g2_decap_4 FILLER_43_1841 ();
 sg13g2_fill_1 FILLER_43_1845 ();
 sg13g2_fill_1 FILLER_43_1896 ();
 sg13g2_fill_2 FILLER_43_1907 ();
 sg13g2_fill_1 FILLER_43_1909 ();
 sg13g2_fill_1 FILLER_43_1921 ();
 sg13g2_decap_4 FILLER_43_1927 ();
 sg13g2_fill_1 FILLER_43_1944 ();
 sg13g2_decap_8 FILLER_43_1950 ();
 sg13g2_fill_1 FILLER_43_1957 ();
 sg13g2_fill_1 FILLER_43_2000 ();
 sg13g2_fill_2 FILLER_43_2005 ();
 sg13g2_fill_2 FILLER_43_2033 ();
 sg13g2_fill_2 FILLER_43_2049 ();
 sg13g2_fill_1 FILLER_43_2051 ();
 sg13g2_fill_1 FILLER_43_2065 ();
 sg13g2_fill_1 FILLER_43_2092 ();
 sg13g2_fill_2 FILLER_43_2103 ();
 sg13g2_fill_2 FILLER_43_2139 ();
 sg13g2_decap_4 FILLER_43_2162 ();
 sg13g2_fill_1 FILLER_43_2170 ();
 sg13g2_fill_2 FILLER_43_2207 ();
 sg13g2_fill_1 FILLER_43_2209 ();
 sg13g2_decap_8 FILLER_43_2214 ();
 sg13g2_decap_8 FILLER_43_2221 ();
 sg13g2_decap_8 FILLER_43_2228 ();
 sg13g2_fill_2 FILLER_43_2235 ();
 sg13g2_fill_2 FILLER_43_2245 ();
 sg13g2_fill_1 FILLER_43_2247 ();
 sg13g2_decap_4 FILLER_43_2281 ();
 sg13g2_decap_8 FILLER_43_2311 ();
 sg13g2_decap_8 FILLER_43_2318 ();
 sg13g2_fill_1 FILLER_43_2325 ();
 sg13g2_fill_2 FILLER_43_2330 ();
 sg13g2_fill_1 FILLER_43_2332 ();
 sg13g2_fill_2 FILLER_43_2337 ();
 sg13g2_fill_1 FILLER_43_2339 ();
 sg13g2_decap_4 FILLER_43_2370 ();
 sg13g2_fill_1 FILLER_43_2374 ();
 sg13g2_decap_4 FILLER_43_2381 ();
 sg13g2_fill_2 FILLER_43_2385 ();
 sg13g2_decap_4 FILLER_43_2413 ();
 sg13g2_fill_2 FILLER_43_2417 ();
 sg13g2_fill_1 FILLER_43_2481 ();
 sg13g2_fill_1 FILLER_43_2492 ();
 sg13g2_fill_2 FILLER_43_2499 ();
 sg13g2_fill_1 FILLER_43_2501 ();
 sg13g2_fill_2 FILLER_43_2631 ();
 sg13g2_decap_4 FILLER_43_2643 ();
 sg13g2_decap_8 FILLER_43_2651 ();
 sg13g2_decap_8 FILLER_43_2658 ();
 sg13g2_decap_4 FILLER_43_2665 ();
 sg13g2_fill_1 FILLER_43_2669 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_28 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_58 ();
 sg13g2_decap_8 FILLER_44_80 ();
 sg13g2_fill_2 FILLER_44_87 ();
 sg13g2_fill_2 FILLER_44_103 ();
 sg13g2_fill_1 FILLER_44_105 ();
 sg13g2_fill_2 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_144 ();
 sg13g2_decap_4 FILLER_44_151 ();
 sg13g2_fill_2 FILLER_44_155 ();
 sg13g2_fill_1 FILLER_44_205 ();
 sg13g2_fill_2 FILLER_44_216 ();
 sg13g2_fill_2 FILLER_44_222 ();
 sg13g2_fill_2 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_232 ();
 sg13g2_fill_2 FILLER_44_244 ();
 sg13g2_fill_1 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_251 ();
 sg13g2_fill_2 FILLER_44_260 ();
 sg13g2_fill_1 FILLER_44_266 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_287 ();
 sg13g2_fill_1 FILLER_44_309 ();
 sg13g2_decap_4 FILLER_44_314 ();
 sg13g2_fill_2 FILLER_44_318 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_fill_2 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_342 ();
 sg13g2_fill_2 FILLER_44_349 ();
 sg13g2_decap_4 FILLER_44_355 ();
 sg13g2_fill_1 FILLER_44_359 ();
 sg13g2_decap_4 FILLER_44_366 ();
 sg13g2_fill_1 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_4 FILLER_44_483 ();
 sg13g2_fill_2 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_493 ();
 sg13g2_decap_8 FILLER_44_500 ();
 sg13g2_decap_8 FILLER_44_507 ();
 sg13g2_fill_2 FILLER_44_514 ();
 sg13g2_fill_2 FILLER_44_533 ();
 sg13g2_fill_1 FILLER_44_535 ();
 sg13g2_fill_2 FILLER_44_540 ();
 sg13g2_fill_1 FILLER_44_542 ();
 sg13g2_decap_4 FILLER_44_557 ();
 sg13g2_fill_1 FILLER_44_567 ();
 sg13g2_fill_1 FILLER_44_620 ();
 sg13g2_fill_1 FILLER_44_624 ();
 sg13g2_decap_4 FILLER_44_643 ();
 sg13g2_fill_1 FILLER_44_647 ();
 sg13g2_fill_2 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_731 ();
 sg13g2_decap_4 FILLER_44_738 ();
 sg13g2_fill_1 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_755 ();
 sg13g2_fill_2 FILLER_44_775 ();
 sg13g2_decap_4 FILLER_44_787 ();
 sg13g2_fill_1 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_860 ();
 sg13g2_decap_4 FILLER_44_867 ();
 sg13g2_fill_1 FILLER_44_871 ();
 sg13g2_decap_4 FILLER_44_915 ();
 sg13g2_fill_1 FILLER_44_919 ();
 sg13g2_decap_8 FILLER_44_928 ();
 sg13g2_fill_2 FILLER_44_935 ();
 sg13g2_fill_1 FILLER_44_937 ();
 sg13g2_fill_2 FILLER_44_951 ();
 sg13g2_fill_1 FILLER_44_953 ();
 sg13g2_decap_4 FILLER_44_967 ();
 sg13g2_fill_2 FILLER_44_971 ();
 sg13g2_fill_1 FILLER_44_977 ();
 sg13g2_fill_1 FILLER_44_983 ();
 sg13g2_fill_1 FILLER_44_988 ();
 sg13g2_fill_2 FILLER_44_1015 ();
 sg13g2_decap_8 FILLER_44_1038 ();
 sg13g2_fill_2 FILLER_44_1045 ();
 sg13g2_decap_4 FILLER_44_1072 ();
 sg13g2_fill_1 FILLER_44_1076 ();
 sg13g2_decap_4 FILLER_44_1127 ();
 sg13g2_decap_4 FILLER_44_1217 ();
 sg13g2_decap_8 FILLER_44_1261 ();
 sg13g2_decap_8 FILLER_44_1268 ();
 sg13g2_decap_8 FILLER_44_1275 ();
 sg13g2_decap_8 FILLER_44_1282 ();
 sg13g2_decap_8 FILLER_44_1289 ();
 sg13g2_decap_8 FILLER_44_1296 ();
 sg13g2_decap_4 FILLER_44_1303 ();
 sg13g2_decap_4 FILLER_44_1311 ();
 sg13g2_decap_4 FILLER_44_1319 ();
 sg13g2_fill_2 FILLER_44_1327 ();
 sg13g2_decap_8 FILLER_44_1334 ();
 sg13g2_decap_4 FILLER_44_1341 ();
 sg13g2_fill_2 FILLER_44_1345 ();
 sg13g2_decap_4 FILLER_44_1366 ();
 sg13g2_fill_1 FILLER_44_1370 ();
 sg13g2_fill_2 FILLER_44_1381 ();
 sg13g2_fill_2 FILLER_44_1387 ();
 sg13g2_fill_2 FILLER_44_1428 ();
 sg13g2_fill_1 FILLER_44_1430 ();
 sg13g2_fill_1 FILLER_44_1450 ();
 sg13g2_fill_2 FILLER_44_1506 ();
 sg13g2_fill_1 FILLER_44_1512 ();
 sg13g2_decap_4 FILLER_44_1516 ();
 sg13g2_fill_1 FILLER_44_1524 ();
 sg13g2_fill_1 FILLER_44_1530 ();
 sg13g2_fill_1 FILLER_44_1557 ();
 sg13g2_fill_2 FILLER_44_1622 ();
 sg13g2_fill_1 FILLER_44_1624 ();
 sg13g2_decap_4 FILLER_44_1670 ();
 sg13g2_fill_1 FILLER_44_1674 ();
 sg13g2_decap_8 FILLER_44_1704 ();
 sg13g2_decap_8 FILLER_44_1711 ();
 sg13g2_fill_2 FILLER_44_1718 ();
 sg13g2_decap_8 FILLER_44_1730 ();
 sg13g2_fill_2 FILLER_44_1737 ();
 sg13g2_fill_1 FILLER_44_1749 ();
 sg13g2_decap_8 FILLER_44_1842 ();
 sg13g2_fill_2 FILLER_44_1849 ();
 sg13g2_fill_1 FILLER_44_1851 ();
 sg13g2_fill_1 FILLER_44_1862 ();
 sg13g2_fill_1 FILLER_44_1905 ();
 sg13g2_fill_1 FILLER_44_1924 ();
 sg13g2_fill_2 FILLER_44_1929 ();
 sg13g2_decap_4 FILLER_44_1934 ();
 sg13g2_fill_2 FILLER_44_1943 ();
 sg13g2_fill_1 FILLER_44_1996 ();
 sg13g2_decap_8 FILLER_44_2002 ();
 sg13g2_decap_4 FILLER_44_2009 ();
 sg13g2_fill_1 FILLER_44_2013 ();
 sg13g2_fill_2 FILLER_44_2022 ();
 sg13g2_decap_4 FILLER_44_2034 ();
 sg13g2_fill_1 FILLER_44_2038 ();
 sg13g2_fill_1 FILLER_44_2080 ();
 sg13g2_decap_4 FILLER_44_2098 ();
 sg13g2_fill_2 FILLER_44_2102 ();
 sg13g2_decap_8 FILLER_44_2150 ();
 sg13g2_fill_2 FILLER_44_2157 ();
 sg13g2_fill_1 FILLER_44_2185 ();
 sg13g2_fill_2 FILLER_44_2212 ();
 sg13g2_fill_1 FILLER_44_2222 ();
 sg13g2_decap_4 FILLER_44_2233 ();
 sg13g2_fill_2 FILLER_44_2263 ();
 sg13g2_fill_1 FILLER_44_2265 ();
 sg13g2_decap_8 FILLER_44_2318 ();
 sg13g2_decap_8 FILLER_44_2325 ();
 sg13g2_decap_4 FILLER_44_2332 ();
 sg13g2_fill_1 FILLER_44_2336 ();
 sg13g2_decap_8 FILLER_44_2367 ();
 sg13g2_decap_8 FILLER_44_2374 ();
 sg13g2_fill_2 FILLER_44_2381 ();
 sg13g2_fill_1 FILLER_44_2383 ();
 sg13g2_decap_4 FILLER_44_2390 ();
 sg13g2_fill_2 FILLER_44_2394 ();
 sg13g2_fill_1 FILLER_44_2400 ();
 sg13g2_fill_2 FILLER_44_2414 ();
 sg13g2_fill_2 FILLER_44_2425 ();
 sg13g2_decap_8 FILLER_44_2431 ();
 sg13g2_decap_4 FILLER_44_2497 ();
 sg13g2_fill_2 FILLER_44_2510 ();
 sg13g2_fill_1 FILLER_44_2512 ();
 sg13g2_decap_4 FILLER_44_2518 ();
 sg13g2_fill_2 FILLER_44_2522 ();
 sg13g2_fill_2 FILLER_44_2545 ();
 sg13g2_fill_1 FILLER_44_2621 ();
 sg13g2_decap_4 FILLER_44_2638 ();
 sg13g2_fill_2 FILLER_44_2668 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_7 ();
 sg13g2_fill_1 FILLER_45_9 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_4 FILLER_45_21 ();
 sg13g2_fill_2 FILLER_45_29 ();
 sg13g2_decap_8 FILLER_45_45 ();
 sg13g2_decap_8 FILLER_45_52 ();
 sg13g2_fill_2 FILLER_45_59 ();
 sg13g2_fill_2 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_120 ();
 sg13g2_fill_2 FILLER_45_139 ();
 sg13g2_fill_1 FILLER_45_141 ();
 sg13g2_fill_1 FILLER_45_150 ();
 sg13g2_decap_8 FILLER_45_164 ();
 sg13g2_fill_2 FILLER_45_171 ();
 sg13g2_fill_1 FILLER_45_173 ();
 sg13g2_fill_1 FILLER_45_178 ();
 sg13g2_fill_2 FILLER_45_185 ();
 sg13g2_fill_1 FILLER_45_187 ();
 sg13g2_decap_8 FILLER_45_202 ();
 sg13g2_decap_4 FILLER_45_209 ();
 sg13g2_fill_1 FILLER_45_213 ();
 sg13g2_fill_2 FILLER_45_229 ();
 sg13g2_decap_4 FILLER_45_235 ();
 sg13g2_decap_4 FILLER_45_247 ();
 sg13g2_decap_4 FILLER_45_256 ();
 sg13g2_decap_4 FILLER_45_265 ();
 sg13g2_fill_2 FILLER_45_269 ();
 sg13g2_fill_2 FILLER_45_291 ();
 sg13g2_decap_4 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_410 ();
 sg13g2_fill_1 FILLER_45_412 ();
 sg13g2_fill_1 FILLER_45_426 ();
 sg13g2_fill_1 FILLER_45_442 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_fill_1 FILLER_45_462 ();
 sg13g2_fill_2 FILLER_45_467 ();
 sg13g2_fill_1 FILLER_45_495 ();
 sg13g2_fill_1 FILLER_45_509 ();
 sg13g2_decap_4 FILLER_45_518 ();
 sg13g2_fill_2 FILLER_45_522 ();
 sg13g2_decap_8 FILLER_45_527 ();
 sg13g2_fill_2 FILLER_45_534 ();
 sg13g2_fill_2 FILLER_45_540 ();
 sg13g2_fill_1 FILLER_45_575 ();
 sg13g2_fill_1 FILLER_45_583 ();
 sg13g2_fill_2 FILLER_45_602 ();
 sg13g2_fill_2 FILLER_45_629 ();
 sg13g2_fill_1 FILLER_45_639 ();
 sg13g2_fill_2 FILLER_45_643 ();
 sg13g2_fill_1 FILLER_45_645 ();
 sg13g2_fill_1 FILLER_45_652 ();
 sg13g2_fill_1 FILLER_45_656 ();
 sg13g2_decap_8 FILLER_45_729 ();
 sg13g2_decap_4 FILLER_45_736 ();
 sg13g2_fill_1 FILLER_45_744 ();
 sg13g2_decap_4 FILLER_45_749 ();
 sg13g2_fill_2 FILLER_45_753 ();
 sg13g2_fill_2 FILLER_45_868 ();
 sg13g2_fill_1 FILLER_45_870 ();
 sg13g2_decap_4 FILLER_45_875 ();
 sg13g2_fill_1 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_926 ();
 sg13g2_decap_8 FILLER_45_933 ();
 sg13g2_fill_2 FILLER_45_997 ();
 sg13g2_fill_1 FILLER_45_1003 ();
 sg13g2_fill_2 FILLER_45_1034 ();
 sg13g2_decap_8 FILLER_45_1045 ();
 sg13g2_decap_4 FILLER_45_1052 ();
 sg13g2_decap_8 FILLER_45_1060 ();
 sg13g2_decap_8 FILLER_45_1067 ();
 sg13g2_decap_8 FILLER_45_1074 ();
 sg13g2_decap_8 FILLER_45_1081 ();
 sg13g2_decap_4 FILLER_45_1092 ();
 sg13g2_fill_1 FILLER_45_1096 ();
 sg13g2_decap_4 FILLER_45_1110 ();
 sg13g2_fill_2 FILLER_45_1114 ();
 sg13g2_fill_2 FILLER_45_1150 ();
 sg13g2_fill_1 FILLER_45_1152 ();
 sg13g2_decap_8 FILLER_45_1158 ();
 sg13g2_decap_8 FILLER_45_1165 ();
 sg13g2_fill_1 FILLER_45_1172 ();
 sg13g2_decap_4 FILLER_45_1177 ();
 sg13g2_decap_4 FILLER_45_1195 ();
 sg13g2_decap_8 FILLER_45_1204 ();
 sg13g2_decap_4 FILLER_45_1211 ();
 sg13g2_fill_1 FILLER_45_1227 ();
 sg13g2_fill_1 FILLER_45_1250 ();
 sg13g2_fill_1 FILLER_45_1257 ();
 sg13g2_fill_2 FILLER_45_1261 ();
 sg13g2_fill_1 FILLER_45_1263 ();
 sg13g2_fill_2 FILLER_45_1278 ();
 sg13g2_fill_1 FILLER_45_1280 ();
 sg13g2_decap_4 FILLER_45_1294 ();
 sg13g2_fill_1 FILLER_45_1298 ();
 sg13g2_decap_8 FILLER_45_1306 ();
 sg13g2_decap_8 FILLER_45_1324 ();
 sg13g2_decap_8 FILLER_45_1331 ();
 sg13g2_fill_2 FILLER_45_1338 ();
 sg13g2_fill_1 FILLER_45_1406 ();
 sg13g2_fill_1 FILLER_45_1439 ();
 sg13g2_fill_1 FILLER_45_1489 ();
 sg13g2_fill_1 FILLER_45_1500 ();
 sg13g2_fill_2 FILLER_45_1530 ();
 sg13g2_fill_1 FILLER_45_1532 ();
 sg13g2_fill_1 FILLER_45_1541 ();
 sg13g2_fill_2 FILLER_45_1570 ();
 sg13g2_decap_8 FILLER_45_1606 ();
 sg13g2_decap_8 FILLER_45_1613 ();
 sg13g2_fill_2 FILLER_45_1620 ();
 sg13g2_fill_2 FILLER_45_1626 ();
 sg13g2_decap_4 FILLER_45_1632 ();
 sg13g2_fill_1 FILLER_45_1640 ();
 sg13g2_fill_2 FILLER_45_1650 ();
 sg13g2_fill_2 FILLER_45_1676 ();
 sg13g2_decap_4 FILLER_45_1721 ();
 sg13g2_fill_2 FILLER_45_1725 ();
 sg13g2_decap_8 FILLER_45_1732 ();
 sg13g2_fill_1 FILLER_45_1739 ();
 sg13g2_decap_4 FILLER_45_1763 ();
 sg13g2_decap_4 FILLER_45_1777 ();
 sg13g2_fill_1 FILLER_45_1781 ();
 sg13g2_decap_4 FILLER_45_1786 ();
 sg13g2_fill_1 FILLER_45_1790 ();
 sg13g2_fill_1 FILLER_45_1820 ();
 sg13g2_fill_2 FILLER_45_1828 ();
 sg13g2_fill_1 FILLER_45_1830 ();
 sg13g2_decap_8 FILLER_45_1838 ();
 sg13g2_decap_4 FILLER_45_1845 ();
 sg13g2_fill_2 FILLER_45_1849 ();
 sg13g2_decap_4 FILLER_45_1869 ();
 sg13g2_fill_1 FILLER_45_1873 ();
 sg13g2_decap_8 FILLER_45_1879 ();
 sg13g2_fill_2 FILLER_45_1886 ();
 sg13g2_fill_1 FILLER_45_1902 ();
 sg13g2_fill_2 FILLER_45_1949 ();
 sg13g2_fill_1 FILLER_45_1951 ();
 sg13g2_decap_8 FILLER_45_2009 ();
 sg13g2_decap_8 FILLER_45_2016 ();
 sg13g2_decap_8 FILLER_45_2023 ();
 sg13g2_decap_8 FILLER_45_2030 ();
 sg13g2_decap_8 FILLER_45_2037 ();
 sg13g2_decap_8 FILLER_45_2044 ();
 sg13g2_decap_8 FILLER_45_2055 ();
 sg13g2_fill_2 FILLER_45_2062 ();
 sg13g2_decap_4 FILLER_45_2103 ();
 sg13g2_fill_2 FILLER_45_2107 ();
 sg13g2_decap_4 FILLER_45_2149 ();
 sg13g2_fill_2 FILLER_45_2153 ();
 sg13g2_decap_8 FILLER_45_2165 ();
 sg13g2_decap_8 FILLER_45_2172 ();
 sg13g2_decap_8 FILLER_45_2179 ();
 sg13g2_decap_8 FILLER_45_2186 ();
 sg13g2_fill_2 FILLER_45_2193 ();
 sg13g2_decap_4 FILLER_45_2272 ();
 sg13g2_decap_8 FILLER_45_2306 ();
 sg13g2_fill_2 FILLER_45_2313 ();
 sg13g2_fill_1 FILLER_45_2315 ();
 sg13g2_fill_2 FILLER_45_2340 ();
 sg13g2_fill_1 FILLER_45_2342 ();
 sg13g2_decap_8 FILLER_45_2347 ();
 sg13g2_fill_2 FILLER_45_2354 ();
 sg13g2_decap_4 FILLER_45_2362 ();
 sg13g2_fill_1 FILLER_45_2366 ();
 sg13g2_fill_1 FILLER_45_2403 ();
 sg13g2_decap_8 FILLER_45_2436 ();
 sg13g2_fill_2 FILLER_45_2443 ();
 sg13g2_decap_8 FILLER_45_2450 ();
 sg13g2_fill_1 FILLER_45_2457 ();
 sg13g2_fill_2 FILLER_45_2468 ();
 sg13g2_fill_1 FILLER_45_2470 ();
 sg13g2_fill_1 FILLER_45_2475 ();
 sg13g2_fill_2 FILLER_45_2514 ();
 sg13g2_fill_1 FILLER_45_2526 ();
 sg13g2_fill_2 FILLER_45_2533 ();
 sg13g2_fill_1 FILLER_45_2583 ();
 sg13g2_decap_8 FILLER_45_2594 ();
 sg13g2_fill_1 FILLER_45_2610 ();
 sg13g2_decap_4 FILLER_45_2647 ();
 sg13g2_decap_8 FILLER_45_2655 ();
 sg13g2_decap_8 FILLER_45_2662 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_2 ();
 sg13g2_decap_8 FILLER_46_29 ();
 sg13g2_fill_1 FILLER_46_36 ();
 sg13g2_decap_4 FILLER_46_77 ();
 sg13g2_fill_2 FILLER_46_81 ();
 sg13g2_decap_8 FILLER_46_103 ();
 sg13g2_decap_8 FILLER_46_110 ();
 sg13g2_decap_4 FILLER_46_117 ();
 sg13g2_fill_2 FILLER_46_121 ();
 sg13g2_fill_1 FILLER_46_153 ();
 sg13g2_decap_8 FILLER_46_178 ();
 sg13g2_decap_4 FILLER_46_185 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_2 FILLER_46_200 ();
 sg13g2_fill_1 FILLER_46_202 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_fill_1 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_230 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_fill_1 FILLER_46_257 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_fill_1 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_279 ();
 sg13g2_fill_1 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_367 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_2 FILLER_46_435 ();
 sg13g2_fill_2 FILLER_46_450 ();
 sg13g2_fill_1 FILLER_46_457 ();
 sg13g2_fill_2 FILLER_46_484 ();
 sg13g2_fill_1 FILLER_46_547 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_fill_2 FILLER_46_591 ();
 sg13g2_fill_1 FILLER_46_610 ();
 sg13g2_fill_1 FILLER_46_622 ();
 sg13g2_fill_1 FILLER_46_633 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_fill_2 FILLER_46_681 ();
 sg13g2_fill_2 FILLER_46_703 ();
 sg13g2_decap_4 FILLER_46_720 ();
 sg13g2_fill_2 FILLER_46_728 ();
 sg13g2_fill_1 FILLER_46_730 ();
 sg13g2_fill_2 FILLER_46_761 ();
 sg13g2_fill_1 FILLER_46_763 ();
 sg13g2_fill_1 FILLER_46_800 ();
 sg13g2_fill_2 FILLER_46_812 ();
 sg13g2_fill_1 FILLER_46_855 ();
 sg13g2_fill_2 FILLER_46_861 ();
 sg13g2_fill_1 FILLER_46_863 ();
 sg13g2_fill_2 FILLER_46_890 ();
 sg13g2_fill_2 FILLER_46_904 ();
 sg13g2_fill_1 FILLER_46_906 ();
 sg13g2_decap_4 FILLER_46_911 ();
 sg13g2_fill_1 FILLER_46_915 ();
 sg13g2_decap_4 FILLER_46_968 ();
 sg13g2_fill_2 FILLER_46_972 ();
 sg13g2_decap_8 FILLER_46_979 ();
 sg13g2_decap_8 FILLER_46_986 ();
 sg13g2_decap_4 FILLER_46_993 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_decap_8 FILLER_46_1090 ();
 sg13g2_decap_8 FILLER_46_1102 ();
 sg13g2_decap_8 FILLER_46_1109 ();
 sg13g2_fill_2 FILLER_46_1116 ();
 sg13g2_fill_1 FILLER_46_1118 ();
 sg13g2_fill_1 FILLER_46_1123 ();
 sg13g2_fill_2 FILLER_46_1129 ();
 sg13g2_fill_2 FILLER_46_1157 ();
 sg13g2_decap_8 FILLER_46_1164 ();
 sg13g2_decap_8 FILLER_46_1171 ();
 sg13g2_fill_2 FILLER_46_1178 ();
 sg13g2_decap_4 FILLER_46_1221 ();
 sg13g2_fill_1 FILLER_46_1225 ();
 sg13g2_fill_1 FILLER_46_1259 ();
 sg13g2_fill_1 FILLER_46_1274 ();
 sg13g2_fill_2 FILLER_46_1311 ();
 sg13g2_decap_8 FILLER_46_1318 ();
 sg13g2_decap_8 FILLER_46_1325 ();
 sg13g2_fill_2 FILLER_46_1372 ();
 sg13g2_decap_8 FILLER_46_1410 ();
 sg13g2_fill_1 FILLER_46_1417 ();
 sg13g2_fill_1 FILLER_46_1427 ();
 sg13g2_fill_2 FILLER_46_1483 ();
 sg13g2_fill_2 FILLER_46_1512 ();
 sg13g2_fill_2 FILLER_46_1519 ();
 sg13g2_fill_1 FILLER_46_1531 ();
 sg13g2_fill_2 FILLER_46_1539 ();
 sg13g2_fill_1 FILLER_46_1547 ();
 sg13g2_fill_2 FILLER_46_1553 ();
 sg13g2_fill_1 FILLER_46_1561 ();
 sg13g2_fill_1 FILLER_46_1579 ();
 sg13g2_fill_2 FILLER_46_1587 ();
 sg13g2_decap_8 FILLER_46_1604 ();
 sg13g2_decap_4 FILLER_46_1611 ();
 sg13g2_fill_2 FILLER_46_1615 ();
 sg13g2_decap_8 FILLER_46_1627 ();
 sg13g2_decap_8 FILLER_46_1634 ();
 sg13g2_fill_1 FILLER_46_1649 ();
 sg13g2_fill_1 FILLER_46_1695 ();
 sg13g2_fill_1 FILLER_46_1716 ();
 sg13g2_fill_1 FILLER_46_1725 ();
 sg13g2_fill_2 FILLER_46_1733 ();
 sg13g2_fill_2 FILLER_46_1743 ();
 sg13g2_fill_2 FILLER_46_1771 ();
 sg13g2_fill_1 FILLER_46_1773 ();
 sg13g2_fill_2 FILLER_46_1811 ();
 sg13g2_decap_4 FILLER_46_1849 ();
 sg13g2_fill_1 FILLER_46_1853 ();
 sg13g2_fill_2 FILLER_46_1879 ();
 sg13g2_fill_1 FILLER_46_1881 ();
 sg13g2_decap_4 FILLER_46_1887 ();
 sg13g2_decap_8 FILLER_46_1895 ();
 sg13g2_fill_1 FILLER_46_1902 ();
 sg13g2_fill_1 FILLER_46_1918 ();
 sg13g2_fill_1 FILLER_46_1925 ();
 sg13g2_fill_1 FILLER_46_1930 ();
 sg13g2_fill_2 FILLER_46_1952 ();
 sg13g2_fill_1 FILLER_46_1954 ();
 sg13g2_fill_2 FILLER_46_1988 ();
 sg13g2_fill_1 FILLER_46_1990 ();
 sg13g2_decap_8 FILLER_46_2013 ();
 sg13g2_decap_8 FILLER_46_2020 ();
 sg13g2_fill_2 FILLER_46_2037 ();
 sg13g2_fill_1 FILLER_46_2039 ();
 sg13g2_decap_8 FILLER_46_2054 ();
 sg13g2_decap_4 FILLER_46_2061 ();
 sg13g2_fill_1 FILLER_46_2065 ();
 sg13g2_decap_8 FILLER_46_2076 ();
 sg13g2_decap_8 FILLER_46_2083 ();
 sg13g2_decap_8 FILLER_46_2090 ();
 sg13g2_decap_8 FILLER_46_2097 ();
 sg13g2_decap_8 FILLER_46_2104 ();
 sg13g2_fill_2 FILLER_46_2111 ();
 sg13g2_decap_8 FILLER_46_2156 ();
 sg13g2_decap_8 FILLER_46_2163 ();
 sg13g2_decap_8 FILLER_46_2170 ();
 sg13g2_decap_8 FILLER_46_2177 ();
 sg13g2_decap_4 FILLER_46_2184 ();
 sg13g2_decap_8 FILLER_46_2192 ();
 sg13g2_fill_1 FILLER_46_2199 ();
 sg13g2_fill_1 FILLER_46_2239 ();
 sg13g2_fill_1 FILLER_46_2266 ();
 sg13g2_fill_2 FILLER_46_2277 ();
 sg13g2_fill_1 FILLER_46_2279 ();
 sg13g2_decap_4 FILLER_46_2306 ();
 sg13g2_decap_4 FILLER_46_2391 ();
 sg13g2_fill_1 FILLER_46_2395 ();
 sg13g2_fill_2 FILLER_46_2401 ();
 sg13g2_decap_8 FILLER_46_2449 ();
 sg13g2_decap_8 FILLER_46_2456 ();
 sg13g2_decap_4 FILLER_46_2463 ();
 sg13g2_fill_1 FILLER_46_2467 ();
 sg13g2_decap_8 FILLER_46_2473 ();
 sg13g2_fill_2 FILLER_46_2486 ();
 sg13g2_fill_2 FILLER_46_2496 ();
 sg13g2_fill_2 FILLER_46_2566 ();
 sg13g2_fill_2 FILLER_46_2629 ();
 sg13g2_fill_1 FILLER_46_2631 ();
 sg13g2_fill_2 FILLER_46_2668 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_13 ();
 sg13g2_decap_4 FILLER_47_45 ();
 sg13g2_fill_2 FILLER_47_49 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_decap_4 FILLER_47_69 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_2 FILLER_47_88 ();
 sg13g2_decap_8 FILLER_47_96 ();
 sg13g2_decap_8 FILLER_47_108 ();
 sg13g2_fill_1 FILLER_47_144 ();
 sg13g2_decap_8 FILLER_47_191 ();
 sg13g2_decap_8 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_47_205 ();
 sg13g2_decap_8 FILLER_47_261 ();
 sg13g2_fill_2 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_296 ();
 sg13g2_fill_1 FILLER_47_298 ();
 sg13g2_decap_4 FILLER_47_305 ();
 sg13g2_decap_8 FILLER_47_317 ();
 sg13g2_decap_8 FILLER_47_324 ();
 sg13g2_decap_8 FILLER_47_335 ();
 sg13g2_decap_8 FILLER_47_342 ();
 sg13g2_fill_2 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_361 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_378 ();
 sg13g2_fill_2 FILLER_47_383 ();
 sg13g2_fill_2 FILLER_47_394 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_433 ();
 sg13g2_fill_1 FILLER_47_439 ();
 sg13g2_fill_1 FILLER_47_445 ();
 sg13g2_fill_2 FILLER_47_486 ();
 sg13g2_fill_1 FILLER_47_501 ();
 sg13g2_fill_2 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_640 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_fill_1 FILLER_47_674 ();
 sg13g2_fill_2 FILLER_47_690 ();
 sg13g2_decap_4 FILLER_47_719 ();
 sg13g2_fill_1 FILLER_47_723 ();
 sg13g2_decap_8 FILLER_47_729 ();
 sg13g2_fill_2 FILLER_47_736 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_4 FILLER_47_749 ();
 sg13g2_fill_2 FILLER_47_753 ();
 sg13g2_decap_4 FILLER_47_767 ();
 sg13g2_fill_2 FILLER_47_783 ();
 sg13g2_fill_1 FILLER_47_802 ();
 sg13g2_fill_1 FILLER_47_806 ();
 sg13g2_fill_1 FILLER_47_835 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_fill_1 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_911 ();
 sg13g2_decap_8 FILLER_47_926 ();
 sg13g2_fill_1 FILLER_47_933 ();
 sg13g2_fill_1 FILLER_47_944 ();
 sg13g2_fill_2 FILLER_47_971 ();
 sg13g2_decap_4 FILLER_47_1025 ();
 sg13g2_decap_8 FILLER_47_1055 ();
 sg13g2_fill_1 FILLER_47_1062 ();
 sg13g2_decap_8 FILLER_47_1088 ();
 sg13g2_decap_8 FILLER_47_1095 ();
 sg13g2_fill_2 FILLER_47_1102 ();
 sg13g2_decap_8 FILLER_47_1150 ();
 sg13g2_decap_8 FILLER_47_1157 ();
 sg13g2_decap_8 FILLER_47_1164 ();
 sg13g2_decap_8 FILLER_47_1171 ();
 sg13g2_fill_1 FILLER_47_1178 ();
 sg13g2_fill_2 FILLER_47_1206 ();
 sg13g2_fill_1 FILLER_47_1208 ();
 sg13g2_fill_2 FILLER_47_1213 ();
 sg13g2_fill_2 FILLER_47_1236 ();
 sg13g2_decap_4 FILLER_47_1283 ();
 sg13g2_decap_4 FILLER_47_1326 ();
 sg13g2_fill_2 FILLER_47_1335 ();
 sg13g2_fill_2 FILLER_47_1341 ();
 sg13g2_fill_1 FILLER_47_1347 ();
 sg13g2_fill_1 FILLER_47_1378 ();
 sg13g2_fill_2 FILLER_47_1406 ();
 sg13g2_fill_2 FILLER_47_1415 ();
 sg13g2_fill_1 FILLER_47_1462 ();
 sg13g2_fill_2 FILLER_47_1472 ();
 sg13g2_fill_1 FILLER_47_1486 ();
 sg13g2_fill_1 FILLER_47_1492 ();
 sg13g2_fill_2 FILLER_47_1497 ();
 sg13g2_fill_1 FILLER_47_1536 ();
 sg13g2_fill_1 FILLER_47_1559 ();
 sg13g2_fill_1 FILLER_47_1592 ();
 sg13g2_fill_2 FILLER_47_1601 ();
 sg13g2_fill_2 FILLER_47_1613 ();
 sg13g2_decap_8 FILLER_47_1619 ();
 sg13g2_fill_1 FILLER_47_1626 ();
 sg13g2_fill_1 FILLER_47_1641 ();
 sg13g2_fill_1 FILLER_47_1656 ();
 sg13g2_fill_2 FILLER_47_1678 ();
 sg13g2_fill_1 FILLER_47_1755 ();
 sg13g2_fill_2 FILLER_47_1772 ();
 sg13g2_decap_4 FILLER_47_1785 ();
 sg13g2_fill_1 FILLER_47_1789 ();
 sg13g2_fill_2 FILLER_47_1797 ();
 sg13g2_fill_1 FILLER_47_1799 ();
 sg13g2_fill_1 FILLER_47_1807 ();
 sg13g2_fill_2 FILLER_47_1838 ();
 sg13g2_fill_1 FILLER_47_1840 ();
 sg13g2_decap_8 FILLER_47_1848 ();
 sg13g2_decap_4 FILLER_47_1855 ();
 sg13g2_fill_1 FILLER_47_1859 ();
 sg13g2_decap_4 FILLER_47_1865 ();
 sg13g2_fill_2 FILLER_47_1869 ();
 sg13g2_decap_4 FILLER_47_1875 ();
 sg13g2_fill_1 FILLER_47_1879 ();
 sg13g2_fill_2 FILLER_47_1885 ();
 sg13g2_fill_2 FILLER_47_1891 ();
 sg13g2_fill_1 FILLER_47_1897 ();
 sg13g2_fill_2 FILLER_47_1911 ();
 sg13g2_fill_1 FILLER_47_1913 ();
 sg13g2_fill_2 FILLER_47_1918 ();
 sg13g2_fill_1 FILLER_47_1920 ();
 sg13g2_fill_2 FILLER_47_1925 ();
 sg13g2_fill_1 FILLER_47_1927 ();
 sg13g2_fill_1 FILLER_47_1938 ();
 sg13g2_fill_2 FILLER_47_1944 ();
 sg13g2_fill_1 FILLER_47_1946 ();
 sg13g2_fill_1 FILLER_47_1956 ();
 sg13g2_fill_2 FILLER_47_1966 ();
 sg13g2_decap_8 FILLER_47_1993 ();
 sg13g2_decap_8 FILLER_47_2000 ();
 sg13g2_decap_4 FILLER_47_2007 ();
 sg13g2_fill_2 FILLER_47_2011 ();
 sg13g2_decap_8 FILLER_47_2073 ();
 sg13g2_decap_8 FILLER_47_2080 ();
 sg13g2_decap_8 FILLER_47_2087 ();
 sg13g2_decap_8 FILLER_47_2094 ();
 sg13g2_decap_4 FILLER_47_2101 ();
 sg13g2_fill_2 FILLER_47_2115 ();
 sg13g2_decap_4 FILLER_47_2138 ();
 sg13g2_fill_2 FILLER_47_2142 ();
 sg13g2_fill_1 FILLER_47_2183 ();
 sg13g2_decap_4 FILLER_47_2216 ();
 sg13g2_fill_1 FILLER_47_2220 ();
 sg13g2_decap_8 FILLER_47_2225 ();
 sg13g2_fill_1 FILLER_47_2232 ();
 sg13g2_fill_2 FILLER_47_2237 ();
 sg13g2_fill_2 FILLER_47_2249 ();
 sg13g2_fill_2 FILLER_47_2255 ();
 sg13g2_fill_1 FILLER_47_2257 ();
 sg13g2_fill_2 FILLER_47_2268 ();
 sg13g2_fill_1 FILLER_47_2270 ();
 sg13g2_fill_2 FILLER_47_2281 ();
 sg13g2_fill_1 FILLER_47_2283 ();
 sg13g2_decap_4 FILLER_47_2292 ();
 sg13g2_fill_2 FILLER_47_2296 ();
 sg13g2_fill_1 FILLER_47_2311 ();
 sg13g2_decap_8 FILLER_47_2349 ();
 sg13g2_fill_2 FILLER_47_2356 ();
 sg13g2_fill_1 FILLER_47_2358 ();
 sg13g2_fill_2 FILLER_47_2368 ();
 sg13g2_fill_1 FILLER_47_2384 ();
 sg13g2_fill_1 FILLER_47_2391 ();
 sg13g2_fill_2 FILLER_47_2398 ();
 sg13g2_fill_2 FILLER_47_2410 ();
 sg13g2_fill_1 FILLER_47_2412 ();
 sg13g2_decap_4 FILLER_47_2417 ();
 sg13g2_fill_2 FILLER_47_2421 ();
 sg13g2_fill_2 FILLER_47_2447 ();
 sg13g2_fill_2 FILLER_47_2483 ();
 sg13g2_fill_1 FILLER_47_2485 ();
 sg13g2_decap_4 FILLER_47_2512 ();
 sg13g2_fill_1 FILLER_47_2526 ();
 sg13g2_fill_2 FILLER_47_2530 ();
 sg13g2_fill_1 FILLER_47_2545 ();
 sg13g2_decap_8 FILLER_47_2610 ();
 sg13g2_fill_1 FILLER_47_2617 ();
 sg13g2_fill_2 FILLER_47_2631 ();
 sg13g2_fill_1 FILLER_47_2633 ();
 sg13g2_fill_1 FILLER_47_2648 ();
 sg13g2_decap_8 FILLER_47_2653 ();
 sg13g2_decap_8 FILLER_47_2660 ();
 sg13g2_fill_2 FILLER_47_2667 ();
 sg13g2_fill_1 FILLER_47_2669 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_33 ();
 sg13g2_fill_1 FILLER_48_93 ();
 sg13g2_fill_1 FILLER_48_99 ();
 sg13g2_decap_4 FILLER_48_114 ();
 sg13g2_fill_2 FILLER_48_118 ();
 sg13g2_decap_4 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_fill_2 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_169 ();
 sg13g2_fill_2 FILLER_48_176 ();
 sg13g2_fill_1 FILLER_48_204 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_fill_2 FILLER_48_217 ();
 sg13g2_fill_2 FILLER_48_223 ();
 sg13g2_fill_1 FILLER_48_225 ();
 sg13g2_fill_1 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_237 ();
 sg13g2_fill_2 FILLER_48_244 ();
 sg13g2_fill_2 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_263 ();
 sg13g2_decap_8 FILLER_48_270 ();
 sg13g2_fill_2 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_283 ();
 sg13g2_decap_4 FILLER_48_299 ();
 sg13g2_fill_2 FILLER_48_303 ();
 sg13g2_fill_1 FILLER_48_309 ();
 sg13g2_decap_4 FILLER_48_315 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_decap_8 FILLER_48_325 ();
 sg13g2_decap_8 FILLER_48_332 ();
 sg13g2_decap_8 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_351 ();
 sg13g2_decap_4 FILLER_48_357 ();
 sg13g2_fill_2 FILLER_48_365 ();
 sg13g2_decap_8 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_383 ();
 sg13g2_decap_4 FILLER_48_390 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_fill_2 FILLER_48_417 ();
 sg13g2_fill_1 FILLER_48_451 ();
 sg13g2_fill_1 FILLER_48_457 ();
 sg13g2_fill_2 FILLER_48_475 ();
 sg13g2_fill_2 FILLER_48_535 ();
 sg13g2_fill_2 FILLER_48_578 ();
 sg13g2_fill_1 FILLER_48_580 ();
 sg13g2_fill_1 FILLER_48_617 ();
 sg13g2_fill_1 FILLER_48_623 ();
 sg13g2_fill_1 FILLER_48_639 ();
 sg13g2_fill_1 FILLER_48_653 ();
 sg13g2_fill_2 FILLER_48_713 ();
 sg13g2_fill_1 FILLER_48_715 ();
 sg13g2_fill_2 FILLER_48_731 ();
 sg13g2_decap_4 FILLER_48_743 ();
 sg13g2_fill_1 FILLER_48_747 ();
 sg13g2_decap_4 FILLER_48_758 ();
 sg13g2_fill_2 FILLER_48_792 ();
 sg13g2_fill_2 FILLER_48_815 ();
 sg13g2_fill_2 FILLER_48_824 ();
 sg13g2_fill_1 FILLER_48_832 ();
 sg13g2_fill_1 FILLER_48_837 ();
 sg13g2_fill_2 FILLER_48_862 ();
 sg13g2_fill_2 FILLER_48_868 ();
 sg13g2_fill_2 FILLER_48_878 ();
 sg13g2_fill_1 FILLER_48_880 ();
 sg13g2_decap_8 FILLER_48_923 ();
 sg13g2_fill_2 FILLER_48_930 ();
 sg13g2_fill_1 FILLER_48_932 ();
 sg13g2_fill_2 FILLER_48_938 ();
 sg13g2_fill_2 FILLER_48_944 ();
 sg13g2_decap_8 FILLER_48_964 ();
 sg13g2_decap_8 FILLER_48_971 ();
 sg13g2_fill_2 FILLER_48_978 ();
 sg13g2_decap_8 FILLER_48_988 ();
 sg13g2_decap_4 FILLER_48_995 ();
 sg13g2_decap_8 FILLER_48_1025 ();
 sg13g2_fill_2 FILLER_48_1072 ();
 sg13g2_fill_1 FILLER_48_1074 ();
 sg13g2_fill_2 FILLER_48_1105 ();
 sg13g2_fill_1 FILLER_48_1107 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_decap_8 FILLER_48_1120 ();
 sg13g2_fill_2 FILLER_48_1140 ();
 sg13g2_fill_2 FILLER_48_1147 ();
 sg13g2_decap_8 FILLER_48_1175 ();
 sg13g2_fill_1 FILLER_48_1182 ();
 sg13g2_fill_1 FILLER_48_1264 ();
 sg13g2_fill_2 FILLER_48_1311 ();
 sg13g2_fill_2 FILLER_48_1324 ();
 sg13g2_fill_2 FILLER_48_1352 ();
 sg13g2_decap_4 FILLER_48_1378 ();
 sg13g2_fill_2 FILLER_48_1388 ();
 sg13g2_fill_1 FILLER_48_1416 ();
 sg13g2_fill_2 FILLER_48_1439 ();
 sg13g2_fill_1 FILLER_48_1497 ();
 sg13g2_fill_1 FILLER_48_1512 ();
 sg13g2_fill_2 FILLER_48_1529 ();
 sg13g2_fill_2 FILLER_48_1562 ();
 sg13g2_fill_1 FILLER_48_1602 ();
 sg13g2_fill_1 FILLER_48_1613 ();
 sg13g2_fill_2 FILLER_48_1627 ();
 sg13g2_fill_1 FILLER_48_1629 ();
 sg13g2_fill_2 FILLER_48_1643 ();
 sg13g2_fill_1 FILLER_48_1645 ();
 sg13g2_fill_2 FILLER_48_1659 ();
 sg13g2_fill_1 FILLER_48_1713 ();
 sg13g2_decap_8 FILLER_48_1719 ();
 sg13g2_fill_1 FILLER_48_1726 ();
 sg13g2_decap_8 FILLER_48_1790 ();
 sg13g2_fill_2 FILLER_48_1797 ();
 sg13g2_decap_8 FILLER_48_1803 ();
 sg13g2_fill_2 FILLER_48_1814 ();
 sg13g2_decap_8 FILLER_48_1846 ();
 sg13g2_fill_1 FILLER_48_1853 ();
 sg13g2_decap_4 FILLER_48_1862 ();
 sg13g2_fill_1 FILLER_48_1866 ();
 sg13g2_fill_2 FILLER_48_1881 ();
 sg13g2_fill_2 FILLER_48_1886 ();
 sg13g2_decap_8 FILLER_48_1896 ();
 sg13g2_decap_4 FILLER_48_1903 ();
 sg13g2_fill_2 FILLER_48_1907 ();
 sg13g2_fill_2 FILLER_48_1914 ();
 sg13g2_fill_1 FILLER_48_1916 ();
 sg13g2_fill_1 FILLER_48_1937 ();
 sg13g2_decap_4 FILLER_48_1944 ();
 sg13g2_fill_1 FILLER_48_1948 ();
 sg13g2_fill_2 FILLER_48_1959 ();
 sg13g2_fill_1 FILLER_48_1961 ();
 sg13g2_decap_8 FILLER_48_1978 ();
 sg13g2_decap_8 FILLER_48_1985 ();
 sg13g2_decap_8 FILLER_48_1992 ();
 sg13g2_decap_8 FILLER_48_1999 ();
 sg13g2_fill_2 FILLER_48_2006 ();
 sg13g2_fill_1 FILLER_48_2008 ();
 sg13g2_decap_8 FILLER_48_2023 ();
 sg13g2_fill_2 FILLER_48_2082 ();
 sg13g2_fill_2 FILLER_48_2118 ();
 sg13g2_decap_4 FILLER_48_2146 ();
 sg13g2_fill_1 FILLER_48_2206 ();
 sg13g2_decap_8 FILLER_48_2227 ();
 sg13g2_decap_8 FILLER_48_2234 ();
 sg13g2_decap_8 FILLER_48_2241 ();
 sg13g2_decap_8 FILLER_48_2248 ();
 sg13g2_decap_4 FILLER_48_2255 ();
 sg13g2_fill_1 FILLER_48_2259 ();
 sg13g2_fill_1 FILLER_48_2311 ();
 sg13g2_fill_2 FILLER_48_2315 ();
 sg13g2_decap_8 FILLER_48_2371 ();
 sg13g2_fill_2 FILLER_48_2378 ();
 sg13g2_fill_1 FILLER_48_2380 ();
 sg13g2_decap_8 FILLER_48_2386 ();
 sg13g2_decap_8 FILLER_48_2393 ();
 sg13g2_decap_4 FILLER_48_2400 ();
 sg13g2_decap_8 FILLER_48_2414 ();
 sg13g2_decap_4 FILLER_48_2421 ();
 sg13g2_fill_1 FILLER_48_2425 ();
 sg13g2_decap_8 FILLER_48_2514 ();
 sg13g2_fill_1 FILLER_48_2521 ();
 sg13g2_fill_2 FILLER_48_2571 ();
 sg13g2_fill_1 FILLER_48_2573 ();
 sg13g2_fill_1 FILLER_48_2588 ();
 sg13g2_fill_1 FILLER_48_2641 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_2 ();
 sg13g2_fill_1 FILLER_49_37 ();
 sg13g2_fill_2 FILLER_49_46 ();
 sg13g2_decap_4 FILLER_49_66 ();
 sg13g2_fill_1 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_fill_1 FILLER_49_130 ();
 sg13g2_fill_2 FILLER_49_139 ();
 sg13g2_fill_1 FILLER_49_150 ();
 sg13g2_fill_2 FILLER_49_159 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_2 FILLER_49_189 ();
 sg13g2_fill_1 FILLER_49_191 ();
 sg13g2_fill_1 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_fill_2 FILLER_49_252 ();
 sg13g2_fill_1 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_fill_2 FILLER_49_280 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_313 ();
 sg13g2_fill_1 FILLER_49_356 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_fill_2 FILLER_49_403 ();
 sg13g2_fill_1 FILLER_49_405 ();
 sg13g2_fill_1 FILLER_49_411 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_fill_2 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_49_431 ();
 sg13g2_fill_1 FILLER_49_436 ();
 sg13g2_fill_1 FILLER_49_449 ();
 sg13g2_fill_1 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_482 ();
 sg13g2_fill_1 FILLER_49_507 ();
 sg13g2_fill_1 FILLER_49_517 ();
 sg13g2_fill_2 FILLER_49_585 ();
 sg13g2_fill_1 FILLER_49_587 ();
 sg13g2_fill_2 FILLER_49_595 ();
 sg13g2_fill_1 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_fill_1 FILLER_49_680 ();
 sg13g2_fill_2 FILLER_49_744 ();
 sg13g2_decap_8 FILLER_49_759 ();
 sg13g2_fill_1 FILLER_49_766 ();
 sg13g2_fill_2 FILLER_49_790 ();
 sg13g2_fill_2 FILLER_49_807 ();
 sg13g2_fill_1 FILLER_49_898 ();
 sg13g2_fill_1 FILLER_49_906 ();
 sg13g2_fill_2 FILLER_49_915 ();
 sg13g2_fill_1 FILLER_49_922 ();
 sg13g2_decap_4 FILLER_49_936 ();
 sg13g2_fill_1 FILLER_49_940 ();
 sg13g2_decap_4 FILLER_49_946 ();
 sg13g2_fill_1 FILLER_49_950 ();
 sg13g2_decap_8 FILLER_49_956 ();
 sg13g2_decap_8 FILLER_49_963 ();
 sg13g2_decap_4 FILLER_49_970 ();
 sg13g2_fill_1 FILLER_49_974 ();
 sg13g2_fill_2 FILLER_49_984 ();
 sg13g2_fill_2 FILLER_49_1025 ();
 sg13g2_decap_8 FILLER_49_1036 ();
 sg13g2_decap_4 FILLER_49_1043 ();
 sg13g2_fill_2 FILLER_49_1047 ();
 sg13g2_fill_2 FILLER_49_1069 ();
 sg13g2_fill_1 FILLER_49_1080 ();
 sg13g2_fill_1 FILLER_49_1084 ();
 sg13g2_fill_1 FILLER_49_1090 ();
 sg13g2_decap_8 FILLER_49_1096 ();
 sg13g2_decap_8 FILLER_49_1103 ();
 sg13g2_fill_2 FILLER_49_1110 ();
 sg13g2_decap_4 FILLER_49_1129 ();
 sg13g2_fill_1 FILLER_49_1133 ();
 sg13g2_fill_2 FILLER_49_1169 ();
 sg13g2_fill_2 FILLER_49_1207 ();
 sg13g2_fill_1 FILLER_49_1223 ();
 sg13g2_fill_1 FILLER_49_1258 ();
 sg13g2_fill_2 FILLER_49_1275 ();
 sg13g2_fill_1 FILLER_49_1288 ();
 sg13g2_decap_4 FILLER_49_1301 ();
 sg13g2_fill_1 FILLER_49_1308 ();
 sg13g2_decap_8 FILLER_49_1313 ();
 sg13g2_fill_1 FILLER_49_1320 ();
 sg13g2_decap_4 FILLER_49_1327 ();
 sg13g2_fill_1 FILLER_49_1336 ();
 sg13g2_fill_2 FILLER_49_1374 ();
 sg13g2_fill_2 FILLER_49_1389 ();
 sg13g2_fill_2 FILLER_49_1417 ();
 sg13g2_fill_2 FILLER_49_1422 ();
 sg13g2_fill_2 FILLER_49_1496 ();
 sg13g2_fill_2 FILLER_49_1502 ();
 sg13g2_fill_2 FILLER_49_1562 ();
 sg13g2_fill_2 FILLER_49_1570 ();
 sg13g2_fill_2 FILLER_49_1610 ();
 sg13g2_fill_1 FILLER_49_1617 ();
 sg13g2_fill_1 FILLER_49_1626 ();
 sg13g2_fill_2 FILLER_49_1631 ();
 sg13g2_fill_1 FILLER_49_1633 ();
 sg13g2_decap_4 FILLER_49_1644 ();
 sg13g2_fill_2 FILLER_49_1667 ();
 sg13g2_fill_1 FILLER_49_1677 ();
 sg13g2_fill_2 FILLER_49_1699 ();
 sg13g2_decap_4 FILLER_49_1727 ();
 sg13g2_fill_2 FILLER_49_1731 ();
 sg13g2_fill_1 FILLER_49_1737 ();
 sg13g2_decap_8 FILLER_49_1788 ();
 sg13g2_fill_2 FILLER_49_1795 ();
 sg13g2_fill_1 FILLER_49_1797 ();
 sg13g2_decap_4 FILLER_49_1855 ();
 sg13g2_fill_1 FILLER_49_1859 ();
 sg13g2_decap_8 FILLER_49_1869 ();
 sg13g2_fill_1 FILLER_49_1876 ();
 sg13g2_fill_2 FILLER_49_1881 ();
 sg13g2_fill_1 FILLER_49_1893 ();
 sg13g2_decap_4 FILLER_49_1899 ();
 sg13g2_fill_1 FILLER_49_1903 ();
 sg13g2_decap_4 FILLER_49_1909 ();
 sg13g2_fill_1 FILLER_49_1913 ();
 sg13g2_decap_8 FILLER_49_1921 ();
 sg13g2_decap_8 FILLER_49_1928 ();
 sg13g2_decap_4 FILLER_49_1935 ();
 sg13g2_fill_2 FILLER_49_1939 ();
 sg13g2_decap_8 FILLER_49_1970 ();
 sg13g2_decap_8 FILLER_49_1977 ();
 sg13g2_decap_8 FILLER_49_1984 ();
 sg13g2_decap_8 FILLER_49_1991 ();
 sg13g2_fill_1 FILLER_49_1998 ();
 sg13g2_fill_2 FILLER_49_2003 ();
 sg13g2_fill_1 FILLER_49_2005 ();
 sg13g2_decap_4 FILLER_49_2032 ();
 sg13g2_fill_2 FILLER_49_2057 ();
 sg13g2_fill_2 FILLER_49_2069 ();
 sg13g2_fill_1 FILLER_49_2071 ();
 sg13g2_decap_8 FILLER_49_2144 ();
 sg13g2_decap_4 FILLER_49_2151 ();
 sg13g2_fill_1 FILLER_49_2165 ();
 sg13g2_fill_1 FILLER_49_2176 ();
 sg13g2_fill_2 FILLER_49_2221 ();
 sg13g2_decap_8 FILLER_49_2233 ();
 sg13g2_fill_2 FILLER_49_2240 ();
 sg13g2_decap_4 FILLER_49_2273 ();
 sg13g2_fill_1 FILLER_49_2277 ();
 sg13g2_decap_8 FILLER_49_2282 ();
 sg13g2_decap_4 FILLER_49_2289 ();
 sg13g2_fill_2 FILLER_49_2310 ();
 sg13g2_decap_8 FILLER_49_2322 ();
 sg13g2_decap_8 FILLER_49_2329 ();
 sg13g2_decap_8 FILLER_49_2336 ();
 sg13g2_decap_8 FILLER_49_2343 ();
 sg13g2_fill_2 FILLER_49_2350 ();
 sg13g2_decap_4 FILLER_49_2356 ();
 sg13g2_fill_2 FILLER_49_2364 ();
 sg13g2_fill_2 FILLER_49_2375 ();
 sg13g2_fill_1 FILLER_49_2377 ();
 sg13g2_fill_2 FILLER_49_2382 ();
 sg13g2_fill_2 FILLER_49_2388 ();
 sg13g2_fill_2 FILLER_49_2425 ();
 sg13g2_fill_1 FILLER_49_2435 ();
 sg13g2_fill_1 FILLER_49_2456 ();
 sg13g2_fill_2 FILLER_49_2461 ();
 sg13g2_fill_1 FILLER_49_2469 ();
 sg13g2_fill_1 FILLER_49_2480 ();
 sg13g2_decap_4 FILLER_49_2498 ();
 sg13g2_fill_2 FILLER_49_2502 ();
 sg13g2_fill_1 FILLER_49_2547 ();
 sg13g2_decap_8 FILLER_49_2563 ();
 sg13g2_fill_1 FILLER_49_2570 ();
 sg13g2_decap_8 FILLER_49_2581 ();
 sg13g2_decap_4 FILLER_49_2588 ();
 sg13g2_fill_2 FILLER_49_2592 ();
 sg13g2_fill_1 FILLER_49_2598 ();
 sg13g2_decap_4 FILLER_49_2606 ();
 sg13g2_fill_2 FILLER_49_2610 ();
 sg13g2_fill_2 FILLER_49_2668 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_55 ();
 sg13g2_decap_8 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_69 ();
 sg13g2_decap_4 FILLER_50_76 ();
 sg13g2_decap_4 FILLER_50_88 ();
 sg13g2_decap_8 FILLER_50_106 ();
 sg13g2_fill_2 FILLER_50_113 ();
 sg13g2_fill_1 FILLER_50_115 ();
 sg13g2_fill_2 FILLER_50_124 ();
 sg13g2_fill_2 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_157 ();
 sg13g2_fill_2 FILLER_50_163 ();
 sg13g2_fill_1 FILLER_50_165 ();
 sg13g2_fill_2 FILLER_50_170 ();
 sg13g2_fill_2 FILLER_50_191 ();
 sg13g2_fill_1 FILLER_50_193 ();
 sg13g2_decap_8 FILLER_50_242 ();
 sg13g2_fill_2 FILLER_50_249 ();
 sg13g2_fill_1 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_278 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_fill_1 FILLER_50_308 ();
 sg13g2_fill_2 FILLER_50_314 ();
 sg13g2_fill_1 FILLER_50_370 ();
 sg13g2_fill_2 FILLER_50_446 ();
 sg13g2_fill_2 FILLER_50_456 ();
 sg13g2_decap_4 FILLER_50_466 ();
 sg13g2_fill_1 FILLER_50_470 ();
 sg13g2_fill_2 FILLER_50_497 ();
 sg13g2_fill_1 FILLER_50_540 ();
 sg13g2_fill_1 FILLER_50_557 ();
 sg13g2_fill_1 FILLER_50_561 ();
 sg13g2_fill_1 FILLER_50_567 ();
 sg13g2_fill_1 FILLER_50_600 ();
 sg13g2_fill_2 FILLER_50_647 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_698 ();
 sg13g2_decap_8 FILLER_50_704 ();
 sg13g2_decap_4 FILLER_50_711 ();
 sg13g2_fill_1 FILLER_50_715 ();
 sg13g2_fill_1 FILLER_50_724 ();
 sg13g2_decap_4 FILLER_50_769 ();
 sg13g2_fill_2 FILLER_50_773 ();
 sg13g2_fill_1 FILLER_50_779 ();
 sg13g2_fill_2 FILLER_50_805 ();
 sg13g2_fill_2 FILLER_50_831 ();
 sg13g2_fill_1 FILLER_50_846 ();
 sg13g2_fill_1 FILLER_50_867 ();
 sg13g2_fill_2 FILLER_50_873 ();
 sg13g2_fill_1 FILLER_50_875 ();
 sg13g2_fill_1 FILLER_50_904 ();
 sg13g2_fill_1 FILLER_50_923 ();
 sg13g2_fill_2 FILLER_50_929 ();
 sg13g2_fill_2 FILLER_50_935 ();
 sg13g2_decap_4 FILLER_50_969 ();
 sg13g2_fill_2 FILLER_50_973 ();
 sg13g2_fill_2 FILLER_50_1004 ();
 sg13g2_fill_1 FILLER_50_1006 ();
 sg13g2_decap_8 FILLER_50_1015 ();
 sg13g2_decap_4 FILLER_50_1022 ();
 sg13g2_fill_2 FILLER_50_1026 ();
 sg13g2_decap_4 FILLER_50_1038 ();
 sg13g2_fill_2 FILLER_50_1042 ();
 sg13g2_fill_1 FILLER_50_1058 ();
 sg13g2_fill_1 FILLER_50_1064 ();
 sg13g2_fill_1 FILLER_50_1070 ();
 sg13g2_fill_2 FILLER_50_1105 ();
 sg13g2_fill_1 FILLER_50_1107 ();
 sg13g2_fill_2 FILLER_50_1143 ();
 sg13g2_fill_1 FILLER_50_1145 ();
 sg13g2_fill_2 FILLER_50_1163 ();
 sg13g2_fill_2 FILLER_50_1186 ();
 sg13g2_fill_1 FILLER_50_1188 ();
 sg13g2_decap_8 FILLER_50_1193 ();
 sg13g2_fill_2 FILLER_50_1200 ();
 sg13g2_fill_1 FILLER_50_1202 ();
 sg13g2_fill_2 FILLER_50_1240 ();
 sg13g2_fill_1 FILLER_50_1253 ();
 sg13g2_fill_2 FILLER_50_1263 ();
 sg13g2_fill_2 FILLER_50_1311 ();
 sg13g2_decap_4 FILLER_50_1316 ();
 sg13g2_decap_4 FILLER_50_1329 ();
 sg13g2_fill_1 FILLER_50_1333 ();
 sg13g2_fill_2 FILLER_50_1339 ();
 sg13g2_fill_1 FILLER_50_1378 ();
 sg13g2_fill_2 FILLER_50_1392 ();
 sg13g2_fill_2 FILLER_50_1400 ();
 sg13g2_fill_1 FILLER_50_1410 ();
 sg13g2_fill_1 FILLER_50_1427 ();
 sg13g2_fill_1 FILLER_50_1455 ();
 sg13g2_fill_2 FILLER_50_1486 ();
 sg13g2_fill_1 FILLER_50_1494 ();
 sg13g2_fill_1 FILLER_50_1528 ();
 sg13g2_fill_2 FILLER_50_1555 ();
 sg13g2_fill_1 FILLER_50_1565 ();
 sg13g2_fill_1 FILLER_50_1586 ();
 sg13g2_fill_1 FILLER_50_1611 ();
 sg13g2_fill_1 FILLER_50_1679 ();
 sg13g2_fill_2 FILLER_50_1715 ();
 sg13g2_fill_2 FILLER_50_1763 ();
 sg13g2_fill_2 FILLER_50_1772 ();
 sg13g2_fill_1 FILLER_50_1790 ();
 sg13g2_fill_2 FILLER_50_1796 ();
 sg13g2_fill_1 FILLER_50_1798 ();
 sg13g2_decap_4 FILLER_50_1803 ();
 sg13g2_fill_1 FILLER_50_1807 ();
 sg13g2_fill_1 FILLER_50_1845 ();
 sg13g2_decap_4 FILLER_50_1850 ();
 sg13g2_fill_1 FILLER_50_1854 ();
 sg13g2_fill_1 FILLER_50_1860 ();
 sg13g2_fill_1 FILLER_50_1867 ();
 sg13g2_fill_1 FILLER_50_1873 ();
 sg13g2_fill_1 FILLER_50_1905 ();
 sg13g2_fill_2 FILLER_50_1910 ();
 sg13g2_fill_1 FILLER_50_1912 ();
 sg13g2_decap_4 FILLER_50_1927 ();
 sg13g2_fill_2 FILLER_50_1931 ();
 sg13g2_decap_8 FILLER_50_1972 ();
 sg13g2_decap_4 FILLER_50_1979 ();
 sg13g2_fill_2 FILLER_50_1983 ();
 sg13g2_decap_4 FILLER_50_1989 ();
 sg13g2_fill_2 FILLER_50_1993 ();
 sg13g2_fill_2 FILLER_50_2005 ();
 sg13g2_fill_1 FILLER_50_2007 ();
 sg13g2_decap_8 FILLER_50_2033 ();
 sg13g2_decap_8 FILLER_50_2040 ();
 sg13g2_decap_4 FILLER_50_2047 ();
 sg13g2_fill_2 FILLER_50_2051 ();
 sg13g2_decap_8 FILLER_50_2063 ();
 sg13g2_decap_8 FILLER_50_2070 ();
 sg13g2_decap_8 FILLER_50_2077 ();
 sg13g2_decap_8 FILLER_50_2146 ();
 sg13g2_decap_8 FILLER_50_2153 ();
 sg13g2_decap_4 FILLER_50_2160 ();
 sg13g2_decap_4 FILLER_50_2168 ();
 sg13g2_decap_4 FILLER_50_2182 ();
 sg13g2_fill_2 FILLER_50_2186 ();
 sg13g2_fill_1 FILLER_50_2198 ();
 sg13g2_fill_1 FILLER_50_2225 ();
 sg13g2_fill_1 FILLER_50_2230 ();
 sg13g2_fill_2 FILLER_50_2257 ();
 sg13g2_fill_2 FILLER_50_2269 ();
 sg13g2_fill_1 FILLER_50_2271 ();
 sg13g2_decap_8 FILLER_50_2306 ();
 sg13g2_decap_4 FILLER_50_2313 ();
 sg13g2_decap_4 FILLER_50_2320 ();
 sg13g2_fill_1 FILLER_50_2324 ();
 sg13g2_decap_8 FILLER_50_2329 ();
 sg13g2_decap_8 FILLER_50_2336 ();
 sg13g2_fill_2 FILLER_50_2343 ();
 sg13g2_fill_1 FILLER_50_2345 ();
 sg13g2_decap_4 FILLER_50_2376 ();
 sg13g2_decap_8 FILLER_50_2384 ();
 sg13g2_decap_4 FILLER_50_2391 ();
 sg13g2_fill_1 FILLER_50_2395 ();
 sg13g2_fill_1 FILLER_50_2420 ();
 sg13g2_fill_2 FILLER_50_2426 ();
 sg13g2_fill_1 FILLER_50_2453 ();
 sg13g2_decap_4 FILLER_50_2458 ();
 sg13g2_fill_2 FILLER_50_2462 ();
 sg13g2_decap_4 FILLER_50_2469 ();
 sg13g2_fill_1 FILLER_50_2473 ();
 sg13g2_decap_4 FILLER_50_2479 ();
 sg13g2_fill_2 FILLER_50_2483 ();
 sg13g2_fill_2 FILLER_50_2493 ();
 sg13g2_decap_4 FILLER_50_2507 ();
 sg13g2_fill_2 FILLER_50_2511 ();
 sg13g2_decap_4 FILLER_50_2517 ();
 sg13g2_fill_2 FILLER_50_2521 ();
 sg13g2_decap_8 FILLER_50_2562 ();
 sg13g2_decap_8 FILLER_50_2569 ();
 sg13g2_decap_8 FILLER_50_2576 ();
 sg13g2_fill_2 FILLER_50_2583 ();
 sg13g2_decap_8 FILLER_50_2620 ();
 sg13g2_decap_8 FILLER_50_2627 ();
 sg13g2_fill_1 FILLER_50_2634 ();
 sg13g2_decap_4 FILLER_50_2643 ();
 sg13g2_fill_1 FILLER_50_2647 ();
 sg13g2_fill_1 FILLER_50_2652 ();
 sg13g2_decap_8 FILLER_50_2657 ();
 sg13g2_decap_4 FILLER_50_2664 ();
 sg13g2_fill_2 FILLER_50_2668 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_4 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_59 ();
 sg13g2_decap_8 FILLER_51_66 ();
 sg13g2_decap_4 FILLER_51_73 ();
 sg13g2_fill_1 FILLER_51_77 ();
 sg13g2_fill_2 FILLER_51_82 ();
 sg13g2_decap_8 FILLER_51_109 ();
 sg13g2_decap_8 FILLER_51_116 ();
 sg13g2_fill_1 FILLER_51_123 ();
 sg13g2_decap_4 FILLER_51_134 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_fill_1 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_170 ();
 sg13g2_decap_4 FILLER_51_177 ();
 sg13g2_fill_1 FILLER_51_181 ();
 sg13g2_decap_4 FILLER_51_192 ();
 sg13g2_decap_8 FILLER_51_240 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_254 ();
 sg13g2_decap_4 FILLER_51_268 ();
 sg13g2_decap_4 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_281 ();
 sg13g2_fill_2 FILLER_51_319 ();
 sg13g2_fill_2 FILLER_51_347 ();
 sg13g2_fill_1 FILLER_51_354 ();
 sg13g2_fill_2 FILLER_51_363 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_4 FILLER_51_392 ();
 sg13g2_fill_1 FILLER_51_396 ();
 sg13g2_fill_2 FILLER_51_412 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_fill_1 FILLER_51_470 ();
 sg13g2_fill_2 FILLER_51_515 ();
 sg13g2_fill_2 FILLER_51_549 ();
 sg13g2_fill_1 FILLER_51_554 ();
 sg13g2_fill_2 FILLER_51_568 ();
 sg13g2_fill_1 FILLER_51_577 ();
 sg13g2_fill_1 FILLER_51_592 ();
 sg13g2_fill_2 FILLER_51_601 ();
 sg13g2_fill_2 FILLER_51_607 ();
 sg13g2_fill_2 FILLER_51_647 ();
 sg13g2_decap_8 FILLER_51_699 ();
 sg13g2_decap_8 FILLER_51_706 ();
 sg13g2_decap_8 FILLER_51_713 ();
 sg13g2_decap_8 FILLER_51_720 ();
 sg13g2_fill_2 FILLER_51_727 ();
 sg13g2_fill_1 FILLER_51_729 ();
 sg13g2_decap_4 FILLER_51_733 ();
 sg13g2_fill_1 FILLER_51_737 ();
 sg13g2_decap_4 FILLER_51_742 ();
 sg13g2_fill_2 FILLER_51_746 ();
 sg13g2_fill_1 FILLER_51_803 ();
 sg13g2_fill_1 FILLER_51_826 ();
 sg13g2_fill_1 FILLER_51_847 ();
 sg13g2_fill_2 FILLER_51_879 ();
 sg13g2_fill_1 FILLER_51_893 ();
 sg13g2_fill_1 FILLER_51_905 ();
 sg13g2_fill_2 FILLER_51_913 ();
 sg13g2_fill_1 FILLER_51_915 ();
 sg13g2_fill_2 FILLER_51_924 ();
 sg13g2_fill_1 FILLER_51_926 ();
 sg13g2_decap_4 FILLER_51_945 ();
 sg13g2_fill_1 FILLER_51_949 ();
 sg13g2_decap_4 FILLER_51_954 ();
 sg13g2_fill_2 FILLER_51_972 ();
 sg13g2_fill_1 FILLER_51_974 ();
 sg13g2_decap_8 FILLER_51_989 ();
 sg13g2_decap_4 FILLER_51_996 ();
 sg13g2_fill_2 FILLER_51_1000 ();
 sg13g2_decap_8 FILLER_51_1007 ();
 sg13g2_decap_8 FILLER_51_1014 ();
 sg13g2_decap_4 FILLER_51_1021 ();
 sg13g2_fill_2 FILLER_51_1059 ();
 sg13g2_fill_1 FILLER_51_1061 ();
 sg13g2_fill_2 FILLER_51_1145 ();
 sg13g2_fill_1 FILLER_51_1147 ();
 sg13g2_fill_2 FILLER_51_1192 ();
 sg13g2_fill_1 FILLER_51_1194 ();
 sg13g2_fill_2 FILLER_51_1221 ();
 sg13g2_fill_1 FILLER_51_1251 ();
 sg13g2_fill_1 FILLER_51_1279 ();
 sg13g2_fill_1 FILLER_51_1310 ();
 sg13g2_fill_1 FILLER_51_1351 ();
 sg13g2_fill_2 FILLER_51_1410 ();
 sg13g2_fill_1 FILLER_51_1420 ();
 sg13g2_fill_1 FILLER_51_1429 ();
 sg13g2_fill_1 FILLER_51_1445 ();
 sg13g2_fill_2 FILLER_51_1467 ();
 sg13g2_fill_1 FILLER_51_1540 ();
 sg13g2_fill_2 FILLER_51_1583 ();
 sg13g2_decap_4 FILLER_51_1627 ();
 sg13g2_fill_1 FILLER_51_1631 ();
 sg13g2_fill_2 FILLER_51_1636 ();
 sg13g2_fill_2 FILLER_51_1679 ();
 sg13g2_fill_2 FILLER_51_1692 ();
 sg13g2_fill_2 FILLER_51_1703 ();
 sg13g2_fill_1 FILLER_51_1715 ();
 sg13g2_fill_1 FILLER_51_1745 ();
 sg13g2_fill_1 FILLER_51_1750 ();
 sg13g2_fill_2 FILLER_51_1777 ();
 sg13g2_decap_8 FILLER_51_1822 ();
 sg13g2_decap_8 FILLER_51_1833 ();
 sg13g2_fill_2 FILLER_51_1840 ();
 sg13g2_fill_2 FILLER_51_1857 ();
 sg13g2_fill_1 FILLER_51_1859 ();
 sg13g2_fill_2 FILLER_51_1872 ();
 sg13g2_fill_1 FILLER_51_1874 ();
 sg13g2_fill_1 FILLER_51_1889 ();
 sg13g2_decap_8 FILLER_51_1905 ();
 sg13g2_decap_8 FILLER_51_1912 ();
 sg13g2_fill_2 FILLER_51_1919 ();
 sg13g2_decap_4 FILLER_51_1931 ();
 sg13g2_fill_1 FILLER_51_1935 ();
 sg13g2_decap_4 FILLER_51_1941 ();
 sg13g2_fill_2 FILLER_51_1974 ();
 sg13g2_fill_2 FILLER_51_2012 ();
 sg13g2_fill_2 FILLER_51_2040 ();
 sg13g2_fill_2 FILLER_51_2045 ();
 sg13g2_decap_8 FILLER_51_2051 ();
 sg13g2_decap_8 FILLER_51_2062 ();
 sg13g2_decap_8 FILLER_51_2069 ();
 sg13g2_fill_2 FILLER_51_2076 ();
 sg13g2_fill_1 FILLER_51_2082 ();
 sg13g2_fill_1 FILLER_51_2096 ();
 sg13g2_fill_1 FILLER_51_2101 ();
 sg13g2_fill_2 FILLER_51_2106 ();
 sg13g2_fill_2 FILLER_51_2116 ();
 sg13g2_fill_1 FILLER_51_2118 ();
 sg13g2_fill_2 FILLER_51_2140 ();
 sg13g2_fill_1 FILLER_51_2142 ();
 sg13g2_fill_2 FILLER_51_2156 ();
 sg13g2_fill_1 FILLER_51_2158 ();
 sg13g2_fill_1 FILLER_51_2189 ();
 sg13g2_decap_8 FILLER_51_2226 ();
 sg13g2_decap_4 FILLER_51_2233 ();
 sg13g2_fill_1 FILLER_51_2267 ();
 sg13g2_decap_4 FILLER_51_2278 ();
 sg13g2_decap_4 FILLER_51_2308 ();
 sg13g2_fill_2 FILLER_51_2312 ();
 sg13g2_decap_8 FILLER_51_2345 ();
 sg13g2_fill_1 FILLER_51_2352 ();
 sg13g2_decap_4 FILLER_51_2383 ();
 sg13g2_fill_1 FILLER_51_2387 ();
 sg13g2_decap_4 FILLER_51_2391 ();
 sg13g2_fill_1 FILLER_51_2395 ();
 sg13g2_decap_8 FILLER_51_2442 ();
 sg13g2_decap_4 FILLER_51_2449 ();
 sg13g2_decap_4 FILLER_51_2457 ();
 sg13g2_decap_8 FILLER_51_2465 ();
 sg13g2_fill_2 FILLER_51_2472 ();
 sg13g2_fill_1 FILLER_51_2474 ();
 sg13g2_decap_8 FILLER_51_2479 ();
 sg13g2_decap_8 FILLER_51_2486 ();
 sg13g2_fill_2 FILLER_51_2493 ();
 sg13g2_decap_8 FILLER_51_2534 ();
 sg13g2_decap_8 FILLER_51_2541 ();
 sg13g2_decap_8 FILLER_51_2548 ();
 sg13g2_fill_2 FILLER_51_2555 ();
 sg13g2_fill_1 FILLER_51_2557 ();
 sg13g2_decap_8 FILLER_51_2572 ();
 sg13g2_fill_2 FILLER_51_2579 ();
 sg13g2_fill_1 FILLER_51_2581 ();
 sg13g2_fill_2 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2652 ();
 sg13g2_decap_8 FILLER_51_2659 ();
 sg13g2_decap_4 FILLER_51_2666 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_1 FILLER_52_9 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_fill_1 FILLER_52_28 ();
 sg13g2_fill_1 FILLER_52_43 ();
 sg13g2_decap_8 FILLER_52_48 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_decap_8 FILLER_52_108 ();
 sg13g2_decap_8 FILLER_52_115 ();
 sg13g2_decap_8 FILLER_52_122 ();
 sg13g2_fill_2 FILLER_52_137 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_173 ();
 sg13g2_fill_2 FILLER_52_178 ();
 sg13g2_fill_1 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_239 ();
 sg13g2_fill_2 FILLER_52_246 ();
 sg13g2_decap_4 FILLER_52_253 ();
 sg13g2_fill_1 FILLER_52_257 ();
 sg13g2_fill_2 FILLER_52_306 ();
 sg13g2_fill_2 FILLER_52_312 ();
 sg13g2_fill_2 FILLER_52_361 ();
 sg13g2_fill_2 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_382 ();
 sg13g2_fill_1 FILLER_52_397 ();
 sg13g2_decap_4 FILLER_52_410 ();
 sg13g2_fill_2 FILLER_52_446 ();
 sg13g2_fill_1 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_459 ();
 sg13g2_decap_8 FILLER_52_466 ();
 sg13g2_fill_1 FILLER_52_473 ();
 sg13g2_fill_2 FILLER_52_512 ();
 sg13g2_fill_2 FILLER_52_521 ();
 sg13g2_fill_1 FILLER_52_532 ();
 sg13g2_fill_1 FILLER_52_560 ();
 sg13g2_fill_2 FILLER_52_578 ();
 sg13g2_fill_2 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_629 ();
 sg13g2_fill_2 FILLER_52_636 ();
 sg13g2_fill_2 FILLER_52_641 ();
 sg13g2_fill_2 FILLER_52_691 ();
 sg13g2_decap_8 FILLER_52_703 ();
 sg13g2_decap_8 FILLER_52_710 ();
 sg13g2_decap_8 FILLER_52_717 ();
 sg13g2_decap_4 FILLER_52_724 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_1 FILLER_52_759 ();
 sg13g2_fill_1 FILLER_52_770 ();
 sg13g2_fill_1 FILLER_52_781 ();
 sg13g2_fill_2 FILLER_52_786 ();
 sg13g2_fill_1 FILLER_52_794 ();
 sg13g2_fill_1 FILLER_52_806 ();
 sg13g2_fill_2 FILLER_52_815 ();
 sg13g2_fill_1 FILLER_52_826 ();
 sg13g2_fill_2 FILLER_52_830 ();
 sg13g2_fill_2 FILLER_52_870 ();
 sg13g2_fill_1 FILLER_52_872 ();
 sg13g2_decap_4 FILLER_52_877 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_fill_2 FILLER_52_889 ();
 sg13g2_fill_2 FILLER_52_981 ();
 sg13g2_decap_8 FILLER_52_1009 ();
 sg13g2_decap_8 FILLER_52_1016 ();
 sg13g2_decap_8 FILLER_52_1023 ();
 sg13g2_fill_2 FILLER_52_1030 ();
 sg13g2_fill_2 FILLER_52_1091 ();
 sg13g2_fill_1 FILLER_52_1093 ();
 sg13g2_fill_1 FILLER_52_1103 ();
 sg13g2_decap_8 FILLER_52_1125 ();
 sg13g2_decap_4 FILLER_52_1179 ();
 sg13g2_fill_2 FILLER_52_1183 ();
 sg13g2_fill_2 FILLER_52_1194 ();
 sg13g2_fill_1 FILLER_52_1196 ();
 sg13g2_fill_2 FILLER_52_1256 ();
 sg13g2_fill_1 FILLER_52_1263 ();
 sg13g2_fill_1 FILLER_52_1293 ();
 sg13g2_fill_1 FILLER_52_1324 ();
 sg13g2_fill_1 FILLER_52_1343 ();
 sg13g2_fill_2 FILLER_52_1409 ();
 sg13g2_fill_1 FILLER_52_1427 ();
 sg13g2_fill_2 FILLER_52_1451 ();
 sg13g2_fill_1 FILLER_52_1495 ();
 sg13g2_fill_1 FILLER_52_1518 ();
 sg13g2_fill_1 FILLER_52_1568 ();
 sg13g2_fill_1 FILLER_52_1593 ();
 sg13g2_fill_1 FILLER_52_1598 ();
 sg13g2_fill_1 FILLER_52_1607 ();
 sg13g2_decap_8 FILLER_52_1615 ();
 sg13g2_decap_4 FILLER_52_1622 ();
 sg13g2_decap_8 FILLER_52_1631 ();
 sg13g2_decap_4 FILLER_52_1638 ();
 sg13g2_fill_1 FILLER_52_1642 ();
 sg13g2_fill_1 FILLER_52_1654 ();
 sg13g2_fill_1 FILLER_52_1669 ();
 sg13g2_fill_2 FILLER_52_1675 ();
 sg13g2_fill_1 FILLER_52_1712 ();
 sg13g2_fill_1 FILLER_52_1718 ();
 sg13g2_decap_8 FILLER_52_1728 ();
 sg13g2_fill_2 FILLER_52_1740 ();
 sg13g2_fill_1 FILLER_52_1742 ();
 sg13g2_fill_1 FILLER_52_1750 ();
 sg13g2_fill_1 FILLER_52_1769 ();
 sg13g2_fill_1 FILLER_52_1775 ();
 sg13g2_fill_1 FILLER_52_1781 ();
 sg13g2_fill_1 FILLER_52_1799 ();
 sg13g2_decap_8 FILLER_52_1856 ();
 sg13g2_decap_4 FILLER_52_1863 ();
 sg13g2_decap_8 FILLER_52_1876 ();
 sg13g2_decap_8 FILLER_52_1883 ();
 sg13g2_decap_8 FILLER_52_1890 ();
 sg13g2_decap_8 FILLER_52_1901 ();
 sg13g2_decap_4 FILLER_52_1908 ();
 sg13g2_fill_1 FILLER_52_1912 ();
 sg13g2_decap_4 FILLER_52_1926 ();
 sg13g2_fill_2 FILLER_52_1930 ();
 sg13g2_fill_2 FILLER_52_1948 ();
 sg13g2_fill_2 FILLER_52_1956 ();
 sg13g2_fill_2 FILLER_52_1988 ();
 sg13g2_fill_1 FILLER_52_1990 ();
 sg13g2_fill_2 FILLER_52_2097 ();
 sg13g2_fill_1 FILLER_52_2099 ();
 sg13g2_decap_4 FILLER_52_2121 ();
 sg13g2_fill_1 FILLER_52_2125 ();
 sg13g2_fill_2 FILLER_52_2130 ();
 sg13g2_fill_1 FILLER_52_2162 ();
 sg13g2_decap_8 FILLER_52_2173 ();
 sg13g2_decap_8 FILLER_52_2180 ();
 sg13g2_decap_8 FILLER_52_2187 ();
 sg13g2_fill_1 FILLER_52_2194 ();
 sg13g2_fill_1 FILLER_52_2272 ();
 sg13g2_fill_2 FILLER_52_2309 ();
 sg13g2_fill_1 FILLER_52_2311 ();
 sg13g2_fill_1 FILLER_52_2338 ();
 sg13g2_decap_8 FILLER_52_2345 ();
 sg13g2_decap_8 FILLER_52_2352 ();
 sg13g2_fill_2 FILLER_52_2359 ();
 sg13g2_fill_1 FILLER_52_2361 ();
 sg13g2_decap_8 FILLER_52_2397 ();
 sg13g2_decap_8 FILLER_52_2404 ();
 sg13g2_decap_8 FILLER_52_2411 ();
 sg13g2_fill_2 FILLER_52_2418 ();
 sg13g2_fill_1 FILLER_52_2420 ();
 sg13g2_decap_8 FILLER_52_2425 ();
 sg13g2_fill_2 FILLER_52_2436 ();
 sg13g2_fill_1 FILLER_52_2469 ();
 sg13g2_decap_4 FILLER_52_2475 ();
 sg13g2_fill_1 FILLER_52_2479 ();
 sg13g2_decap_8 FILLER_52_2484 ();
 sg13g2_fill_2 FILLER_52_2491 ();
 sg13g2_decap_4 FILLER_52_2502 ();
 sg13g2_decap_8 FILLER_52_2510 ();
 sg13g2_decap_4 FILLER_52_2517 ();
 sg13g2_fill_2 FILLER_52_2521 ();
 sg13g2_decap_8 FILLER_52_2549 ();
 sg13g2_fill_2 FILLER_52_2556 ();
 sg13g2_fill_1 FILLER_52_2588 ();
 sg13g2_fill_1 FILLER_52_2619 ();
 sg13g2_fill_2 FILLER_52_2624 ();
 sg13g2_fill_2 FILLER_52_2630 ();
 sg13g2_fill_2 FILLER_52_2636 ();
 sg13g2_decap_4 FILLER_52_2664 ();
 sg13g2_fill_2 FILLER_52_2668 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_decap_4 FILLER_53_33 ();
 sg13g2_fill_1 FILLER_53_37 ();
 sg13g2_fill_1 FILLER_53_43 ();
 sg13g2_fill_1 FILLER_53_61 ();
 sg13g2_fill_1 FILLER_53_76 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_decap_4 FILLER_53_108 ();
 sg13g2_decap_8 FILLER_53_116 ();
 sg13g2_decap_4 FILLER_53_123 ();
 sg13g2_fill_2 FILLER_53_127 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_150 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_2 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_187 ();
 sg13g2_fill_2 FILLER_53_192 ();
 sg13g2_fill_1 FILLER_53_194 ();
 sg13g2_decap_4 FILLER_53_199 ();
 sg13g2_fill_1 FILLER_53_203 ();
 sg13g2_decap_4 FILLER_53_212 ();
 sg13g2_fill_2 FILLER_53_271 ();
 sg13g2_fill_1 FILLER_53_273 ();
 sg13g2_fill_1 FILLER_53_279 ();
 sg13g2_fill_2 FILLER_53_293 ();
 sg13g2_decap_4 FILLER_53_304 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_346 ();
 sg13g2_fill_1 FILLER_53_352 ();
 sg13g2_fill_2 FILLER_53_358 ();
 sg13g2_fill_2 FILLER_53_365 ();
 sg13g2_decap_8 FILLER_53_370 ();
 sg13g2_fill_2 FILLER_53_377 ();
 sg13g2_fill_1 FILLER_53_379 ();
 sg13g2_fill_2 FILLER_53_389 ();
 sg13g2_fill_1 FILLER_53_391 ();
 sg13g2_fill_2 FILLER_53_403 ();
 sg13g2_decap_4 FILLER_53_415 ();
 sg13g2_fill_1 FILLER_53_419 ();
 sg13g2_fill_1 FILLER_53_424 ();
 sg13g2_fill_2 FILLER_53_462 ();
 sg13g2_fill_1 FILLER_53_479 ();
 sg13g2_decap_4 FILLER_53_484 ();
 sg13g2_fill_2 FILLER_53_488 ();
 sg13g2_fill_1 FILLER_53_494 ();
 sg13g2_fill_1 FILLER_53_551 ();
 sg13g2_fill_1 FILLER_53_568 ();
 sg13g2_fill_1 FILLER_53_575 ();
 sg13g2_fill_1 FILLER_53_584 ();
 sg13g2_fill_1 FILLER_53_590 ();
 sg13g2_fill_1 FILLER_53_596 ();
 sg13g2_fill_1 FILLER_53_609 ();
 sg13g2_fill_1 FILLER_53_618 ();
 sg13g2_fill_2 FILLER_53_697 ();
 sg13g2_fill_1 FILLER_53_699 ();
 sg13g2_decap_4 FILLER_53_726 ();
 sg13g2_fill_2 FILLER_53_730 ();
 sg13g2_fill_1 FILLER_53_770 ();
 sg13g2_fill_1 FILLER_53_800 ();
 sg13g2_fill_2 FILLER_53_827 ();
 sg13g2_fill_1 FILLER_53_863 ();
 sg13g2_fill_2 FILLER_53_868 ();
 sg13g2_fill_1 FILLER_53_874 ();
 sg13g2_fill_1 FILLER_53_883 ();
 sg13g2_decap_4 FILLER_53_898 ();
 sg13g2_fill_1 FILLER_53_909 ();
 sg13g2_fill_2 FILLER_53_941 ();
 sg13g2_fill_1 FILLER_53_943 ();
 sg13g2_decap_4 FILLER_53_948 ();
 sg13g2_fill_2 FILLER_53_987 ();
 sg13g2_decap_8 FILLER_53_1022 ();
 sg13g2_fill_1 FILLER_53_1029 ();
 sg13g2_fill_1 FILLER_53_1092 ();
 sg13g2_decap_8 FILLER_53_1182 ();
 sg13g2_fill_2 FILLER_53_1189 ();
 sg13g2_fill_1 FILLER_53_1191 ();
 sg13g2_decap_8 FILLER_53_1205 ();
 sg13g2_fill_1 FILLER_53_1212 ();
 sg13g2_fill_2 FILLER_53_1351 ();
 sg13g2_fill_2 FILLER_53_1361 ();
 sg13g2_fill_1 FILLER_53_1372 ();
 sg13g2_fill_1 FILLER_53_1385 ();
 sg13g2_fill_1 FILLER_53_1400 ();
 sg13g2_fill_2 FILLER_53_1420 ();
 sg13g2_fill_2 FILLER_53_1452 ();
 sg13g2_fill_2 FILLER_53_1462 ();
 sg13g2_fill_1 FILLER_53_1487 ();
 sg13g2_fill_1 FILLER_53_1541 ();
 sg13g2_fill_1 FILLER_53_1567 ();
 sg13g2_fill_1 FILLER_53_1596 ();
 sg13g2_fill_2 FILLER_53_1627 ();
 sg13g2_fill_1 FILLER_53_1639 ();
 sg13g2_decap_8 FILLER_53_1644 ();
 sg13g2_fill_2 FILLER_53_1651 ();
 sg13g2_fill_1 FILLER_53_1653 ();
 sg13g2_fill_2 FILLER_53_1672 ();
 sg13g2_fill_2 FILLER_53_1696 ();
 sg13g2_decap_4 FILLER_53_1728 ();
 sg13g2_fill_2 FILLER_53_1799 ();
 sg13g2_fill_2 FILLER_53_1808 ();
 sg13g2_fill_1 FILLER_53_1810 ();
 sg13g2_decap_8 FILLER_53_1815 ();
 sg13g2_decap_4 FILLER_53_1822 ();
 sg13g2_decap_4 FILLER_53_1831 ();
 sg13g2_decap_4 FILLER_53_1845 ();
 sg13g2_decap_8 FILLER_53_1853 ();
 sg13g2_fill_2 FILLER_53_1860 ();
 sg13g2_decap_4 FILLER_53_1867 ();
 sg13g2_fill_1 FILLER_53_1901 ();
 sg13g2_fill_1 FILLER_53_1906 ();
 sg13g2_fill_1 FILLER_53_1936 ();
 sg13g2_fill_1 FILLER_53_1953 ();
 sg13g2_decap_8 FILLER_53_1980 ();
 sg13g2_decap_4 FILLER_53_1987 ();
 sg13g2_decap_4 FILLER_53_1995 ();
 sg13g2_decap_4 FILLER_53_2003 ();
 sg13g2_fill_2 FILLER_53_2007 ();
 sg13g2_fill_1 FILLER_53_2044 ();
 sg13g2_fill_1 FILLER_53_2076 ();
 sg13g2_fill_1 FILLER_53_2087 ();
 sg13g2_fill_1 FILLER_53_2114 ();
 sg13g2_fill_1 FILLER_53_2125 ();
 sg13g2_decap_4 FILLER_53_2152 ();
 sg13g2_fill_2 FILLER_53_2186 ();
 sg13g2_fill_2 FILLER_53_2192 ();
 sg13g2_fill_1 FILLER_53_2194 ();
 sg13g2_fill_1 FILLER_53_2225 ();
 sg13g2_decap_8 FILLER_53_2230 ();
 sg13g2_decap_8 FILLER_53_2237 ();
 sg13g2_decap_8 FILLER_53_2244 ();
 sg13g2_decap_4 FILLER_53_2255 ();
 sg13g2_fill_1 FILLER_53_2259 ();
 sg13g2_decap_4 FILLER_53_2270 ();
 sg13g2_fill_1 FILLER_53_2274 ();
 sg13g2_fill_2 FILLER_53_2315 ();
 sg13g2_fill_1 FILLER_53_2317 ();
 sg13g2_fill_2 FILLER_53_2351 ();
 sg13g2_decap_4 FILLER_53_2358 ();
 sg13g2_fill_1 FILLER_53_2362 ();
 sg13g2_decap_8 FILLER_53_2367 ();
 sg13g2_decap_4 FILLER_53_2374 ();
 sg13g2_fill_2 FILLER_53_2378 ();
 sg13g2_fill_1 FILLER_53_2390 ();
 sg13g2_decap_8 FILLER_53_2395 ();
 sg13g2_decap_4 FILLER_53_2410 ();
 sg13g2_fill_2 FILLER_53_2414 ();
 sg13g2_fill_1 FILLER_53_2420 ();
 sg13g2_fill_2 FILLER_53_2426 ();
 sg13g2_fill_1 FILLER_53_2428 ();
 sg13g2_fill_2 FILLER_53_2433 ();
 sg13g2_fill_1 FILLER_53_2539 ();
 sg13g2_fill_2 FILLER_53_2606 ();
 sg13g2_fill_2 FILLER_53_2668 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_32 ();
 sg13g2_fill_1 FILLER_54_34 ();
 sg13g2_fill_2 FILLER_54_40 ();
 sg13g2_fill_2 FILLER_54_59 ();
 sg13g2_fill_2 FILLER_54_87 ();
 sg13g2_fill_1 FILLER_54_89 ();
 sg13g2_decap_4 FILLER_54_116 ();
 sg13g2_fill_1 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_147 ();
 sg13g2_fill_2 FILLER_54_153 ();
 sg13g2_fill_2 FILLER_54_159 ();
 sg13g2_fill_2 FILLER_54_169 ();
 sg13g2_decap_4 FILLER_54_175 ();
 sg13g2_fill_2 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_4 FILLER_54_210 ();
 sg13g2_fill_1 FILLER_54_214 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_261 ();
 sg13g2_fill_1 FILLER_54_266 ();
 sg13g2_fill_2 FILLER_54_290 ();
 sg13g2_fill_1 FILLER_54_296 ();
 sg13g2_decap_8 FILLER_54_309 ();
 sg13g2_decap_8 FILLER_54_316 ();
 sg13g2_decap_8 FILLER_54_323 ();
 sg13g2_decap_8 FILLER_54_338 ();
 sg13g2_decap_8 FILLER_54_345 ();
 sg13g2_fill_1 FILLER_54_352 ();
 sg13g2_decap_8 FILLER_54_361 ();
 sg13g2_decap_8 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_375 ();
 sg13g2_fill_2 FILLER_54_386 ();
 sg13g2_fill_1 FILLER_54_388 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_fill_1 FILLER_54_404 ();
 sg13g2_fill_1 FILLER_54_424 ();
 sg13g2_fill_1 FILLER_54_448 ();
 sg13g2_fill_1 FILLER_54_489 ();
 sg13g2_fill_1 FILLER_54_558 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_2 FILLER_54_592 ();
 sg13g2_fill_1 FILLER_54_639 ();
 sg13g2_fill_2 FILLER_54_670 ();
 sg13g2_fill_2 FILLER_54_698 ();
 sg13g2_fill_1 FILLER_54_700 ();
 sg13g2_fill_2 FILLER_54_751 ();
 sg13g2_fill_2 FILLER_54_761 ();
 sg13g2_fill_1 FILLER_54_763 ();
 sg13g2_fill_2 FILLER_54_779 ();
 sg13g2_fill_1 FILLER_54_781 ();
 sg13g2_fill_1 FILLER_54_786 ();
 sg13g2_fill_1 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_818 ();
 sg13g2_fill_2 FILLER_54_823 ();
 sg13g2_decap_4 FILLER_54_859 ();
 sg13g2_fill_1 FILLER_54_863 ();
 sg13g2_decap_8 FILLER_54_874 ();
 sg13g2_decap_4 FILLER_54_881 ();
 sg13g2_fill_1 FILLER_54_885 ();
 sg13g2_fill_1 FILLER_54_895 ();
 sg13g2_fill_2 FILLER_54_901 ();
 sg13g2_fill_1 FILLER_54_903 ();
 sg13g2_decap_8 FILLER_54_908 ();
 sg13g2_fill_2 FILLER_54_922 ();
 sg13g2_fill_1 FILLER_54_924 ();
 sg13g2_fill_1 FILLER_54_929 ();
 sg13g2_decap_8 FILLER_54_940 ();
 sg13g2_decap_8 FILLER_54_947 ();
 sg13g2_decap_8 FILLER_54_954 ();
 sg13g2_decap_4 FILLER_54_965 ();
 sg13g2_decap_4 FILLER_54_977 ();
 sg13g2_decap_8 FILLER_54_986 ();
 sg13g2_fill_1 FILLER_54_993 ();
 sg13g2_fill_1 FILLER_54_999 ();
 sg13g2_fill_1 FILLER_54_1005 ();
 sg13g2_fill_2 FILLER_54_1027 ();
 sg13g2_fill_2 FILLER_54_1038 ();
 sg13g2_fill_1 FILLER_54_1040 ();
 sg13g2_decap_8 FILLER_54_1045 ();
 sg13g2_fill_1 FILLER_54_1056 ();
 sg13g2_fill_1 FILLER_54_1066 ();
 sg13g2_fill_1 FILLER_54_1086 ();
 sg13g2_fill_2 FILLER_54_1098 ();
 sg13g2_fill_1 FILLER_54_1100 ();
 sg13g2_fill_2 FILLER_54_1118 ();
 sg13g2_fill_1 FILLER_54_1132 ();
 sg13g2_decap_8 FILLER_54_1138 ();
 sg13g2_fill_2 FILLER_54_1145 ();
 sg13g2_fill_1 FILLER_54_1194 ();
 sg13g2_decap_8 FILLER_54_1200 ();
 sg13g2_decap_8 FILLER_54_1207 ();
 sg13g2_decap_4 FILLER_54_1214 ();
 sg13g2_fill_2 FILLER_54_1222 ();
 sg13g2_fill_1 FILLER_54_1244 ();
 sg13g2_fill_1 FILLER_54_1274 ();
 sg13g2_fill_2 FILLER_54_1282 ();
 sg13g2_fill_1 FILLER_54_1303 ();
 sg13g2_fill_2 FILLER_54_1315 ();
 sg13g2_fill_1 FILLER_54_1320 ();
 sg13g2_decap_4 FILLER_54_1333 ();
 sg13g2_decap_8 FILLER_54_1349 ();
 sg13g2_decap_8 FILLER_54_1356 ();
 sg13g2_decap_8 FILLER_54_1363 ();
 sg13g2_fill_2 FILLER_54_1370 ();
 sg13g2_fill_1 FILLER_54_1372 ();
 sg13g2_fill_2 FILLER_54_1392 ();
 sg13g2_fill_2 FILLER_54_1485 ();
 sg13g2_fill_1 FILLER_54_1521 ();
 sg13g2_fill_1 FILLER_54_1527 ();
 sg13g2_fill_2 FILLER_54_1536 ();
 sg13g2_fill_1 FILLER_54_1547 ();
 sg13g2_fill_2 FILLER_54_1573 ();
 sg13g2_fill_2 FILLER_54_1583 ();
 sg13g2_fill_1 FILLER_54_1626 ();
 sg13g2_fill_2 FILLER_54_1636 ();
 sg13g2_fill_2 FILLER_54_1642 ();
 sg13g2_fill_2 FILLER_54_1650 ();
 sg13g2_decap_4 FILLER_54_1660 ();
 sg13g2_fill_2 FILLER_54_1664 ();
 sg13g2_fill_2 FILLER_54_1695 ();
 sg13g2_decap_4 FILLER_54_1738 ();
 sg13g2_fill_1 FILLER_54_1742 ();
 sg13g2_fill_2 FILLER_54_1786 ();
 sg13g2_fill_1 FILLER_54_1788 ();
 sg13g2_fill_2 FILLER_54_1793 ();
 sg13g2_fill_1 FILLER_54_1795 ();
 sg13g2_decap_8 FILLER_54_1804 ();
 sg13g2_fill_2 FILLER_54_1811 ();
 sg13g2_decap_8 FILLER_54_1839 ();
 sg13g2_decap_8 FILLER_54_1846 ();
 sg13g2_decap_4 FILLER_54_1853 ();
 sg13g2_decap_8 FILLER_54_1864 ();
 sg13g2_decap_4 FILLER_54_1871 ();
 sg13g2_fill_1 FILLER_54_1875 ();
 sg13g2_decap_8 FILLER_54_1880 ();
 sg13g2_fill_2 FILLER_54_1887 ();
 sg13g2_fill_1 FILLER_54_1919 ();
 sg13g2_fill_2 FILLER_54_1926 ();
 sg13g2_decap_8 FILLER_54_1971 ();
 sg13g2_decap_8 FILLER_54_1978 ();
 sg13g2_decap_4 FILLER_54_1985 ();
 sg13g2_fill_2 FILLER_54_1989 ();
 sg13g2_fill_1 FILLER_54_2003 ();
 sg13g2_fill_2 FILLER_54_2013 ();
 sg13g2_fill_1 FILLER_54_2073 ();
 sg13g2_fill_1 FILLER_54_2095 ();
 sg13g2_fill_1 FILLER_54_2106 ();
 sg13g2_decap_4 FILLER_54_2142 ();
 sg13g2_fill_2 FILLER_54_2194 ();
 sg13g2_fill_1 FILLER_54_2196 ();
 sg13g2_decap_8 FILLER_54_2235 ();
 sg13g2_decap_8 FILLER_54_2242 ();
 sg13g2_decap_8 FILLER_54_2249 ();
 sg13g2_decap_8 FILLER_54_2256 ();
 sg13g2_decap_8 FILLER_54_2263 ();
 sg13g2_fill_1 FILLER_54_2270 ();
 sg13g2_fill_2 FILLER_54_2292 ();
 sg13g2_fill_1 FILLER_54_2294 ();
 sg13g2_decap_8 FILLER_54_2299 ();
 sg13g2_decap_4 FILLER_54_2306 ();
 sg13g2_fill_2 FILLER_54_2310 ();
 sg13g2_fill_1 FILLER_54_2315 ();
 sg13g2_fill_1 FILLER_54_2346 ();
 sg13g2_fill_1 FILLER_54_2372 ();
 sg13g2_fill_1 FILLER_54_2413 ();
 sg13g2_fill_2 FILLER_54_2422 ();
 sg13g2_fill_1 FILLER_54_2443 ();
 sg13g2_fill_2 FILLER_54_2452 ();
 sg13g2_fill_1 FILLER_54_2510 ();
 sg13g2_fill_1 FILLER_54_2524 ();
 sg13g2_fill_1 FILLER_54_2529 ();
 sg13g2_fill_2 FILLER_54_2561 ();
 sg13g2_decap_4 FILLER_54_2574 ();
 sg13g2_decap_8 FILLER_54_2582 ();
 sg13g2_decap_8 FILLER_54_2589 ();
 sg13g2_decap_8 FILLER_54_2600 ();
 sg13g2_decap_4 FILLER_54_2607 ();
 sg13g2_decap_8 FILLER_54_2624 ();
 sg13g2_fill_1 FILLER_54_2631 ();
 sg13g2_fill_2 FILLER_54_2640 ();
 sg13g2_fill_2 FILLER_54_2668 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_43 ();
 sg13g2_fill_2 FILLER_55_62 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_78 ();
 sg13g2_fill_2 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_decap_8 FILLER_55_122 ();
 sg13g2_decap_8 FILLER_55_136 ();
 sg13g2_decap_4 FILLER_55_143 ();
 sg13g2_fill_2 FILLER_55_147 ();
 sg13g2_decap_4 FILLER_55_153 ();
 sg13g2_fill_2 FILLER_55_157 ();
 sg13g2_decap_8 FILLER_55_170 ();
 sg13g2_fill_2 FILLER_55_177 ();
 sg13g2_fill_2 FILLER_55_204 ();
 sg13g2_fill_1 FILLER_55_235 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_decap_4 FILLER_55_253 ();
 sg13g2_fill_2 FILLER_55_257 ();
 sg13g2_decap_8 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_309 ();
 sg13g2_fill_1 FILLER_55_311 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_323 ();
 sg13g2_fill_1 FILLER_55_325 ();
 sg13g2_fill_2 FILLER_55_330 ();
 sg13g2_decap_8 FILLER_55_362 ();
 sg13g2_decap_8 FILLER_55_369 ();
 sg13g2_fill_2 FILLER_55_376 ();
 sg13g2_fill_1 FILLER_55_378 ();
 sg13g2_fill_2 FILLER_55_389 ();
 sg13g2_fill_1 FILLER_55_391 ();
 sg13g2_fill_2 FILLER_55_434 ();
 sg13g2_fill_1 FILLER_55_436 ();
 sg13g2_fill_2 FILLER_55_442 ();
 sg13g2_fill_1 FILLER_55_453 ();
 sg13g2_fill_2 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_465 ();
 sg13g2_fill_2 FILLER_55_470 ();
 sg13g2_fill_2 FILLER_55_476 ();
 sg13g2_decap_8 FILLER_55_483 ();
 sg13g2_fill_2 FILLER_55_490 ();
 sg13g2_fill_1 FILLER_55_492 ();
 sg13g2_fill_1 FILLER_55_506 ();
 sg13g2_fill_1 FILLER_55_533 ();
 sg13g2_fill_1 FILLER_55_537 ();
 sg13g2_fill_1 FILLER_55_551 ();
 sg13g2_fill_1 FILLER_55_561 ();
 sg13g2_fill_1 FILLER_55_580 ();
 sg13g2_fill_1 FILLER_55_601 ();
 sg13g2_fill_1 FILLER_55_607 ();
 sg13g2_fill_1 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_649 ();
 sg13g2_fill_2 FILLER_55_663 ();
 sg13g2_decap_4 FILLER_55_669 ();
 sg13g2_fill_1 FILLER_55_693 ();
 sg13g2_decap_8 FILLER_55_725 ();
 sg13g2_fill_2 FILLER_55_765 ();
 sg13g2_fill_1 FILLER_55_767 ();
 sg13g2_decap_4 FILLER_55_865 ();
 sg13g2_fill_1 FILLER_55_869 ();
 sg13g2_fill_1 FILLER_55_899 ();
 sg13g2_fill_2 FILLER_55_904 ();
 sg13g2_fill_1 FILLER_55_906 ();
 sg13g2_fill_2 FILLER_55_913 ();
 sg13g2_fill_1 FILLER_55_915 ();
 sg13g2_decap_8 FILLER_55_930 ();
 sg13g2_decap_8 FILLER_55_937 ();
 sg13g2_fill_2 FILLER_55_944 ();
 sg13g2_fill_1 FILLER_55_946 ();
 sg13g2_decap_4 FILLER_55_950 ();
 sg13g2_fill_1 FILLER_55_954 ();
 sg13g2_decap_8 FILLER_55_959 ();
 sg13g2_decap_8 FILLER_55_966 ();
 sg13g2_fill_2 FILLER_55_973 ();
 sg13g2_fill_1 FILLER_55_975 ();
 sg13g2_fill_2 FILLER_55_1002 ();
 sg13g2_fill_1 FILLER_55_1004 ();
 sg13g2_fill_1 FILLER_55_1009 ();
 sg13g2_decap_8 FILLER_55_1056 ();
 sg13g2_decap_4 FILLER_55_1063 ();
 sg13g2_fill_1 FILLER_55_1112 ();
 sg13g2_fill_2 FILLER_55_1116 ();
 sg13g2_decap_4 FILLER_55_1144 ();
 sg13g2_fill_1 FILLER_55_1148 ();
 sg13g2_fill_1 FILLER_55_1154 ();
 sg13g2_fill_2 FILLER_55_1159 ();
 sg13g2_fill_2 FILLER_55_1166 ();
 sg13g2_decap_8 FILLER_55_1211 ();
 sg13g2_decap_4 FILLER_55_1218 ();
 sg13g2_fill_2 FILLER_55_1222 ();
 sg13g2_fill_1 FILLER_55_1251 ();
 sg13g2_fill_2 FILLER_55_1256 ();
 sg13g2_fill_2 FILLER_55_1274 ();
 sg13g2_fill_2 FILLER_55_1280 ();
 sg13g2_fill_1 FILLER_55_1285 ();
 sg13g2_fill_1 FILLER_55_1315 ();
 sg13g2_fill_2 FILLER_55_1319 ();
 sg13g2_decap_4 FILLER_55_1330 ();
 sg13g2_decap_8 FILLER_55_1364 ();
 sg13g2_decap_8 FILLER_55_1371 ();
 sg13g2_decap_4 FILLER_55_1378 ();
 sg13g2_fill_2 FILLER_55_1412 ();
 sg13g2_fill_1 FILLER_55_1420 ();
 sg13g2_fill_2 FILLER_55_1466 ();
 sg13g2_fill_2 FILLER_55_1509 ();
 sg13g2_fill_2 FILLER_55_1518 ();
 sg13g2_fill_1 FILLER_55_1544 ();
 sg13g2_fill_1 FILLER_55_1554 ();
 sg13g2_fill_2 FILLER_55_1560 ();
 sg13g2_fill_1 FILLER_55_1584 ();
 sg13g2_fill_1 FILLER_55_1595 ();
 sg13g2_fill_1 FILLER_55_1601 ();
 sg13g2_fill_1 FILLER_55_1605 ();
 sg13g2_fill_1 FILLER_55_1635 ();
 sg13g2_decap_4 FILLER_55_1655 ();
 sg13g2_decap_8 FILLER_55_1685 ();
 sg13g2_fill_2 FILLER_55_1692 ();
 sg13g2_decap_8 FILLER_55_1704 ();
 sg13g2_decap_8 FILLER_55_1711 ();
 sg13g2_fill_1 FILLER_55_1718 ();
 sg13g2_decap_8 FILLER_55_1726 ();
 sg13g2_decap_8 FILLER_55_1733 ();
 sg13g2_decap_8 FILLER_55_1740 ();
 sg13g2_decap_8 FILLER_55_1751 ();
 sg13g2_fill_2 FILLER_55_1758 ();
 sg13g2_fill_1 FILLER_55_1760 ();
 sg13g2_fill_1 FILLER_55_1765 ();
 sg13g2_fill_1 FILLER_55_1771 ();
 sg13g2_decap_8 FILLER_55_1780 ();
 sg13g2_decap_8 FILLER_55_1795 ();
 sg13g2_decap_8 FILLER_55_1802 ();
 sg13g2_decap_8 FILLER_55_1809 ();
 sg13g2_decap_4 FILLER_55_1816 ();
 sg13g2_fill_1 FILLER_55_1824 ();
 sg13g2_fill_2 FILLER_55_1855 ();
 sg13g2_decap_4 FILLER_55_1888 ();
 sg13g2_fill_1 FILLER_55_1892 ();
 sg13g2_decap_8 FILLER_55_1898 ();
 sg13g2_fill_2 FILLER_55_1905 ();
 sg13g2_decap_8 FILLER_55_1965 ();
 sg13g2_decap_8 FILLER_55_1972 ();
 sg13g2_fill_2 FILLER_55_1979 ();
 sg13g2_fill_2 FILLER_55_2001 ();
 sg13g2_fill_1 FILLER_55_2003 ();
 sg13g2_fill_2 FILLER_55_2102 ();
 sg13g2_decap_8 FILLER_55_2114 ();
 sg13g2_decap_8 FILLER_55_2121 ();
 sg13g2_decap_8 FILLER_55_2128 ();
 sg13g2_decap_8 FILLER_55_2135 ();
 sg13g2_decap_8 FILLER_55_2142 ();
 sg13g2_decap_4 FILLER_55_2149 ();
 sg13g2_fill_2 FILLER_55_2153 ();
 sg13g2_decap_4 FILLER_55_2170 ();
 sg13g2_fill_1 FILLER_55_2174 ();
 sg13g2_fill_1 FILLER_55_2203 ();
 sg13g2_fill_2 FILLER_55_2247 ();
 sg13g2_fill_1 FILLER_55_2249 ();
 sg13g2_decap_4 FILLER_55_2254 ();
 sg13g2_fill_1 FILLER_55_2258 ();
 sg13g2_decap_8 FILLER_55_2290 ();
 sg13g2_decap_4 FILLER_55_2297 ();
 sg13g2_fill_2 FILLER_55_2301 ();
 sg13g2_fill_1 FILLER_55_2319 ();
 sg13g2_fill_1 FILLER_55_2335 ();
 sg13g2_fill_2 FILLER_55_2385 ();
 sg13g2_fill_1 FILLER_55_2447 ();
 sg13g2_fill_2 FILLER_55_2483 ();
 sg13g2_fill_1 FILLER_55_2485 ();
 sg13g2_decap_8 FILLER_55_2490 ();
 sg13g2_fill_1 FILLER_55_2497 ();
 sg13g2_decap_4 FILLER_55_2503 ();
 sg13g2_fill_2 FILLER_55_2507 ();
 sg13g2_decap_8 FILLER_55_2513 ();
 sg13g2_fill_2 FILLER_55_2520 ();
 sg13g2_fill_2 FILLER_55_2533 ();
 sg13g2_fill_2 FILLER_55_2544 ();
 sg13g2_fill_1 FILLER_55_2546 ();
 sg13g2_fill_2 FILLER_55_2552 ();
 sg13g2_decap_8 FILLER_55_2592 ();
 sg13g2_decap_8 FILLER_55_2599 ();
 sg13g2_decap_8 FILLER_55_2606 ();
 sg13g2_decap_8 FILLER_55_2613 ();
 sg13g2_decap_8 FILLER_55_2620 ();
 sg13g2_decap_8 FILLER_55_2627 ();
 sg13g2_fill_2 FILLER_55_2634 ();
 sg13g2_fill_1 FILLER_55_2636 ();
 sg13g2_decap_4 FILLER_55_2641 ();
 sg13g2_fill_1 FILLER_55_2645 ();
 sg13g2_decap_8 FILLER_55_2658 ();
 sg13g2_decap_4 FILLER_55_2665 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_decap_4 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_4 ();
 sg13g2_fill_1 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_59 ();
 sg13g2_fill_2 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_93 ();
 sg13g2_fill_1 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_138 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_1 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_217 ();
 sg13g2_fill_1 FILLER_56_219 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_fill_2 FILLER_56_231 ();
 sg13g2_fill_1 FILLER_56_233 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_250 ();
 sg13g2_decap_8 FILLER_56_255 ();
 sg13g2_decap_8 FILLER_56_262 ();
 sg13g2_decap_4 FILLER_56_269 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_314 ();
 sg13g2_fill_2 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_322 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_fill_1 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_339 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_2 FILLER_56_356 ();
 sg13g2_fill_1 FILLER_56_362 ();
 sg13g2_fill_2 FILLER_56_411 ();
 sg13g2_fill_1 FILLER_56_434 ();
 sg13g2_decap_4 FILLER_56_474 ();
 sg13g2_fill_2 FILLER_56_478 ();
 sg13g2_decap_8 FILLER_56_486 ();
 sg13g2_fill_1 FILLER_56_493 ();
 sg13g2_fill_1 FILLER_56_498 ();
 sg13g2_fill_1 FILLER_56_548 ();
 sg13g2_fill_1 FILLER_56_558 ();
 sg13g2_fill_2 FILLER_56_573 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_fill_2 FILLER_56_615 ();
 sg13g2_fill_2 FILLER_56_629 ();
 sg13g2_decap_8 FILLER_56_669 ();
 sg13g2_fill_2 FILLER_56_676 ();
 sg13g2_decap_4 FILLER_56_701 ();
 sg13g2_fill_2 FILLER_56_705 ();
 sg13g2_fill_2 FILLER_56_715 ();
 sg13g2_fill_1 FILLER_56_743 ();
 sg13g2_decap_4 FILLER_56_784 ();
 sg13g2_fill_2 FILLER_56_788 ();
 sg13g2_fill_1 FILLER_56_799 ();
 sg13g2_fill_2 FILLER_56_807 ();
 sg13g2_fill_1 FILLER_56_829 ();
 sg13g2_fill_2 FILLER_56_835 ();
 sg13g2_fill_1 FILLER_56_837 ();
 sg13g2_decap_8 FILLER_56_854 ();
 sg13g2_decap_8 FILLER_56_861 ();
 sg13g2_fill_2 FILLER_56_868 ();
 sg13g2_fill_1 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_886 ();
 sg13g2_fill_2 FILLER_56_931 ();
 sg13g2_fill_1 FILLER_56_940 ();
 sg13g2_fill_2 FILLER_56_944 ();
 sg13g2_fill_1 FILLER_56_964 ();
 sg13g2_fill_2 FILLER_56_981 ();
 sg13g2_fill_1 FILLER_56_987 ();
 sg13g2_fill_1 FILLER_56_992 ();
 sg13g2_decap_4 FILLER_56_1012 ();
 sg13g2_fill_1 FILLER_56_1016 ();
 sg13g2_decap_8 FILLER_56_1027 ();
 sg13g2_decap_4 FILLER_56_1034 ();
 sg13g2_decap_8 FILLER_56_1042 ();
 sg13g2_decap_4 FILLER_56_1049 ();
 sg13g2_fill_2 FILLER_56_1053 ();
 sg13g2_decap_4 FILLER_56_1068 ();
 sg13g2_fill_1 FILLER_56_1086 ();
 sg13g2_fill_2 FILLER_56_1120 ();
 sg13g2_fill_1 FILLER_56_1129 ();
 sg13g2_fill_1 FILLER_56_1139 ();
 sg13g2_decap_8 FILLER_56_1170 ();
 sg13g2_decap_8 FILLER_56_1177 ();
 sg13g2_fill_1 FILLER_56_1184 ();
 sg13g2_fill_2 FILLER_56_1206 ();
 sg13g2_fill_1 FILLER_56_1234 ();
 sg13g2_decap_4 FILLER_56_1256 ();
 sg13g2_fill_1 FILLER_56_1260 ();
 sg13g2_decap_8 FILLER_56_1329 ();
 sg13g2_fill_1 FILLER_56_1345 ();
 sg13g2_fill_1 FILLER_56_1402 ();
 sg13g2_fill_1 FILLER_56_1418 ();
 sg13g2_fill_2 FILLER_56_1428 ();
 sg13g2_fill_1 FILLER_56_1471 ();
 sg13g2_fill_1 FILLER_56_1482 ();
 sg13g2_fill_2 FILLER_56_1496 ();
 sg13g2_fill_1 FILLER_56_1514 ();
 sg13g2_fill_2 FILLER_56_1518 ();
 sg13g2_fill_1 FILLER_56_1530 ();
 sg13g2_fill_2 FILLER_56_1537 ();
 sg13g2_fill_1 FILLER_56_1560 ();
 sg13g2_fill_1 FILLER_56_1593 ();
 sg13g2_fill_2 FILLER_56_1623 ();
 sg13g2_fill_2 FILLER_56_1656 ();
 sg13g2_fill_1 FILLER_56_1658 ();
 sg13g2_fill_2 FILLER_56_1685 ();
 sg13g2_fill_1 FILLER_56_1687 ();
 sg13g2_fill_1 FILLER_56_1722 ();
 sg13g2_fill_2 FILLER_56_1733 ();
 sg13g2_decap_8 FILLER_56_1748 ();
 sg13g2_decap_4 FILLER_56_1755 ();
 sg13g2_decap_8 FILLER_56_1764 ();
 sg13g2_decap_8 FILLER_56_1771 ();
 sg13g2_fill_1 FILLER_56_1778 ();
 sg13g2_decap_8 FILLER_56_1783 ();
 sg13g2_decap_4 FILLER_56_1790 ();
 sg13g2_fill_2 FILLER_56_1804 ();
 sg13g2_decap_8 FILLER_56_1812 ();
 sg13g2_decap_8 FILLER_56_1819 ();
 sg13g2_fill_2 FILLER_56_1826 ();
 sg13g2_fill_1 FILLER_56_1828 ();
 sg13g2_decap_4 FILLER_56_1841 ();
 sg13g2_fill_2 FILLER_56_1845 ();
 sg13g2_fill_1 FILLER_56_1851 ();
 sg13g2_fill_2 FILLER_56_1878 ();
 sg13g2_fill_2 FILLER_56_1910 ();
 sg13g2_fill_1 FILLER_56_1912 ();
 sg13g2_decap_8 FILLER_56_1917 ();
 sg13g2_fill_1 FILLER_56_1946 ();
 sg13g2_fill_2 FILLER_56_1955 ();
 sg13g2_decap_8 FILLER_56_1961 ();
 sg13g2_decap_4 FILLER_56_1968 ();
 sg13g2_fill_1 FILLER_56_1972 ();
 sg13g2_fill_2 FILLER_56_2011 ();
 sg13g2_fill_1 FILLER_56_2013 ();
 sg13g2_fill_1 FILLER_56_2040 ();
 sg13g2_fill_2 FILLER_56_2066 ();
 sg13g2_fill_1 FILLER_56_2097 ();
 sg13g2_fill_2 FILLER_56_2134 ();
 sg13g2_decap_8 FILLER_56_2140 ();
 sg13g2_fill_2 FILLER_56_2147 ();
 sg13g2_decap_8 FILLER_56_2153 ();
 sg13g2_fill_1 FILLER_56_2160 ();
 sg13g2_fill_1 FILLER_56_2187 ();
 sg13g2_fill_2 FILLER_56_2210 ();
 sg13g2_decap_4 FILLER_56_2238 ();
 sg13g2_fill_2 FILLER_56_2242 ();
 sg13g2_decap_4 FILLER_56_2270 ();
 sg13g2_fill_1 FILLER_56_2274 ();
 sg13g2_decap_8 FILLER_56_2301 ();
 sg13g2_fill_2 FILLER_56_2308 ();
 sg13g2_fill_2 FILLER_56_2369 ();
 sg13g2_fill_1 FILLER_56_2397 ();
 sg13g2_fill_1 FILLER_56_2411 ();
 sg13g2_fill_1 FILLER_56_2438 ();
 sg13g2_fill_1 FILLER_56_2444 ();
 sg13g2_fill_1 FILLER_56_2471 ();
 sg13g2_fill_1 FILLER_56_2476 ();
 sg13g2_fill_2 FILLER_56_2485 ();
 sg13g2_fill_1 FILLER_56_2491 ();
 sg13g2_fill_1 FILLER_56_2547 ();
 sg13g2_decap_4 FILLER_56_2589 ();
 sg13g2_decap_8 FILLER_56_2633 ();
 sg13g2_decap_8 FILLER_56_2640 ();
 sg13g2_fill_2 FILLER_56_2647 ();
 sg13g2_decap_8 FILLER_56_2653 ();
 sg13g2_decap_8 FILLER_56_2660 ();
 sg13g2_fill_2 FILLER_56_2667 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_4 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_30 ();
 sg13g2_fill_1 FILLER_57_36 ();
 sg13g2_fill_2 FILLER_57_65 ();
 sg13g2_fill_2 FILLER_57_85 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_166 ();
 sg13g2_decap_4 FILLER_57_176 ();
 sg13g2_fill_2 FILLER_57_180 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_210 ();
 sg13g2_fill_1 FILLER_57_212 ();
 sg13g2_fill_2 FILLER_57_227 ();
 sg13g2_fill_1 FILLER_57_229 ();
 sg13g2_decap_4 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_decap_4 FILLER_57_279 ();
 sg13g2_fill_2 FILLER_57_283 ();
 sg13g2_decap_8 FILLER_57_290 ();
 sg13g2_decap_4 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_305 ();
 sg13g2_fill_2 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_348 ();
 sg13g2_decap_4 FILLER_57_364 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_2 FILLER_57_373 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_fill_2 FILLER_57_390 ();
 sg13g2_fill_1 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_398 ();
 sg13g2_fill_2 FILLER_57_409 ();
 sg13g2_fill_2 FILLER_57_416 ();
 sg13g2_decap_4 FILLER_57_422 ();
 sg13g2_fill_2 FILLER_57_435 ();
 sg13g2_fill_1 FILLER_57_437 ();
 sg13g2_fill_2 FILLER_57_455 ();
 sg13g2_fill_1 FILLER_57_457 ();
 sg13g2_fill_2 FILLER_57_508 ();
 sg13g2_fill_2 FILLER_57_560 ();
 sg13g2_fill_1 FILLER_57_588 ();
 sg13g2_fill_1 FILLER_57_619 ();
 sg13g2_fill_1 FILLER_57_623 ();
 sg13g2_fill_1 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_652 ();
 sg13g2_decap_8 FILLER_57_692 ();
 sg13g2_decap_8 FILLER_57_699 ();
 sg13g2_decap_8 FILLER_57_706 ();
 sg13g2_decap_8 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_720 ();
 sg13g2_fill_1 FILLER_57_749 ();
 sg13g2_fill_1 FILLER_57_759 ();
 sg13g2_fill_2 FILLER_57_773 ();
 sg13g2_fill_1 FILLER_57_775 ();
 sg13g2_fill_2 FILLER_57_780 ();
 sg13g2_fill_1 FILLER_57_818 ();
 sg13g2_fill_2 FILLER_57_825 ();
 sg13g2_fill_2 FILLER_57_863 ();
 sg13g2_fill_1 FILLER_57_865 ();
 sg13g2_fill_1 FILLER_57_879 ();
 sg13g2_fill_2 FILLER_57_890 ();
 sg13g2_fill_1 FILLER_57_897 ();
 sg13g2_fill_2 FILLER_57_907 ();
 sg13g2_fill_1 FILLER_57_920 ();
 sg13g2_fill_1 FILLER_57_982 ();
 sg13g2_fill_1 FILLER_57_992 ();
 sg13g2_fill_1 FILLER_57_1008 ();
 sg13g2_fill_1 FILLER_57_1022 ();
 sg13g2_fill_2 FILLER_57_1026 ();
 sg13g2_fill_2 FILLER_57_1070 ();
 sg13g2_fill_1 FILLER_57_1072 ();
 sg13g2_decap_8 FILLER_57_1146 ();
 sg13g2_decap_8 FILLER_57_1153 ();
 sg13g2_decap_4 FILLER_57_1160 ();
 sg13g2_fill_1 FILLER_57_1164 ();
 sg13g2_fill_1 FILLER_57_1191 ();
 sg13g2_fill_1 FILLER_57_1202 ();
 sg13g2_fill_1 FILLER_57_1229 ();
 sg13g2_fill_2 FILLER_57_1240 ();
 sg13g2_decap_8 FILLER_57_1246 ();
 sg13g2_decap_4 FILLER_57_1282 ();
 sg13g2_fill_2 FILLER_57_1293 ();
 sg13g2_decap_4 FILLER_57_1324 ();
 sg13g2_fill_1 FILLER_57_1328 ();
 sg13g2_fill_1 FILLER_57_1338 ();
 sg13g2_fill_1 FILLER_57_1342 ();
 sg13g2_decap_4 FILLER_57_1365 ();
 sg13g2_fill_1 FILLER_57_1369 ();
 sg13g2_fill_2 FILLER_57_1453 ();
 sg13g2_fill_2 FILLER_57_1511 ();
 sg13g2_fill_2 FILLER_57_1530 ();
 sg13g2_fill_2 FILLER_57_1605 ();
 sg13g2_fill_2 FILLER_57_1628 ();
 sg13g2_fill_1 FILLER_57_1640 ();
 sg13g2_fill_1 FILLER_57_1645 ();
 sg13g2_fill_1 FILLER_57_1666 ();
 sg13g2_fill_2 FILLER_57_1671 ();
 sg13g2_fill_1 FILLER_57_1673 ();
 sg13g2_fill_1 FILLER_57_1725 ();
 sg13g2_decap_8 FILLER_57_1730 ();
 sg13g2_decap_8 FILLER_57_1741 ();
 sg13g2_decap_8 FILLER_57_1748 ();
 sg13g2_decap_8 FILLER_57_1755 ();
 sg13g2_decap_8 FILLER_57_1762 ();
 sg13g2_decap_8 FILLER_57_1769 ();
 sg13g2_fill_2 FILLER_57_1776 ();
 sg13g2_fill_1 FILLER_57_1783 ();
 sg13g2_fill_1 FILLER_57_1804 ();
 sg13g2_fill_2 FILLER_57_1810 ();
 sg13g2_fill_1 FILLER_57_1812 ();
 sg13g2_decap_8 FILLER_57_1828 ();
 sg13g2_fill_1 FILLER_57_1835 ();
 sg13g2_fill_1 FILLER_57_1840 ();
 sg13g2_fill_1 FILLER_57_1867 ();
 sg13g2_decap_8 FILLER_57_1872 ();
 sg13g2_fill_2 FILLER_57_1886 ();
 sg13g2_fill_2 FILLER_57_1892 ();
 sg13g2_fill_2 FILLER_57_1927 ();
 sg13g2_fill_1 FILLER_57_1935 ();
 sg13g2_fill_1 FILLER_57_1943 ();
 sg13g2_fill_1 FILLER_57_1970 ();
 sg13g2_fill_2 FILLER_57_1997 ();
 sg13g2_fill_1 FILLER_57_1999 ();
 sg13g2_decap_4 FILLER_57_2034 ();
 sg13g2_decap_8 FILLER_57_2048 ();
 sg13g2_fill_1 FILLER_57_2081 ();
 sg13g2_fill_1 FILLER_57_2087 ();
 sg13g2_decap_4 FILLER_57_2121 ();
 sg13g2_decap_8 FILLER_57_2233 ();
 sg13g2_decap_4 FILLER_57_2240 ();
 sg13g2_fill_2 FILLER_57_2244 ();
 sg13g2_decap_4 FILLER_57_2256 ();
 sg13g2_fill_2 FILLER_57_2260 ();
 sg13g2_decap_8 FILLER_57_2309 ();
 sg13g2_fill_1 FILLER_57_2325 ();
 sg13g2_fill_2 FILLER_57_2386 ();
 sg13g2_fill_1 FILLER_57_2388 ();
 sg13g2_fill_2 FILLER_57_2394 ();
 sg13g2_fill_1 FILLER_57_2396 ();
 sg13g2_decap_4 FILLER_57_2407 ();
 sg13g2_decap_8 FILLER_57_2424 ();
 sg13g2_fill_2 FILLER_57_2431 ();
 sg13g2_fill_1 FILLER_57_2439 ();
 sg13g2_fill_2 FILLER_57_2449 ();
 sg13g2_fill_1 FILLER_57_2451 ();
 sg13g2_fill_1 FILLER_57_2524 ();
 sg13g2_fill_1 FILLER_57_2641 ();
 sg13g2_fill_2 FILLER_57_2668 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_13 ();
 sg13g2_fill_2 FILLER_58_20 ();
 sg13g2_fill_1 FILLER_58_22 ();
 sg13g2_fill_2 FILLER_58_26 ();
 sg13g2_fill_1 FILLER_58_28 ();
 sg13g2_fill_2 FILLER_58_89 ();
 sg13g2_fill_2 FILLER_58_97 ();
 sg13g2_fill_2 FILLER_58_108 ();
 sg13g2_fill_1 FILLER_58_110 ();
 sg13g2_fill_2 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_190 ();
 sg13g2_fill_1 FILLER_58_197 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_fill_1 FILLER_58_218 ();
 sg13g2_fill_1 FILLER_58_231 ();
 sg13g2_decap_4 FILLER_58_263 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_decap_8 FILLER_58_272 ();
 sg13g2_decap_4 FILLER_58_279 ();
 sg13g2_fill_1 FILLER_58_283 ();
 sg13g2_decap_8 FILLER_58_289 ();
 sg13g2_decap_4 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_300 ();
 sg13g2_decap_4 FILLER_58_342 ();
 sg13g2_fill_1 FILLER_58_346 ();
 sg13g2_decap_8 FILLER_58_387 ();
 sg13g2_fill_2 FILLER_58_450 ();
 sg13g2_fill_2 FILLER_58_471 ();
 sg13g2_fill_1 FILLER_58_477 ();
 sg13g2_decap_8 FILLER_58_486 ();
 sg13g2_fill_1 FILLER_58_523 ();
 sg13g2_fill_1 FILLER_58_529 ();
 sg13g2_fill_1 FILLER_58_535 ();
 sg13g2_fill_1 FILLER_58_570 ();
 sg13g2_decap_4 FILLER_58_582 ();
 sg13g2_fill_1 FILLER_58_590 ();
 sg13g2_fill_1 FILLER_58_595 ();
 sg13g2_fill_1 FILLER_58_604 ();
 sg13g2_fill_2 FILLER_58_620 ();
 sg13g2_decap_8 FILLER_58_655 ();
 sg13g2_fill_1 FILLER_58_662 ();
 sg13g2_decap_8 FILLER_58_666 ();
 sg13g2_decap_4 FILLER_58_677 ();
 sg13g2_fill_1 FILLER_58_681 ();
 sg13g2_decap_8 FILLER_58_688 ();
 sg13g2_decap_4 FILLER_58_695 ();
 sg13g2_decap_8 FILLER_58_703 ();
 sg13g2_decap_4 FILLER_58_710 ();
 sg13g2_fill_2 FILLER_58_714 ();
 sg13g2_fill_2 FILLER_58_742 ();
 sg13g2_fill_2 FILLER_58_759 ();
 sg13g2_fill_1 FILLER_58_761 ();
 sg13g2_fill_2 FILLER_58_766 ();
 sg13g2_fill_2 FILLER_58_778 ();
 sg13g2_fill_1 FILLER_58_780 ();
 sg13g2_fill_2 FILLER_58_817 ();
 sg13g2_fill_1 FILLER_58_819 ();
 sg13g2_fill_1 FILLER_58_826 ();
 sg13g2_fill_2 FILLER_58_831 ();
 sg13g2_fill_1 FILLER_58_833 ();
 sg13g2_fill_2 FILLER_58_870 ();
 sg13g2_fill_1 FILLER_58_904 ();
 sg13g2_fill_1 FILLER_58_919 ();
 sg13g2_fill_1 FILLER_58_950 ();
 sg13g2_fill_2 FILLER_58_954 ();
 sg13g2_fill_2 FILLER_58_1005 ();
 sg13g2_decap_8 FILLER_58_1066 ();
 sg13g2_decap_4 FILLER_58_1073 ();
 sg13g2_fill_2 FILLER_58_1124 ();
 sg13g2_fill_1 FILLER_58_1166 ();
 sg13g2_decap_8 FILLER_58_1197 ();
 sg13g2_fill_2 FILLER_58_1204 ();
 sg13g2_fill_1 FILLER_58_1206 ();
 sg13g2_fill_2 FILLER_58_1211 ();
 sg13g2_fill_1 FILLER_58_1213 ();
 sg13g2_decap_8 FILLER_58_1218 ();
 sg13g2_decap_8 FILLER_58_1265 ();
 sg13g2_decap_8 FILLER_58_1272 ();
 sg13g2_fill_1 FILLER_58_1279 ();
 sg13g2_fill_1 FILLER_58_1293 ();
 sg13g2_fill_1 FILLER_58_1304 ();
 sg13g2_fill_2 FILLER_58_1342 ();
 sg13g2_fill_1 FILLER_58_1360 ();
 sg13g2_fill_1 FILLER_58_1370 ();
 sg13g2_fill_1 FILLER_58_1376 ();
 sg13g2_decap_8 FILLER_58_1387 ();
 sg13g2_fill_1 FILLER_58_1394 ();
 sg13g2_fill_1 FILLER_58_1440 ();
 sg13g2_fill_1 FILLER_58_1474 ();
 sg13g2_fill_1 FILLER_58_1485 ();
 sg13g2_fill_2 FILLER_58_1502 ();
 sg13g2_fill_2 FILLER_58_1545 ();
 sg13g2_fill_2 FILLER_58_1554 ();
 sg13g2_decap_4 FILLER_58_1561 ();
 sg13g2_fill_1 FILLER_58_1565 ();
 sg13g2_fill_1 FILLER_58_1571 ();
 sg13g2_fill_1 FILLER_58_1580 ();
 sg13g2_fill_2 FILLER_58_1610 ();
 sg13g2_fill_2 FILLER_58_1643 ();
 sg13g2_fill_1 FILLER_58_1658 ();
 sg13g2_fill_1 FILLER_58_1701 ();
 sg13g2_fill_2 FILLER_58_1707 ();
 sg13g2_fill_1 FILLER_58_1709 ();
 sg13g2_decap_8 FILLER_58_1745 ();
 sg13g2_decap_8 FILLER_58_1752 ();
 sg13g2_decap_8 FILLER_58_1759 ();
 sg13g2_fill_2 FILLER_58_1766 ();
 sg13g2_decap_4 FILLER_58_1781 ();
 sg13g2_fill_1 FILLER_58_1828 ();
 sg13g2_decap_4 FILLER_58_1834 ();
 sg13g2_fill_1 FILLER_58_1838 ();
 sg13g2_decap_4 FILLER_58_1854 ();
 sg13g2_decap_8 FILLER_58_1871 ();
 sg13g2_decap_4 FILLER_58_1878 ();
 sg13g2_fill_2 FILLER_58_1893 ();
 sg13g2_decap_8 FILLER_58_1921 ();
 sg13g2_fill_1 FILLER_58_1928 ();
 sg13g2_fill_2 FILLER_58_1936 ();
 sg13g2_fill_1 FILLER_58_1938 ();
 sg13g2_decap_8 FILLER_58_1965 ();
 sg13g2_decap_8 FILLER_58_1972 ();
 sg13g2_fill_1 FILLER_58_1979 ();
 sg13g2_decap_4 FILLER_58_2016 ();
 sg13g2_fill_1 FILLER_58_2020 ();
 sg13g2_fill_1 FILLER_58_2025 ();
 sg13g2_decap_4 FILLER_58_2035 ();
 sg13g2_decap_8 FILLER_58_2069 ();
 sg13g2_fill_2 FILLER_58_2130 ();
 sg13g2_fill_1 FILLER_58_2132 ();
 sg13g2_decap_4 FILLER_58_2164 ();
 sg13g2_fill_1 FILLER_58_2168 ();
 sg13g2_decap_8 FILLER_58_2173 ();
 sg13g2_fill_2 FILLER_58_2180 ();
 sg13g2_fill_1 FILLER_58_2182 ();
 sg13g2_fill_1 FILLER_58_2223 ();
 sg13g2_decap_8 FILLER_58_2234 ();
 sg13g2_fill_2 FILLER_58_2241 ();
 sg13g2_fill_1 FILLER_58_2243 ();
 sg13g2_fill_2 FILLER_58_2270 ();
 sg13g2_fill_1 FILLER_58_2303 ();
 sg13g2_fill_2 FILLER_58_2314 ();
 sg13g2_fill_1 FILLER_58_2316 ();
 sg13g2_fill_1 FILLER_58_2363 ();
 sg13g2_fill_1 FILLER_58_2378 ();
 sg13g2_fill_1 FILLER_58_2394 ();
 sg13g2_decap_8 FILLER_58_2402 ();
 sg13g2_decap_4 FILLER_58_2409 ();
 sg13g2_fill_2 FILLER_58_2413 ();
 sg13g2_decap_8 FILLER_58_2420 ();
 sg13g2_decap_4 FILLER_58_2427 ();
 sg13g2_decap_8 FILLER_58_2435 ();
 sg13g2_decap_8 FILLER_58_2442 ();
 sg13g2_fill_2 FILLER_58_2449 ();
 sg13g2_fill_1 FILLER_58_2451 ();
 sg13g2_fill_2 FILLER_58_2491 ();
 sg13g2_fill_1 FILLER_58_2597 ();
 sg13g2_fill_2 FILLER_58_2604 ();
 sg13g2_fill_2 FILLER_58_2668 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_34 ();
 sg13g2_fill_2 FILLER_59_41 ();
 sg13g2_fill_2 FILLER_59_48 ();
 sg13g2_fill_2 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_135 ();
 sg13g2_fill_1 FILLER_59_140 ();
 sg13g2_fill_1 FILLER_59_146 ();
 sg13g2_fill_1 FILLER_59_162 ();
 sg13g2_fill_1 FILLER_59_179 ();
 sg13g2_fill_2 FILLER_59_184 ();
 sg13g2_fill_1 FILLER_59_193 ();
 sg13g2_fill_2 FILLER_59_207 ();
 sg13g2_fill_2 FILLER_59_221 ();
 sg13g2_fill_1 FILLER_59_223 ();
 sg13g2_fill_2 FILLER_59_237 ();
 sg13g2_fill_1 FILLER_59_239 ();
 sg13g2_decap_8 FILLER_59_248 ();
 sg13g2_decap_8 FILLER_59_255 ();
 sg13g2_decap_4 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_270 ();
 sg13g2_fill_1 FILLER_59_274 ();
 sg13g2_fill_1 FILLER_59_279 ();
 sg13g2_fill_2 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_290 ();
 sg13g2_fill_2 FILLER_59_305 ();
 sg13g2_decap_4 FILLER_59_311 ();
 sg13g2_decap_4 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_decap_4 FILLER_59_341 ();
 sg13g2_fill_1 FILLER_59_371 ();
 sg13g2_fill_2 FILLER_59_376 ();
 sg13g2_fill_1 FILLER_59_378 ();
 sg13g2_fill_2 FILLER_59_391 ();
 sg13g2_fill_1 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_419 ();
 sg13g2_fill_2 FILLER_59_449 ();
 sg13g2_decap_8 FILLER_59_477 ();
 sg13g2_decap_8 FILLER_59_484 ();
 sg13g2_decap_4 FILLER_59_491 ();
 sg13g2_fill_1 FILLER_59_495 ();
 sg13g2_fill_2 FILLER_59_501 ();
 sg13g2_fill_1 FILLER_59_503 ();
 sg13g2_fill_1 FILLER_59_516 ();
 sg13g2_fill_1 FILLER_59_522 ();
 sg13g2_fill_1 FILLER_59_554 ();
 sg13g2_fill_2 FILLER_59_559 ();
 sg13g2_fill_1 FILLER_59_568 ();
 sg13g2_fill_2 FILLER_59_586 ();
 sg13g2_fill_2 FILLER_59_592 ();
 sg13g2_fill_1 FILLER_59_606 ();
 sg13g2_fill_1 FILLER_59_650 ();
 sg13g2_fill_1 FILLER_59_654 ();
 sg13g2_fill_1 FILLER_59_658 ();
 sg13g2_fill_2 FILLER_59_664 ();
 sg13g2_fill_1 FILLER_59_692 ();
 sg13g2_decap_8 FILLER_59_699 ();
 sg13g2_fill_1 FILLER_59_706 ();
 sg13g2_fill_2 FILLER_59_713 ();
 sg13g2_fill_2 FILLER_59_719 ();
 sg13g2_decap_4 FILLER_59_763 ();
 sg13g2_fill_1 FILLER_59_767 ();
 sg13g2_fill_2 FILLER_59_772 ();
 sg13g2_decap_8 FILLER_59_779 ();
 sg13g2_fill_2 FILLER_59_790 ();
 sg13g2_fill_1 FILLER_59_792 ();
 sg13g2_fill_1 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_fill_2 FILLER_59_841 ();
 sg13g2_fill_1 FILLER_59_843 ();
 sg13g2_decap_4 FILLER_59_848 ();
 sg13g2_fill_1 FILLER_59_868 ();
 sg13g2_fill_1 FILLER_59_874 ();
 sg13g2_fill_2 FILLER_59_891 ();
 sg13g2_fill_1 FILLER_59_935 ();
 sg13g2_fill_1 FILLER_59_940 ();
 sg13g2_fill_1 FILLER_59_962 ();
 sg13g2_fill_2 FILLER_59_968 ();
 sg13g2_fill_1 FILLER_59_984 ();
 sg13g2_fill_1 FILLER_59_992 ();
 sg13g2_fill_2 FILLER_59_1073 ();
 sg13g2_fill_1 FILLER_59_1075 ();
 sg13g2_fill_2 FILLER_59_1129 ();
 sg13g2_fill_1 FILLER_59_1157 ();
 sg13g2_fill_1 FILLER_59_1163 ();
 sg13g2_fill_2 FILLER_59_1169 ();
 sg13g2_fill_1 FILLER_59_1175 ();
 sg13g2_decap_4 FILLER_59_1180 ();
 sg13g2_fill_2 FILLER_59_1184 ();
 sg13g2_fill_2 FILLER_59_1190 ();
 sg13g2_fill_1 FILLER_59_1192 ();
 sg13g2_decap_8 FILLER_59_1233 ();
 sg13g2_decap_4 FILLER_59_1240 ();
 sg13g2_decap_8 FILLER_59_1257 ();
 sg13g2_decap_8 FILLER_59_1264 ();
 sg13g2_decap_8 FILLER_59_1271 ();
 sg13g2_fill_1 FILLER_59_1278 ();
 sg13g2_fill_1 FILLER_59_1332 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_fill_1 FILLER_59_1377 ();
 sg13g2_decap_8 FILLER_59_1390 ();
 sg13g2_fill_2 FILLER_59_1402 ();
 sg13g2_fill_2 FILLER_59_1477 ();
 sg13g2_fill_2 FILLER_59_1485 ();
 sg13g2_fill_1 FILLER_59_1487 ();
 sg13g2_fill_2 FILLER_59_1518 ();
 sg13g2_fill_1 FILLER_59_1524 ();
 sg13g2_fill_2 FILLER_59_1530 ();
 sg13g2_decap_8 FILLER_59_1539 ();
 sg13g2_decap_4 FILLER_59_1546 ();
 sg13g2_fill_1 FILLER_59_1604 ();
 sg13g2_fill_1 FILLER_59_1610 ();
 sg13g2_fill_2 FILLER_59_1637 ();
 sg13g2_fill_1 FILLER_59_1667 ();
 sg13g2_fill_2 FILLER_59_1672 ();
 sg13g2_decap_8 FILLER_59_1686 ();
 sg13g2_fill_1 FILLER_59_1693 ();
 sg13g2_fill_2 FILLER_59_1703 ();
 sg13g2_fill_1 FILLER_59_1705 ();
 sg13g2_decap_8 FILLER_59_1758 ();
 sg13g2_decap_8 FILLER_59_1765 ();
 sg13g2_decap_8 FILLER_59_1772 ();
 sg13g2_decap_4 FILLER_59_1779 ();
 sg13g2_fill_1 FILLER_59_1783 ();
 sg13g2_fill_1 FILLER_59_1797 ();
 sg13g2_decap_4 FILLER_59_1803 ();
 sg13g2_fill_1 FILLER_59_1807 ();
 sg13g2_fill_2 FILLER_59_1813 ();
 sg13g2_fill_1 FILLER_59_1815 ();
 sg13g2_decap_8 FILLER_59_1836 ();
 sg13g2_fill_2 FILLER_59_1843 ();
 sg13g2_fill_1 FILLER_59_1845 ();
 sg13g2_fill_2 FILLER_59_1857 ();
 sg13g2_decap_4 FILLER_59_1863 ();
 sg13g2_fill_1 FILLER_59_1867 ();
 sg13g2_fill_1 FILLER_59_1872 ();
 sg13g2_fill_2 FILLER_59_1877 ();
 sg13g2_fill_2 FILLER_59_1884 ();
 sg13g2_decap_8 FILLER_59_1916 ();
 sg13g2_decap_8 FILLER_59_1923 ();
 sg13g2_fill_1 FILLER_59_1930 ();
 sg13g2_decap_8 FILLER_59_1962 ();
 sg13g2_decap_8 FILLER_59_1969 ();
 sg13g2_decap_8 FILLER_59_1976 ();
 sg13g2_fill_1 FILLER_59_1983 ();
 sg13g2_decap_8 FILLER_59_1988 ();
 sg13g2_decap_8 FILLER_59_1995 ();
 sg13g2_decap_8 FILLER_59_2002 ();
 sg13g2_decap_8 FILLER_59_2009 ();
 sg13g2_decap_8 FILLER_59_2016 ();
 sg13g2_decap_8 FILLER_59_2023 ();
 sg13g2_decap_8 FILLER_59_2030 ();
 sg13g2_decap_8 FILLER_59_2037 ();
 sg13g2_fill_2 FILLER_59_2044 ();
 sg13g2_fill_1 FILLER_59_2046 ();
 sg13g2_decap_4 FILLER_59_2061 ();
 sg13g2_fill_2 FILLER_59_2065 ();
 sg13g2_fill_2 FILLER_59_2103 ();
 sg13g2_fill_2 FILLER_59_2124 ();
 sg13g2_decap_8 FILLER_59_2162 ();
 sg13g2_decap_8 FILLER_59_2169 ();
 sg13g2_decap_8 FILLER_59_2176 ();
 sg13g2_decap_8 FILLER_59_2183 ();
 sg13g2_decap_8 FILLER_59_2190 ();
 sg13g2_decap_8 FILLER_59_2197 ();
 sg13g2_decap_4 FILLER_59_2204 ();
 sg13g2_decap_8 FILLER_59_2212 ();
 sg13g2_decap_8 FILLER_59_2219 ();
 sg13g2_decap_4 FILLER_59_2226 ();
 sg13g2_fill_2 FILLER_59_2230 ();
 sg13g2_decap_4 FILLER_59_2258 ();
 sg13g2_fill_2 FILLER_59_2266 ();
 sg13g2_fill_1 FILLER_59_2268 ();
 sg13g2_fill_2 FILLER_59_2295 ();
 sg13g2_fill_2 FILLER_59_2349 ();
 sg13g2_fill_1 FILLER_59_2394 ();
 sg13g2_fill_1 FILLER_59_2400 ();
 sg13g2_decap_8 FILLER_59_2407 ();
 sg13g2_fill_1 FILLER_59_2440 ();
 sg13g2_fill_1 FILLER_59_2446 ();
 sg13g2_decap_4 FILLER_59_2483 ();
 sg13g2_fill_2 FILLER_59_2487 ();
 sg13g2_fill_1 FILLER_59_2493 ();
 sg13g2_fill_2 FILLER_59_2528 ();
 sg13g2_fill_2 FILLER_59_2539 ();
 sg13g2_decap_4 FILLER_59_2545 ();
 sg13g2_fill_1 FILLER_59_2549 ();
 sg13g2_fill_1 FILLER_59_2558 ();
 sg13g2_fill_1 FILLER_59_2563 ();
 sg13g2_fill_1 FILLER_59_2568 ();
 sg13g2_fill_1 FILLER_59_2578 ();
 sg13g2_fill_1 FILLER_59_2595 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_39 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_decap_4 FILLER_60_121 ();
 sg13g2_fill_1 FILLER_60_125 ();
 sg13g2_fill_2 FILLER_60_130 ();
 sg13g2_fill_1 FILLER_60_132 ();
 sg13g2_decap_4 FILLER_60_137 ();
 sg13g2_fill_1 FILLER_60_171 ();
 sg13g2_fill_1 FILLER_60_198 ();
 sg13g2_fill_2 FILLER_60_207 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_decap_4 FILLER_60_254 ();
 sg13g2_fill_2 FILLER_60_258 ();
 sg13g2_decap_4 FILLER_60_264 ();
 sg13g2_fill_1 FILLER_60_268 ();
 sg13g2_fill_1 FILLER_60_273 ();
 sg13g2_fill_2 FILLER_60_305 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_fill_2 FILLER_60_354 ();
 sg13g2_decap_8 FILLER_60_370 ();
 sg13g2_decap_4 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_401 ();
 sg13g2_decap_8 FILLER_60_411 ();
 sg13g2_decap_8 FILLER_60_418 ();
 sg13g2_decap_4 FILLER_60_425 ();
 sg13g2_fill_1 FILLER_60_460 ();
 sg13g2_decap_8 FILLER_60_465 ();
 sg13g2_fill_1 FILLER_60_472 ();
 sg13g2_fill_1 FILLER_60_523 ();
 sg13g2_fill_2 FILLER_60_550 ();
 sg13g2_fill_1 FILLER_60_561 ();
 sg13g2_fill_1 FILLER_60_605 ();
 sg13g2_fill_2 FILLER_60_610 ();
 sg13g2_fill_2 FILLER_60_616 ();
 sg13g2_fill_1 FILLER_60_628 ();
 sg13g2_fill_1 FILLER_60_640 ();
 sg13g2_fill_1 FILLER_60_649 ();
 sg13g2_fill_2 FILLER_60_655 ();
 sg13g2_fill_1 FILLER_60_657 ();
 sg13g2_fill_1 FILLER_60_667 ();
 sg13g2_fill_2 FILLER_60_682 ();
 sg13g2_fill_1 FILLER_60_684 ();
 sg13g2_fill_1 FILLER_60_724 ();
 sg13g2_decap_4 FILLER_60_769 ();
 sg13g2_fill_1 FILLER_60_783 ();
 sg13g2_decap_8 FILLER_60_826 ();
 sg13g2_fill_1 FILLER_60_833 ();
 sg13g2_fill_2 FILLER_60_878 ();
 sg13g2_fill_1 FILLER_60_897 ();
 sg13g2_fill_2 FILLER_60_966 ();
 sg13g2_fill_1 FILLER_60_978 ();
 sg13g2_fill_2 FILLER_60_990 ();
 sg13g2_fill_2 FILLER_60_1011 ();
 sg13g2_fill_1 FILLER_60_1027 ();
 sg13g2_fill_1 FILLER_60_1060 ();
 sg13g2_decap_8 FILLER_60_1071 ();
 sg13g2_decap_8 FILLER_60_1078 ();
 sg13g2_decap_8 FILLER_60_1085 ();
 sg13g2_fill_2 FILLER_60_1092 ();
 sg13g2_fill_1 FILLER_60_1094 ();
 sg13g2_fill_1 FILLER_60_1099 ();
 sg13g2_fill_2 FILLER_60_1110 ();
 sg13g2_fill_2 FILLER_60_1127 ();
 sg13g2_decap_8 FILLER_60_1159 ();
 sg13g2_decap_8 FILLER_60_1166 ();
 sg13g2_decap_8 FILLER_60_1173 ();
 sg13g2_decap_4 FILLER_60_1180 ();
 sg13g2_decap_4 FILLER_60_1188 ();
 sg13g2_fill_2 FILLER_60_1192 ();
 sg13g2_decap_4 FILLER_60_1198 ();
 sg13g2_fill_2 FILLER_60_1202 ();
 sg13g2_decap_8 FILLER_60_1234 ();
 sg13g2_decap_8 FILLER_60_1241 ();
 sg13g2_decap_8 FILLER_60_1248 ();
 sg13g2_fill_2 FILLER_60_1255 ();
 sg13g2_fill_2 FILLER_60_1261 ();
 sg13g2_fill_1 FILLER_60_1268 ();
 sg13g2_fill_2 FILLER_60_1273 ();
 sg13g2_fill_2 FILLER_60_1291 ();
 sg13g2_fill_2 FILLER_60_1324 ();
 sg13g2_fill_1 FILLER_60_1343 ();
 sg13g2_decap_4 FILLER_60_1367 ();
 sg13g2_fill_2 FILLER_60_1371 ();
 sg13g2_fill_1 FILLER_60_1376 ();
 sg13g2_fill_1 FILLER_60_1381 ();
 sg13g2_decap_8 FILLER_60_1423 ();
 sg13g2_decap_4 FILLER_60_1430 ();
 sg13g2_fill_2 FILLER_60_1450 ();
 sg13g2_fill_1 FILLER_60_1456 ();
 sg13g2_fill_1 FILLER_60_1462 ();
 sg13g2_fill_1 FILLER_60_1473 ();
 sg13g2_decap_4 FILLER_60_1479 ();
 sg13g2_decap_8 FILLER_60_1487 ();
 sg13g2_decap_4 FILLER_60_1494 ();
 sg13g2_fill_2 FILLER_60_1502 ();
 sg13g2_fill_1 FILLER_60_1504 ();
 sg13g2_fill_2 FILLER_60_1514 ();
 sg13g2_fill_1 FILLER_60_1516 ();
 sg13g2_fill_1 FILLER_60_1527 ();
 sg13g2_fill_1 FILLER_60_1535 ();
 sg13g2_decap_8 FILLER_60_1566 ();
 sg13g2_fill_2 FILLER_60_1609 ();
 sg13g2_fill_1 FILLER_60_1627 ();
 sg13g2_fill_2 FILLER_60_1682 ();
 sg13g2_fill_2 FILLER_60_1695 ();
 sg13g2_fill_1 FILLER_60_1716 ();
 sg13g2_fill_2 FILLER_60_1738 ();
 sg13g2_decap_4 FILLER_60_1770 ();
 sg13g2_fill_2 FILLER_60_1774 ();
 sg13g2_decap_8 FILLER_60_1780 ();
 sg13g2_decap_8 FILLER_60_1791 ();
 sg13g2_decap_4 FILLER_60_1802 ();
 sg13g2_fill_1 FILLER_60_1806 ();
 sg13g2_decap_8 FILLER_60_1812 ();
 sg13g2_decap_4 FILLER_60_1855 ();
 sg13g2_fill_1 FILLER_60_1864 ();
 sg13g2_fill_1 FILLER_60_1875 ();
 sg13g2_decap_8 FILLER_60_1883 ();
 sg13g2_decap_8 FILLER_60_1890 ();
 sg13g2_decap_8 FILLER_60_1897 ();
 sg13g2_decap_8 FILLER_60_1904 ();
 sg13g2_decap_8 FILLER_60_1911 ();
 sg13g2_decap_8 FILLER_60_1918 ();
 sg13g2_decap_8 FILLER_60_1925 ();
 sg13g2_decap_4 FILLER_60_1932 ();
 sg13g2_fill_1 FILLER_60_1936 ();
 sg13g2_fill_1 FILLER_60_1941 ();
 sg13g2_decap_4 FILLER_60_1951 ();
 sg13g2_fill_1 FILLER_60_1955 ();
 sg13g2_decap_8 FILLER_60_1964 ();
 sg13g2_decap_8 FILLER_60_1971 ();
 sg13g2_decap_4 FILLER_60_1978 ();
 sg13g2_fill_2 FILLER_60_1982 ();
 sg13g2_decap_8 FILLER_60_2056 ();
 sg13g2_decap_8 FILLER_60_2063 ();
 sg13g2_fill_2 FILLER_60_2070 ();
 sg13g2_decap_8 FILLER_60_2082 ();
 sg13g2_fill_2 FILLER_60_2125 ();
 sg13g2_fill_1 FILLER_60_2127 ();
 sg13g2_decap_8 FILLER_60_2132 ();
 sg13g2_decap_8 FILLER_60_2139 ();
 sg13g2_decap_8 FILLER_60_2146 ();
 sg13g2_fill_1 FILLER_60_2153 ();
 sg13g2_fill_2 FILLER_60_2164 ();
 sg13g2_fill_1 FILLER_60_2166 ();
 sg13g2_decap_8 FILLER_60_2193 ();
 sg13g2_decap_8 FILLER_60_2200 ();
 sg13g2_decap_8 FILLER_60_2211 ();
 sg13g2_decap_8 FILLER_60_2218 ();
 sg13g2_fill_2 FILLER_60_2225 ();
 sg13g2_fill_1 FILLER_60_2279 ();
 sg13g2_decap_8 FILLER_60_2310 ();
 sg13g2_fill_2 FILLER_60_2348 ();
 sg13g2_fill_1 FILLER_60_2350 ();
 sg13g2_fill_1 FILLER_60_2370 ();
 sg13g2_fill_2 FILLER_60_2397 ();
 sg13g2_fill_1 FILLER_60_2431 ();
 sg13g2_fill_1 FILLER_60_2448 ();
 sg13g2_fill_1 FILLER_60_2471 ();
 sg13g2_decap_8 FILLER_60_2478 ();
 sg13g2_fill_2 FILLER_60_2485 ();
 sg13g2_decap_8 FILLER_60_2491 ();
 sg13g2_decap_4 FILLER_60_2498 ();
 sg13g2_fill_1 FILLER_60_2507 ();
 sg13g2_fill_2 FILLER_60_2528 ();
 sg13g2_fill_1 FILLER_60_2530 ();
 sg13g2_fill_2 FILLER_60_2536 ();
 sg13g2_decap_8 FILLER_60_2543 ();
 sg13g2_decap_4 FILLER_60_2550 ();
 sg13g2_fill_1 FILLER_60_2554 ();
 sg13g2_fill_1 FILLER_60_2565 ();
 sg13g2_fill_1 FILLER_60_2586 ();
 sg13g2_fill_1 FILLER_60_2595 ();
 sg13g2_fill_2 FILLER_60_2601 ();
 sg13g2_decap_8 FILLER_60_2663 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_decap_4 FILLER_61_29 ();
 sg13g2_fill_1 FILLER_61_33 ();
 sg13g2_fill_2 FILLER_61_39 ();
 sg13g2_fill_1 FILLER_61_41 ();
 sg13g2_decap_8 FILLER_61_46 ();
 sg13g2_decap_8 FILLER_61_61 ();
 sg13g2_fill_1 FILLER_61_108 ();
 sg13g2_decap_8 FILLER_61_135 ();
 sg13g2_decap_8 FILLER_61_142 ();
 sg13g2_fill_1 FILLER_61_153 ();
 sg13g2_decap_4 FILLER_61_158 ();
 sg13g2_fill_1 FILLER_61_162 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_175 ();
 sg13g2_fill_1 FILLER_61_177 ();
 sg13g2_decap_8 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_207 ();
 sg13g2_fill_1 FILLER_61_209 ();
 sg13g2_decap_8 FILLER_61_233 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_2 FILLER_61_252 ();
 sg13g2_fill_1 FILLER_61_258 ();
 sg13g2_fill_2 FILLER_61_299 ();
 sg13g2_fill_1 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_307 ();
 sg13g2_fill_2 FILLER_61_314 ();
 sg13g2_decap_4 FILLER_61_320 ();
 sg13g2_fill_1 FILLER_61_369 ();
 sg13g2_fill_2 FILLER_61_374 ();
 sg13g2_fill_1 FILLER_61_376 ();
 sg13g2_decap_8 FILLER_61_389 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_fill_2 FILLER_61_403 ();
 sg13g2_fill_1 FILLER_61_412 ();
 sg13g2_decap_8 FILLER_61_419 ();
 sg13g2_decap_8 FILLER_61_426 ();
 sg13g2_decap_4 FILLER_61_433 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_fill_2 FILLER_61_448 ();
 sg13g2_decap_8 FILLER_61_455 ();
 sg13g2_fill_1 FILLER_61_462 ();
 sg13g2_decap_8 FILLER_61_473 ();
 sg13g2_fill_2 FILLER_61_480 ();
 sg13g2_fill_2 FILLER_61_525 ();
 sg13g2_fill_1 FILLER_61_527 ();
 sg13g2_decap_4 FILLER_61_560 ();
 sg13g2_fill_1 FILLER_61_564 ();
 sg13g2_decap_4 FILLER_61_582 ();
 sg13g2_fill_1 FILLER_61_586 ();
 sg13g2_decap_8 FILLER_61_638 ();
 sg13g2_decap_8 FILLER_61_645 ();
 sg13g2_decap_8 FILLER_61_656 ();
 sg13g2_decap_4 FILLER_61_663 ();
 sg13g2_fill_1 FILLER_61_672 ();
 sg13g2_fill_2 FILLER_61_677 ();
 sg13g2_fill_1 FILLER_61_679 ();
 sg13g2_decap_4 FILLER_61_685 ();
 sg13g2_fill_1 FILLER_61_689 ();
 sg13g2_fill_1 FILLER_61_698 ();
 sg13g2_fill_2 FILLER_61_704 ();
 sg13g2_fill_2 FILLER_61_720 ();
 sg13g2_fill_2 FILLER_61_730 ();
 sg13g2_fill_2 FILLER_61_742 ();
 sg13g2_decap_4 FILLER_61_770 ();
 sg13g2_fill_2 FILLER_61_787 ();
 sg13g2_fill_1 FILLER_61_789 ();
 sg13g2_decap_8 FILLER_61_800 ();
 sg13g2_decap_8 FILLER_61_807 ();
 sg13g2_decap_8 FILLER_61_814 ();
 sg13g2_decap_8 FILLER_61_821 ();
 sg13g2_decap_4 FILLER_61_828 ();
 sg13g2_fill_1 FILLER_61_850 ();
 sg13g2_fill_1 FILLER_61_897 ();
 sg13g2_fill_2 FILLER_61_916 ();
 sg13g2_fill_1 FILLER_61_952 ();
 sg13g2_fill_2 FILLER_61_1005 ();
 sg13g2_fill_1 FILLER_61_1034 ();
 sg13g2_fill_2 FILLER_61_1081 ();
 sg13g2_decap_8 FILLER_61_1087 ();
 sg13g2_decap_8 FILLER_61_1094 ();
 sg13g2_decap_8 FILLER_61_1101 ();
 sg13g2_fill_2 FILLER_61_1108 ();
 sg13g2_fill_1 FILLER_61_1110 ();
 sg13g2_fill_2 FILLER_61_1132 ();
 sg13g2_fill_1 FILLER_61_1134 ();
 sg13g2_decap_8 FILLER_61_1139 ();
 sg13g2_decap_8 FILLER_61_1146 ();
 sg13g2_decap_4 FILLER_61_1153 ();
 sg13g2_fill_1 FILLER_61_1157 ();
 sg13g2_decap_4 FILLER_61_1162 ();
 sg13g2_fill_1 FILLER_61_1166 ();
 sg13g2_fill_1 FILLER_61_1176 ();
 sg13g2_fill_2 FILLER_61_1186 ();
 sg13g2_decap_4 FILLER_61_1192 ();
 sg13g2_fill_1 FILLER_61_1196 ();
 sg13g2_decap_8 FILLER_61_1232 ();
 sg13g2_decap_8 FILLER_61_1239 ();
 sg13g2_decap_4 FILLER_61_1252 ();
 sg13g2_fill_2 FILLER_61_1256 ();
 sg13g2_fill_2 FILLER_61_1262 ();
 sg13g2_fill_2 FILLER_61_1295 ();
 sg13g2_decap_8 FILLER_61_1324 ();
 sg13g2_decap_8 FILLER_61_1331 ();
 sg13g2_fill_1 FILLER_61_1338 ();
 sg13g2_fill_1 FILLER_61_1352 ();
 sg13g2_fill_2 FILLER_61_1358 ();
 sg13g2_fill_1 FILLER_61_1368 ();
 sg13g2_fill_1 FILLER_61_1379 ();
 sg13g2_fill_1 FILLER_61_1385 ();
 sg13g2_fill_1 FILLER_61_1417 ();
 sg13g2_fill_1 FILLER_61_1448 ();
 sg13g2_fill_2 FILLER_61_1453 ();
 sg13g2_fill_1 FILLER_61_1455 ();
 sg13g2_decap_4 FILLER_61_1460 ();
 sg13g2_fill_1 FILLER_61_1464 ();
 sg13g2_fill_1 FILLER_61_1469 ();
 sg13g2_decap_8 FILLER_61_1490 ();
 sg13g2_decap_8 FILLER_61_1497 ();
 sg13g2_decap_8 FILLER_61_1504 ();
 sg13g2_fill_1 FILLER_61_1511 ();
 sg13g2_fill_1 FILLER_61_1516 ();
 sg13g2_decap_8 FILLER_61_1521 ();
 sg13g2_fill_1 FILLER_61_1528 ();
 sg13g2_fill_1 FILLER_61_1537 ();
 sg13g2_fill_1 FILLER_61_1542 ();
 sg13g2_fill_1 FILLER_61_1547 ();
 sg13g2_decap_8 FILLER_61_1556 ();
 sg13g2_fill_2 FILLER_61_1563 ();
 sg13g2_fill_1 FILLER_61_1565 ();
 sg13g2_fill_2 FILLER_61_1578 ();
 sg13g2_fill_2 FILLER_61_1634 ();
 sg13g2_fill_1 FILLER_61_1679 ();
 sg13g2_fill_1 FILLER_61_1693 ();
 sg13g2_fill_1 FILLER_61_1726 ();
 sg13g2_fill_2 FILLER_61_1741 ();
 sg13g2_decap_8 FILLER_61_1758 ();
 sg13g2_decap_8 FILLER_61_1765 ();
 sg13g2_decap_4 FILLER_61_1772 ();
 sg13g2_fill_2 FILLER_61_1776 ();
 sg13g2_fill_2 FILLER_61_1782 ();
 sg13g2_fill_2 FILLER_61_1833 ();
 sg13g2_fill_1 FILLER_61_1835 ();
 sg13g2_fill_1 FILLER_61_1844 ();
 sg13g2_fill_2 FILLER_61_1858 ();
 sg13g2_fill_2 FILLER_61_1874 ();
 sg13g2_fill_1 FILLER_61_1876 ();
 sg13g2_fill_2 FILLER_61_1886 ();
 sg13g2_fill_1 FILLER_61_1888 ();
 sg13g2_decap_4 FILLER_61_1898 ();
 sg13g2_fill_2 FILLER_61_1902 ();
 sg13g2_decap_4 FILLER_61_1908 ();
 sg13g2_fill_1 FILLER_61_1912 ();
 sg13g2_decap_8 FILLER_61_1921 ();
 sg13g2_decap_8 FILLER_61_1928 ();
 sg13g2_decap_8 FILLER_61_1935 ();
 sg13g2_decap_8 FILLER_61_1942 ();
 sg13g2_decap_8 FILLER_61_1949 ();
 sg13g2_decap_8 FILLER_61_1956 ();
 sg13g2_fill_2 FILLER_61_1963 ();
 sg13g2_fill_2 FILLER_61_2062 ();
 sg13g2_decap_8 FILLER_61_2068 ();
 sg13g2_decap_4 FILLER_61_2075 ();
 sg13g2_fill_2 FILLER_61_2079 ();
 sg13g2_fill_1 FILLER_61_2117 ();
 sg13g2_fill_1 FILLER_61_2144 ();
 sg13g2_fill_2 FILLER_61_2228 ();
 sg13g2_fill_1 FILLER_61_2238 ();
 sg13g2_fill_2 FILLER_61_2249 ();
 sg13g2_fill_1 FILLER_61_2292 ();
 sg13g2_fill_1 FILLER_61_2319 ();
 sg13g2_fill_1 FILLER_61_2324 ();
 sg13g2_fill_2 FILLER_61_2329 ();
 sg13g2_fill_2 FILLER_61_2336 ();
 sg13g2_fill_1 FILLER_61_2342 ();
 sg13g2_decap_4 FILLER_61_2357 ();
 sg13g2_fill_1 FILLER_61_2361 ();
 sg13g2_decap_8 FILLER_61_2366 ();
 sg13g2_fill_1 FILLER_61_2373 ();
 sg13g2_fill_1 FILLER_61_2413 ();
 sg13g2_fill_2 FILLER_61_2448 ();
 sg13g2_fill_1 FILLER_61_2450 ();
 sg13g2_fill_2 FILLER_61_2460 ();
 sg13g2_fill_1 FILLER_61_2462 ();
 sg13g2_fill_2 FILLER_61_2468 ();
 sg13g2_decap_8 FILLER_61_2479 ();
 sg13g2_fill_2 FILLER_61_2486 ();
 sg13g2_fill_1 FILLER_61_2488 ();
 sg13g2_fill_1 FILLER_61_2497 ();
 sg13g2_fill_2 FILLER_61_2510 ();
 sg13g2_fill_2 FILLER_61_2555 ();
 sg13g2_fill_1 FILLER_61_2586 ();
 sg13g2_fill_2 FILLER_61_2597 ();
 sg13g2_decap_4 FILLER_61_2658 ();
 sg13g2_fill_2 FILLER_61_2668 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_7 ();
 sg13g2_decap_4 FILLER_62_12 ();
 sg13g2_fill_1 FILLER_62_16 ();
 sg13g2_fill_2 FILLER_62_21 ();
 sg13g2_fill_1 FILLER_62_23 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_46 ();
 sg13g2_decap_4 FILLER_62_53 ();
 sg13g2_fill_1 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_68 ();
 sg13g2_fill_2 FILLER_62_79 ();
 sg13g2_decap_8 FILLER_62_89 ();
 sg13g2_fill_1 FILLER_62_96 ();
 sg13g2_decap_8 FILLER_62_102 ();
 sg13g2_decap_4 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_113 ();
 sg13g2_decap_4 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_fill_1 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_222 ();
 sg13g2_fill_1 FILLER_62_229 ();
 sg13g2_fill_1 FILLER_62_256 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_fill_1 FILLER_62_293 ();
 sg13g2_decap_8 FILLER_62_299 ();
 sg13g2_fill_2 FILLER_62_306 ();
 sg13g2_decap_8 FILLER_62_320 ();
 sg13g2_decap_4 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_340 ();
 sg13g2_fill_1 FILLER_62_345 ();
 sg13g2_fill_2 FILLER_62_377 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_fill_2 FILLER_62_394 ();
 sg13g2_decap_4 FILLER_62_437 ();
 sg13g2_fill_1 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_446 ();
 sg13g2_fill_2 FILLER_62_453 ();
 sg13g2_fill_1 FILLER_62_459 ();
 sg13g2_decap_8 FILLER_62_491 ();
 sg13g2_fill_1 FILLER_62_503 ();
 sg13g2_fill_1 FILLER_62_508 ();
 sg13g2_fill_1 FILLER_62_513 ();
 sg13g2_fill_2 FILLER_62_519 ();
 sg13g2_fill_2 FILLER_62_530 ();
 sg13g2_fill_2 FILLER_62_540 ();
 sg13g2_decap_8 FILLER_62_547 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_fill_1 FILLER_62_556 ();
 sg13g2_decap_8 FILLER_62_566 ();
 sg13g2_fill_2 FILLER_62_573 ();
 sg13g2_fill_1 FILLER_62_575 ();
 sg13g2_decap_8 FILLER_62_580 ();
 sg13g2_decap_4 FILLER_62_587 ();
 sg13g2_fill_1 FILLER_62_601 ();
 sg13g2_decap_4 FILLER_62_637 ();
 sg13g2_decap_4 FILLER_62_676 ();
 sg13g2_fill_1 FILLER_62_680 ();
 sg13g2_fill_1 FILLER_62_686 ();
 sg13g2_fill_1 FILLER_62_693 ();
 sg13g2_fill_2 FILLER_62_711 ();
 sg13g2_fill_1 FILLER_62_752 ();
 sg13g2_fill_1 FILLER_62_840 ();
 sg13g2_fill_2 FILLER_62_849 ();
 sg13g2_fill_2 FILLER_62_961 ();
 sg13g2_fill_2 FILLER_62_1001 ();
 sg13g2_fill_2 FILLER_62_1033 ();
 sg13g2_fill_2 FILLER_62_1095 ();
 sg13g2_fill_1 FILLER_62_1105 ();
 sg13g2_decap_8 FILLER_62_1132 ();
 sg13g2_decap_8 FILLER_62_1139 ();
 sg13g2_fill_2 FILLER_62_1177 ();
 sg13g2_fill_1 FILLER_62_1179 ();
 sg13g2_fill_1 FILLER_62_1253 ();
 sg13g2_fill_1 FILLER_62_1280 ();
 sg13g2_fill_1 FILLER_62_1288 ();
 sg13g2_fill_1 FILLER_62_1299 ();
 sg13g2_fill_2 FILLER_62_1312 ();
 sg13g2_fill_1 FILLER_62_1314 ();
 sg13g2_fill_2 FILLER_62_1323 ();
 sg13g2_fill_1 FILLER_62_1325 ();
 sg13g2_fill_1 FILLER_62_1330 ();
 sg13g2_decap_8 FILLER_62_1336 ();
 sg13g2_decap_8 FILLER_62_1343 ();
 sg13g2_fill_2 FILLER_62_1350 ();
 sg13g2_fill_1 FILLER_62_1352 ();
 sg13g2_decap_8 FILLER_62_1366 ();
 sg13g2_decap_8 FILLER_62_1373 ();
 sg13g2_fill_2 FILLER_62_1398 ();
 sg13g2_fill_1 FILLER_62_1400 ();
 sg13g2_fill_1 FILLER_62_1416 ();
 sg13g2_fill_2 FILLER_62_1452 ();
 sg13g2_decap_4 FILLER_62_1459 ();
 sg13g2_fill_2 FILLER_62_1472 ();
 sg13g2_decap_8 FILLER_62_1491 ();
 sg13g2_decap_4 FILLER_62_1498 ();
 sg13g2_fill_1 FILLER_62_1502 ();
 sg13g2_fill_2 FILLER_62_1566 ();
 sg13g2_fill_1 FILLER_62_1568 ();
 sg13g2_decap_4 FILLER_62_1611 ();
 sg13g2_fill_1 FILLER_62_1615 ();
 sg13g2_fill_2 FILLER_62_1625 ();
 sg13g2_fill_2 FILLER_62_1638 ();
 sg13g2_fill_2 FILLER_62_1689 ();
 sg13g2_decap_8 FILLER_62_1751 ();
 sg13g2_fill_1 FILLER_62_1758 ();
 sg13g2_decap_4 FILLER_62_1763 ();
 sg13g2_fill_1 FILLER_62_1772 ();
 sg13g2_fill_2 FILLER_62_1783 ();
 sg13g2_fill_1 FILLER_62_1818 ();
 sg13g2_fill_2 FILLER_62_1834 ();
 sg13g2_decap_4 FILLER_62_1856 ();
 sg13g2_decap_4 FILLER_62_1870 ();
 sg13g2_fill_1 FILLER_62_1874 ();
 sg13g2_fill_1 FILLER_62_1884 ();
 sg13g2_fill_2 FILLER_62_1902 ();
 sg13g2_decap_4 FILLER_62_1909 ();
 sg13g2_fill_1 FILLER_62_1913 ();
 sg13g2_fill_1 FILLER_62_1938 ();
 sg13g2_decap_4 FILLER_62_1949 ();
 sg13g2_fill_2 FILLER_62_1953 ();
 sg13g2_decap_8 FILLER_62_1959 ();
 sg13g2_decap_8 FILLER_62_1966 ();
 sg13g2_fill_2 FILLER_62_2032 ();
 sg13g2_fill_2 FILLER_62_2092 ();
 sg13g2_fill_1 FILLER_62_2269 ();
 sg13g2_decap_8 FILLER_62_2280 ();
 sg13g2_decap_8 FILLER_62_2287 ();
 sg13g2_decap_8 FILLER_62_2294 ();
 sg13g2_fill_1 FILLER_62_2301 ();
 sg13g2_fill_2 FILLER_62_2306 ();
 sg13g2_fill_1 FILLER_62_2308 ();
 sg13g2_fill_1 FILLER_62_2331 ();
 sg13g2_fill_2 FILLER_62_2341 ();
 sg13g2_fill_1 FILLER_62_2383 ();
 sg13g2_fill_1 FILLER_62_2390 ();
 sg13g2_fill_1 FILLER_62_2401 ();
 sg13g2_fill_1 FILLER_62_2415 ();
 sg13g2_decap_4 FILLER_62_2425 ();
 sg13g2_fill_2 FILLER_62_2433 ();
 sg13g2_fill_1 FILLER_62_2435 ();
 sg13g2_fill_2 FILLER_62_2441 ();
 sg13g2_fill_2 FILLER_62_2448 ();
 sg13g2_fill_1 FILLER_62_2450 ();
 sg13g2_fill_2 FILLER_62_2455 ();
 sg13g2_fill_1 FILLER_62_2457 ();
 sg13g2_fill_2 FILLER_62_2469 ();
 sg13g2_fill_1 FILLER_62_2471 ();
 sg13g2_fill_1 FILLER_62_2519 ();
 sg13g2_fill_2 FILLER_62_2537 ();
 sg13g2_decap_8 FILLER_62_2544 ();
 sg13g2_fill_2 FILLER_62_2551 ();
 sg13g2_fill_1 FILLER_62_2553 ();
 sg13g2_fill_1 FILLER_62_2570 ();
 sg13g2_fill_1 FILLER_62_2586 ();
 sg13g2_fill_1 FILLER_62_2596 ();
 sg13g2_fill_1 FILLER_62_2611 ();
 sg13g2_fill_2 FILLER_62_2668 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_61 ();
 sg13g2_fill_2 FILLER_63_68 ();
 sg13g2_fill_2 FILLER_63_83 ();
 sg13g2_fill_1 FILLER_63_85 ();
 sg13g2_fill_1 FILLER_63_95 ();
 sg13g2_decap_4 FILLER_63_101 ();
 sg13g2_fill_2 FILLER_63_105 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_fill_1 FILLER_63_164 ();
 sg13g2_fill_2 FILLER_63_191 ();
 sg13g2_decap_8 FILLER_63_227 ();
 sg13g2_decap_8 FILLER_63_234 ();
 sg13g2_decap_8 FILLER_63_241 ();
 sg13g2_fill_1 FILLER_63_251 ();
 sg13g2_decap_4 FILLER_63_272 ();
 sg13g2_fill_2 FILLER_63_281 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_1 FILLER_63_289 ();
 sg13g2_fill_1 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_decap_8 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_337 ();
 sg13g2_decap_8 FILLER_63_344 ();
 sg13g2_decap_4 FILLER_63_351 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_decap_4 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_376 ();
 sg13g2_decap_4 FILLER_63_418 ();
 sg13g2_fill_1 FILLER_63_422 ();
 sg13g2_fill_2 FILLER_63_455 ();
 sg13g2_fill_1 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_decap_8 FILLER_63_483 ();
 sg13g2_fill_2 FILLER_63_490 ();
 sg13g2_fill_1 FILLER_63_492 ();
 sg13g2_fill_1 FILLER_63_499 ();
 sg13g2_fill_2 FILLER_63_509 ();
 sg13g2_decap_4 FILLER_63_515 ();
 sg13g2_fill_1 FILLER_63_519 ();
 sg13g2_decap_8 FILLER_63_546 ();
 sg13g2_decap_4 FILLER_63_553 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_fill_2 FILLER_63_588 ();
 sg13g2_fill_2 FILLER_63_616 ();
 sg13g2_fill_2 FILLER_63_622 ();
 sg13g2_decap_4 FILLER_63_650 ();
 sg13g2_decap_8 FILLER_63_666 ();
 sg13g2_decap_8 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_680 ();
 sg13g2_fill_1 FILLER_63_682 ();
 sg13g2_fill_2 FILLER_63_689 ();
 sg13g2_fill_1 FILLER_63_704 ();
 sg13g2_fill_2 FILLER_63_753 ();
 sg13g2_fill_2 FILLER_63_759 ();
 sg13g2_fill_1 FILLER_63_761 ();
 sg13g2_fill_2 FILLER_63_844 ();
 sg13g2_fill_1 FILLER_63_853 ();
 sg13g2_fill_1 FILLER_63_910 ();
 sg13g2_fill_1 FILLER_63_953 ();
 sg13g2_fill_2 FILLER_63_975 ();
 sg13g2_fill_1 FILLER_63_987 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_fill_2 FILLER_63_1039 ();
 sg13g2_decap_8 FILLER_63_1054 ();
 sg13g2_fill_2 FILLER_63_1061 ();
 sg13g2_fill_2 FILLER_63_1068 ();
 sg13g2_decap_8 FILLER_63_1080 ();
 sg13g2_decap_4 FILLER_63_1087 ();
 sg13g2_fill_1 FILLER_63_1096 ();
 sg13g2_fill_1 FILLER_63_1115 ();
 sg13g2_decap_4 FILLER_63_1146 ();
 sg13g2_fill_1 FILLER_63_1181 ();
 sg13g2_fill_2 FILLER_63_1190 ();
 sg13g2_fill_1 FILLER_63_1192 ();
 sg13g2_decap_8 FILLER_63_1232 ();
 sg13g2_decap_8 FILLER_63_1239 ();
 sg13g2_fill_1 FILLER_63_1267 ();
 sg13g2_fill_2 FILLER_63_1273 ();
 sg13g2_fill_2 FILLER_63_1322 ();
 sg13g2_fill_1 FILLER_63_1324 ();
 sg13g2_decap_8 FILLER_63_1328 ();
 sg13g2_fill_2 FILLER_63_1335 ();
 sg13g2_fill_2 FILLER_63_1346 ();
 sg13g2_fill_1 FILLER_63_1348 ();
 sg13g2_fill_2 FILLER_63_1372 ();
 sg13g2_fill_1 FILLER_63_1374 ();
 sg13g2_fill_1 FILLER_63_1396 ();
 sg13g2_fill_2 FILLER_63_1431 ();
 sg13g2_fill_2 FILLER_63_1463 ();
 sg13g2_fill_1 FILLER_63_1465 ();
 sg13g2_fill_2 FILLER_63_1476 ();
 sg13g2_fill_1 FILLER_63_1478 ();
 sg13g2_decap_4 FILLER_63_1483 ();
 sg13g2_fill_2 FILLER_63_1487 ();
 sg13g2_fill_1 FILLER_63_1494 ();
 sg13g2_fill_2 FILLER_63_1504 ();
 sg13g2_fill_2 FILLER_63_1511 ();
 sg13g2_fill_2 FILLER_63_1533 ();
 sg13g2_fill_1 FILLER_63_1535 ();
 sg13g2_decap_4 FILLER_63_1541 ();
 sg13g2_fill_1 FILLER_63_1545 ();
 sg13g2_decap_8 FILLER_63_1550 ();
 sg13g2_fill_1 FILLER_63_1557 ();
 sg13g2_decap_8 FILLER_63_1567 ();
 sg13g2_fill_2 FILLER_63_1574 ();
 sg13g2_fill_1 FILLER_63_1576 ();
 sg13g2_fill_1 FILLER_63_1581 ();
 sg13g2_fill_1 FILLER_63_1597 ();
 sg13g2_fill_1 FILLER_63_1601 ();
 sg13g2_fill_1 FILLER_63_1626 ();
 sg13g2_fill_1 FILLER_63_1643 ();
 sg13g2_fill_1 FILLER_63_1658 ();
 sg13g2_fill_1 FILLER_63_1666 ();
 sg13g2_decap_8 FILLER_63_1677 ();
 sg13g2_decap_4 FILLER_63_1684 ();
 sg13g2_fill_1 FILLER_63_1688 ();
 sg13g2_fill_1 FILLER_63_1693 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_fill_1 FILLER_63_1772 ();
 sg13g2_fill_2 FILLER_63_1781 ();
 sg13g2_fill_2 FILLER_63_1826 ();
 sg13g2_fill_1 FILLER_63_1828 ();
 sg13g2_decap_8 FILLER_63_1835 ();
 sg13g2_decap_8 FILLER_63_1847 ();
 sg13g2_fill_2 FILLER_63_1854 ();
 sg13g2_fill_2 FILLER_63_1905 ();
 sg13g2_fill_1 FILLER_63_1920 ();
 sg13g2_fill_2 FILLER_63_1926 ();
 sg13g2_fill_1 FILLER_63_1928 ();
 sg13g2_fill_2 FILLER_63_1952 ();
 sg13g2_fill_1 FILLER_63_1954 ();
 sg13g2_decap_8 FILLER_63_1963 ();
 sg13g2_decap_8 FILLER_63_1970 ();
 sg13g2_decap_8 FILLER_63_1977 ();
 sg13g2_fill_2 FILLER_63_1984 ();
 sg13g2_fill_2 FILLER_63_1995 ();
 sg13g2_fill_1 FILLER_63_1997 ();
 sg13g2_decap_4 FILLER_63_2008 ();
 sg13g2_decap_8 FILLER_63_2016 ();
 sg13g2_decap_8 FILLER_63_2076 ();
 sg13g2_decap_8 FILLER_63_2083 ();
 sg13g2_decap_8 FILLER_63_2090 ();
 sg13g2_fill_2 FILLER_63_2097 ();
 sg13g2_fill_1 FILLER_63_2099 ();
 sg13g2_decap_8 FILLER_63_2114 ();
 sg13g2_decap_4 FILLER_63_2121 ();
 sg13g2_fill_2 FILLER_63_2125 ();
 sg13g2_fill_2 FILLER_63_2131 ();
 sg13g2_fill_2 FILLER_63_2159 ();
 sg13g2_fill_1 FILLER_63_2161 ();
 sg13g2_fill_2 FILLER_63_2172 ();
 sg13g2_decap_8 FILLER_63_2233 ();
 sg13g2_fill_1 FILLER_63_2240 ();
 sg13g2_decap_4 FILLER_63_2247 ();
 sg13g2_fill_1 FILLER_63_2251 ();
 sg13g2_decap_8 FILLER_63_2278 ();
 sg13g2_decap_4 FILLER_63_2285 ();
 sg13g2_fill_1 FILLER_63_2289 ();
 sg13g2_fill_1 FILLER_63_2333 ();
 sg13g2_fill_2 FILLER_63_2356 ();
 sg13g2_fill_1 FILLER_63_2358 ();
 sg13g2_fill_2 FILLER_63_2373 ();
 sg13g2_fill_1 FILLER_63_2398 ();
 sg13g2_fill_2 FILLER_63_2436 ();
 sg13g2_fill_1 FILLER_63_2490 ();
 sg13g2_fill_1 FILLER_63_2566 ();
 sg13g2_fill_1 FILLER_63_2571 ();
 sg13g2_fill_1 FILLER_63_2616 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_4 FILLER_64_21 ();
 sg13g2_fill_1 FILLER_64_25 ();
 sg13g2_fill_1 FILLER_64_82 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_fill_1 FILLER_64_99 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_4 FILLER_64_119 ();
 sg13g2_fill_2 FILLER_64_123 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_4 FILLER_64_151 ();
 sg13g2_fill_2 FILLER_64_155 ();
 sg13g2_decap_8 FILLER_64_167 ();
 sg13g2_decap_4 FILLER_64_178 ();
 sg13g2_fill_2 FILLER_64_182 ();
 sg13g2_fill_1 FILLER_64_189 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_fill_1 FILLER_64_205 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_216 ();
 sg13g2_fill_1 FILLER_64_222 ();
 sg13g2_fill_1 FILLER_64_233 ();
 sg13g2_fill_1 FILLER_64_247 ();
 sg13g2_fill_2 FILLER_64_252 ();
 sg13g2_fill_2 FILLER_64_285 ();
 sg13g2_fill_2 FILLER_64_301 ();
 sg13g2_fill_1 FILLER_64_303 ();
 sg13g2_fill_2 FILLER_64_335 ();
 sg13g2_fill_1 FILLER_64_337 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_fill_2 FILLER_64_371 ();
 sg13g2_fill_1 FILLER_64_387 ();
 sg13g2_decap_8 FILLER_64_431 ();
 sg13g2_fill_2 FILLER_64_442 ();
 sg13g2_fill_1 FILLER_64_492 ();
 sg13g2_fill_2 FILLER_64_529 ();
 sg13g2_decap_8 FILLER_64_535 ();
 sg13g2_decap_4 FILLER_64_542 ();
 sg13g2_fill_2 FILLER_64_576 ();
 sg13g2_fill_1 FILLER_64_592 ();
 sg13g2_fill_2 FILLER_64_611 ();
 sg13g2_decap_8 FILLER_64_623 ();
 sg13g2_decap_8 FILLER_64_630 ();
 sg13g2_decap_8 FILLER_64_637 ();
 sg13g2_decap_4 FILLER_64_644 ();
 sg13g2_decap_4 FILLER_64_652 ();
 sg13g2_decap_8 FILLER_64_664 ();
 sg13g2_decap_8 FILLER_64_671 ();
 sg13g2_decap_4 FILLER_64_678 ();
 sg13g2_fill_2 FILLER_64_682 ();
 sg13g2_fill_2 FILLER_64_716 ();
 sg13g2_fill_1 FILLER_64_722 ();
 sg13g2_decap_8 FILLER_64_727 ();
 sg13g2_fill_2 FILLER_64_734 ();
 sg13g2_fill_1 FILLER_64_736 ();
 sg13g2_decap_4 FILLER_64_772 ();
 sg13g2_fill_1 FILLER_64_776 ();
 sg13g2_fill_2 FILLER_64_795 ();
 sg13g2_fill_1 FILLER_64_797 ();
 sg13g2_fill_1 FILLER_64_802 ();
 sg13g2_fill_1 FILLER_64_813 ();
 sg13g2_fill_1 FILLER_64_859 ();
 sg13g2_fill_2 FILLER_64_879 ();
 sg13g2_fill_2 FILLER_64_910 ();
 sg13g2_fill_1 FILLER_64_922 ();
 sg13g2_fill_2 FILLER_64_945 ();
 sg13g2_fill_1 FILLER_64_976 ();
 sg13g2_fill_2 FILLER_64_987 ();
 sg13g2_fill_1 FILLER_64_997 ();
 sg13g2_fill_2 FILLER_64_1013 ();
 sg13g2_fill_1 FILLER_64_1033 ();
 sg13g2_decap_8 FILLER_64_1060 ();
 sg13g2_decap_4 FILLER_64_1124 ();
 sg13g2_fill_1 FILLER_64_1189 ();
 sg13g2_fill_2 FILLER_64_1214 ();
 sg13g2_fill_1 FILLER_64_1216 ();
 sg13g2_decap_8 FILLER_64_1243 ();
 sg13g2_decap_8 FILLER_64_1250 ();
 sg13g2_fill_2 FILLER_64_1257 ();
 sg13g2_fill_1 FILLER_64_1259 ();
 sg13g2_fill_2 FILLER_64_1264 ();
 sg13g2_fill_1 FILLER_64_1276 ();
 sg13g2_fill_2 FILLER_64_1285 ();
 sg13g2_fill_1 FILLER_64_1292 ();
 sg13g2_fill_1 FILLER_64_1298 ();
 sg13g2_fill_2 FILLER_64_1304 ();
 sg13g2_fill_1 FILLER_64_1314 ();
 sg13g2_fill_2 FILLER_64_1320 ();
 sg13g2_fill_2 FILLER_64_1327 ();
 sg13g2_fill_1 FILLER_64_1329 ();
 sg13g2_fill_1 FILLER_64_1347 ();
 sg13g2_fill_2 FILLER_64_1397 ();
 sg13g2_fill_2 FILLER_64_1407 ();
 sg13g2_fill_2 FILLER_64_1414 ();
 sg13g2_fill_2 FILLER_64_1463 ();
 sg13g2_fill_1 FILLER_64_1465 ();
 sg13g2_decap_4 FILLER_64_1483 ();
 sg13g2_fill_1 FILLER_64_1487 ();
 sg13g2_fill_2 FILLER_64_1510 ();
 sg13g2_fill_2 FILLER_64_1526 ();
 sg13g2_decap_8 FILLER_64_1532 ();
 sg13g2_fill_1 FILLER_64_1539 ();
 sg13g2_fill_2 FILLER_64_1546 ();
 sg13g2_fill_1 FILLER_64_1548 ();
 sg13g2_decap_8 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1560 ();
 sg13g2_decap_8 FILLER_64_1567 ();
 sg13g2_fill_2 FILLER_64_1574 ();
 sg13g2_fill_1 FILLER_64_1576 ();
 sg13g2_fill_2 FILLER_64_1582 ();
 sg13g2_decap_8 FILLER_64_1588 ();
 sg13g2_fill_2 FILLER_64_1595 ();
 sg13g2_fill_1 FILLER_64_1597 ();
 sg13g2_fill_2 FILLER_64_1606 ();
 sg13g2_fill_1 FILLER_64_1608 ();
 sg13g2_fill_1 FILLER_64_1617 ();
 sg13g2_fill_2 FILLER_64_1650 ();
 sg13g2_decap_4 FILLER_64_1666 ();
 sg13g2_fill_1 FILLER_64_1695 ();
 sg13g2_fill_2 FILLER_64_1700 ();
 sg13g2_fill_2 FILLER_64_1716 ();
 sg13g2_decap_8 FILLER_64_1728 ();
 sg13g2_decap_8 FILLER_64_1735 ();
 sg13g2_fill_1 FILLER_64_1794 ();
 sg13g2_fill_2 FILLER_64_1799 ();
 sg13g2_fill_1 FILLER_64_1809 ();
 sg13g2_decap_8 FILLER_64_1832 ();
 sg13g2_decap_4 FILLER_64_1839 ();
 sg13g2_decap_4 FILLER_64_1854 ();
 sg13g2_fill_2 FILLER_64_1862 ();
 sg13g2_fill_1 FILLER_64_1874 ();
 sg13g2_fill_2 FILLER_64_1890 ();
 sg13g2_fill_1 FILLER_64_1927 ();
 sg13g2_fill_2 FILLER_64_1953 ();
 sg13g2_decap_8 FILLER_64_1963 ();
 sg13g2_decap_8 FILLER_64_1970 ();
 sg13g2_decap_4 FILLER_64_1977 ();
 sg13g2_fill_2 FILLER_64_1981 ();
 sg13g2_decap_4 FILLER_64_1993 ();
 sg13g2_fill_1 FILLER_64_1997 ();
 sg13g2_decap_8 FILLER_64_2026 ();
 sg13g2_decap_8 FILLER_64_2033 ();
 sg13g2_decap_8 FILLER_64_2040 ();
 sg13g2_decap_4 FILLER_64_2047 ();
 sg13g2_fill_1 FILLER_64_2051 ();
 sg13g2_fill_2 FILLER_64_2078 ();
 sg13g2_fill_1 FILLER_64_2080 ();
 sg13g2_decap_8 FILLER_64_2152 ();
 sg13g2_fill_2 FILLER_64_2159 ();
 sg13g2_fill_1 FILLER_64_2161 ();
 sg13g2_fill_2 FILLER_64_2239 ();
 sg13g2_fill_1 FILLER_64_2266 ();
 sg13g2_fill_2 FILLER_64_2322 ();
 sg13g2_fill_2 FILLER_64_2332 ();
 sg13g2_fill_1 FILLER_64_2374 ();
 sg13g2_fill_1 FILLER_64_2385 ();
 sg13g2_decap_4 FILLER_64_2442 ();
 sg13g2_fill_1 FILLER_64_2446 ();
 sg13g2_fill_1 FILLER_64_2455 ();
 sg13g2_fill_2 FILLER_64_2461 ();
 sg13g2_fill_1 FILLER_64_2467 ();
 sg13g2_fill_1 FILLER_64_2475 ();
 sg13g2_fill_2 FILLER_64_2519 ();
 sg13g2_fill_2 FILLER_64_2526 ();
 sg13g2_fill_2 FILLER_64_2532 ();
 sg13g2_decap_8 FILLER_64_2542 ();
 sg13g2_decap_4 FILLER_64_2549 ();
 sg13g2_fill_1 FILLER_64_2553 ();
 sg13g2_fill_2 FILLER_64_2558 ();
 sg13g2_decap_8 FILLER_64_2565 ();
 sg13g2_fill_1 FILLER_64_2572 ();
 sg13g2_fill_2 FILLER_64_2630 ();
 sg13g2_fill_2 FILLER_64_2642 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_33 ();
 sg13g2_fill_2 FILLER_65_38 ();
 sg13g2_fill_2 FILLER_65_45 ();
 sg13g2_decap_8 FILLER_65_51 ();
 sg13g2_fill_1 FILLER_65_58 ();
 sg13g2_fill_2 FILLER_65_64 ();
 sg13g2_fill_2 FILLER_65_70 ();
 sg13g2_fill_1 FILLER_65_72 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_1 FILLER_65_88 ();
 sg13g2_fill_1 FILLER_65_136 ();
 sg13g2_decap_4 FILLER_65_152 ();
 sg13g2_fill_2 FILLER_65_177 ();
 sg13g2_fill_1 FILLER_65_179 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_decap_8 FILLER_65_209 ();
 sg13g2_fill_2 FILLER_65_216 ();
 sg13g2_fill_1 FILLER_65_218 ();
 sg13g2_decap_8 FILLER_65_225 ();
 sg13g2_fill_2 FILLER_65_232 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_decap_4 FILLER_65_301 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_fill_1 FILLER_65_311 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_1 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_355 ();
 sg13g2_fill_2 FILLER_65_362 ();
 sg13g2_fill_2 FILLER_65_379 ();
 sg13g2_fill_1 FILLER_65_404 ();
 sg13g2_decap_8 FILLER_65_431 ();
 sg13g2_decap_4 FILLER_65_438 ();
 sg13g2_fill_1 FILLER_65_442 ();
 sg13g2_fill_1 FILLER_65_478 ();
 sg13g2_fill_2 FILLER_65_495 ();
 sg13g2_fill_1 FILLER_65_512 ();
 sg13g2_fill_1 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_531 ();
 sg13g2_decap_4 FILLER_65_538 ();
 sg13g2_fill_1 FILLER_65_542 ();
 sg13g2_fill_2 FILLER_65_552 ();
 sg13g2_fill_1 FILLER_65_575 ();
 sg13g2_decap_4 FILLER_65_584 ();
 sg13g2_fill_2 FILLER_65_588 ();
 sg13g2_decap_8 FILLER_65_594 ();
 sg13g2_decap_8 FILLER_65_601 ();
 sg13g2_decap_8 FILLER_65_608 ();
 sg13g2_decap_8 FILLER_65_615 ();
 sg13g2_decap_8 FILLER_65_622 ();
 sg13g2_fill_2 FILLER_65_629 ();
 sg13g2_fill_2 FILLER_65_664 ();
 sg13g2_fill_2 FILLER_65_676 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_fill_1 FILLER_65_684 ();
 sg13g2_fill_2 FILLER_65_711 ();
 sg13g2_fill_1 FILLER_65_713 ();
 sg13g2_decap_8 FILLER_65_718 ();
 sg13g2_decap_8 FILLER_65_725 ();
 sg13g2_decap_4 FILLER_65_732 ();
 sg13g2_decap_8 FILLER_65_767 ();
 sg13g2_decap_8 FILLER_65_774 ();
 sg13g2_decap_8 FILLER_65_781 ();
 sg13g2_fill_2 FILLER_65_788 ();
 sg13g2_decap_4 FILLER_65_795 ();
 sg13g2_fill_1 FILLER_65_799 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_4 FILLER_65_812 ();
 sg13g2_fill_2 FILLER_65_872 ();
 sg13g2_fill_1 FILLER_65_904 ();
 sg13g2_fill_2 FILLER_65_911 ();
 sg13g2_fill_1 FILLER_65_930 ();
 sg13g2_fill_1 FILLER_65_971 ();
 sg13g2_fill_1 FILLER_65_1017 ();
 sg13g2_decap_4 FILLER_65_1054 ();
 sg13g2_fill_2 FILLER_65_1078 ();
 sg13g2_fill_2 FILLER_65_1106 ();
 sg13g2_decap_8 FILLER_65_1120 ();
 sg13g2_decap_8 FILLER_65_1127 ();
 sg13g2_fill_1 FILLER_65_1173 ();
 sg13g2_decap_8 FILLER_65_1178 ();
 sg13g2_fill_1 FILLER_65_1185 ();
 sg13g2_decap_4 FILLER_65_1190 ();
 sg13g2_decap_8 FILLER_65_1225 ();
 sg13g2_decap_8 FILLER_65_1232 ();
 sg13g2_decap_4 FILLER_65_1239 ();
 sg13g2_fill_2 FILLER_65_1243 ();
 sg13g2_fill_2 FILLER_65_1255 ();
 sg13g2_decap_8 FILLER_65_1280 ();
 sg13g2_decap_4 FILLER_65_1287 ();
 sg13g2_fill_2 FILLER_65_1299 ();
 sg13g2_fill_1 FILLER_65_1305 ();
 sg13g2_fill_1 FILLER_65_1311 ();
 sg13g2_fill_1 FILLER_65_1319 ();
 sg13g2_fill_1 FILLER_65_1328 ();
 sg13g2_fill_1 FILLER_65_1337 ();
 sg13g2_fill_2 FILLER_65_1342 ();
 sg13g2_fill_1 FILLER_65_1369 ();
 sg13g2_fill_1 FILLER_65_1383 ();
 sg13g2_decap_4 FILLER_65_1417 ();
 sg13g2_fill_2 FILLER_65_1426 ();
 sg13g2_fill_2 FILLER_65_1447 ();
 sg13g2_fill_1 FILLER_65_1460 ();
 sg13g2_fill_2 FILLER_65_1470 ();
 sg13g2_fill_2 FILLER_65_1482 ();
 sg13g2_decap_8 FILLER_65_1489 ();
 sg13g2_decap_8 FILLER_65_1500 ();
 sg13g2_fill_1 FILLER_65_1507 ();
 sg13g2_decap_4 FILLER_65_1520 ();
 sg13g2_fill_2 FILLER_65_1524 ();
 sg13g2_fill_2 FILLER_65_1569 ();
 sg13g2_fill_1 FILLER_65_1575 ();
 sg13g2_decap_4 FILLER_65_1602 ();
 sg13g2_fill_2 FILLER_65_1606 ();
 sg13g2_fill_2 FILLER_65_1625 ();
 sg13g2_fill_1 FILLER_65_1627 ();
 sg13g2_fill_1 FILLER_65_1640 ();
 sg13g2_fill_1 FILLER_65_1653 ();
 sg13g2_fill_2 FILLER_65_1666 ();
 sg13g2_fill_2 FILLER_65_1682 ();
 sg13g2_fill_1 FILLER_65_1688 ();
 sg13g2_fill_2 FILLER_65_1710 ();
 sg13g2_fill_2 FILLER_65_1734 ();
 sg13g2_fill_1 FILLER_65_1736 ();
 sg13g2_decap_8 FILLER_65_1742 ();
 sg13g2_decap_4 FILLER_65_1749 ();
 sg13g2_fill_2 FILLER_65_1792 ();
 sg13g2_fill_2 FILLER_65_1798 ();
 sg13g2_decap_4 FILLER_65_1831 ();
 sg13g2_fill_2 FILLER_65_1835 ();
 sg13g2_decap_4 FILLER_65_1847 ();
 sg13g2_fill_2 FILLER_65_1851 ();
 sg13g2_fill_2 FILLER_65_1881 ();
 sg13g2_fill_1 FILLER_65_1924 ();
 sg13g2_fill_1 FILLER_65_1930 ();
 sg13g2_fill_1 FILLER_65_1940 ();
 sg13g2_decap_4 FILLER_65_1968 ();
 sg13g2_fill_2 FILLER_65_2006 ();
 sg13g2_decap_8 FILLER_65_2041 ();
 sg13g2_fill_2 FILLER_65_2048 ();
 sg13g2_decap_8 FILLER_65_2055 ();
 sg13g2_decap_8 FILLER_65_2062 ();
 sg13g2_fill_2 FILLER_65_2069 ();
 sg13g2_decap_8 FILLER_65_2081 ();
 sg13g2_decap_4 FILLER_65_2114 ();
 sg13g2_fill_1 FILLER_65_2118 ();
 sg13g2_decap_4 FILLER_65_2138 ();
 sg13g2_fill_2 FILLER_65_2163 ();
 sg13g2_decap_8 FILLER_65_2223 ();
 sg13g2_fill_1 FILLER_65_2230 ();
 sg13g2_fill_1 FILLER_65_2267 ();
 sg13g2_fill_1 FILLER_65_2289 ();
 sg13g2_fill_2 FILLER_65_2307 ();
 sg13g2_fill_1 FILLER_65_2309 ();
 sg13g2_fill_1 FILLER_65_2349 ();
 sg13g2_fill_2 FILLER_65_2475 ();
 sg13g2_fill_1 FILLER_65_2486 ();
 sg13g2_fill_2 FILLER_65_2495 ();
 sg13g2_fill_1 FILLER_65_2515 ();
 sg13g2_fill_2 FILLER_65_2520 ();
 sg13g2_fill_1 FILLER_65_2526 ();
 sg13g2_fill_1 FILLER_65_2579 ();
 sg13g2_fill_2 FILLER_65_2625 ();
 sg13g2_decap_4 FILLER_65_2666 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_12 ();
 sg13g2_decap_8 FILLER_66_18 ();
 sg13g2_decap_4 FILLER_66_25 ();
 sg13g2_fill_2 FILLER_66_29 ();
 sg13g2_fill_2 FILLER_66_41 ();
 sg13g2_fill_1 FILLER_66_43 ();
 sg13g2_fill_2 FILLER_66_54 ();
 sg13g2_fill_2 FILLER_66_86 ();
 sg13g2_fill_1 FILLER_66_88 ();
 sg13g2_fill_2 FILLER_66_97 ();
 sg13g2_fill_1 FILLER_66_104 ();
 sg13g2_decap_4 FILLER_66_115 ();
 sg13g2_decap_4 FILLER_66_145 ();
 sg13g2_fill_2 FILLER_66_149 ();
 sg13g2_fill_1 FILLER_66_177 ();
 sg13g2_fill_2 FILLER_66_188 ();
 sg13g2_fill_2 FILLER_66_230 ();
 sg13g2_fill_1 FILLER_66_232 ();
 sg13g2_fill_1 FILLER_66_247 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_2 FILLER_66_264 ();
 sg13g2_decap_4 FILLER_66_271 ();
 sg13g2_decap_8 FILLER_66_279 ();
 sg13g2_decap_4 FILLER_66_286 ();
 sg13g2_fill_2 FILLER_66_294 ();
 sg13g2_decap_4 FILLER_66_301 ();
 sg13g2_fill_1 FILLER_66_305 ();
 sg13g2_fill_2 FILLER_66_311 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_376 ();
 sg13g2_fill_2 FILLER_66_408 ();
 sg13g2_fill_2 FILLER_66_413 ();
 sg13g2_fill_2 FILLER_66_430 ();
 sg13g2_fill_1 FILLER_66_441 ();
 sg13g2_fill_1 FILLER_66_462 ();
 sg13g2_fill_1 FILLER_66_468 ();
 sg13g2_fill_1 FILLER_66_491 ();
 sg13g2_decap_8 FILLER_66_521 ();
 sg13g2_decap_8 FILLER_66_528 ();
 sg13g2_fill_1 FILLER_66_535 ();
 sg13g2_fill_2 FILLER_66_598 ();
 sg13g2_fill_1 FILLER_66_600 ();
 sg13g2_decap_8 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_630 ();
 sg13g2_fill_2 FILLER_66_637 ();
 sg13g2_fill_1 FILLER_66_639 ();
 sg13g2_fill_2 FILLER_66_644 ();
 sg13g2_fill_1 FILLER_66_651 ();
 sg13g2_fill_1 FILLER_66_667 ();
 sg13g2_fill_1 FILLER_66_674 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_decap_8 FILLER_66_710 ();
 sg13g2_decap_8 FILLER_66_717 ();
 sg13g2_decap_8 FILLER_66_724 ();
 sg13g2_fill_1 FILLER_66_741 ();
 sg13g2_fill_1 FILLER_66_774 ();
 sg13g2_fill_2 FILLER_66_780 ();
 sg13g2_fill_1 FILLER_66_782 ();
 sg13g2_decap_8 FILLER_66_809 ();
 sg13g2_decap_8 FILLER_66_816 ();
 sg13g2_decap_8 FILLER_66_823 ();
 sg13g2_decap_4 FILLER_66_834 ();
 sg13g2_fill_2 FILLER_66_864 ();
 sg13g2_fill_1 FILLER_66_895 ();
 sg13g2_fill_2 FILLER_66_913 ();
 sg13g2_fill_2 FILLER_66_928 ();
 sg13g2_decap_8 FILLER_66_985 ();
 sg13g2_decap_8 FILLER_66_992 ();
 sg13g2_decap_4 FILLER_66_999 ();
 sg13g2_fill_1 FILLER_66_1003 ();
 sg13g2_fill_1 FILLER_66_1035 ();
 sg13g2_fill_1 FILLER_66_1049 ();
 sg13g2_decap_8 FILLER_66_1058 ();
 sg13g2_decap_8 FILLER_66_1065 ();
 sg13g2_fill_2 FILLER_66_1072 ();
 sg13g2_fill_1 FILLER_66_1074 ();
 sg13g2_decap_8 FILLER_66_1079 ();
 sg13g2_fill_2 FILLER_66_1086 ();
 sg13g2_fill_1 FILLER_66_1088 ();
 sg13g2_decap_8 FILLER_66_1097 ();
 sg13g2_decap_8 FILLER_66_1104 ();
 sg13g2_fill_2 FILLER_66_1111 ();
 sg13g2_fill_2 FILLER_66_1118 ();
 sg13g2_decap_8 FILLER_66_1128 ();
 sg13g2_decap_4 FILLER_66_1140 ();
 sg13g2_fill_2 FILLER_66_1144 ();
 sg13g2_fill_1 FILLER_66_1154 ();
 sg13g2_decap_4 FILLER_66_1173 ();
 sg13g2_fill_2 FILLER_66_1203 ();
 sg13g2_fill_2 FILLER_66_1235 ();
 sg13g2_fill_1 FILLER_66_1237 ();
 sg13g2_decap_8 FILLER_66_1301 ();
 sg13g2_decap_4 FILLER_66_1308 ();
 sg13g2_fill_2 FILLER_66_1312 ();
 sg13g2_fill_2 FILLER_66_1324 ();
 sg13g2_fill_2 FILLER_66_1338 ();
 sg13g2_decap_4 FILLER_66_1357 ();
 sg13g2_fill_1 FILLER_66_1361 ();
 sg13g2_fill_2 FILLER_66_1372 ();
 sg13g2_decap_8 FILLER_66_1386 ();
 sg13g2_decap_4 FILLER_66_1393 ();
 sg13g2_fill_2 FILLER_66_1397 ();
 sg13g2_decap_8 FILLER_66_1409 ();
 sg13g2_decap_8 FILLER_66_1416 ();
 sg13g2_decap_8 FILLER_66_1423 ();
 sg13g2_fill_1 FILLER_66_1430 ();
 sg13g2_fill_2 FILLER_66_1434 ();
 sg13g2_fill_1 FILLER_66_1436 ();
 sg13g2_decap_4 FILLER_66_1441 ();
 sg13g2_decap_4 FILLER_66_1450 ();
 sg13g2_fill_2 FILLER_66_1470 ();
 sg13g2_fill_2 FILLER_66_1490 ();
 sg13g2_fill_2 FILLER_66_1497 ();
 sg13g2_fill_1 FILLER_66_1499 ();
 sg13g2_fill_2 FILLER_66_1504 ();
 sg13g2_fill_1 FILLER_66_1506 ();
 sg13g2_fill_2 FILLER_66_1512 ();
 sg13g2_decap_8 FILLER_66_1522 ();
 sg13g2_fill_2 FILLER_66_1529 ();
 sg13g2_fill_1 FILLER_66_1555 ();
 sg13g2_fill_2 FILLER_66_1561 ();
 sg13g2_fill_1 FILLER_66_1563 ();
 sg13g2_fill_1 FILLER_66_1569 ();
 sg13g2_fill_1 FILLER_66_1577 ();
 sg13g2_fill_2 FILLER_66_1586 ();
 sg13g2_fill_1 FILLER_66_1609 ();
 sg13g2_decap_8 FILLER_66_1618 ();
 sg13g2_fill_1 FILLER_66_1625 ();
 sg13g2_decap_8 FILLER_66_1660 ();
 sg13g2_decap_4 FILLER_66_1667 ();
 sg13g2_fill_2 FILLER_66_1700 ();
 sg13g2_fill_1 FILLER_66_1707 ();
 sg13g2_fill_1 FILLER_66_1721 ();
 sg13g2_decap_8 FILLER_66_1733 ();
 sg13g2_decap_8 FILLER_66_1745 ();
 sg13g2_decap_4 FILLER_66_1752 ();
 sg13g2_fill_1 FILLER_66_1765 ();
 sg13g2_fill_2 FILLER_66_1771 ();
 sg13g2_fill_1 FILLER_66_1800 ();
 sg13g2_fill_1 FILLER_66_1817 ();
 sg13g2_decap_8 FILLER_66_1836 ();
 sg13g2_decap_8 FILLER_66_1843 ();
 sg13g2_fill_1 FILLER_66_1850 ();
 sg13g2_fill_2 FILLER_66_1884 ();
 sg13g2_fill_1 FILLER_66_1886 ();
 sg13g2_fill_1 FILLER_66_1892 ();
 sg13g2_fill_1 FILLER_66_1906 ();
 sg13g2_fill_1 FILLER_66_1911 ();
 sg13g2_fill_2 FILLER_66_1917 ();
 sg13g2_fill_1 FILLER_66_1919 ();
 sg13g2_fill_2 FILLER_66_1947 ();
 sg13g2_fill_1 FILLER_66_1949 ();
 sg13g2_decap_8 FILLER_66_1966 ();
 sg13g2_decap_8 FILLER_66_1973 ();
 sg13g2_decap_4 FILLER_66_1980 ();
 sg13g2_fill_1 FILLER_66_1984 ();
 sg13g2_decap_8 FILLER_66_2046 ();
 sg13g2_decap_8 FILLER_66_2063 ();
 sg13g2_decap_8 FILLER_66_2148 ();
 sg13g2_decap_8 FILLER_66_2155 ();
 sg13g2_decap_4 FILLER_66_2162 ();
 sg13g2_fill_2 FILLER_66_2166 ();
 sg13g2_decap_8 FILLER_66_2234 ();
 sg13g2_decap_4 FILLER_66_2241 ();
 sg13g2_fill_1 FILLER_66_2245 ();
 sg13g2_decap_8 FILLER_66_2260 ();
 sg13g2_decap_8 FILLER_66_2267 ();
 sg13g2_fill_2 FILLER_66_2274 ();
 sg13g2_fill_1 FILLER_66_2280 ();
 sg13g2_decap_8 FILLER_66_2285 ();
 sg13g2_fill_1 FILLER_66_2292 ();
 sg13g2_fill_2 FILLER_66_2296 ();
 sg13g2_fill_1 FILLER_66_2304 ();
 sg13g2_decap_4 FILLER_66_2316 ();
 sg13g2_fill_1 FILLER_66_2320 ();
 sg13g2_decap_4 FILLER_66_2325 ();
 sg13g2_fill_2 FILLER_66_2329 ();
 sg13g2_fill_1 FILLER_66_2363 ();
 sg13g2_fill_2 FILLER_66_2395 ();
 sg13g2_fill_2 FILLER_66_2401 ();
 sg13g2_fill_1 FILLER_66_2408 ();
 sg13g2_fill_2 FILLER_66_2414 ();
 sg13g2_fill_2 FILLER_66_2424 ();
 sg13g2_decap_4 FILLER_66_2434 ();
 sg13g2_fill_2 FILLER_66_2442 ();
 sg13g2_fill_1 FILLER_66_2444 ();
 sg13g2_fill_2 FILLER_66_2454 ();
 sg13g2_fill_2 FILLER_66_2490 ();
 sg13g2_fill_1 FILLER_66_2496 ();
 sg13g2_fill_1 FILLER_66_2523 ();
 sg13g2_fill_2 FILLER_66_2548 ();
 sg13g2_fill_2 FILLER_66_2555 ();
 sg13g2_fill_1 FILLER_66_2557 ();
 sg13g2_fill_1 FILLER_66_2587 ();
 sg13g2_decap_8 FILLER_66_2651 ();
 sg13g2_decap_8 FILLER_66_2658 ();
 sg13g2_decap_4 FILLER_66_2665 ();
 sg13g2_fill_1 FILLER_66_2669 ();
 sg13g2_decap_4 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_30 ();
 sg13g2_decap_4 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_60 ();
 sg13g2_decap_8 FILLER_67_66 ();
 sg13g2_decap_8 FILLER_67_73 ();
 sg13g2_fill_1 FILLER_67_80 ();
 sg13g2_fill_2 FILLER_67_107 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_157 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_4 FILLER_67_203 ();
 sg13g2_fill_1 FILLER_67_207 ();
 sg13g2_fill_1 FILLER_67_216 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_229 ();
 sg13g2_fill_2 FILLER_67_234 ();
 sg13g2_fill_1 FILLER_67_267 ();
 sg13g2_decap_4 FILLER_67_273 ();
 sg13g2_fill_2 FILLER_67_277 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_fill_2 FILLER_67_289 ();
 sg13g2_fill_1 FILLER_67_296 ();
 sg13g2_fill_2 FILLER_67_312 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_1 FILLER_67_325 ();
 sg13g2_decap_4 FILLER_67_352 ();
 sg13g2_fill_1 FILLER_67_356 ();
 sg13g2_decap_8 FILLER_67_361 ();
 sg13g2_fill_2 FILLER_67_368 ();
 sg13g2_fill_1 FILLER_67_370 ();
 sg13g2_decap_4 FILLER_67_375 ();
 sg13g2_fill_1 FILLER_67_379 ();
 sg13g2_fill_1 FILLER_67_409 ();
 sg13g2_fill_1 FILLER_67_424 ();
 sg13g2_fill_1 FILLER_67_451 ();
 sg13g2_fill_2 FILLER_67_482 ();
 sg13g2_fill_2 FILLER_67_526 ();
 sg13g2_fill_1 FILLER_67_528 ();
 sg13g2_fill_2 FILLER_67_581 ();
 sg13g2_fill_1 FILLER_67_623 ();
 sg13g2_fill_1 FILLER_67_629 ();
 sg13g2_fill_2 FILLER_67_638 ();
 sg13g2_fill_1 FILLER_67_764 ();
 sg13g2_fill_2 FILLER_67_796 ();
 sg13g2_decap_4 FILLER_67_824 ();
 sg13g2_fill_2 FILLER_67_828 ();
 sg13g2_decap_8 FILLER_67_835 ();
 sg13g2_fill_2 FILLER_67_842 ();
 sg13g2_fill_1 FILLER_67_851 ();
 sg13g2_decap_8 FILLER_67_950 ();
 sg13g2_fill_2 FILLER_67_957 ();
 sg13g2_fill_2 FILLER_67_964 ();
 sg13g2_fill_1 FILLER_67_971 ();
 sg13g2_fill_2 FILLER_67_996 ();
 sg13g2_fill_2 FILLER_67_1005 ();
 sg13g2_decap_4 FILLER_67_1069 ();
 sg13g2_decap_8 FILLER_67_1103 ();
 sg13g2_fill_1 FILLER_67_1110 ();
 sg13g2_decap_8 FILLER_67_1150 ();
 sg13g2_decap_8 FILLER_67_1157 ();
 sg13g2_decap_4 FILLER_67_1164 ();
 sg13g2_fill_1 FILLER_67_1168 ();
 sg13g2_decap_8 FILLER_67_1225 ();
 sg13g2_fill_2 FILLER_67_1241 ();
 sg13g2_fill_1 FILLER_67_1276 ();
 sg13g2_decap_4 FILLER_67_1285 ();
 sg13g2_fill_1 FILLER_67_1289 ();
 sg13g2_fill_2 FILLER_67_1295 ();
 sg13g2_fill_1 FILLER_67_1297 ();
 sg13g2_decap_4 FILLER_67_1310 ();
 sg13g2_fill_1 FILLER_67_1314 ();
 sg13g2_decap_8 FILLER_67_1322 ();
 sg13g2_decap_8 FILLER_67_1329 ();
 sg13g2_decap_4 FILLER_67_1336 ();
 sg13g2_fill_2 FILLER_67_1340 ();
 sg13g2_fill_1 FILLER_67_1380 ();
 sg13g2_decap_4 FILLER_67_1387 ();
 sg13g2_fill_2 FILLER_67_1391 ();
 sg13g2_decap_8 FILLER_67_1413 ();
 sg13g2_decap_8 FILLER_67_1420 ();
 sg13g2_decap_4 FILLER_67_1427 ();
 sg13g2_fill_2 FILLER_67_1431 ();
 sg13g2_decap_8 FILLER_67_1437 ();
 sg13g2_decap_8 FILLER_67_1444 ();
 sg13g2_decap_8 FILLER_67_1451 ();
 sg13g2_fill_1 FILLER_67_1458 ();
 sg13g2_fill_1 FILLER_67_1468 ();
 sg13g2_fill_2 FILLER_67_1494 ();
 sg13g2_fill_1 FILLER_67_1496 ();
 sg13g2_fill_1 FILLER_67_1500 ();
 sg13g2_decap_8 FILLER_67_1511 ();
 sg13g2_decap_4 FILLER_67_1518 ();
 sg13g2_decap_4 FILLER_67_1526 ();
 sg13g2_fill_1 FILLER_67_1530 ();
 sg13g2_fill_1 FILLER_67_1562 ();
 sg13g2_fill_1 FILLER_67_1585 ();
 sg13g2_fill_1 FILLER_67_1612 ();
 sg13g2_fill_2 FILLER_67_1643 ();
 sg13g2_decap_8 FILLER_67_1650 ();
 sg13g2_decap_4 FILLER_67_1657 ();
 sg13g2_fill_1 FILLER_67_1661 ();
 sg13g2_fill_2 FILLER_67_1667 ();
 sg13g2_fill_1 FILLER_67_1669 ();
 sg13g2_fill_2 FILLER_67_1680 ();
 sg13g2_fill_1 FILLER_67_1687 ();
 sg13g2_decap_4 FILLER_67_1693 ();
 sg13g2_fill_1 FILLER_67_1697 ();
 sg13g2_fill_2 FILLER_67_1708 ();
 sg13g2_decap_8 FILLER_67_1727 ();
 sg13g2_decap_8 FILLER_67_1734 ();
 sg13g2_decap_8 FILLER_67_1741 ();
 sg13g2_decap_8 FILLER_67_1748 ();
 sg13g2_decap_4 FILLER_67_1755 ();
 sg13g2_fill_1 FILLER_67_1759 ();
 sg13g2_fill_1 FILLER_67_1781 ();
 sg13g2_fill_1 FILLER_67_1790 ();
 sg13g2_fill_1 FILLER_67_1796 ();
 sg13g2_decap_8 FILLER_67_1820 ();
 sg13g2_fill_2 FILLER_67_1827 ();
 sg13g2_fill_1 FILLER_67_1829 ();
 sg13g2_decap_8 FILLER_67_1835 ();
 sg13g2_decap_8 FILLER_67_1842 ();
 sg13g2_decap_8 FILLER_67_1849 ();
 sg13g2_decap_4 FILLER_67_1856 ();
 sg13g2_fill_1 FILLER_67_1860 ();
 sg13g2_decap_4 FILLER_67_1866 ();
 sg13g2_fill_1 FILLER_67_1870 ();
 sg13g2_fill_1 FILLER_67_1890 ();
 sg13g2_fill_1 FILLER_67_1919 ();
 sg13g2_fill_1 FILLER_67_1926 ();
 sg13g2_decap_8 FILLER_67_1962 ();
 sg13g2_decap_8 FILLER_67_1969 ();
 sg13g2_fill_2 FILLER_67_1976 ();
 sg13g2_fill_1 FILLER_67_1978 ();
 sg13g2_fill_1 FILLER_67_2005 ();
 sg13g2_fill_2 FILLER_67_2009 ();
 sg13g2_fill_2 FILLER_67_2107 ();
 sg13g2_fill_1 FILLER_67_2119 ();
 sg13g2_decap_4 FILLER_67_2124 ();
 sg13g2_fill_1 FILLER_67_2128 ();
 sg13g2_decap_8 FILLER_67_2133 ();
 sg13g2_decap_8 FILLER_67_2140 ();
 sg13g2_fill_2 FILLER_67_2147 ();
 sg13g2_fill_1 FILLER_67_2191 ();
 sg13g2_fill_2 FILLER_67_2212 ();
 sg13g2_decap_8 FILLER_67_2246 ();
 sg13g2_decap_8 FILLER_67_2253 ();
 sg13g2_fill_2 FILLER_67_2260 ();
 sg13g2_fill_2 FILLER_67_2308 ();
 sg13g2_decap_8 FILLER_67_2345 ();
 sg13g2_fill_1 FILLER_67_2352 ();
 sg13g2_fill_1 FILLER_67_2358 ();
 sg13g2_decap_8 FILLER_67_2363 ();
 sg13g2_fill_2 FILLER_67_2370 ();
 sg13g2_decap_8 FILLER_67_2396 ();
 sg13g2_decap_8 FILLER_67_2403 ();
 sg13g2_decap_8 FILLER_67_2410 ();
 sg13g2_decap_8 FILLER_67_2417 ();
 sg13g2_fill_1 FILLER_67_2424 ();
 sg13g2_decap_4 FILLER_67_2429 ();
 sg13g2_fill_1 FILLER_67_2433 ();
 sg13g2_decap_4 FILLER_67_2439 ();
 sg13g2_fill_1 FILLER_67_2443 ();
 sg13g2_fill_2 FILLER_67_2451 ();
 sg13g2_fill_1 FILLER_67_2496 ();
 sg13g2_fill_1 FILLER_67_2549 ();
 sg13g2_fill_2 FILLER_67_2582 ();
 sg13g2_fill_2 FILLER_67_2624 ();
 sg13g2_decap_8 FILLER_67_2658 ();
 sg13g2_decap_4 FILLER_67_2665 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_2 ();
 sg13g2_decap_8 FILLER_68_38 ();
 sg13g2_decap_8 FILLER_68_45 ();
 sg13g2_fill_2 FILLER_68_52 ();
 sg13g2_decap_4 FILLER_68_75 ();
 sg13g2_fill_2 FILLER_68_79 ();
 sg13g2_fill_1 FILLER_68_106 ();
 sg13g2_decap_4 FILLER_68_112 ();
 sg13g2_decap_4 FILLER_68_120 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_fill_2 FILLER_68_137 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_174 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_decap_4 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_266 ();
 sg13g2_fill_1 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_331 ();
 sg13g2_fill_2 FILLER_68_338 ();
 sg13g2_fill_1 FILLER_68_340 ();
 sg13g2_decap_8 FILLER_68_345 ();
 sg13g2_decap_8 FILLER_68_352 ();
 sg13g2_decap_4 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_363 ();
 sg13g2_decap_8 FILLER_68_447 ();
 sg13g2_decap_8 FILLER_68_454 ();
 sg13g2_fill_1 FILLER_68_500 ();
 sg13g2_fill_1 FILLER_68_505 ();
 sg13g2_fill_1 FILLER_68_515 ();
 sg13g2_decap_4 FILLER_68_520 ();
 sg13g2_fill_1 FILLER_68_524 ();
 sg13g2_fill_2 FILLER_68_532 ();
 sg13g2_fill_2 FILLER_68_576 ();
 sg13g2_fill_1 FILLER_68_578 ();
 sg13g2_fill_1 FILLER_68_605 ();
 sg13g2_decap_4 FILLER_68_632 ();
 sg13g2_fill_2 FILLER_68_636 ();
 sg13g2_fill_1 FILLER_68_662 ();
 sg13g2_fill_2 FILLER_68_667 ();
 sg13g2_fill_2 FILLER_68_689 ();
 sg13g2_fill_1 FILLER_68_773 ();
 sg13g2_fill_2 FILLER_68_796 ();
 sg13g2_fill_2 FILLER_68_834 ();
 sg13g2_fill_1 FILLER_68_836 ();
 sg13g2_fill_1 FILLER_68_842 ();
 sg13g2_fill_2 FILLER_68_851 ();
 sg13g2_fill_1 FILLER_68_853 ();
 sg13g2_fill_1 FILLER_68_918 ();
 sg13g2_decap_8 FILLER_68_945 ();
 sg13g2_decap_8 FILLER_68_952 ();
 sg13g2_decap_8 FILLER_68_959 ();
 sg13g2_decap_8 FILLER_68_966 ();
 sg13g2_decap_4 FILLER_68_973 ();
 sg13g2_fill_1 FILLER_68_977 ();
 sg13g2_fill_1 FILLER_68_1008 ();
 sg13g2_fill_1 FILLER_68_1037 ();
 sg13g2_fill_2 FILLER_68_1048 ();
 sg13g2_fill_1 FILLER_68_1050 ();
 sg13g2_fill_1 FILLER_68_1077 ();
 sg13g2_decap_4 FILLER_68_1130 ();
 sg13g2_fill_2 FILLER_68_1160 ();
 sg13g2_fill_1 FILLER_68_1162 ();
 sg13g2_fill_2 FILLER_68_1172 ();
 sg13g2_fill_1 FILLER_68_1174 ();
 sg13g2_decap_4 FILLER_68_1179 ();
 sg13g2_fill_1 FILLER_68_1183 ();
 sg13g2_decap_4 FILLER_68_1188 ();
 sg13g2_fill_2 FILLER_68_1222 ();
 sg13g2_fill_1 FILLER_68_1224 ();
 sg13g2_fill_2 FILLER_68_1251 ();
 sg13g2_fill_2 FILLER_68_1258 ();
 sg13g2_fill_2 FILLER_68_1291 ();
 sg13g2_fill_1 FILLER_68_1293 ();
 sg13g2_fill_2 FILLER_68_1305 ();
 sg13g2_fill_1 FILLER_68_1307 ();
 sg13g2_fill_1 FILLER_68_1324 ();
 sg13g2_fill_2 FILLER_68_1333 ();
 sg13g2_fill_1 FILLER_68_1335 ();
 sg13g2_decap_8 FILLER_68_1341 ();
 sg13g2_fill_1 FILLER_68_1385 ();
 sg13g2_fill_1 FILLER_68_1415 ();
 sg13g2_decap_8 FILLER_68_1430 ();
 sg13g2_fill_2 FILLER_68_1437 ();
 sg13g2_fill_1 FILLER_68_1447 ();
 sg13g2_fill_1 FILLER_68_1474 ();
 sg13g2_decap_8 FILLER_68_1489 ();
 sg13g2_fill_2 FILLER_68_1496 ();
 sg13g2_fill_1 FILLER_68_1498 ();
 sg13g2_decap_8 FILLER_68_1512 ();
 sg13g2_fill_2 FILLER_68_1519 ();
 sg13g2_fill_1 FILLER_68_1564 ();
 sg13g2_fill_2 FILLER_68_1570 ();
 sg13g2_fill_2 FILLER_68_1578 ();
 sg13g2_fill_2 FILLER_68_1584 ();
 sg13g2_decap_8 FILLER_68_1632 ();
 sg13g2_fill_1 FILLER_68_1639 ();
 sg13g2_fill_2 FILLER_68_1644 ();
 sg13g2_fill_1 FILLER_68_1646 ();
 sg13g2_decap_8 FILLER_68_1677 ();
 sg13g2_decap_4 FILLER_68_1684 ();
 sg13g2_fill_1 FILLER_68_1688 ();
 sg13g2_decap_8 FILLER_68_1694 ();
 sg13g2_decap_8 FILLER_68_1701 ();
 sg13g2_fill_2 FILLER_68_1721 ();
 sg13g2_fill_1 FILLER_68_1723 ();
 sg13g2_fill_1 FILLER_68_1729 ();
 sg13g2_fill_1 FILLER_68_1737 ();
 sg13g2_fill_1 FILLER_68_1746 ();
 sg13g2_decap_4 FILLER_68_1758 ();
 sg13g2_fill_2 FILLER_68_1762 ();
 sg13g2_decap_4 FILLER_68_1773 ();
 sg13g2_decap_4 FILLER_68_1814 ();
 sg13g2_decap_8 FILLER_68_1821 ();
 sg13g2_decap_8 FILLER_68_1828 ();
 sg13g2_decap_8 FILLER_68_1835 ();
 sg13g2_decap_8 FILLER_68_1842 ();
 sg13g2_decap_8 FILLER_68_1849 ();
 sg13g2_fill_2 FILLER_68_1856 ();
 sg13g2_fill_1 FILLER_68_1881 ();
 sg13g2_fill_1 FILLER_68_1886 ();
 sg13g2_fill_1 FILLER_68_1901 ();
 sg13g2_fill_2 FILLER_68_1917 ();
 sg13g2_fill_1 FILLER_68_1919 ();
 sg13g2_fill_2 FILLER_68_1943 ();
 sg13g2_fill_1 FILLER_68_1945 ();
 sg13g2_fill_1 FILLER_68_1955 ();
 sg13g2_decap_8 FILLER_68_1966 ();
 sg13g2_decap_8 FILLER_68_1973 ();
 sg13g2_decap_4 FILLER_68_1980 ();
 sg13g2_fill_2 FILLER_68_1984 ();
 sg13g2_fill_2 FILLER_68_1990 ();
 sg13g2_fill_1 FILLER_68_2005 ();
 sg13g2_fill_2 FILLER_68_2009 ();
 sg13g2_fill_1 FILLER_68_2030 ();
 sg13g2_fill_2 FILLER_68_2052 ();
 sg13g2_fill_1 FILLER_68_2087 ();
 sg13g2_decap_8 FILLER_68_2098 ();
 sg13g2_decap_8 FILLER_68_2105 ();
 sg13g2_fill_2 FILLER_68_2142 ();
 sg13g2_fill_1 FILLER_68_2144 ();
 sg13g2_decap_8 FILLER_68_2171 ();
 sg13g2_fill_1 FILLER_68_2178 ();
 sg13g2_fill_1 FILLER_68_2195 ();
 sg13g2_fill_1 FILLER_68_2217 ();
 sg13g2_fill_2 FILLER_68_2278 ();
 sg13g2_fill_1 FILLER_68_2280 ();
 sg13g2_fill_1 FILLER_68_2311 ();
 sg13g2_fill_2 FILLER_68_2329 ();
 sg13g2_fill_1 FILLER_68_2331 ();
 sg13g2_decap_4 FILLER_68_2337 ();
 sg13g2_fill_1 FILLER_68_2341 ();
 sg13g2_fill_2 FILLER_68_2350 ();
 sg13g2_decap_8 FILLER_68_2361 ();
 sg13g2_decap_4 FILLER_68_2368 ();
 sg13g2_fill_2 FILLER_68_2381 ();
 sg13g2_fill_1 FILLER_68_2383 ();
 sg13g2_fill_1 FILLER_68_2408 ();
 sg13g2_fill_2 FILLER_68_2413 ();
 sg13g2_fill_1 FILLER_68_2415 ();
 sg13g2_fill_1 FILLER_68_2447 ();
 sg13g2_fill_2 FILLER_68_2456 ();
 sg13g2_fill_2 FILLER_68_2488 ();
 sg13g2_fill_1 FILLER_68_2511 ();
 sg13g2_decap_4 FILLER_68_2517 ();
 sg13g2_fill_2 FILLER_68_2534 ();
 sg13g2_decap_8 FILLER_68_2540 ();
 sg13g2_decap_4 FILLER_68_2547 ();
 sg13g2_fill_2 FILLER_68_2551 ();
 sg13g2_fill_2 FILLER_68_2556 ();
 sg13g2_fill_1 FILLER_68_2581 ();
 sg13g2_fill_1 FILLER_68_2626 ();
 sg13g2_fill_2 FILLER_68_2668 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_12 ();
 sg13g2_fill_1 FILLER_69_17 ();
 sg13g2_fill_1 FILLER_69_44 ();
 sg13g2_fill_1 FILLER_69_71 ();
 sg13g2_decap_8 FILLER_69_92 ();
 sg13g2_decap_4 FILLER_69_104 ();
 sg13g2_decap_8 FILLER_69_123 ();
 sg13g2_decap_4 FILLER_69_130 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_decap_8 FILLER_69_174 ();
 sg13g2_decap_8 FILLER_69_181 ();
 sg13g2_decap_4 FILLER_69_188 ();
 sg13g2_decap_8 FILLER_69_207 ();
 sg13g2_fill_2 FILLER_69_214 ();
 sg13g2_fill_1 FILLER_69_216 ();
 sg13g2_fill_2 FILLER_69_230 ();
 sg13g2_fill_2 FILLER_69_237 ();
 sg13g2_fill_1 FILLER_69_239 ();
 sg13g2_fill_2 FILLER_69_250 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_258 ();
 sg13g2_fill_2 FILLER_69_271 ();
 sg13g2_fill_1 FILLER_69_291 ();
 sg13g2_decap_4 FILLER_69_335 ();
 sg13g2_fill_1 FILLER_69_339 ();
 sg13g2_decap_4 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_354 ();
 sg13g2_decap_4 FILLER_69_390 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_fill_2 FILLER_69_423 ();
 sg13g2_fill_1 FILLER_69_425 ();
 sg13g2_decap_4 FILLER_69_430 ();
 sg13g2_decap_4 FILLER_69_438 ();
 sg13g2_fill_2 FILLER_69_442 ();
 sg13g2_decap_8 FILLER_69_448 ();
 sg13g2_fill_2 FILLER_69_482 ();
 sg13g2_fill_1 FILLER_69_484 ();
 sg13g2_fill_1 FILLER_69_492 ();
 sg13g2_decap_8 FILLER_69_497 ();
 sg13g2_fill_2 FILLER_69_504 ();
 sg13g2_decap_8 FILLER_69_511 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_fill_2 FILLER_69_525 ();
 sg13g2_fill_1 FILLER_69_527 ();
 sg13g2_fill_2 FILLER_69_596 ();
 sg13g2_decap_8 FILLER_69_616 ();
 sg13g2_fill_2 FILLER_69_623 ();
 sg13g2_decap_8 FILLER_69_628 ();
 sg13g2_decap_4 FILLER_69_635 ();
 sg13g2_fill_2 FILLER_69_639 ();
 sg13g2_fill_2 FILLER_69_648 ();
 sg13g2_fill_2 FILLER_69_659 ();
 sg13g2_fill_1 FILLER_69_665 ();
 sg13g2_fill_2 FILLER_69_692 ();
 sg13g2_fill_2 FILLER_69_701 ();
 sg13g2_fill_2 FILLER_69_729 ();
 sg13g2_fill_1 FILLER_69_731 ();
 sg13g2_fill_1 FILLER_69_763 ();
 sg13g2_fill_2 FILLER_69_777 ();
 sg13g2_fill_1 FILLER_69_779 ();
 sg13g2_fill_1 FILLER_69_794 ();
 sg13g2_fill_2 FILLER_69_822 ();
 sg13g2_decap_8 FILLER_69_830 ();
 sg13g2_decap_8 FILLER_69_927 ();
 sg13g2_fill_1 FILLER_69_934 ();
 sg13g2_decap_4 FILLER_69_972 ();
 sg13g2_fill_2 FILLER_69_976 ();
 sg13g2_fill_2 FILLER_69_982 ();
 sg13g2_fill_1 FILLER_69_984 ();
 sg13g2_decap_4 FILLER_69_998 ();
 sg13g2_fill_1 FILLER_69_1002 ();
 sg13g2_decap_4 FILLER_69_1035 ();
 sg13g2_fill_2 FILLER_69_1059 ();
 sg13g2_fill_1 FILLER_69_1061 ();
 sg13g2_decap_4 FILLER_69_1066 ();
 sg13g2_fill_1 FILLER_69_1070 ();
 sg13g2_fill_2 FILLER_69_1084 ();
 sg13g2_fill_1 FILLER_69_1091 ();
 sg13g2_fill_1 FILLER_69_1117 ();
 sg13g2_fill_2 FILLER_69_1122 ();
 sg13g2_decap_8 FILLER_69_1184 ();
 sg13g2_decap_8 FILLER_69_1191 ();
 sg13g2_decap_8 FILLER_69_1198 ();
 sg13g2_decap_8 FILLER_69_1205 ();
 sg13g2_decap_8 FILLER_69_1212 ();
 sg13g2_fill_2 FILLER_69_1228 ();
 sg13g2_fill_1 FILLER_69_1230 ();
 sg13g2_fill_1 FILLER_69_1239 ();
 sg13g2_fill_2 FILLER_69_1243 ();
 sg13g2_fill_2 FILLER_69_1252 ();
 sg13g2_decap_8 FILLER_69_1262 ();
 sg13g2_fill_2 FILLER_69_1273 ();
 sg13g2_decap_8 FILLER_69_1333 ();
 sg13g2_fill_1 FILLER_69_1391 ();
 sg13g2_fill_1 FILLER_69_1419 ();
 sg13g2_decap_4 FILLER_69_1424 ();
 sg13g2_decap_8 FILLER_69_1433 ();
 sg13g2_fill_1 FILLER_69_1440 ();
 sg13g2_decap_4 FILLER_69_1445 ();
 sg13g2_fill_2 FILLER_69_1449 ();
 sg13g2_decap_4 FILLER_69_1456 ();
 sg13g2_fill_1 FILLER_69_1465 ();
 sg13g2_fill_2 FILLER_69_1476 ();
 sg13g2_decap_8 FILLER_69_1483 ();
 sg13g2_decap_4 FILLER_69_1490 ();
 sg13g2_fill_2 FILLER_69_1498 ();
 sg13g2_fill_1 FILLER_69_1500 ();
 sg13g2_decap_8 FILLER_69_1510 ();
 sg13g2_decap_4 FILLER_69_1517 ();
 sg13g2_fill_2 FILLER_69_1521 ();
 sg13g2_decap_4 FILLER_69_1535 ();
 sg13g2_fill_1 FILLER_69_1552 ();
 sg13g2_decap_8 FILLER_69_1558 ();
 sg13g2_fill_2 FILLER_69_1565 ();
 sg13g2_decap_8 FILLER_69_1574 ();
 sg13g2_fill_2 FILLER_69_1586 ();
 sg13g2_fill_1 FILLER_69_1593 ();
 sg13g2_decap_8 FILLER_69_1598 ();
 sg13g2_fill_2 FILLER_69_1605 ();
 sg13g2_fill_1 FILLER_69_1607 ();
 sg13g2_decap_8 FILLER_69_1612 ();
 sg13g2_decap_4 FILLER_69_1619 ();
 sg13g2_fill_1 FILLER_69_1631 ();
 sg13g2_decap_8 FILLER_69_1639 ();
 sg13g2_decap_8 FILLER_69_1646 ();
 sg13g2_decap_4 FILLER_69_1653 ();
 sg13g2_decap_8 FILLER_69_1661 ();
 sg13g2_decap_8 FILLER_69_1668 ();
 sg13g2_decap_4 FILLER_69_1675 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_decap_8 FILLER_69_1692 ();
 sg13g2_decap_8 FILLER_69_1699 ();
 sg13g2_decap_8 FILLER_69_1706 ();
 sg13g2_decap_4 FILLER_69_1713 ();
 sg13g2_fill_1 FILLER_69_1717 ();
 sg13g2_decap_4 FILLER_69_1726 ();
 sg13g2_fill_1 FILLER_69_1730 ();
 sg13g2_fill_1 FILLER_69_1735 ();
 sg13g2_fill_2 FILLER_69_1746 ();
 sg13g2_fill_2 FILLER_69_1776 ();
 sg13g2_fill_1 FILLER_69_1778 ();
 sg13g2_fill_2 FILLER_69_1793 ();
 sg13g2_fill_2 FILLER_69_1824 ();
 sg13g2_fill_2 FILLER_69_1835 ();
 sg13g2_fill_2 FILLER_69_1842 ();
 sg13g2_decap_8 FILLER_69_1849 ();
 sg13g2_fill_2 FILLER_69_1856 ();
 sg13g2_decap_8 FILLER_69_1863 ();
 sg13g2_fill_2 FILLER_69_1879 ();
 sg13g2_fill_1 FILLER_69_1908 ();
 sg13g2_fill_1 FILLER_69_1919 ();
 sg13g2_fill_2 FILLER_69_1925 ();
 sg13g2_fill_2 FILLER_69_1970 ();
 sg13g2_fill_1 FILLER_69_1972 ();
 sg13g2_decap_4 FILLER_69_1977 ();
 sg13g2_fill_2 FILLER_69_1981 ();
 sg13g2_fill_2 FILLER_69_1987 ();
 sg13g2_fill_1 FILLER_69_1989 ();
 sg13g2_fill_1 FILLER_69_1995 ();
 sg13g2_fill_1 FILLER_69_2037 ();
 sg13g2_fill_2 FILLER_69_2074 ();
 sg13g2_fill_1 FILLER_69_2076 ();
 sg13g2_decap_8 FILLER_69_2123 ();
 sg13g2_fill_1 FILLER_69_2130 ();
 sg13g2_decap_4 FILLER_69_2167 ();
 sg13g2_decap_8 FILLER_69_2175 ();
 sg13g2_decap_8 FILLER_69_2182 ();
 sg13g2_fill_1 FILLER_69_2240 ();
 sg13g2_decap_4 FILLER_69_2255 ();
 sg13g2_fill_1 FILLER_69_2259 ();
 sg13g2_decap_4 FILLER_69_2270 ();
 sg13g2_decap_8 FILLER_69_2288 ();
 sg13g2_decap_8 FILLER_69_2295 ();
 sg13g2_decap_4 FILLER_69_2302 ();
 sg13g2_fill_1 FILLER_69_2306 ();
 sg13g2_fill_2 FILLER_69_2341 ();
 sg13g2_fill_1 FILLER_69_2343 ();
 sg13g2_fill_1 FILLER_69_2349 ();
 sg13g2_fill_2 FILLER_69_2376 ();
 sg13g2_fill_1 FILLER_69_2423 ();
 sg13g2_decap_4 FILLER_69_2443 ();
 sg13g2_fill_1 FILLER_69_2471 ();
 sg13g2_decap_4 FILLER_69_2502 ();
 sg13g2_fill_1 FILLER_69_2506 ();
 sg13g2_fill_1 FILLER_69_2512 ();
 sg13g2_decap_8 FILLER_69_2522 ();
 sg13g2_fill_1 FILLER_69_2529 ();
 sg13g2_fill_2 FILLER_69_2534 ();
 sg13g2_fill_1 FILLER_69_2536 ();
 sg13g2_decap_4 FILLER_69_2560 ();
 sg13g2_fill_1 FILLER_69_2567 ();
 sg13g2_fill_2 FILLER_69_2592 ();
 sg13g2_fill_1 FILLER_69_2636 ();
 sg13g2_fill_1 FILLER_69_2647 ();
 sg13g2_decap_8 FILLER_69_2655 ();
 sg13g2_decap_8 FILLER_69_2662 ();
 sg13g2_fill_1 FILLER_69_2669 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_1 FILLER_70_37 ();
 sg13g2_fill_1 FILLER_70_48 ();
 sg13g2_fill_2 FILLER_70_79 ();
 sg13g2_decap_4 FILLER_70_85 ();
 sg13g2_fill_1 FILLER_70_115 ();
 sg13g2_fill_2 FILLER_70_121 ();
 sg13g2_fill_1 FILLER_70_123 ();
 sg13g2_fill_1 FILLER_70_142 ();
 sg13g2_decap_4 FILLER_70_148 ();
 sg13g2_fill_1 FILLER_70_152 ();
 sg13g2_fill_1 FILLER_70_206 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_4 FILLER_70_238 ();
 sg13g2_fill_2 FILLER_70_242 ();
 sg13g2_fill_1 FILLER_70_249 ();
 sg13g2_decap_4 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_258 ();
 sg13g2_fill_2 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_283 ();
 sg13g2_decap_8 FILLER_70_290 ();
 sg13g2_decap_4 FILLER_70_297 ();
 sg13g2_fill_1 FILLER_70_301 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_318 ();
 sg13g2_fill_1 FILLER_70_324 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_1 FILLER_70_337 ();
 sg13g2_fill_2 FILLER_70_343 ();
 sg13g2_decap_4 FILLER_70_349 ();
 sg13g2_fill_2 FILLER_70_353 ();
 sg13g2_decap_4 FILLER_70_359 ();
 sg13g2_fill_1 FILLER_70_363 ();
 sg13g2_fill_2 FILLER_70_372 ();
 sg13g2_decap_4 FILLER_70_378 ();
 sg13g2_decap_4 FILLER_70_386 ();
 sg13g2_decap_8 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_70_426 ();
 sg13g2_decap_4 FILLER_70_433 ();
 sg13g2_fill_1 FILLER_70_509 ();
 sg13g2_fill_1 FILLER_70_546 ();
 sg13g2_fill_1 FILLER_70_550 ();
 sg13g2_fill_2 FILLER_70_555 ();
 sg13g2_fill_1 FILLER_70_557 ();
 sg13g2_fill_2 FILLER_70_563 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_604 ();
 sg13g2_fill_2 FILLER_70_618 ();
 sg13g2_fill_2 FILLER_70_624 ();
 sg13g2_fill_2 FILLER_70_678 ();
 sg13g2_decap_8 FILLER_70_702 ();
 sg13g2_fill_1 FILLER_70_709 ();
 sg13g2_fill_2 FILLER_70_718 ();
 sg13g2_fill_1 FILLER_70_763 ();
 sg13g2_fill_2 FILLER_70_768 ();
 sg13g2_fill_2 FILLER_70_784 ();
 sg13g2_fill_2 FILLER_70_795 ();
 sg13g2_decap_4 FILLER_70_807 ();
 sg13g2_decap_4 FILLER_70_815 ();
 sg13g2_decap_8 FILLER_70_831 ();
 sg13g2_decap_4 FILLER_70_842 ();
 sg13g2_fill_2 FILLER_70_851 ();
 sg13g2_decap_8 FILLER_70_865 ();
 sg13g2_fill_1 FILLER_70_872 ();
 sg13g2_decap_8 FILLER_70_879 ();
 sg13g2_fill_2 FILLER_70_890 ();
 sg13g2_fill_2 FILLER_70_895 ();
 sg13g2_fill_1 FILLER_70_897 ();
 sg13g2_decap_8 FILLER_70_928 ();
 sg13g2_decap_8 FILLER_70_935 ();
 sg13g2_decap_4 FILLER_70_942 ();
 sg13g2_decap_4 FILLER_70_951 ();
 sg13g2_fill_1 FILLER_70_969 ();
 sg13g2_decap_4 FILLER_70_975 ();
 sg13g2_fill_1 FILLER_70_979 ();
 sg13g2_decap_8 FILLER_70_1063 ();
 sg13g2_decap_4 FILLER_70_1070 ();
 sg13g2_fill_2 FILLER_70_1074 ();
 sg13g2_decap_8 FILLER_70_1114 ();
 sg13g2_fill_1 FILLER_70_1121 ();
 sg13g2_fill_2 FILLER_70_1132 ();
 sg13g2_fill_1 FILLER_70_1134 ();
 sg13g2_fill_1 FILLER_70_1148 ();
 sg13g2_fill_1 FILLER_70_1157 ();
 sg13g2_fill_2 FILLER_70_1161 ();
 sg13g2_fill_1 FILLER_70_1163 ();
 sg13g2_decap_8 FILLER_70_1167 ();
 sg13g2_decap_8 FILLER_70_1174 ();
 sg13g2_fill_2 FILLER_70_1181 ();
 sg13g2_decap_4 FILLER_70_1208 ();
 sg13g2_fill_2 FILLER_70_1212 ();
 sg13g2_fill_1 FILLER_70_1263 ();
 sg13g2_decap_4 FILLER_70_1289 ();
 sg13g2_fill_2 FILLER_70_1304 ();
 sg13g2_fill_1 FILLER_70_1310 ();
 sg13g2_fill_2 FILLER_70_1318 ();
 sg13g2_fill_1 FILLER_70_1325 ();
 sg13g2_fill_2 FILLER_70_1364 ();
 sg13g2_decap_4 FILLER_70_1376 ();
 sg13g2_fill_2 FILLER_70_1380 ();
 sg13g2_decap_4 FILLER_70_1400 ();
 sg13g2_fill_2 FILLER_70_1404 ();
 sg13g2_fill_1 FILLER_70_1423 ();
 sg13g2_decap_4 FILLER_70_1440 ();
 sg13g2_decap_8 FILLER_70_1449 ();
 sg13g2_fill_1 FILLER_70_1456 ();
 sg13g2_fill_1 FILLER_70_1461 ();
 sg13g2_decap_4 FILLER_70_1483 ();
 sg13g2_fill_2 FILLER_70_1492 ();
 sg13g2_fill_1 FILLER_70_1494 ();
 sg13g2_decap_4 FILLER_70_1535 ();
 sg13g2_decap_4 FILLER_70_1553 ();
 sg13g2_fill_1 FILLER_70_1557 ();
 sg13g2_decap_4 FILLER_70_1580 ();
 sg13g2_fill_1 FILLER_70_1589 ();
 sg13g2_fill_1 FILLER_70_1595 ();
 sg13g2_decap_8 FILLER_70_1601 ();
 sg13g2_decap_4 FILLER_70_1608 ();
 sg13g2_decap_4 FILLER_70_1617 ();
 sg13g2_fill_1 FILLER_70_1621 ();
 sg13g2_fill_2 FILLER_70_1629 ();
 sg13g2_fill_2 FILLER_70_1652 ();
 sg13g2_fill_1 FILLER_70_1654 ();
 sg13g2_decap_8 FILLER_70_1662 ();
 sg13g2_decap_8 FILLER_70_1669 ();
 sg13g2_fill_2 FILLER_70_1676 ();
 sg13g2_fill_1 FILLER_70_1678 ();
 sg13g2_decap_4 FILLER_70_1683 ();
 sg13g2_decap_8 FILLER_70_1691 ();
 sg13g2_decap_4 FILLER_70_1698 ();
 sg13g2_fill_2 FILLER_70_1702 ();
 sg13g2_decap_4 FILLER_70_1708 ();
 sg13g2_fill_2 FILLER_70_1712 ();
 sg13g2_decap_8 FILLER_70_1719 ();
 sg13g2_fill_2 FILLER_70_1726 ();
 sg13g2_fill_1 FILLER_70_1740 ();
 sg13g2_fill_1 FILLER_70_1744 ();
 sg13g2_fill_1 FILLER_70_1750 ();
 sg13g2_fill_2 FILLER_70_1775 ();
 sg13g2_fill_1 FILLER_70_1798 ();
 sg13g2_fill_1 FILLER_70_1817 ();
 sg13g2_fill_2 FILLER_70_1823 ();
 sg13g2_fill_1 FILLER_70_1830 ();
 sg13g2_fill_2 FILLER_70_1839 ();
 sg13g2_fill_1 FILLER_70_1850 ();
 sg13g2_decap_8 FILLER_70_1861 ();
 sg13g2_decap_8 FILLER_70_1868 ();
 sg13g2_decap_4 FILLER_70_1875 ();
 sg13g2_fill_2 FILLER_70_1885 ();
 sg13g2_decap_4 FILLER_70_1900 ();
 sg13g2_fill_1 FILLER_70_1904 ();
 sg13g2_fill_2 FILLER_70_1917 ();
 sg13g2_fill_1 FILLER_70_1943 ();
 sg13g2_fill_2 FILLER_70_1948 ();
 sg13g2_decap_8 FILLER_70_1971 ();
 sg13g2_decap_8 FILLER_70_1978 ();
 sg13g2_decap_4 FILLER_70_1985 ();
 sg13g2_fill_2 FILLER_70_1993 ();
 sg13g2_fill_2 FILLER_70_2011 ();
 sg13g2_decap_4 FILLER_70_2047 ();
 sg13g2_fill_2 FILLER_70_2051 ();
 sg13g2_fill_1 FILLER_70_2057 ();
 sg13g2_decap_8 FILLER_70_2111 ();
 sg13g2_decap_4 FILLER_70_2118 ();
 sg13g2_decap_8 FILLER_70_2132 ();
 sg13g2_fill_2 FILLER_70_2139 ();
 sg13g2_decap_4 FILLER_70_2158 ();
 sg13g2_fill_2 FILLER_70_2162 ();
 sg13g2_decap_8 FILLER_70_2190 ();
 sg13g2_decap_4 FILLER_70_2234 ();
 sg13g2_fill_2 FILLER_70_2238 ();
 sg13g2_decap_8 FILLER_70_2266 ();
 sg13g2_fill_2 FILLER_70_2273 ();
 sg13g2_fill_1 FILLER_70_2275 ();
 sg13g2_fill_2 FILLER_70_2302 ();
 sg13g2_fill_1 FILLER_70_2304 ();
 sg13g2_decap_4 FILLER_70_2309 ();
 sg13g2_fill_2 FILLER_70_2313 ();
 sg13g2_fill_2 FILLER_70_2361 ();
 sg13g2_fill_1 FILLER_70_2363 ();
 sg13g2_fill_1 FILLER_70_2426 ();
 sg13g2_fill_2 FILLER_70_2456 ();
 sg13g2_decap_8 FILLER_70_2496 ();
 sg13g2_fill_2 FILLER_70_2503 ();
 sg13g2_fill_1 FILLER_70_2505 ();
 sg13g2_decap_4 FILLER_70_2511 ();
 sg13g2_decap_8 FILLER_70_2546 ();
 sg13g2_decap_8 FILLER_70_2553 ();
 sg13g2_decap_4 FILLER_70_2560 ();
 sg13g2_fill_1 FILLER_70_2593 ();
 sg13g2_fill_1 FILLER_70_2599 ();
 sg13g2_fill_2 FILLER_70_2618 ();
 sg13g2_decap_4 FILLER_70_2666 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_decap_8 FILLER_71_48 ();
 sg13g2_decap_4 FILLER_71_69 ();
 sg13g2_fill_2 FILLER_71_94 ();
 sg13g2_fill_1 FILLER_71_96 ();
 sg13g2_fill_1 FILLER_71_128 ();
 sg13g2_fill_2 FILLER_71_181 ();
 sg13g2_fill_1 FILLER_71_183 ();
 sg13g2_decap_4 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_234 ();
 sg13g2_fill_2 FILLER_71_245 ();
 sg13g2_fill_1 FILLER_71_247 ();
 sg13g2_fill_2 FILLER_71_251 ();
 sg13g2_fill_1 FILLER_71_253 ();
 sg13g2_fill_2 FILLER_71_267 ();
 sg13g2_fill_1 FILLER_71_269 ();
 sg13g2_decap_4 FILLER_71_275 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_fill_2 FILLER_71_301 ();
 sg13g2_fill_1 FILLER_71_303 ();
 sg13g2_decap_4 FILLER_71_309 ();
 sg13g2_fill_1 FILLER_71_313 ();
 sg13g2_decap_8 FILLER_71_326 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_335 ();
 sg13g2_fill_2 FILLER_71_346 ();
 sg13g2_fill_1 FILLER_71_348 ();
 sg13g2_decap_4 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_393 ();
 sg13g2_fill_2 FILLER_71_400 ();
 sg13g2_decap_4 FILLER_71_419 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_fill_2 FILLER_71_450 ();
 sg13g2_fill_1 FILLER_71_452 ();
 sg13g2_fill_1 FILLER_71_530 ();
 sg13g2_fill_2 FILLER_71_544 ();
 sg13g2_fill_1 FILLER_71_546 ();
 sg13g2_fill_2 FILLER_71_560 ();
 sg13g2_fill_1 FILLER_71_562 ();
 sg13g2_fill_2 FILLER_71_567 ();
 sg13g2_fill_1 FILLER_71_588 ();
 sg13g2_fill_1 FILLER_71_595 ();
 sg13g2_fill_2 FILLER_71_675 ();
 sg13g2_decap_4 FILLER_71_689 ();
 sg13g2_fill_1 FILLER_71_693 ();
 sg13g2_fill_1 FILLER_71_699 ();
 sg13g2_decap_8 FILLER_71_708 ();
 sg13g2_decap_8 FILLER_71_715 ();
 sg13g2_decap_4 FILLER_71_722 ();
 sg13g2_fill_2 FILLER_71_726 ();
 sg13g2_fill_1 FILLER_71_754 ();
 sg13g2_fill_2 FILLER_71_781 ();
 sg13g2_fill_2 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_829 ();
 sg13g2_decap_8 FILLER_71_836 ();
 sg13g2_decap_4 FILLER_71_843 ();
 sg13g2_fill_1 FILLER_71_847 ();
 sg13g2_decap_4 FILLER_71_872 ();
 sg13g2_fill_1 FILLER_71_876 ();
 sg13g2_decap_4 FILLER_71_882 ();
 sg13g2_fill_2 FILLER_71_886 ();
 sg13g2_fill_1 FILLER_71_970 ();
 sg13g2_fill_1 FILLER_71_997 ();
 sg13g2_fill_1 FILLER_71_1003 ();
 sg13g2_fill_1 FILLER_71_1008 ();
 sg13g2_fill_2 FILLER_71_1017 ();
 sg13g2_decap_8 FILLER_71_1036 ();
 sg13g2_decap_8 FILLER_71_1043 ();
 sg13g2_decap_8 FILLER_71_1050 ();
 sg13g2_decap_8 FILLER_71_1057 ();
 sg13g2_decap_8 FILLER_71_1064 ();
 sg13g2_decap_8 FILLER_71_1071 ();
 sg13g2_decap_4 FILLER_71_1078 ();
 sg13g2_fill_1 FILLER_71_1082 ();
 sg13g2_fill_1 FILLER_71_1092 ();
 sg13g2_fill_1 FILLER_71_1097 ();
 sg13g2_decap_8 FILLER_71_1107 ();
 sg13g2_decap_4 FILLER_71_1114 ();
 sg13g2_fill_1 FILLER_71_1157 ();
 sg13g2_fill_2 FILLER_71_1171 ();
 sg13g2_fill_1 FILLER_71_1173 ();
 sg13g2_fill_1 FILLER_71_1193 ();
 sg13g2_decap_4 FILLER_71_1220 ();
 sg13g2_fill_2 FILLER_71_1236 ();
 sg13g2_fill_1 FILLER_71_1238 ();
 sg13g2_fill_1 FILLER_71_1243 ();
 sg13g2_fill_2 FILLER_71_1255 ();
 sg13g2_fill_2 FILLER_71_1262 ();
 sg13g2_fill_1 FILLER_71_1264 ();
 sg13g2_fill_1 FILLER_71_1273 ();
 sg13g2_fill_1 FILLER_71_1278 ();
 sg13g2_fill_1 FILLER_71_1283 ();
 sg13g2_fill_1 FILLER_71_1306 ();
 sg13g2_decap_8 FILLER_71_1312 ();
 sg13g2_decap_8 FILLER_71_1319 ();
 sg13g2_decap_4 FILLER_71_1326 ();
 sg13g2_fill_2 FILLER_71_1330 ();
 sg13g2_decap_8 FILLER_71_1340 ();
 sg13g2_decap_4 FILLER_71_1347 ();
 sg13g2_decap_8 FILLER_71_1369 ();
 sg13g2_decap_8 FILLER_71_1376 ();
 sg13g2_decap_8 FILLER_71_1383 ();
 sg13g2_decap_8 FILLER_71_1390 ();
 sg13g2_fill_2 FILLER_71_1397 ();
 sg13g2_fill_1 FILLER_71_1399 ();
 sg13g2_fill_1 FILLER_71_1420 ();
 sg13g2_fill_2 FILLER_71_1436 ();
 sg13g2_fill_1 FILLER_71_1443 ();
 sg13g2_fill_1 FILLER_71_1453 ();
 sg13g2_fill_1 FILLER_71_1458 ();
 sg13g2_fill_1 FILLER_71_1471 ();
 sg13g2_fill_2 FILLER_71_1484 ();
 sg13g2_fill_1 FILLER_71_1491 ();
 sg13g2_fill_2 FILLER_71_1501 ();
 sg13g2_fill_1 FILLER_71_1511 ();
 sg13g2_fill_1 FILLER_71_1526 ();
 sg13g2_decap_4 FILLER_71_1535 ();
 sg13g2_fill_2 FILLER_71_1539 ();
 sg13g2_fill_2 FILLER_71_1593 ();
 sg13g2_fill_2 FILLER_71_1600 ();
 sg13g2_fill_1 FILLER_71_1606 ();
 sg13g2_fill_2 FILLER_71_1612 ();
 sg13g2_fill_1 FILLER_71_1614 ();
 sg13g2_fill_2 FILLER_71_1620 ();
 sg13g2_fill_1 FILLER_71_1622 ();
 sg13g2_fill_2 FILLER_71_1628 ();
 sg13g2_fill_2 FILLER_71_1656 ();
 sg13g2_fill_1 FILLER_71_1658 ();
 sg13g2_decap_4 FILLER_71_1668 ();
 sg13g2_fill_2 FILLER_71_1672 ();
 sg13g2_fill_2 FILLER_71_1683 ();
 sg13g2_fill_1 FILLER_71_1685 ();
 sg13g2_fill_2 FILLER_71_1692 ();
 sg13g2_fill_1 FILLER_71_1694 ();
 sg13g2_decap_4 FILLER_71_1703 ();
 sg13g2_decap_8 FILLER_71_1712 ();
 sg13g2_decap_4 FILLER_71_1719 ();
 sg13g2_fill_2 FILLER_71_1723 ();
 sg13g2_fill_2 FILLER_71_1729 ();
 sg13g2_fill_1 FILLER_71_1748 ();
 sg13g2_fill_1 FILLER_71_1755 ();
 sg13g2_fill_1 FILLER_71_1761 ();
 sg13g2_fill_1 FILLER_71_1767 ();
 sg13g2_fill_1 FILLER_71_1782 ();
 sg13g2_fill_1 FILLER_71_1787 ();
 sg13g2_fill_1 FILLER_71_1814 ();
 sg13g2_fill_2 FILLER_71_1823 ();
 sg13g2_fill_1 FILLER_71_1825 ();
 sg13g2_fill_2 FILLER_71_1831 ();
 sg13g2_fill_1 FILLER_71_1833 ();
 sg13g2_decap_8 FILLER_71_1839 ();
 sg13g2_fill_1 FILLER_71_1846 ();
 sg13g2_fill_2 FILLER_71_1863 ();
 sg13g2_fill_1 FILLER_71_1871 ();
 sg13g2_fill_1 FILLER_71_1881 ();
 sg13g2_fill_1 FILLER_71_1892 ();
 sg13g2_fill_2 FILLER_71_1902 ();
 sg13g2_fill_1 FILLER_71_1912 ();
 sg13g2_fill_1 FILLER_71_1937 ();
 sg13g2_fill_1 FILLER_71_1956 ();
 sg13g2_decap_8 FILLER_71_1976 ();
 sg13g2_fill_1 FILLER_71_1983 ();
 sg13g2_fill_1 FILLER_71_2090 ();
 sg13g2_fill_2 FILLER_71_2112 ();
 sg13g2_decap_8 FILLER_71_2190 ();
 sg13g2_decap_8 FILLER_71_2197 ();
 sg13g2_fill_2 FILLER_71_2204 ();
 sg13g2_decap_4 FILLER_71_2216 ();
 sg13g2_fill_2 FILLER_71_2220 ();
 sg13g2_decap_8 FILLER_71_2227 ();
 sg13g2_decap_4 FILLER_71_2234 ();
 sg13g2_decap_4 FILLER_71_2251 ();
 sg13g2_fill_1 FILLER_71_2255 ();
 sg13g2_decap_8 FILLER_71_2282 ();
 sg13g2_fill_1 FILLER_71_2289 ();
 sg13g2_fill_1 FILLER_71_2329 ();
 sg13g2_fill_1 FILLER_71_2338 ();
 sg13g2_decap_4 FILLER_71_2343 ();
 sg13g2_fill_2 FILLER_71_2397 ();
 sg13g2_fill_1 FILLER_71_2450 ();
 sg13g2_fill_2 FILLER_71_2464 ();
 sg13g2_decap_8 FILLER_71_2484 ();
 sg13g2_fill_1 FILLER_71_2491 ();
 sg13g2_fill_1 FILLER_71_2497 ();
 sg13g2_fill_1 FILLER_71_2502 ();
 sg13g2_fill_1 FILLER_71_2509 ();
 sg13g2_fill_2 FILLER_71_2515 ();
 sg13g2_decap_4 FILLER_71_2521 ();
 sg13g2_fill_1 FILLER_71_2525 ();
 sg13g2_decap_8 FILLER_71_2612 ();
 sg13g2_fill_1 FILLER_71_2619 ();
 sg13g2_decap_4 FILLER_71_2666 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_11 ();
 sg13g2_fill_2 FILLER_72_17 ();
 sg13g2_fill_1 FILLER_72_19 ();
 sg13g2_decap_8 FILLER_72_72 ();
 sg13g2_decap_8 FILLER_72_79 ();
 sg13g2_decap_8 FILLER_72_86 ();
 sg13g2_decap_8 FILLER_72_93 ();
 sg13g2_decap_8 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_107 ();
 sg13g2_fill_2 FILLER_72_114 ();
 sg13g2_decap_4 FILLER_72_134 ();
 sg13g2_fill_2 FILLER_72_138 ();
 sg13g2_fill_2 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_156 ();
 sg13g2_fill_1 FILLER_72_160 ();
 sg13g2_fill_2 FILLER_72_166 ();
 sg13g2_fill_1 FILLER_72_168 ();
 sg13g2_decap_4 FILLER_72_172 ();
 sg13g2_fill_2 FILLER_72_176 ();
 sg13g2_fill_2 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_183 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_253 ();
 sg13g2_fill_2 FILLER_72_270 ();
 sg13g2_fill_1 FILLER_72_277 ();
 sg13g2_decap_4 FILLER_72_283 ();
 sg13g2_fill_1 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_354 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_366 ();
 sg13g2_fill_1 FILLER_72_398 ();
 sg13g2_fill_1 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_452 ();
 sg13g2_fill_1 FILLER_72_483 ();
 sg13g2_fill_1 FILLER_72_510 ();
 sg13g2_fill_2 FILLER_72_537 ();
 sg13g2_fill_1 FILLER_72_565 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_fill_2 FILLER_72_582 ();
 sg13g2_fill_1 FILLER_72_597 ();
 sg13g2_fill_2 FILLER_72_608 ();
 sg13g2_fill_1 FILLER_72_620 ();
 sg13g2_fill_1 FILLER_72_640 ();
 sg13g2_fill_1 FILLER_72_645 ();
 sg13g2_fill_1 FILLER_72_658 ();
 sg13g2_fill_1 FILLER_72_667 ();
 sg13g2_fill_2 FILLER_72_677 ();
 sg13g2_fill_1 FILLER_72_687 ();
 sg13g2_fill_1 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_719 ();
 sg13g2_fill_2 FILLER_72_726 ();
 sg13g2_fill_1 FILLER_72_728 ();
 sg13g2_fill_1 FILLER_72_795 ();
 sg13g2_decap_8 FILLER_72_827 ();
 sg13g2_fill_1 FILLER_72_834 ();
 sg13g2_fill_2 FILLER_72_839 ();
 sg13g2_fill_1 FILLER_72_841 ();
 sg13g2_decap_4 FILLER_72_879 ();
 sg13g2_fill_2 FILLER_72_883 ();
 sg13g2_fill_1 FILLER_72_922 ();
 sg13g2_fill_1 FILLER_72_927 ();
 sg13g2_fill_1 FILLER_72_933 ();
 sg13g2_fill_1 FILLER_72_938 ();
 sg13g2_decap_8 FILLER_72_958 ();
 sg13g2_decap_4 FILLER_72_965 ();
 sg13g2_fill_2 FILLER_72_969 ();
 sg13g2_fill_1 FILLER_72_976 ();
 sg13g2_decap_8 FILLER_72_981 ();
 sg13g2_fill_2 FILLER_72_991 ();
 sg13g2_fill_1 FILLER_72_993 ();
 sg13g2_decap_4 FILLER_72_1025 ();
 sg13g2_fill_1 FILLER_72_1029 ();
 sg13g2_decap_8 FILLER_72_1076 ();
 sg13g2_decap_8 FILLER_72_1083 ();
 sg13g2_fill_2 FILLER_72_1099 ();
 sg13g2_fill_1 FILLER_72_1101 ();
 sg13g2_fill_2 FILLER_72_1128 ();
 sg13g2_fill_2 FILLER_72_1160 ();
 sg13g2_fill_2 FILLER_72_1188 ();
 sg13g2_fill_1 FILLER_72_1190 ();
 sg13g2_fill_2 FILLER_72_1195 ();
 sg13g2_fill_1 FILLER_72_1197 ();
 sg13g2_fill_2 FILLER_72_1224 ();
 sg13g2_fill_1 FILLER_72_1226 ();
 sg13g2_fill_1 FILLER_72_1242 ();
 sg13g2_fill_2 FILLER_72_1267 ();
 sg13g2_decap_4 FILLER_72_1295 ();
 sg13g2_fill_2 FILLER_72_1303 ();
 sg13g2_decap_8 FILLER_72_1313 ();
 sg13g2_decap_4 FILLER_72_1320 ();
 sg13g2_fill_1 FILLER_72_1324 ();
 sg13g2_decap_4 FILLER_72_1329 ();
 sg13g2_fill_2 FILLER_72_1333 ();
 sg13g2_decap_8 FILLER_72_1339 ();
 sg13g2_decap_8 FILLER_72_1346 ();
 sg13g2_decap_8 FILLER_72_1353 ();
 sg13g2_fill_2 FILLER_72_1374 ();
 sg13g2_fill_1 FILLER_72_1376 ();
 sg13g2_decap_4 FILLER_72_1381 ();
 sg13g2_fill_1 FILLER_72_1388 ();
 sg13g2_decap_8 FILLER_72_1393 ();
 sg13g2_fill_2 FILLER_72_1405 ();
 sg13g2_fill_1 FILLER_72_1420 ();
 sg13g2_fill_2 FILLER_72_1426 ();
 sg13g2_fill_2 FILLER_72_1447 ();
 sg13g2_fill_1 FILLER_72_1449 ();
 sg13g2_fill_2 FILLER_72_1459 ();
 sg13g2_fill_2 FILLER_72_1464 ();
 sg13g2_fill_2 FILLER_72_1479 ();
 sg13g2_decap_8 FILLER_72_1485 ();
 sg13g2_fill_2 FILLER_72_1492 ();
 sg13g2_fill_1 FILLER_72_1499 ();
 sg13g2_fill_1 FILLER_72_1572 ();
 sg13g2_decap_4 FILLER_72_1580 ();
 sg13g2_fill_2 FILLER_72_1593 ();
 sg13g2_fill_1 FILLER_72_1601 ();
 sg13g2_fill_2 FILLER_72_1661 ();
 sg13g2_fill_1 FILLER_72_1663 ();
 sg13g2_decap_4 FILLER_72_1672 ();
 sg13g2_fill_1 FILLER_72_1681 ();
 sg13g2_fill_1 FILLER_72_1709 ();
 sg13g2_decap_4 FILLER_72_1724 ();
 sg13g2_fill_2 FILLER_72_1728 ();
 sg13g2_fill_1 FILLER_72_1735 ();
 sg13g2_decap_8 FILLER_72_1746 ();
 sg13g2_fill_2 FILLER_72_1753 ();
 sg13g2_fill_1 FILLER_72_1755 ();
 sg13g2_fill_2 FILLER_72_1793 ();
 sg13g2_decap_4 FILLER_72_1809 ();
 sg13g2_fill_2 FILLER_72_1813 ();
 sg13g2_fill_1 FILLER_72_1833 ();
 sg13g2_decap_8 FILLER_72_1849 ();
 sg13g2_decap_8 FILLER_72_1856 ();
 sg13g2_fill_2 FILLER_72_1880 ();
 sg13g2_decap_4 FILLER_72_1889 ();
 sg13g2_fill_1 FILLER_72_1897 ();
 sg13g2_decap_4 FILLER_72_1904 ();
 sg13g2_fill_1 FILLER_72_1930 ();
 sg13g2_decap_8 FILLER_72_1978 ();
 sg13g2_fill_2 FILLER_72_1985 ();
 sg13g2_fill_1 FILLER_72_1987 ();
 sg13g2_fill_2 FILLER_72_2040 ();
 sg13g2_decap_4 FILLER_72_2097 ();
 sg13g2_fill_2 FILLER_72_2101 ();
 sg13g2_fill_2 FILLER_72_2126 ();
 sg13g2_fill_1 FILLER_72_2128 ();
 sg13g2_fill_2 FILLER_72_2175 ();
 sg13g2_decap_8 FILLER_72_2239 ();
 sg13g2_decap_8 FILLER_72_2281 ();
 sg13g2_decap_8 FILLER_72_2288 ();
 sg13g2_fill_2 FILLER_72_2295 ();
 sg13g2_decap_8 FILLER_72_2301 ();
 sg13g2_decap_4 FILLER_72_2308 ();
 sg13g2_fill_1 FILLER_72_2312 ();
 sg13g2_decap_4 FILLER_72_2321 ();
 sg13g2_fill_2 FILLER_72_2325 ();
 sg13g2_decap_8 FILLER_72_2338 ();
 sg13g2_decap_8 FILLER_72_2345 ();
 sg13g2_fill_2 FILLER_72_2352 ();
 sg13g2_fill_1 FILLER_72_2362 ();
 sg13g2_fill_1 FILLER_72_2368 ();
 sg13g2_fill_2 FILLER_72_2377 ();
 sg13g2_decap_8 FILLER_72_2383 ();
 sg13g2_decap_8 FILLER_72_2390 ();
 sg13g2_fill_1 FILLER_72_2397 ();
 sg13g2_decap_4 FILLER_72_2415 ();
 sg13g2_decap_4 FILLER_72_2537 ();
 sg13g2_fill_1 FILLER_72_2551 ();
 sg13g2_fill_1 FILLER_72_2556 ();
 sg13g2_fill_2 FILLER_72_2567 ();
 sg13g2_fill_2 FILLER_72_2624 ();
 sg13g2_fill_2 FILLER_72_2635 ();
 sg13g2_fill_2 FILLER_72_2643 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_fill_2 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_23 ();
 sg13g2_fill_1 FILLER_73_28 ();
 sg13g2_fill_2 FILLER_73_49 ();
 sg13g2_fill_1 FILLER_73_51 ();
 sg13g2_fill_2 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_58 ();
 sg13g2_decap_4 FILLER_73_80 ();
 sg13g2_decap_8 FILLER_73_89 ();
 sg13g2_decap_8 FILLER_73_96 ();
 sg13g2_decap_8 FILLER_73_103 ();
 sg13g2_decap_4 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_118 ();
 sg13g2_decap_8 FILLER_73_125 ();
 sg13g2_fill_1 FILLER_73_132 ();
 sg13g2_decap_4 FILLER_73_143 ();
 sg13g2_fill_1 FILLER_73_147 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_179 ();
 sg13g2_decap_4 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_190 ();
 sg13g2_fill_1 FILLER_73_208 ();
 sg13g2_decap_4 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_238 ();
 sg13g2_fill_2 FILLER_73_259 ();
 sg13g2_fill_1 FILLER_73_266 ();
 sg13g2_fill_1 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_311 ();
 sg13g2_decap_4 FILLER_73_318 ();
 sg13g2_decap_8 FILLER_73_332 ();
 sg13g2_decap_8 FILLER_73_339 ();
 sg13g2_decap_4 FILLER_73_346 ();
 sg13g2_fill_2 FILLER_73_350 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_388 ();
 sg13g2_fill_2 FILLER_73_416 ();
 sg13g2_decap_4 FILLER_73_423 ();
 sg13g2_fill_2 FILLER_73_471 ();
 sg13g2_fill_1 FILLER_73_473 ();
 sg13g2_decap_4 FILLER_73_498 ();
 sg13g2_fill_2 FILLER_73_512 ();
 sg13g2_fill_2 FILLER_73_518 ();
 sg13g2_fill_1 FILLER_73_520 ();
 sg13g2_decap_8 FILLER_73_525 ();
 sg13g2_decap_4 FILLER_73_532 ();
 sg13g2_fill_2 FILLER_73_536 ();
 sg13g2_fill_1 FILLER_73_560 ();
 sg13g2_fill_2 FILLER_73_565 ();
 sg13g2_fill_1 FILLER_73_567 ();
 sg13g2_fill_2 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_648 ();
 sg13g2_decap_8 FILLER_73_655 ();
 sg13g2_fill_2 FILLER_73_662 ();
 sg13g2_fill_1 FILLER_73_664 ();
 sg13g2_decap_4 FILLER_73_668 ();
 sg13g2_fill_1 FILLER_73_672 ();
 sg13g2_fill_2 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_694 ();
 sg13g2_decap_8 FILLER_73_721 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_8 FILLER_73_742 ();
 sg13g2_decap_4 FILLER_73_749 ();
 sg13g2_fill_1 FILLER_73_753 ();
 sg13g2_fill_2 FILLER_73_757 ();
 sg13g2_decap_4 FILLER_73_763 ();
 sg13g2_fill_2 FILLER_73_777 ();
 sg13g2_fill_2 FILLER_73_783 ();
 sg13g2_fill_1 FILLER_73_785 ();
 sg13g2_fill_1 FILLER_73_789 ();
 sg13g2_decap_8 FILLER_73_832 ();
 sg13g2_fill_2 FILLER_73_839 ();
 sg13g2_fill_1 FILLER_73_841 ();
 sg13g2_decap_4 FILLER_73_852 ();
 sg13g2_fill_2 FILLER_73_856 ();
 sg13g2_decap_8 FILLER_73_890 ();
 sg13g2_decap_8 FILLER_73_897 ();
 sg13g2_decap_8 FILLER_73_904 ();
 sg13g2_decap_8 FILLER_73_911 ();
 sg13g2_decap_8 FILLER_73_918 ();
 sg13g2_decap_4 FILLER_73_925 ();
 sg13g2_decap_4 FILLER_73_959 ();
 sg13g2_fill_1 FILLER_73_963 ();
 sg13g2_fill_1 FILLER_73_967 ();
 sg13g2_fill_1 FILLER_73_984 ();
 sg13g2_decap_4 FILLER_73_989 ();
 sg13g2_fill_2 FILLER_73_998 ();
 sg13g2_fill_1 FILLER_73_1000 ();
 sg13g2_fill_1 FILLER_73_1005 ();
 sg13g2_fill_2 FILLER_73_1041 ();
 sg13g2_decap_8 FILLER_73_1047 ();
 sg13g2_decap_4 FILLER_73_1054 ();
 sg13g2_fill_1 FILLER_73_1058 ();
 sg13g2_decap_8 FILLER_73_1063 ();
 sg13g2_decap_8 FILLER_73_1070 ();
 sg13g2_fill_1 FILLER_73_1077 ();
 sg13g2_decap_4 FILLER_73_1135 ();
 sg13g2_fill_1 FILLER_73_1143 ();
 sg13g2_fill_1 FILLER_73_1148 ();
 sg13g2_fill_2 FILLER_73_1154 ();
 sg13g2_decap_4 FILLER_73_1160 ();
 sg13g2_fill_2 FILLER_73_1164 ();
 sg13g2_decap_4 FILLER_73_1187 ();
 sg13g2_fill_2 FILLER_73_1191 ();
 sg13g2_fill_2 FILLER_73_1201 ();
 sg13g2_fill_1 FILLER_73_1203 ();
 sg13g2_decap_8 FILLER_73_1208 ();
 sg13g2_decap_8 FILLER_73_1215 ();
 sg13g2_fill_2 FILLER_73_1222 ();
 sg13g2_fill_1 FILLER_73_1224 ();
 sg13g2_fill_1 FILLER_73_1230 ();
 sg13g2_fill_1 FILLER_73_1245 ();
 sg13g2_fill_1 FILLER_73_1260 ();
 sg13g2_fill_2 FILLER_73_1268 ();
 sg13g2_fill_2 FILLER_73_1288 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_fill_2 FILLER_73_1305 ();
 sg13g2_decap_8 FILLER_73_1318 ();
 sg13g2_fill_2 FILLER_73_1344 ();
 sg13g2_fill_1 FILLER_73_1346 ();
 sg13g2_decap_8 FILLER_73_1353 ();
 sg13g2_fill_2 FILLER_73_1360 ();
 sg13g2_decap_8 FILLER_73_1367 ();
 sg13g2_decap_4 FILLER_73_1374 ();
 sg13g2_decap_4 FILLER_73_1386 ();
 sg13g2_fill_1 FILLER_73_1390 ();
 sg13g2_fill_1 FILLER_73_1396 ();
 sg13g2_fill_1 FILLER_73_1420 ();
 sg13g2_fill_1 FILLER_73_1425 ();
 sg13g2_fill_1 FILLER_73_1432 ();
 sg13g2_fill_1 FILLER_73_1452 ();
 sg13g2_fill_1 FILLER_73_1485 ();
 sg13g2_fill_2 FILLER_73_1493 ();
 sg13g2_fill_1 FILLER_73_1495 ();
 sg13g2_fill_1 FILLER_73_1510 ();
 sg13g2_decap_8 FILLER_73_1518 ();
 sg13g2_fill_2 FILLER_73_1525 ();
 sg13g2_fill_1 FILLER_73_1532 ();
 sg13g2_fill_1 FILLER_73_1540 ();
 sg13g2_decap_4 FILLER_73_1560 ();
 sg13g2_fill_1 FILLER_73_1564 ();
 sg13g2_decap_8 FILLER_73_1584 ();
 sg13g2_decap_8 FILLER_73_1591 ();
 sg13g2_fill_2 FILLER_73_1598 ();
 sg13g2_fill_1 FILLER_73_1600 ();
 sg13g2_decap_4 FILLER_73_1631 ();
 sg13g2_decap_8 FILLER_73_1665 ();
 sg13g2_fill_1 FILLER_73_1676 ();
 sg13g2_fill_1 FILLER_73_1701 ();
 sg13g2_fill_1 FILLER_73_1705 ();
 sg13g2_fill_1 FILLER_73_1710 ();
 sg13g2_fill_1 FILLER_73_1731 ();
 sg13g2_decap_8 FILLER_73_1737 ();
 sg13g2_fill_2 FILLER_73_1744 ();
 sg13g2_decap_8 FILLER_73_1751 ();
 sg13g2_decap_4 FILLER_73_1758 ();
 sg13g2_fill_1 FILLER_73_1762 ();
 sg13g2_decap_4 FILLER_73_1778 ();
 sg13g2_fill_2 FILLER_73_1782 ();
 sg13g2_fill_1 FILLER_73_1797 ();
 sg13g2_decap_8 FILLER_73_1802 ();
 sg13g2_decap_8 FILLER_73_1809 ();
 sg13g2_decap_8 FILLER_73_1816 ();
 sg13g2_decap_8 FILLER_73_1823 ();
 sg13g2_decap_4 FILLER_73_1848 ();
 sg13g2_fill_2 FILLER_73_1888 ();
 sg13g2_decap_4 FILLER_73_1895 ();
 sg13g2_fill_1 FILLER_73_1899 ();
 sg13g2_fill_2 FILLER_73_1915 ();
 sg13g2_fill_1 FILLER_73_1917 ();
 sg13g2_fill_1 FILLER_73_1924 ();
 sg13g2_fill_2 FILLER_73_1929 ();
 sg13g2_fill_1 FILLER_73_1931 ();
 sg13g2_fill_1 FILLER_73_1969 ();
 sg13g2_decap_8 FILLER_73_1974 ();
 sg13g2_decap_8 FILLER_73_1981 ();
 sg13g2_fill_1 FILLER_73_2014 ();
 sg13g2_decap_8 FILLER_73_2040 ();
 sg13g2_decap_4 FILLER_73_2047 ();
 sg13g2_decap_8 FILLER_73_2090 ();
 sg13g2_decap_4 FILLER_73_2097 ();
 sg13g2_fill_2 FILLER_73_2101 ();
 sg13g2_fill_1 FILLER_73_2139 ();
 sg13g2_decap_8 FILLER_73_2149 ();
 sg13g2_decap_8 FILLER_73_2156 ();
 sg13g2_decap_4 FILLER_73_2214 ();
 sg13g2_fill_2 FILLER_73_2218 ();
 sg13g2_decap_4 FILLER_73_2224 ();
 sg13g2_decap_4 FILLER_73_2304 ();
 sg13g2_decap_8 FILLER_73_2313 ();
 sg13g2_fill_1 FILLER_73_2320 ();
 sg13g2_fill_1 FILLER_73_2329 ();
 sg13g2_decap_8 FILLER_73_2335 ();
 sg13g2_fill_1 FILLER_73_2346 ();
 sg13g2_decap_8 FILLER_73_2366 ();
 sg13g2_decap_8 FILLER_73_2373 ();
 sg13g2_fill_2 FILLER_73_2380 ();
 sg13g2_fill_1 FILLER_73_2382 ();
 sg13g2_fill_1 FILLER_73_2387 ();
 sg13g2_decap_4 FILLER_73_2418 ();
 sg13g2_fill_1 FILLER_73_2510 ();
 sg13g2_fill_1 FILLER_73_2516 ();
 sg13g2_fill_1 FILLER_73_2547 ();
 sg13g2_decap_8 FILLER_73_2554 ();
 sg13g2_decap_8 FILLER_73_2561 ();
 sg13g2_decap_8 FILLER_73_2663 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_4 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_44 ();
 sg13g2_fill_2 FILLER_74_51 ();
 sg13g2_fill_1 FILLER_74_53 ();
 sg13g2_decap_4 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_79 ();
 sg13g2_decap_4 FILLER_74_109 ();
 sg13g2_decap_8 FILLER_74_134 ();
 sg13g2_fill_1 FILLER_74_177 ();
 sg13g2_fill_2 FILLER_74_187 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_223 ();
 sg13g2_fill_2 FILLER_74_235 ();
 sg13g2_fill_1 FILLER_74_242 ();
 sg13g2_fill_1 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_252 ();
 sg13g2_fill_2 FILLER_74_263 ();
 sg13g2_fill_2 FILLER_74_305 ();
 sg13g2_decap_8 FILLER_74_313 ();
 sg13g2_decap_4 FILLER_74_320 ();
 sg13g2_fill_1 FILLER_74_324 ();
 sg13g2_decap_4 FILLER_74_350 ();
 sg13g2_fill_2 FILLER_74_354 ();
 sg13g2_fill_1 FILLER_74_360 ();
 sg13g2_fill_2 FILLER_74_378 ();
 sg13g2_fill_1 FILLER_74_380 ();
 sg13g2_decap_8 FILLER_74_394 ();
 sg13g2_fill_2 FILLER_74_401 ();
 sg13g2_fill_1 FILLER_74_403 ();
 sg13g2_decap_8 FILLER_74_430 ();
 sg13g2_decap_8 FILLER_74_437 ();
 sg13g2_fill_2 FILLER_74_444 ();
 sg13g2_fill_1 FILLER_74_446 ();
 sg13g2_fill_1 FILLER_74_458 ();
 sg13g2_decap_4 FILLER_74_468 ();
 sg13g2_fill_1 FILLER_74_472 ();
 sg13g2_decap_8 FILLER_74_478 ();
 sg13g2_fill_1 FILLER_74_485 ();
 sg13g2_decap_8 FILLER_74_505 ();
 sg13g2_decap_8 FILLER_74_512 ();
 sg13g2_decap_8 FILLER_74_519 ();
 sg13g2_decap_8 FILLER_74_526 ();
 sg13g2_decap_8 FILLER_74_533 ();
 sg13g2_fill_2 FILLER_74_540 ();
 sg13g2_decap_8 FILLER_74_576 ();
 sg13g2_fill_1 FILLER_74_583 ();
 sg13g2_fill_1 FILLER_74_603 ();
 sg13g2_decap_8 FILLER_74_626 ();
 sg13g2_decap_4 FILLER_74_633 ();
 sg13g2_fill_1 FILLER_74_637 ();
 sg13g2_fill_1 FILLER_74_647 ();
 sg13g2_fill_1 FILLER_74_656 ();
 sg13g2_fill_1 FILLER_74_671 ();
 sg13g2_fill_2 FILLER_74_705 ();
 sg13g2_decap_4 FILLER_74_711 ();
 sg13g2_fill_2 FILLER_74_715 ();
 sg13g2_fill_2 FILLER_74_791 ();
 sg13g2_fill_1 FILLER_74_793 ();
 sg13g2_fill_1 FILLER_74_800 ();
 sg13g2_decap_4 FILLER_74_815 ();
 sg13g2_fill_2 FILLER_74_819 ();
 sg13g2_fill_2 FILLER_74_908 ();
 sg13g2_decap_8 FILLER_74_921 ();
 sg13g2_decap_8 FILLER_74_928 ();
 sg13g2_decap_8 FILLER_74_945 ();
 sg13g2_fill_2 FILLER_74_952 ();
 sg13g2_fill_1 FILLER_74_954 ();
 sg13g2_fill_2 FILLER_74_972 ();
 sg13g2_fill_2 FILLER_74_1026 ();
 sg13g2_fill_1 FILLER_74_1028 ();
 sg13g2_decap_8 FILLER_74_1055 ();
 sg13g2_decap_8 FILLER_74_1062 ();
 sg13g2_decap_8 FILLER_74_1069 ();
 sg13g2_fill_1 FILLER_74_1127 ();
 sg13g2_decap_8 FILLER_74_1137 ();
 sg13g2_decap_8 FILLER_74_1144 ();
 sg13g2_decap_8 FILLER_74_1151 ();
 sg13g2_fill_1 FILLER_74_1158 ();
 sg13g2_decap_8 FILLER_74_1164 ();
 sg13g2_fill_2 FILLER_74_1171 ();
 sg13g2_fill_1 FILLER_74_1173 ();
 sg13g2_fill_2 FILLER_74_1203 ();
 sg13g2_fill_1 FILLER_74_1205 ();
 sg13g2_decap_8 FILLER_74_1214 ();
 sg13g2_fill_1 FILLER_74_1221 ();
 sg13g2_fill_1 FILLER_74_1243 ();
 sg13g2_fill_1 FILLER_74_1258 ();
 sg13g2_decap_8 FILLER_74_1281 ();
 sg13g2_fill_2 FILLER_74_1288 ();
 sg13g2_fill_1 FILLER_74_1295 ();
 sg13g2_fill_2 FILLER_74_1305 ();
 sg13g2_decap_4 FILLER_74_1316 ();
 sg13g2_decap_8 FILLER_74_1324 ();
 sg13g2_decap_4 FILLER_74_1331 ();
 sg13g2_fill_1 FILLER_74_1335 ();
 sg13g2_decap_4 FILLER_74_1343 ();
 sg13g2_fill_2 FILLER_74_1347 ();
 sg13g2_decap_8 FILLER_74_1354 ();
 sg13g2_decap_8 FILLER_74_1361 ();
 sg13g2_decap_4 FILLER_74_1368 ();
 sg13g2_fill_2 FILLER_74_1372 ();
 sg13g2_fill_2 FILLER_74_1383 ();
 sg13g2_decap_4 FILLER_74_1392 ();
 sg13g2_fill_2 FILLER_74_1396 ();
 sg13g2_fill_2 FILLER_74_1416 ();
 sg13g2_decap_8 FILLER_74_1424 ();
 sg13g2_fill_2 FILLER_74_1436 ();
 sg13g2_fill_1 FILLER_74_1441 ();
 sg13g2_fill_1 FILLER_74_1469 ();
 sg13g2_decap_8 FILLER_74_1489 ();
 sg13g2_fill_2 FILLER_74_1496 ();
 sg13g2_decap_8 FILLER_74_1518 ();
 sg13g2_fill_1 FILLER_74_1525 ();
 sg13g2_fill_2 FILLER_74_1531 ();
 sg13g2_fill_2 FILLER_74_1566 ();
 sg13g2_fill_2 FILLER_74_1590 ();
 sg13g2_fill_1 FILLER_74_1592 ();
 sg13g2_decap_8 FILLER_74_1598 ();
 sg13g2_decap_4 FILLER_74_1605 ();
 sg13g2_fill_2 FILLER_74_1622 ();
 sg13g2_fill_1 FILLER_74_1624 ();
 sg13g2_decap_8 FILLER_74_1629 ();
 sg13g2_decap_8 FILLER_74_1636 ();
 sg13g2_fill_2 FILLER_74_1643 ();
 sg13g2_fill_2 FILLER_74_1658 ();
 sg13g2_fill_1 FILLER_74_1660 ();
 sg13g2_decap_4 FILLER_74_1665 ();
 sg13g2_fill_1 FILLER_74_1692 ();
 sg13g2_fill_1 FILLER_74_1696 ();
 sg13g2_decap_4 FILLER_74_1702 ();
 sg13g2_fill_2 FILLER_74_1710 ();
 sg13g2_fill_1 FILLER_74_1728 ();
 sg13g2_fill_1 FILLER_74_1737 ();
 sg13g2_fill_1 FILLER_74_1743 ();
 sg13g2_fill_2 FILLER_74_1748 ();
 sg13g2_decap_4 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1764 ();
 sg13g2_fill_1 FILLER_74_1766 ();
 sg13g2_decap_4 FILLER_74_1771 ();
 sg13g2_fill_2 FILLER_74_1775 ();
 sg13g2_decap_4 FILLER_74_1785 ();
 sg13g2_decap_8 FILLER_74_1794 ();
 sg13g2_decap_8 FILLER_74_1801 ();
 sg13g2_decap_4 FILLER_74_1808 ();
 sg13g2_fill_1 FILLER_74_1812 ();
 sg13g2_decap_4 FILLER_74_1818 ();
 sg13g2_fill_1 FILLER_74_1822 ();
 sg13g2_decap_4 FILLER_74_1827 ();
 sg13g2_decap_4 FILLER_74_1834 ();
 sg13g2_decap_4 FILLER_74_1842 ();
 sg13g2_decap_8 FILLER_74_1856 ();
 sg13g2_fill_1 FILLER_74_1881 ();
 sg13g2_fill_2 FILLER_74_1888 ();
 sg13g2_fill_1 FILLER_74_1902 ();
 sg13g2_fill_1 FILLER_74_1911 ();
 sg13g2_fill_2 FILLER_74_1940 ();
 sg13g2_fill_2 FILLER_74_1946 ();
 sg13g2_fill_2 FILLER_74_1959 ();
 sg13g2_decap_8 FILLER_74_1971 ();
 sg13g2_decap_4 FILLER_74_1978 ();
 sg13g2_fill_1 FILLER_74_1982 ();
 sg13g2_decap_8 FILLER_74_2004 ();
 sg13g2_fill_2 FILLER_74_2011 ();
 sg13g2_fill_1 FILLER_74_2013 ();
 sg13g2_decap_4 FILLER_74_2054 ();
 sg13g2_fill_1 FILLER_74_2068 ();
 sg13g2_decap_8 FILLER_74_2105 ();
 sg13g2_decap_4 FILLER_74_2112 ();
 sg13g2_fill_1 FILLER_74_2116 ();
 sg13g2_decap_4 FILLER_74_2125 ();
 sg13g2_fill_2 FILLER_74_2129 ();
 sg13g2_decap_8 FILLER_74_2135 ();
 sg13g2_decap_8 FILLER_74_2142 ();
 sg13g2_decap_8 FILLER_74_2149 ();
 sg13g2_decap_4 FILLER_74_2156 ();
 sg13g2_fill_1 FILLER_74_2160 ();
 sg13g2_decap_8 FILLER_74_2171 ();
 sg13g2_decap_8 FILLER_74_2178 ();
 sg13g2_decap_8 FILLER_74_2185 ();
 sg13g2_decap_4 FILLER_74_2192 ();
 sg13g2_decap_8 FILLER_74_2200 ();
 sg13g2_fill_2 FILLER_74_2207 ();
 sg13g2_fill_1 FILLER_74_2209 ();
 sg13g2_decap_8 FILLER_74_2214 ();
 sg13g2_decap_8 FILLER_74_2221 ();
 sg13g2_fill_2 FILLER_74_2228 ();
 sg13g2_fill_1 FILLER_74_2230 ();
 sg13g2_fill_1 FILLER_74_2297 ();
 sg13g2_fill_1 FILLER_74_2302 ();
 sg13g2_fill_1 FILLER_74_2313 ();
 sg13g2_fill_2 FILLER_74_2319 ();
 sg13g2_fill_1 FILLER_74_2321 ();
 sg13g2_decap_4 FILLER_74_2327 ();
 sg13g2_fill_1 FILLER_74_2331 ();
 sg13g2_fill_2 FILLER_74_2337 ();
 sg13g2_fill_1 FILLER_74_2339 ();
 sg13g2_fill_2 FILLER_74_2357 ();
 sg13g2_fill_1 FILLER_74_2359 ();
 sg13g2_decap_8 FILLER_74_2369 ();
 sg13g2_fill_2 FILLER_74_2376 ();
 sg13g2_fill_1 FILLER_74_2378 ();
 sg13g2_decap_8 FILLER_74_2416 ();
 sg13g2_decap_8 FILLER_74_2438 ();
 sg13g2_decap_8 FILLER_74_2445 ();
 sg13g2_decap_4 FILLER_74_2452 ();
 sg13g2_fill_1 FILLER_74_2480 ();
 sg13g2_fill_1 FILLER_74_2486 ();
 sg13g2_fill_1 FILLER_74_2491 ();
 sg13g2_fill_1 FILLER_74_2496 ();
 sg13g2_decap_8 FILLER_74_2501 ();
 sg13g2_decap_8 FILLER_74_2508 ();
 sg13g2_fill_2 FILLER_74_2515 ();
 sg13g2_decap_8 FILLER_74_2560 ();
 sg13g2_fill_2 FILLER_74_2567 ();
 sg13g2_fill_1 FILLER_74_2569 ();
 sg13g2_fill_1 FILLER_74_2576 ();
 sg13g2_decap_8 FILLER_74_2617 ();
 sg13g2_fill_2 FILLER_74_2634 ();
 sg13g2_fill_2 FILLER_74_2646 ();
 sg13g2_decap_8 FILLER_74_2652 ();
 sg13g2_decap_8 FILLER_74_2659 ();
 sg13g2_decap_4 FILLER_74_2666 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_4 ();
 sg13g2_fill_2 FILLER_75_41 ();
 sg13g2_fill_1 FILLER_75_43 ();
 sg13g2_decap_4 FILLER_75_54 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_decap_4 FILLER_75_73 ();
 sg13g2_fill_2 FILLER_75_103 ();
 sg13g2_decap_4 FILLER_75_110 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_200 ();
 sg13g2_fill_1 FILLER_75_202 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_decap_8 FILLER_75_220 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_4 FILLER_75_238 ();
 sg13g2_fill_1 FILLER_75_242 ();
 sg13g2_decap_4 FILLER_75_246 ();
 sg13g2_fill_2 FILLER_75_250 ();
 sg13g2_fill_1 FILLER_75_277 ();
 sg13g2_fill_1 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_289 ();
 sg13g2_fill_2 FILLER_75_293 ();
 sg13g2_decap_4 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_325 ();
 sg13g2_fill_1 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_340 ();
 sg13g2_decap_8 FILLER_75_347 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_391 ();
 sg13g2_decap_8 FILLER_75_398 ();
 sg13g2_decap_4 FILLER_75_405 ();
 sg13g2_fill_1 FILLER_75_409 ();
 sg13g2_decap_8 FILLER_75_414 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_8 FILLER_75_428 ();
 sg13g2_fill_2 FILLER_75_454 ();
 sg13g2_fill_2 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_471 ();
 sg13g2_fill_2 FILLER_75_492 ();
 sg13g2_fill_1 FILLER_75_494 ();
 sg13g2_fill_2 FILLER_75_535 ();
 sg13g2_fill_1 FILLER_75_537 ();
 sg13g2_fill_1 FILLER_75_570 ();
 sg13g2_fill_2 FILLER_75_585 ();
 sg13g2_fill_2 FILLER_75_592 ();
 sg13g2_decap_4 FILLER_75_598 ();
 sg13g2_decap_4 FILLER_75_609 ();
 sg13g2_fill_1 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_618 ();
 sg13g2_decap_8 FILLER_75_625 ();
 sg13g2_fill_2 FILLER_75_632 ();
 sg13g2_fill_1 FILLER_75_634 ();
 sg13g2_fill_2 FILLER_75_644 ();
 sg13g2_fill_1 FILLER_75_646 ();
 sg13g2_fill_2 FILLER_75_655 ();
 sg13g2_fill_1 FILLER_75_657 ();
 sg13g2_fill_2 FILLER_75_685 ();
 sg13g2_decap_8 FILLER_75_713 ();
 sg13g2_decap_4 FILLER_75_720 ();
 sg13g2_fill_2 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_fill_1 FILLER_75_768 ();
 sg13g2_fill_2 FILLER_75_785 ();
 sg13g2_fill_1 FILLER_75_793 ();
 sg13g2_fill_2 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_fill_2 FILLER_75_824 ();
 sg13g2_fill_1 FILLER_75_826 ();
 sg13g2_decap_4 FILLER_75_837 ();
 sg13g2_decap_4 FILLER_75_845 ();
 sg13g2_fill_1 FILLER_75_849 ();
 sg13g2_decap_8 FILLER_75_860 ();
 sg13g2_fill_2 FILLER_75_867 ();
 sg13g2_fill_1 FILLER_75_869 ();
 sg13g2_fill_2 FILLER_75_874 ();
 sg13g2_fill_1 FILLER_75_888 ();
 sg13g2_decap_4 FILLER_75_931 ();
 sg13g2_decap_4 FILLER_75_975 ();
 sg13g2_fill_2 FILLER_75_979 ();
 sg13g2_decap_8 FILLER_75_993 ();
 sg13g2_decap_8 FILLER_75_1000 ();
 sg13g2_fill_2 FILLER_75_1007 ();
 sg13g2_decap_4 FILLER_75_1035 ();
 sg13g2_fill_1 FILLER_75_1039 ();
 sg13g2_decap_8 FILLER_75_1050 ();
 sg13g2_fill_2 FILLER_75_1057 ();
 sg13g2_decap_8 FILLER_75_1063 ();
 sg13g2_decap_8 FILLER_75_1070 ();
 sg13g2_decap_8 FILLER_75_1077 ();
 sg13g2_decap_4 FILLER_75_1088 ();
 sg13g2_fill_2 FILLER_75_1092 ();
 sg13g2_fill_1 FILLER_75_1098 ();
 sg13g2_fill_2 FILLER_75_1134 ();
 sg13g2_fill_2 FILLER_75_1167 ();
 sg13g2_fill_1 FILLER_75_1173 ();
 sg13g2_fill_1 FILLER_75_1187 ();
 sg13g2_decap_4 FILLER_75_1219 ();
 sg13g2_fill_2 FILLER_75_1223 ();
 sg13g2_fill_1 FILLER_75_1233 ();
 sg13g2_fill_1 FILLER_75_1238 ();
 sg13g2_fill_1 FILLER_75_1249 ();
 sg13g2_decap_4 FILLER_75_1255 ();
 sg13g2_fill_2 FILLER_75_1259 ();
 sg13g2_decap_4 FILLER_75_1267 ();
 sg13g2_fill_1 FILLER_75_1271 ();
 sg13g2_fill_1 FILLER_75_1290 ();
 sg13g2_decap_8 FILLER_75_1304 ();
 sg13g2_fill_2 FILLER_75_1316 ();
 sg13g2_decap_8 FILLER_75_1323 ();
 sg13g2_decap_8 FILLER_75_1330 ();
 sg13g2_decap_8 FILLER_75_1337 ();
 sg13g2_decap_8 FILLER_75_1344 ();
 sg13g2_fill_1 FILLER_75_1351 ();
 sg13g2_fill_2 FILLER_75_1361 ();
 sg13g2_fill_1 FILLER_75_1363 ();
 sg13g2_decap_4 FILLER_75_1377 ();
 sg13g2_fill_1 FILLER_75_1381 ();
 sg13g2_decap_8 FILLER_75_1394 ();
 sg13g2_decap_8 FILLER_75_1401 ();
 sg13g2_decap_4 FILLER_75_1408 ();
 sg13g2_fill_2 FILLER_75_1428 ();
 sg13g2_decap_8 FILLER_75_1440 ();
 sg13g2_fill_1 FILLER_75_1447 ();
 sg13g2_fill_1 FILLER_75_1477 ();
 sg13g2_fill_2 FILLER_75_1496 ();
 sg13g2_fill_1 FILLER_75_1498 ();
 sg13g2_fill_2 FILLER_75_1515 ();
 sg13g2_decap_4 FILLER_75_1526 ();
 sg13g2_fill_2 FILLER_75_1530 ();
 sg13g2_decap_4 FILLER_75_1541 ();
 sg13g2_fill_2 FILLER_75_1545 ();
 sg13g2_fill_1 FILLER_75_1552 ();
 sg13g2_fill_1 FILLER_75_1559 ();
 sg13g2_fill_1 FILLER_75_1565 ();
 sg13g2_fill_2 FILLER_75_1582 ();
 sg13g2_fill_2 FILLER_75_1589 ();
 sg13g2_fill_2 FILLER_75_1596 ();
 sg13g2_decap_8 FILLER_75_1606 ();
 sg13g2_decap_8 FILLER_75_1613 ();
 sg13g2_decap_8 FILLER_75_1620 ();
 sg13g2_fill_2 FILLER_75_1627 ();
 sg13g2_decap_8 FILLER_75_1633 ();
 sg13g2_decap_8 FILLER_75_1640 ();
 sg13g2_decap_4 FILLER_75_1647 ();
 sg13g2_fill_1 FILLER_75_1651 ();
 sg13g2_fill_1 FILLER_75_1665 ();
 sg13g2_decap_8 FILLER_75_1691 ();
 sg13g2_fill_1 FILLER_75_1698 ();
 sg13g2_fill_1 FILLER_75_1709 ();
 sg13g2_fill_1 FILLER_75_1726 ();
 sg13g2_fill_1 FILLER_75_1736 ();
 sg13g2_fill_2 FILLER_75_1755 ();
 sg13g2_decap_4 FILLER_75_1766 ();
 sg13g2_fill_2 FILLER_75_1790 ();
 sg13g2_decap_4 FILLER_75_1797 ();
 sg13g2_fill_1 FILLER_75_1801 ();
 sg13g2_decap_4 FILLER_75_1840 ();
 sg13g2_decap_4 FILLER_75_1849 ();
 sg13g2_fill_2 FILLER_75_1853 ();
 sg13g2_fill_2 FILLER_75_1859 ();
 sg13g2_fill_1 FILLER_75_1861 ();
 sg13g2_fill_2 FILLER_75_1867 ();
 sg13g2_fill_1 FILLER_75_1869 ();
 sg13g2_fill_2 FILLER_75_1873 ();
 sg13g2_fill_1 FILLER_75_1875 ();
 sg13g2_fill_2 FILLER_75_1881 ();
 sg13g2_fill_1 FILLER_75_1883 ();
 sg13g2_fill_1 FILLER_75_1897 ();
 sg13g2_decap_4 FILLER_75_1904 ();
 sg13g2_fill_2 FILLER_75_1908 ();
 sg13g2_decap_4 FILLER_75_1933 ();
 sg13g2_fill_2 FILLER_75_1947 ();
 sg13g2_decap_8 FILLER_75_1968 ();
 sg13g2_decap_8 FILLER_75_1975 ();
 sg13g2_decap_4 FILLER_75_1982 ();
 sg13g2_decap_8 FILLER_75_2022 ();
 sg13g2_fill_2 FILLER_75_2029 ();
 sg13g2_fill_1 FILLER_75_2031 ();
 sg13g2_fill_1 FILLER_75_2042 ();
 sg13g2_decap_8 FILLER_75_2053 ();
 sg13g2_decap_8 FILLER_75_2060 ();
 sg13g2_decap_4 FILLER_75_2067 ();
 sg13g2_fill_1 FILLER_75_2071 ();
 sg13g2_fill_2 FILLER_75_2089 ();
 sg13g2_fill_2 FILLER_75_2112 ();
 sg13g2_decap_8 FILLER_75_2150 ();
 sg13g2_fill_2 FILLER_75_2157 ();
 sg13g2_decap_4 FILLER_75_2172 ();
 sg13g2_fill_1 FILLER_75_2176 ();
 sg13g2_fill_2 FILLER_75_2211 ();
 sg13g2_fill_1 FILLER_75_2213 ();
 sg13g2_decap_4 FILLER_75_2235 ();
 sg13g2_fill_1 FILLER_75_2239 ();
 sg13g2_decap_8 FILLER_75_2244 ();
 sg13g2_decap_4 FILLER_75_2251 ();
 sg13g2_decap_8 FILLER_75_2282 ();
 sg13g2_fill_2 FILLER_75_2289 ();
 sg13g2_fill_1 FILLER_75_2317 ();
 sg13g2_fill_2 FILLER_75_2322 ();
 sg13g2_fill_1 FILLER_75_2324 ();
 sg13g2_fill_2 FILLER_75_2356 ();
 sg13g2_fill_1 FILLER_75_2364 ();
 sg13g2_fill_1 FILLER_75_2369 ();
 sg13g2_fill_2 FILLER_75_2375 ();
 sg13g2_fill_2 FILLER_75_2381 ();
 sg13g2_fill_1 FILLER_75_2383 ();
 sg13g2_fill_2 FILLER_75_2398 ();
 sg13g2_fill_1 FILLER_75_2400 ();
 sg13g2_fill_2 FILLER_75_2407 ();
 sg13g2_fill_1 FILLER_75_2409 ();
 sg13g2_decap_8 FILLER_75_2425 ();
 sg13g2_fill_2 FILLER_75_2432 ();
 sg13g2_fill_1 FILLER_75_2434 ();
 sg13g2_decap_8 FILLER_75_2439 ();
 sg13g2_decap_4 FILLER_75_2446 ();
 sg13g2_fill_1 FILLER_75_2450 ();
 sg13g2_fill_2 FILLER_75_2455 ();
 sg13g2_fill_1 FILLER_75_2457 ();
 sg13g2_fill_2 FILLER_75_2467 ();
 sg13g2_fill_1 FILLER_75_2469 ();
 sg13g2_decap_8 FILLER_75_2474 ();
 sg13g2_decap_8 FILLER_75_2481 ();
 sg13g2_decap_4 FILLER_75_2488 ();
 sg13g2_fill_2 FILLER_75_2492 ();
 sg13g2_decap_8 FILLER_75_2503 ();
 sg13g2_decap_4 FILLER_75_2510 ();
 sg13g2_fill_2 FILLER_75_2514 ();
 sg13g2_decap_8 FILLER_75_2521 ();
 sg13g2_decap_4 FILLER_75_2528 ();
 sg13g2_fill_2 FILLER_75_2538 ();
 sg13g2_fill_1 FILLER_75_2540 ();
 sg13g2_fill_2 FILLER_75_2545 ();
 sg13g2_fill_1 FILLER_75_2547 ();
 sg13g2_fill_2 FILLER_75_2554 ();
 sg13g2_decap_8 FILLER_75_2560 ();
 sg13g2_decap_8 FILLER_75_2567 ();
 sg13g2_fill_1 FILLER_75_2574 ();
 sg13g2_fill_1 FILLER_75_2583 ();
 sg13g2_fill_1 FILLER_75_2588 ();
 sg13g2_fill_2 FILLER_75_2599 ();
 sg13g2_fill_1 FILLER_75_2611 ();
 sg13g2_fill_2 FILLER_75_2638 ();
 sg13g2_decap_4 FILLER_75_2666 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_4 FILLER_76_18 ();
 sg13g2_fill_1 FILLER_76_22 ();
 sg13g2_fill_1 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_38 ();
 sg13g2_fill_1 FILLER_76_69 ();
 sg13g2_decap_8 FILLER_76_113 ();
 sg13g2_fill_2 FILLER_76_120 ();
 sg13g2_fill_2 FILLER_76_126 ();
 sg13g2_fill_1 FILLER_76_216 ();
 sg13g2_fill_2 FILLER_76_222 ();
 sg13g2_fill_2 FILLER_76_229 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_2 FILLER_76_268 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_fill_1 FILLER_76_294 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_decap_4 FILLER_76_340 ();
 sg13g2_fill_2 FILLER_76_344 ();
 sg13g2_fill_1 FILLER_76_367 ();
 sg13g2_decap_8 FILLER_76_372 ();
 sg13g2_decap_4 FILLER_76_379 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_fill_1 FILLER_76_441 ();
 sg13g2_fill_1 FILLER_76_449 ();
 sg13g2_fill_1 FILLER_76_455 ();
 sg13g2_fill_1 FILLER_76_491 ();
 sg13g2_fill_2 FILLER_76_496 ();
 sg13g2_fill_1 FILLER_76_498 ();
 sg13g2_decap_8 FILLER_76_509 ();
 sg13g2_fill_2 FILLER_76_520 ();
 sg13g2_fill_1 FILLER_76_522 ();
 sg13g2_fill_2 FILLER_76_526 ();
 sg13g2_fill_1 FILLER_76_528 ();
 sg13g2_decap_8 FILLER_76_533 ();
 sg13g2_decap_8 FILLER_76_540 ();
 sg13g2_decap_4 FILLER_76_547 ();
 sg13g2_fill_1 FILLER_76_551 ();
 sg13g2_fill_2 FILLER_76_556 ();
 sg13g2_fill_1 FILLER_76_558 ();
 sg13g2_decap_8 FILLER_76_604 ();
 sg13g2_fill_2 FILLER_76_628 ();
 sg13g2_fill_1 FILLER_76_634 ();
 sg13g2_fill_1 FILLER_76_640 ();
 sg13g2_fill_2 FILLER_76_663 ();
 sg13g2_fill_2 FILLER_76_689 ();
 sg13g2_decap_8 FILLER_76_719 ();
 sg13g2_fill_2 FILLER_76_726 ();
 sg13g2_fill_1 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_fill_1 FILLER_76_749 ();
 sg13g2_fill_1 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_fill_2 FILLER_76_819 ();
 sg13g2_fill_1 FILLER_76_821 ();
 sg13g2_decap_8 FILLER_76_828 ();
 sg13g2_decap_8 FILLER_76_879 ();
 sg13g2_fill_1 FILLER_76_896 ();
 sg13g2_decap_8 FILLER_76_959 ();
 sg13g2_decap_8 FILLER_76_966 ();
 sg13g2_decap_4 FILLER_76_973 ();
 sg13g2_fill_2 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_985 ();
 sg13g2_fill_1 FILLER_76_992 ();
 sg13g2_decap_8 FILLER_76_997 ();
 sg13g2_decap_8 FILLER_76_1004 ();
 sg13g2_fill_2 FILLER_76_1011 ();
 sg13g2_decap_4 FILLER_76_1023 ();
 sg13g2_fill_1 FILLER_76_1027 ();
 sg13g2_decap_8 FILLER_76_1033 ();
 sg13g2_fill_2 FILLER_76_1040 ();
 sg13g2_fill_2 FILLER_76_1078 ();
 sg13g2_fill_1 FILLER_76_1080 ();
 sg13g2_decap_4 FILLER_76_1091 ();
 sg13g2_fill_2 FILLER_76_1095 ();
 sg13g2_fill_2 FILLER_76_1118 ();
 sg13g2_fill_1 FILLER_76_1120 ();
 sg13g2_decap_4 FILLER_76_1137 ();
 sg13g2_decap_4 FILLER_76_1149 ();
 sg13g2_fill_1 FILLER_76_1153 ();
 sg13g2_fill_2 FILLER_76_1180 ();
 sg13g2_fill_1 FILLER_76_1182 ();
 sg13g2_decap_8 FILLER_76_1217 ();
 sg13g2_decap_4 FILLER_76_1224 ();
 sg13g2_fill_1 FILLER_76_1239 ();
 sg13g2_decap_4 FILLER_76_1258 ();
 sg13g2_decap_4 FILLER_76_1284 ();
 sg13g2_fill_2 FILLER_76_1288 ();
 sg13g2_fill_2 FILLER_76_1295 ();
 sg13g2_fill_1 FILLER_76_1297 ();
 sg13g2_decap_4 FILLER_76_1345 ();
 sg13g2_fill_2 FILLER_76_1394 ();
 sg13g2_fill_2 FILLER_76_1404 ();
 sg13g2_fill_1 FILLER_76_1406 ();
 sg13g2_fill_2 FILLER_76_1421 ();
 sg13g2_fill_2 FILLER_76_1431 ();
 sg13g2_fill_2 FILLER_76_1466 ();
 sg13g2_fill_1 FILLER_76_1473 ();
 sg13g2_fill_2 FILLER_76_1483 ();
 sg13g2_fill_1 FILLER_76_1485 ();
 sg13g2_fill_2 FILLER_76_1505 ();
 sg13g2_decap_4 FILLER_76_1520 ();
 sg13g2_fill_1 FILLER_76_1524 ();
 sg13g2_decap_4 FILLER_76_1529 ();
 sg13g2_fill_1 FILLER_76_1571 ();
 sg13g2_decap_4 FILLER_76_1576 ();
 sg13g2_fill_1 FILLER_76_1588 ();
 sg13g2_fill_1 FILLER_76_1601 ();
 sg13g2_fill_2 FILLER_76_1615 ();
 sg13g2_fill_2 FILLER_76_1621 ();
 sg13g2_fill_1 FILLER_76_1623 ();
 sg13g2_fill_2 FILLER_76_1629 ();
 sg13g2_fill_1 FILLER_76_1631 ();
 sg13g2_fill_2 FILLER_76_1636 ();
 sg13g2_fill_1 FILLER_76_1638 ();
 sg13g2_fill_2 FILLER_76_1660 ();
 sg13g2_fill_1 FILLER_76_1700 ();
 sg13g2_fill_2 FILLER_76_1706 ();
 sg13g2_fill_1 FILLER_76_1738 ();
 sg13g2_fill_1 FILLER_76_1745 ();
 sg13g2_decap_4 FILLER_76_1758 ();
 sg13g2_fill_1 FILLER_76_1762 ();
 sg13g2_fill_2 FILLER_76_1767 ();
 sg13g2_fill_1 FILLER_76_1769 ();
 sg13g2_decap_4 FILLER_76_1789 ();
 sg13g2_fill_1 FILLER_76_1793 ();
 sg13g2_fill_2 FILLER_76_1813 ();
 sg13g2_fill_2 FILLER_76_1819 ();
 sg13g2_fill_1 FILLER_76_1825 ();
 sg13g2_fill_2 FILLER_76_1831 ();
 sg13g2_fill_1 FILLER_76_1853 ();
 sg13g2_fill_2 FILLER_76_1862 ();
 sg13g2_fill_1 FILLER_76_1897 ();
 sg13g2_fill_2 FILLER_76_1938 ();
 sg13g2_decap_8 FILLER_76_1964 ();
 sg13g2_decap_8 FILLER_76_1971 ();
 sg13g2_decap_8 FILLER_76_1982 ();
 sg13g2_decap_8 FILLER_76_1989 ();
 sg13g2_decap_4 FILLER_76_1996 ();
 sg13g2_decap_8 FILLER_76_2010 ();
 sg13g2_decap_8 FILLER_76_2017 ();
 sg13g2_decap_8 FILLER_76_2024 ();
 sg13g2_decap_8 FILLER_76_2036 ();
 sg13g2_decap_4 FILLER_76_2043 ();
 sg13g2_fill_2 FILLER_76_2073 ();
 sg13g2_fill_1 FILLER_76_2075 ();
 sg13g2_decap_4 FILLER_76_2112 ();
 sg13g2_fill_1 FILLER_76_2116 ();
 sg13g2_fill_1 FILLER_76_2127 ();
 sg13g2_fill_2 FILLER_76_2157 ();
 sg13g2_fill_2 FILLER_76_2195 ();
 sg13g2_decap_4 FILLER_76_2233 ();
 sg13g2_fill_2 FILLER_76_2237 ();
 sg13g2_decap_8 FILLER_76_2249 ();
 sg13g2_decap_8 FILLER_76_2256 ();
 sg13g2_fill_2 FILLER_76_2263 ();
 sg13g2_fill_1 FILLER_76_2265 ();
 sg13g2_decap_8 FILLER_76_2276 ();
 sg13g2_decap_8 FILLER_76_2283 ();
 sg13g2_fill_1 FILLER_76_2290 ();
 sg13g2_fill_2 FILLER_76_2341 ();
 sg13g2_fill_2 FILLER_76_2356 ();
 sg13g2_fill_1 FILLER_76_2401 ();
 sg13g2_fill_2 FILLER_76_2415 ();
 sg13g2_fill_1 FILLER_76_2417 ();
 sg13g2_decap_4 FILLER_76_2429 ();
 sg13g2_fill_1 FILLER_76_2441 ();
 sg13g2_fill_2 FILLER_76_2460 ();
 sg13g2_fill_2 FILLER_76_2466 ();
 sg13g2_fill_1 FILLER_76_2468 ();
 sg13g2_decap_8 FILLER_76_2482 ();
 sg13g2_fill_1 FILLER_76_2489 ();
 sg13g2_fill_1 FILLER_76_2521 ();
 sg13g2_decap_4 FILLER_76_2548 ();
 sg13g2_fill_2 FILLER_76_2565 ();
 sg13g2_fill_1 FILLER_76_2567 ();
 sg13g2_decap_4 FILLER_76_2577 ();
 sg13g2_fill_1 FILLER_76_2581 ();
 sg13g2_fill_2 FILLER_76_2592 ();
 sg13g2_fill_1 FILLER_76_2594 ();
 sg13g2_decap_8 FILLER_76_2605 ();
 sg13g2_decap_8 FILLER_76_2612 ();
 sg13g2_fill_1 FILLER_76_2619 ();
 sg13g2_decap_4 FILLER_76_2624 ();
 sg13g2_fill_1 FILLER_76_2628 ();
 sg13g2_decap_4 FILLER_76_2665 ();
 sg13g2_fill_1 FILLER_76_2669 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_2 ();
 sg13g2_fill_2 FILLER_77_29 ();
 sg13g2_fill_1 FILLER_77_84 ();
 sg13g2_fill_1 FILLER_77_90 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_1 FILLER_77_215 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_4 FILLER_77_266 ();
 sg13g2_decap_4 FILLER_77_275 ();
 sg13g2_fill_1 FILLER_77_288 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_fill_1 FILLER_77_301 ();
 sg13g2_fill_1 FILLER_77_311 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_decap_8 FILLER_77_332 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_2 FILLER_77_364 ();
 sg13g2_fill_2 FILLER_77_392 ();
 sg13g2_fill_1 FILLER_77_394 ();
 sg13g2_decap_8 FILLER_77_403 ();
 sg13g2_decap_8 FILLER_77_410 ();
 sg13g2_decap_8 FILLER_77_417 ();
 sg13g2_decap_8 FILLER_77_424 ();
 sg13g2_fill_2 FILLER_77_431 ();
 sg13g2_fill_1 FILLER_77_433 ();
 sg13g2_fill_2 FILLER_77_484 ();
 sg13g2_fill_1 FILLER_77_491 ();
 sg13g2_fill_2 FILLER_77_511 ();
 sg13g2_fill_1 FILLER_77_538 ();
 sg13g2_decap_8 FILLER_77_543 ();
 sg13g2_decap_4 FILLER_77_550 ();
 sg13g2_fill_2 FILLER_77_580 ();
 sg13g2_fill_1 FILLER_77_582 ();
 sg13g2_decap_4 FILLER_77_590 ();
 sg13g2_fill_2 FILLER_77_594 ();
 sg13g2_fill_1 FILLER_77_689 ();
 sg13g2_fill_2 FILLER_77_702 ();
 sg13g2_fill_2 FILLER_77_730 ();
 sg13g2_fill_2 FILLER_77_736 ();
 sg13g2_fill_1 FILLER_77_738 ();
 sg13g2_fill_2 FILLER_77_765 ();
 sg13g2_fill_1 FILLER_77_767 ();
 sg13g2_fill_2 FILLER_77_772 ();
 sg13g2_fill_1 FILLER_77_774 ();
 sg13g2_fill_2 FILLER_77_795 ();
 sg13g2_decap_8 FILLER_77_853 ();
 sg13g2_decap_8 FILLER_77_919 ();
 sg13g2_fill_1 FILLER_77_957 ();
 sg13g2_fill_2 FILLER_77_972 ();
 sg13g2_decap_4 FILLER_77_1010 ();
 sg13g2_fill_2 FILLER_77_1044 ();
 sg13g2_decap_4 FILLER_77_1085 ();
 sg13g2_fill_1 FILLER_77_1089 ();
 sg13g2_decap_8 FILLER_77_1134 ();
 sg13g2_fill_1 FILLER_77_1141 ();
 sg13g2_fill_1 FILLER_77_1152 ();
 sg13g2_fill_1 FILLER_77_1157 ();
 sg13g2_fill_2 FILLER_77_1184 ();
 sg13g2_fill_1 FILLER_77_1191 ();
 sg13g2_decap_4 FILLER_77_1222 ();
 sg13g2_fill_2 FILLER_77_1226 ();
 sg13g2_fill_2 FILLER_77_1265 ();
 sg13g2_fill_1 FILLER_77_1267 ();
 sg13g2_fill_2 FILLER_77_1293 ();
 sg13g2_fill_1 FILLER_77_1310 ();
 sg13g2_fill_2 FILLER_77_1316 ();
 sg13g2_fill_1 FILLER_77_1324 ();
 sg13g2_fill_1 FILLER_77_1334 ();
 sg13g2_fill_1 FILLER_77_1360 ();
 sg13g2_fill_1 FILLER_77_1399 ();
 sg13g2_fill_2 FILLER_77_1409 ();
 sg13g2_fill_1 FILLER_77_1445 ();
 sg13g2_fill_1 FILLER_77_1451 ();
 sg13g2_decap_8 FILLER_77_1456 ();
 sg13g2_fill_1 FILLER_77_1463 ();
 sg13g2_fill_2 FILLER_77_1473 ();
 sg13g2_fill_1 FILLER_77_1495 ();
 sg13g2_fill_1 FILLER_77_1505 ();
 sg13g2_fill_1 FILLER_77_1526 ();
 sg13g2_fill_2 FILLER_77_1553 ();
 sg13g2_fill_1 FILLER_77_1572 ();
 sg13g2_decap_4 FILLER_77_1687 ();
 sg13g2_fill_1 FILLER_77_1709 ();
 sg13g2_decap_4 FILLER_77_1732 ();
 sg13g2_fill_2 FILLER_77_1780 ();
 sg13g2_fill_2 FILLER_77_1785 ();
 sg13g2_fill_1 FILLER_77_1787 ();
 sg13g2_decap_4 FILLER_77_1793 ();
 sg13g2_fill_2 FILLER_77_1814 ();
 sg13g2_fill_1 FILLER_77_1816 ();
 sg13g2_fill_1 FILLER_77_1835 ();
 sg13g2_fill_1 FILLER_77_1841 ();
 sg13g2_decap_4 FILLER_77_1871 ();
 sg13g2_fill_1 FILLER_77_1880 ();
 sg13g2_fill_2 FILLER_77_1889 ();
 sg13g2_fill_1 FILLER_77_1891 ();
 sg13g2_fill_2 FILLER_77_1897 ();
 sg13g2_fill_2 FILLER_77_1925 ();
 sg13g2_fill_2 FILLER_77_1949 ();
 sg13g2_fill_2 FILLER_77_1978 ();
 sg13g2_decap_4 FILLER_77_2016 ();
 sg13g2_fill_1 FILLER_77_2030 ();
 sg13g2_decap_8 FILLER_77_2108 ();
 sg13g2_fill_1 FILLER_77_2115 ();
 sg13g2_fill_2 FILLER_77_2126 ();
 sg13g2_fill_1 FILLER_77_2128 ();
 sg13g2_decap_8 FILLER_77_2155 ();
 sg13g2_decap_4 FILLER_77_2162 ();
 sg13g2_fill_2 FILLER_77_2166 ();
 sg13g2_decap_8 FILLER_77_2189 ();
 sg13g2_fill_2 FILLER_77_2196 ();
 sg13g2_fill_2 FILLER_77_2211 ();
 sg13g2_fill_1 FILLER_77_2213 ();
 sg13g2_decap_4 FILLER_77_2240 ();
 sg13g2_fill_1 FILLER_77_2244 ();
 sg13g2_decap_4 FILLER_77_2271 ();
 sg13g2_fill_1 FILLER_77_2357 ();
 sg13g2_fill_1 FILLER_77_2362 ();
 sg13g2_fill_2 FILLER_77_2368 ();
 sg13g2_fill_2 FILLER_77_2401 ();
 sg13g2_fill_1 FILLER_77_2403 ();
 sg13g2_fill_1 FILLER_77_2430 ();
 sg13g2_fill_1 FILLER_77_2462 ();
 sg13g2_fill_1 FILLER_77_2489 ();
 sg13g2_fill_2 FILLER_77_2516 ();
 sg13g2_fill_2 FILLER_77_2534 ();
 sg13g2_decap_8 FILLER_77_2562 ();
 sg13g2_decap_4 FILLER_77_2585 ();
 sg13g2_decap_8 FILLER_77_2628 ();
 sg13g2_decap_8 FILLER_77_2635 ();
 sg13g2_fill_1 FILLER_77_2642 ();
 sg13g2_decap_8 FILLER_77_2651 ();
 sg13g2_decap_8 FILLER_77_2658 ();
 sg13g2_decap_4 FILLER_77_2665 ();
 sg13g2_fill_1 FILLER_77_2669 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_32 ();
 sg13g2_fill_1 FILLER_78_38 ();
 sg13g2_fill_1 FILLER_78_75 ();
 sg13g2_fill_1 FILLER_78_116 ();
 sg13g2_fill_1 FILLER_78_126 ();
 sg13g2_fill_1 FILLER_78_194 ();
 sg13g2_decap_4 FILLER_78_259 ();
 sg13g2_fill_1 FILLER_78_263 ();
 sg13g2_decap_8 FILLER_78_269 ();
 sg13g2_decap_4 FILLER_78_276 ();
 sg13g2_decap_4 FILLER_78_288 ();
 sg13g2_fill_1 FILLER_78_332 ();
 sg13g2_decap_4 FILLER_78_337 ();
 sg13g2_fill_2 FILLER_78_341 ();
 sg13g2_fill_2 FILLER_78_352 ();
 sg13g2_fill_1 FILLER_78_359 ();
 sg13g2_fill_1 FILLER_78_374 ();
 sg13g2_fill_1 FILLER_78_410 ();
 sg13g2_fill_1 FILLER_78_477 ();
 sg13g2_fill_2 FILLER_78_483 ();
 sg13g2_fill_1 FILLER_78_495 ();
 sg13g2_fill_2 FILLER_78_511 ();
 sg13g2_fill_1 FILLER_78_544 ();
 sg13g2_fill_2 FILLER_78_571 ();
 sg13g2_fill_1 FILLER_78_573 ();
 sg13g2_fill_1 FILLER_78_639 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_fill_2 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_719 ();
 sg13g2_fill_1 FILLER_78_726 ();
 sg13g2_decap_8 FILLER_78_753 ();
 sg13g2_decap_8 FILLER_78_760 ();
 sg13g2_fill_1 FILLER_78_767 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_fill_1 FILLER_78_801 ();
 sg13g2_fill_2 FILLER_78_828 ();
 sg13g2_fill_1 FILLER_78_856 ();
 sg13g2_fill_1 FILLER_78_871 ();
 sg13g2_decap_4 FILLER_78_960 ();
 sg13g2_fill_1 FILLER_78_964 ();
 sg13g2_fill_1 FILLER_78_1001 ();
 sg13g2_fill_1 FILLER_78_1038 ();
 sg13g2_fill_1 FILLER_78_1085 ();
 sg13g2_fill_1 FILLER_78_1112 ();
 sg13g2_fill_2 FILLER_78_1169 ();
 sg13g2_fill_1 FILLER_78_1171 ();
 sg13g2_fill_1 FILLER_78_1207 ();
 sg13g2_decap_8 FILLER_78_1212 ();
 sg13g2_decap_8 FILLER_78_1219 ();
 sg13g2_decap_8 FILLER_78_1226 ();
 sg13g2_decap_4 FILLER_78_1233 ();
 sg13g2_fill_2 FILLER_78_1256 ();
 sg13g2_fill_1 FILLER_78_1258 ();
 sg13g2_fill_1 FILLER_78_1271 ();
 sg13g2_fill_2 FILLER_78_1282 ();
 sg13g2_fill_1 FILLER_78_1284 ();
 sg13g2_fill_1 FILLER_78_1293 ();
 sg13g2_fill_2 FILLER_78_1336 ();
 sg13g2_fill_1 FILLER_78_1343 ();
 sg13g2_fill_1 FILLER_78_1358 ();
 sg13g2_decap_8 FILLER_78_1381 ();
 sg13g2_decap_8 FILLER_78_1388 ();
 sg13g2_fill_2 FILLER_78_1462 ();
 sg13g2_fill_1 FILLER_78_1464 ();
 sg13g2_fill_1 FILLER_78_1477 ();
 sg13g2_fill_2 FILLER_78_1499 ();
 sg13g2_fill_1 FILLER_78_1501 ();
 sg13g2_decap_8 FILLER_78_1642 ();
 sg13g2_decap_8 FILLER_78_1649 ();
 sg13g2_decap_4 FILLER_78_1662 ();
 sg13g2_fill_1 FILLER_78_1677 ();
 sg13g2_fill_1 FILLER_78_1690 ();
 sg13g2_fill_2 FILLER_78_1706 ();
 sg13g2_fill_1 FILLER_78_1708 ();
 sg13g2_fill_2 FILLER_78_1732 ();
 sg13g2_fill_1 FILLER_78_1734 ();
 sg13g2_decap_4 FILLER_78_1760 ();
 sg13g2_fill_2 FILLER_78_1764 ();
 sg13g2_decap_4 FILLER_78_1775 ();
 sg13g2_fill_1 FILLER_78_1789 ();
 sg13g2_fill_1 FILLER_78_1800 ();
 sg13g2_fill_1 FILLER_78_1809 ();
 sg13g2_fill_2 FILLER_78_1819 ();
 sg13g2_decap_4 FILLER_78_1844 ();
 sg13g2_fill_1 FILLER_78_1848 ();
 sg13g2_fill_1 FILLER_78_1861 ();
 sg13g2_fill_1 FILLER_78_1867 ();
 sg13g2_fill_1 FILLER_78_1872 ();
 sg13g2_fill_2 FILLER_78_1893 ();
 sg13g2_fill_1 FILLER_78_1908 ();
 sg13g2_fill_1 FILLER_78_1920 ();
 sg13g2_decap_4 FILLER_78_1932 ();
 sg13g2_decap_8 FILLER_78_1966 ();
 sg13g2_decap_4 FILLER_78_1973 ();
 sg13g2_fill_1 FILLER_78_1977 ();
 sg13g2_fill_2 FILLER_78_2004 ();
 sg13g2_fill_2 FILLER_78_2027 ();
 sg13g2_fill_2 FILLER_78_2055 ();
 sg13g2_decap_8 FILLER_78_2067 ();
 sg13g2_decap_8 FILLER_78_2074 ();
 sg13g2_fill_1 FILLER_78_2081 ();
 sg13g2_fill_1 FILLER_78_2086 ();
 sg13g2_fill_2 FILLER_78_2091 ();
 sg13g2_fill_1 FILLER_78_2093 ();
 sg13g2_fill_2 FILLER_78_2160 ();
 sg13g2_fill_1 FILLER_78_2162 ();
 sg13g2_fill_1 FILLER_78_2167 ();
 sg13g2_decap_8 FILLER_78_2194 ();
 sg13g2_fill_2 FILLER_78_2237 ();
 sg13g2_fill_1 FILLER_78_2239 ();
 sg13g2_fill_2 FILLER_78_2301 ();
 sg13g2_fill_1 FILLER_78_2303 ();
 sg13g2_fill_2 FILLER_78_2334 ();
 sg13g2_fill_1 FILLER_78_2393 ();
 sg13g2_fill_1 FILLER_78_2398 ();
 sg13g2_fill_2 FILLER_78_2486 ();
 sg13g2_fill_1 FILLER_78_2488 ();
 sg13g2_decap_4 FILLER_78_2520 ();
 sg13g2_fill_2 FILLER_78_2563 ();
 sg13g2_fill_1 FILLER_78_2601 ();
 sg13g2_decap_8 FILLER_78_2628 ();
 sg13g2_decap_8 FILLER_78_2635 ();
 sg13g2_decap_8 FILLER_78_2642 ();
 sg13g2_decap_8 FILLER_78_2649 ();
 sg13g2_decap_8 FILLER_78_2656 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_4 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_4 ();
 sg13g2_fill_1 FILLER_79_36 ();
 sg13g2_fill_1 FILLER_79_42 ();
 sg13g2_fill_1 FILLER_79_53 ();
 sg13g2_fill_1 FILLER_79_76 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_fill_1 FILLER_79_117 ();
 sg13g2_fill_1 FILLER_79_144 ();
 sg13g2_fill_2 FILLER_79_150 ();
 sg13g2_fill_1 FILLER_79_156 ();
 sg13g2_fill_1 FILLER_79_163 ();
 sg13g2_fill_1 FILLER_79_181 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_fill_1 FILLER_79_200 ();
 sg13g2_fill_2 FILLER_79_208 ();
 sg13g2_fill_1 FILLER_79_242 ();
 sg13g2_fill_2 FILLER_79_269 ();
 sg13g2_fill_1 FILLER_79_275 ();
 sg13g2_fill_1 FILLER_79_354 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_fill_1 FILLER_79_409 ();
 sg13g2_fill_2 FILLER_79_436 ();
 sg13g2_fill_2 FILLER_79_493 ();
 sg13g2_fill_1 FILLER_79_555 ();
 sg13g2_fill_2 FILLER_79_573 ();
 sg13g2_fill_2 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_723 ();
 sg13g2_fill_2 FILLER_79_730 ();
 sg13g2_fill_1 FILLER_79_732 ();
 sg13g2_decap_4 FILLER_79_737 ();
 sg13g2_fill_1 FILLER_79_751 ();
 sg13g2_decap_4 FILLER_79_762 ();
 sg13g2_fill_2 FILLER_79_766 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_fill_2 FILLER_79_809 ();
 sg13g2_fill_1 FILLER_79_811 ();
 sg13g2_fill_1 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_857 ();
 sg13g2_fill_1 FILLER_79_864 ();
 sg13g2_decap_8 FILLER_79_891 ();
 sg13g2_fill_1 FILLER_79_934 ();
 sg13g2_fill_2 FILLER_79_945 ();
 sg13g2_fill_2 FILLER_79_951 ();
 sg13g2_fill_2 FILLER_79_979 ();
 sg13g2_fill_1 FILLER_79_981 ();
 sg13g2_fill_2 FILLER_79_996 ();
 sg13g2_fill_1 FILLER_79_998 ();
 sg13g2_fill_2 FILLER_79_1047 ();
 sg13g2_decap_8 FILLER_79_1125 ();
 sg13g2_decap_8 FILLER_79_1132 ();
 sg13g2_fill_2 FILLER_79_1143 ();
 sg13g2_fill_1 FILLER_79_1145 ();
 sg13g2_decap_8 FILLER_79_1172 ();
 sg13g2_fill_2 FILLER_79_1179 ();
 sg13g2_fill_1 FILLER_79_1181 ();
 sg13g2_fill_2 FILLER_79_1186 ();
 sg13g2_decap_8 FILLER_79_1214 ();
 sg13g2_fill_2 FILLER_79_1221 ();
 sg13g2_decap_4 FILLER_79_1254 ();
 sg13g2_decap_8 FILLER_79_1270 ();
 sg13g2_fill_2 FILLER_79_1277 ();
 sg13g2_fill_2 FILLER_79_1284 ();
 sg13g2_fill_1 FILLER_79_1322 ();
 sg13g2_decap_8 FILLER_79_1333 ();
 sg13g2_decap_8 FILLER_79_1340 ();
 sg13g2_decap_4 FILLER_79_1354 ();
 sg13g2_fill_1 FILLER_79_1364 ();
 sg13g2_fill_2 FILLER_79_1371 ();
 sg13g2_fill_1 FILLER_79_1373 ();
 sg13g2_decap_8 FILLER_79_1404 ();
 sg13g2_fill_1 FILLER_79_1411 ();
 sg13g2_decap_4 FILLER_79_1439 ();
 sg13g2_fill_2 FILLER_79_1447 ();
 sg13g2_fill_1 FILLER_79_1449 ();
 sg13g2_decap_8 FILLER_79_1457 ();
 sg13g2_decap_8 FILLER_79_1464 ();
 sg13g2_decap_8 FILLER_79_1480 ();
 sg13g2_fill_2 FILLER_79_1487 ();
 sg13g2_decap_4 FILLER_79_1493 ();
 sg13g2_decap_4 FILLER_79_1511 ();
 sg13g2_decap_8 FILLER_79_1529 ();
 sg13g2_decap_4 FILLER_79_1536 ();
 sg13g2_fill_1 FILLER_79_1540 ();
 sg13g2_fill_2 FILLER_79_1546 ();
 sg13g2_fill_2 FILLER_79_1553 ();
 sg13g2_fill_2 FILLER_79_1587 ();
 sg13g2_fill_2 FILLER_79_1623 ();
 sg13g2_decap_8 FILLER_79_1651 ();
 sg13g2_decap_8 FILLER_79_1658 ();
 sg13g2_decap_8 FILLER_79_1665 ();
 sg13g2_decap_4 FILLER_79_1672 ();
 sg13g2_fill_2 FILLER_79_1681 ();
 sg13g2_fill_2 FILLER_79_1688 ();
 sg13g2_fill_1 FILLER_79_1690 ();
 sg13g2_decap_8 FILLER_79_1714 ();
 sg13g2_fill_1 FILLER_79_1721 ();
 sg13g2_decap_8 FILLER_79_1727 ();
 sg13g2_decap_8 FILLER_79_1734 ();
 sg13g2_decap_8 FILLER_79_1741 ();
 sg13g2_decap_4 FILLER_79_1782 ();
 sg13g2_fill_1 FILLER_79_1795 ();
 sg13g2_fill_1 FILLER_79_1805 ();
 sg13g2_fill_1 FILLER_79_1816 ();
 sg13g2_decap_8 FILLER_79_1834 ();
 sg13g2_decap_8 FILLER_79_1841 ();
 sg13g2_decap_4 FILLER_79_1848 ();
 sg13g2_fill_2 FILLER_79_1852 ();
 sg13g2_fill_1 FILLER_79_1874 ();
 sg13g2_decap_8 FILLER_79_1879 ();
 sg13g2_decap_8 FILLER_79_1886 ();
 sg13g2_decap_8 FILLER_79_1893 ();
 sg13g2_fill_2 FILLER_79_1909 ();
 sg13g2_fill_2 FILLER_79_1916 ();
 sg13g2_fill_1 FILLER_79_1918 ();
 sg13g2_fill_2 FILLER_79_1923 ();
 sg13g2_fill_1 FILLER_79_1925 ();
 sg13g2_fill_2 FILLER_79_1931 ();
 sg13g2_fill_1 FILLER_79_1933 ();
 sg13g2_decap_4 FILLER_79_1943 ();
 sg13g2_fill_1 FILLER_79_1947 ();
 sg13g2_fill_1 FILLER_79_1954 ();
 sg13g2_decap_8 FILLER_79_1960 ();
 sg13g2_decap_4 FILLER_79_1967 ();
 sg13g2_fill_2 FILLER_79_1971 ();
 sg13g2_fill_2 FILLER_79_1999 ();
 sg13g2_fill_1 FILLER_79_2001 ();
 sg13g2_fill_2 FILLER_79_2028 ();
 sg13g2_decap_8 FILLER_79_2113 ();
 sg13g2_decap_8 FILLER_79_2120 ();
 sg13g2_decap_4 FILLER_79_2127 ();
 sg13g2_fill_1 FILLER_79_2131 ();
 sg13g2_fill_1 FILLER_79_2136 ();
 sg13g2_fill_2 FILLER_79_2141 ();
 sg13g2_fill_2 FILLER_79_2169 ();
 sg13g2_fill_1 FILLER_79_2197 ();
 sg13g2_fill_2 FILLER_79_2208 ();
 sg13g2_fill_1 FILLER_79_2214 ();
 sg13g2_fill_1 FILLER_79_2241 ();
 sg13g2_fill_1 FILLER_79_2256 ();
 sg13g2_fill_1 FILLER_79_2278 ();
 sg13g2_fill_2 FILLER_79_2283 ();
 sg13g2_fill_1 FILLER_79_2285 ();
 sg13g2_decap_4 FILLER_79_2290 ();
 sg13g2_fill_1 FILLER_79_2294 ();
 sg13g2_fill_1 FILLER_79_2321 ();
 sg13g2_decap_4 FILLER_79_2352 ();
 sg13g2_fill_2 FILLER_79_2356 ();
 sg13g2_fill_2 FILLER_79_2362 ();
 sg13g2_fill_1 FILLER_79_2364 ();
 sg13g2_fill_2 FILLER_79_2370 ();
 sg13g2_fill_1 FILLER_79_2372 ();
 sg13g2_fill_2 FILLER_79_2377 ();
 sg13g2_fill_1 FILLER_79_2379 ();
 sg13g2_fill_2 FILLER_79_2410 ();
 sg13g2_fill_2 FILLER_79_2417 ();
 sg13g2_fill_1 FILLER_79_2419 ();
 sg13g2_decap_8 FILLER_79_2424 ();
 sg13g2_fill_2 FILLER_79_2435 ();
 sg13g2_decap_4 FILLER_79_2489 ();
 sg13g2_fill_1 FILLER_79_2513 ();
 sg13g2_decap_4 FILLER_79_2566 ();
 sg13g2_fill_2 FILLER_79_2596 ();
 sg13g2_fill_1 FILLER_79_2598 ();
 sg13g2_fill_2 FILLER_79_2609 ();
 sg13g2_decap_8 FILLER_79_2637 ();
 sg13g2_decap_8 FILLER_79_2644 ();
 sg13g2_decap_8 FILLER_79_2651 ();
 sg13g2_decap_8 FILLER_79_2658 ();
 sg13g2_decap_4 FILLER_79_2665 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_2 FILLER_80_14 ();
 sg13g2_fill_1 FILLER_80_16 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_77 ();
 sg13g2_fill_2 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_2 FILLER_80_196 ();
 sg13g2_fill_2 FILLER_80_268 ();
 sg13g2_decap_4 FILLER_80_290 ();
 sg13g2_fill_1 FILLER_80_294 ();
 sg13g2_fill_1 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_312 ();
 sg13g2_decap_8 FILLER_80_319 ();
 sg13g2_decap_8 FILLER_80_326 ();
 sg13g2_fill_1 FILLER_80_333 ();
 sg13g2_decap_8 FILLER_80_339 ();
 sg13g2_fill_1 FILLER_80_351 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_fill_2 FILLER_80_360 ();
 sg13g2_decap_8 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_4 FILLER_80_380 ();
 sg13g2_fill_2 FILLER_80_384 ();
 sg13g2_decap_4 FILLER_80_414 ();
 sg13g2_fill_2 FILLER_80_430 ();
 sg13g2_decap_4 FILLER_80_442 ();
 sg13g2_fill_1 FILLER_80_446 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_4 FILLER_80_469 ();
 sg13g2_fill_1 FILLER_80_473 ();
 sg13g2_decap_8 FILLER_80_484 ();
 sg13g2_decap_4 FILLER_80_491 ();
 sg13g2_fill_2 FILLER_80_499 ();
 sg13g2_decap_8 FILLER_80_505 ();
 sg13g2_decap_8 FILLER_80_512 ();
 sg13g2_decap_8 FILLER_80_519 ();
 sg13g2_fill_1 FILLER_80_526 ();
 sg13g2_decap_4 FILLER_80_531 ();
 sg13g2_fill_2 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_541 ();
 sg13g2_decap_8 FILLER_80_548 ();
 sg13g2_fill_1 FILLER_80_555 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_572 ();
 sg13g2_fill_1 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_4 FILLER_80_602 ();
 sg13g2_fill_2 FILLER_80_606 ();
 sg13g2_decap_8 FILLER_80_612 ();
 sg13g2_decap_8 FILLER_80_619 ();
 sg13g2_decap_8 FILLER_80_626 ();
 sg13g2_decap_4 FILLER_80_633 ();
 sg13g2_fill_2 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_643 ();
 sg13g2_decap_4 FILLER_80_654 ();
 sg13g2_fill_2 FILLER_80_658 ();
 sg13g2_fill_2 FILLER_80_664 ();
 sg13g2_fill_1 FILLER_80_666 ();
 sg13g2_decap_8 FILLER_80_671 ();
 sg13g2_decap_4 FILLER_80_678 ();
 sg13g2_fill_1 FILLER_80_682 ();
 sg13g2_decap_4 FILLER_80_686 ();
 sg13g2_fill_1 FILLER_80_690 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_fill_2 FILLER_80_735 ();
 sg13g2_fill_1 FILLER_80_737 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_4 FILLER_80_775 ();
 sg13g2_decap_4 FILLER_80_783 ();
 sg13g2_fill_2 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_828 ();
 sg13g2_fill_2 FILLER_80_835 ();
 sg13g2_decap_8 FILLER_80_841 ();
 sg13g2_decap_8 FILLER_80_848 ();
 sg13g2_decap_8 FILLER_80_855 ();
 sg13g2_fill_2 FILLER_80_862 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_4 FILLER_80_910 ();
 sg13g2_fill_1 FILLER_80_914 ();
 sg13g2_decap_8 FILLER_80_923 ();
 sg13g2_decap_8 FILLER_80_930 ();
 sg13g2_decap_8 FILLER_80_937 ();
 sg13g2_decap_8 FILLER_80_944 ();
 sg13g2_decap_8 FILLER_80_951 ();
 sg13g2_fill_1 FILLER_80_958 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_977 ();
 sg13g2_decap_8 FILLER_80_984 ();
 sg13g2_fill_1 FILLER_80_991 ();
 sg13g2_decap_8 FILLER_80_1018 ();
 sg13g2_fill_1 FILLER_80_1025 ();
 sg13g2_decap_4 FILLER_80_1030 ();
 sg13g2_fill_2 FILLER_80_1034 ();
 sg13g2_decap_8 FILLER_80_1062 ();
 sg13g2_decap_8 FILLER_80_1069 ();
 sg13g2_decap_8 FILLER_80_1076 ();
 sg13g2_decap_8 FILLER_80_1083 ();
 sg13g2_decap_8 FILLER_80_1090 ();
 sg13g2_decap_4 FILLER_80_1101 ();
 sg13g2_fill_1 FILLER_80_1105 ();
 sg13g2_decap_8 FILLER_80_1119 ();
 sg13g2_decap_8 FILLER_80_1126 ();
 sg13g2_decap_8 FILLER_80_1133 ();
 sg13g2_decap_8 FILLER_80_1140 ();
 sg13g2_decap_8 FILLER_80_1147 ();
 sg13g2_decap_8 FILLER_80_1158 ();
 sg13g2_decap_8 FILLER_80_1165 ();
 sg13g2_decap_8 FILLER_80_1172 ();
 sg13g2_decap_8 FILLER_80_1179 ();
 sg13g2_decap_8 FILLER_80_1186 ();
 sg13g2_fill_2 FILLER_80_1193 ();
 sg13g2_fill_1 FILLER_80_1195 ();
 sg13g2_decap_8 FILLER_80_1200 ();
 sg13g2_decap_8 FILLER_80_1207 ();
 sg13g2_decap_8 FILLER_80_1214 ();
 sg13g2_decap_8 FILLER_80_1221 ();
 sg13g2_fill_2 FILLER_80_1228 ();
 sg13g2_decap_8 FILLER_80_1234 ();
 sg13g2_decap_8 FILLER_80_1241 ();
 sg13g2_decap_8 FILLER_80_1248 ();
 sg13g2_decap_8 FILLER_80_1255 ();
 sg13g2_decap_8 FILLER_80_1262 ();
 sg13g2_decap_8 FILLER_80_1269 ();
 sg13g2_decap_8 FILLER_80_1276 ();
 sg13g2_decap_8 FILLER_80_1283 ();
 sg13g2_decap_8 FILLER_80_1290 ();
 sg13g2_fill_1 FILLER_80_1297 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_8 FILLER_80_1310 ();
 sg13g2_fill_1 FILLER_80_1317 ();
 sg13g2_fill_1 FILLER_80_1323 ();
 sg13g2_decap_8 FILLER_80_1329 ();
 sg13g2_decap_8 FILLER_80_1336 ();
 sg13g2_decap_8 FILLER_80_1343 ();
 sg13g2_decap_8 FILLER_80_1350 ();
 sg13g2_decap_8 FILLER_80_1357 ();
 sg13g2_decap_8 FILLER_80_1364 ();
 sg13g2_decap_8 FILLER_80_1371 ();
 sg13g2_decap_4 FILLER_80_1378 ();
 sg13g2_fill_2 FILLER_80_1382 ();
 sg13g2_decap_8 FILLER_80_1388 ();
 sg13g2_decap_8 FILLER_80_1395 ();
 sg13g2_decap_4 FILLER_80_1402 ();
 sg13g2_fill_1 FILLER_80_1406 ();
 sg13g2_decap_8 FILLER_80_1412 ();
 sg13g2_decap_8 FILLER_80_1419 ();
 sg13g2_decap_8 FILLER_80_1426 ();
 sg13g2_decap_8 FILLER_80_1433 ();
 sg13g2_decap_8 FILLER_80_1440 ();
 sg13g2_decap_8 FILLER_80_1447 ();
 sg13g2_decap_8 FILLER_80_1454 ();
 sg13g2_decap_4 FILLER_80_1461 ();
 sg13g2_fill_2 FILLER_80_1465 ();
 sg13g2_decap_8 FILLER_80_1493 ();
 sg13g2_decap_8 FILLER_80_1500 ();
 sg13g2_decap_8 FILLER_80_1507 ();
 sg13g2_decap_8 FILLER_80_1514 ();
 sg13g2_decap_8 FILLER_80_1521 ();
 sg13g2_decap_8 FILLER_80_1528 ();
 sg13g2_decap_8 FILLER_80_1535 ();
 sg13g2_decap_8 FILLER_80_1542 ();
 sg13g2_decap_8 FILLER_80_1549 ();
 sg13g2_fill_2 FILLER_80_1556 ();
 sg13g2_fill_1 FILLER_80_1558 ();
 sg13g2_decap_8 FILLER_80_1563 ();
 sg13g2_fill_2 FILLER_80_1574 ();
 sg13g2_decap_4 FILLER_80_1580 ();
 sg13g2_decap_8 FILLER_80_1588 ();
 sg13g2_fill_1 FILLER_80_1595 ();
 sg13g2_decap_8 FILLER_80_1600 ();
 sg13g2_decap_8 FILLER_80_1607 ();
 sg13g2_decap_8 FILLER_80_1614 ();
 sg13g2_decap_8 FILLER_80_1621 ();
 sg13g2_decap_8 FILLER_80_1628 ();
 sg13g2_decap_8 FILLER_80_1635 ();
 sg13g2_decap_8 FILLER_80_1642 ();
 sg13g2_decap_8 FILLER_80_1649 ();
 sg13g2_decap_8 FILLER_80_1656 ();
 sg13g2_decap_8 FILLER_80_1663 ();
 sg13g2_decap_4 FILLER_80_1670 ();
 sg13g2_fill_2 FILLER_80_1674 ();
 sg13g2_fill_1 FILLER_80_1681 ();
 sg13g2_decap_8 FILLER_80_1690 ();
 sg13g2_fill_1 FILLER_80_1697 ();
 sg13g2_decap_8 FILLER_80_1702 ();
 sg13g2_decap_8 FILLER_80_1709 ();
 sg13g2_decap_8 FILLER_80_1716 ();
 sg13g2_decap_8 FILLER_80_1723 ();
 sg13g2_decap_8 FILLER_80_1730 ();
 sg13g2_decap_8 FILLER_80_1737 ();
 sg13g2_decap_8 FILLER_80_1744 ();
 sg13g2_decap_8 FILLER_80_1751 ();
 sg13g2_decap_8 FILLER_80_1758 ();
 sg13g2_decap_8 FILLER_80_1765 ();
 sg13g2_decap_8 FILLER_80_1772 ();
 sg13g2_decap_8 FILLER_80_1779 ();
 sg13g2_decap_8 FILLER_80_1786 ();
 sg13g2_decap_4 FILLER_80_1793 ();
 sg13g2_fill_2 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1815 ();
 sg13g2_decap_8 FILLER_80_1827 ();
 sg13g2_decap_8 FILLER_80_1834 ();
 sg13g2_decap_8 FILLER_80_1841 ();
 sg13g2_decap_8 FILLER_80_1848 ();
 sg13g2_decap_8 FILLER_80_1855 ();
 sg13g2_decap_4 FILLER_80_1862 ();
 sg13g2_fill_2 FILLER_80_1866 ();
 sg13g2_decap_8 FILLER_80_1872 ();
 sg13g2_decap_8 FILLER_80_1879 ();
 sg13g2_decap_8 FILLER_80_1886 ();
 sg13g2_decap_8 FILLER_80_1893 ();
 sg13g2_decap_8 FILLER_80_1900 ();
 sg13g2_decap_8 FILLER_80_1907 ();
 sg13g2_decap_8 FILLER_80_1914 ();
 sg13g2_decap_8 FILLER_80_1921 ();
 sg13g2_decap_8 FILLER_80_1928 ();
 sg13g2_decap_8 FILLER_80_1935 ();
 sg13g2_decap_4 FILLER_80_1942 ();
 sg13g2_fill_1 FILLER_80_1946 ();
 sg13g2_decap_8 FILLER_80_1951 ();
 sg13g2_decap_8 FILLER_80_1958 ();
 sg13g2_decap_8 FILLER_80_1965 ();
 sg13g2_decap_8 FILLER_80_1972 ();
 sg13g2_fill_2 FILLER_80_1979 ();
 sg13g2_decap_8 FILLER_80_1989 ();
 sg13g2_fill_2 FILLER_80_1996 ();
 sg13g2_fill_1 FILLER_80_1998 ();
 sg13g2_fill_2 FILLER_80_2009 ();
 sg13g2_fill_1 FILLER_80_2011 ();
 sg13g2_decap_8 FILLER_80_2016 ();
 sg13g2_decap_8 FILLER_80_2023 ();
 sg13g2_decap_8 FILLER_80_2030 ();
 sg13g2_decap_4 FILLER_80_2037 ();
 sg13g2_fill_1 FILLER_80_2041 ();
 sg13g2_decap_8 FILLER_80_2060 ();
 sg13g2_fill_1 FILLER_80_2067 ();
 sg13g2_decap_8 FILLER_80_2072 ();
 sg13g2_decap_8 FILLER_80_2079 ();
 sg13g2_fill_2 FILLER_80_2086 ();
 sg13g2_decap_8 FILLER_80_2124 ();
 sg13g2_decap_8 FILLER_80_2131 ();
 sg13g2_decap_8 FILLER_80_2138 ();
 sg13g2_decap_4 FILLER_80_2145 ();
 sg13g2_fill_2 FILLER_80_2149 ();
 sg13g2_decap_4 FILLER_80_2175 ();
 sg13g2_fill_1 FILLER_80_2179 ();
 sg13g2_decap_8 FILLER_80_2184 ();
 sg13g2_decap_8 FILLER_80_2191 ();
 sg13g2_decap_8 FILLER_80_2198 ();
 sg13g2_fill_2 FILLER_80_2205 ();
 sg13g2_decap_4 FILLER_80_2211 ();
 sg13g2_fill_1 FILLER_80_2215 ();
 sg13g2_decap_8 FILLER_80_2230 ();
 sg13g2_decap_8 FILLER_80_2237 ();
 sg13g2_decap_8 FILLER_80_2244 ();
 sg13g2_decap_8 FILLER_80_2251 ();
 sg13g2_decap_8 FILLER_80_2268 ();
 sg13g2_decap_8 FILLER_80_2275 ();
 sg13g2_decap_8 FILLER_80_2282 ();
 sg13g2_decap_8 FILLER_80_2289 ();
 sg13g2_decap_8 FILLER_80_2296 ();
 sg13g2_fill_2 FILLER_80_2311 ();
 sg13g2_fill_1 FILLER_80_2313 ();
 sg13g2_decap_8 FILLER_80_2318 ();
 sg13g2_decap_4 FILLER_80_2325 ();
 sg13g2_fill_1 FILLER_80_2329 ();
 sg13g2_fill_2 FILLER_80_2334 ();
 sg13g2_fill_1 FILLER_80_2336 ();
 sg13g2_fill_2 FILLER_80_2341 ();
 sg13g2_fill_1 FILLER_80_2343 ();
 sg13g2_decap_8 FILLER_80_2348 ();
 sg13g2_decap_8 FILLER_80_2355 ();
 sg13g2_decap_8 FILLER_80_2362 ();
 sg13g2_decap_4 FILLER_80_2373 ();
 sg13g2_fill_1 FILLER_80_2377 ();
 sg13g2_decap_4 FILLER_80_2382 ();
 sg13g2_fill_1 FILLER_80_2386 ();
 sg13g2_decap_8 FILLER_80_2391 ();
 sg13g2_decap_8 FILLER_80_2398 ();
 sg13g2_decap_8 FILLER_80_2405 ();
 sg13g2_decap_8 FILLER_80_2412 ();
 sg13g2_decap_8 FILLER_80_2419 ();
 sg13g2_decap_8 FILLER_80_2426 ();
 sg13g2_decap_4 FILLER_80_2433 ();
 sg13g2_fill_2 FILLER_80_2437 ();
 sg13g2_decap_4 FILLER_80_2456 ();
 sg13g2_fill_1 FILLER_80_2460 ();
 sg13g2_fill_1 FILLER_80_2466 ();
 sg13g2_fill_2 FILLER_80_2479 ();
 sg13g2_decap_8 FILLER_80_2485 ();
 sg13g2_decap_8 FILLER_80_2492 ();
 sg13g2_decap_8 FILLER_80_2499 ();
 sg13g2_decap_8 FILLER_80_2506 ();
 sg13g2_decap_8 FILLER_80_2513 ();
 sg13g2_fill_1 FILLER_80_2520 ();
 sg13g2_fill_2 FILLER_80_2529 ();
 sg13g2_fill_1 FILLER_80_2531 ();
 sg13g2_decap_4 FILLER_80_2541 ();
 sg13g2_fill_2 FILLER_80_2549 ();
 sg13g2_fill_1 FILLER_80_2551 ();
 sg13g2_decap_8 FILLER_80_2556 ();
 sg13g2_decap_8 FILLER_80_2563 ();
 sg13g2_decap_8 FILLER_80_2570 ();
 sg13g2_fill_1 FILLER_80_2577 ();
 sg13g2_decap_8 FILLER_80_2586 ();
 sg13g2_decap_4 FILLER_80_2593 ();
 sg13g2_decap_8 FILLER_80_2601 ();
 sg13g2_fill_2 FILLER_80_2608 ();
 sg13g2_fill_1 FILLER_80_2610 ();
 sg13g2_fill_2 FILLER_80_2615 ();
 sg13g2_decap_8 FILLER_80_2621 ();
 sg13g2_decap_8 FILLER_80_2628 ();
 sg13g2_decap_8 FILLER_80_2635 ();
 sg13g2_decap_8 FILLER_80_2642 ();
 sg13g2_decap_8 FILLER_80_2649 ();
 sg13g2_decap_8 FILLER_80_2656 ();
 sg13g2_decap_8 FILLER_80_2663 ();
endmodule
