module tt_um_rebeccargb_vga_pride (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire clknet_0_clk;
 wire net333;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire counter_clk;
 wire \flag.flag_abrosexual_inst.pix_x[0] ;
 wire \flag.flag_abrosexual_inst.pix_x[1] ;
 wire \flag.flag_abrosexual_inst.pix_x[2] ;
 wire \flag.flag_abrosexual_inst.pix_x[3] ;
 wire \flag.flag_abrosexual_inst.pix_x[4] ;
 wire \flag.flag_abrosexual_inst.pix_x[5] ;
 wire \flag.flag_abrosexual_inst.pix_x[6] ;
 wire \flag.flag_abrosexual_inst.pix_x[7] ;
 wire \flag.flag_abrosexual_inst.pix_x[8] ;
 wire \flag.flag_abrosexual_inst.pix_x[9] ;
 wire \flag.flag_abrosexual_inst.pix_y[0] ;
 wire \flag.flag_abrosexual_inst.pix_y[1] ;
 wire \flag.flag_abrosexual_inst.pix_y[2] ;
 wire \flag.flag_abrosexual_inst.pix_y[3] ;
 wire \flag.flag_abrosexual_inst.pix_y[4] ;
 wire \flag.flag_abrosexual_inst.pix_y[5] ;
 wire \flag.flag_abrosexual_inst.pix_y[6] ;
 wire \flag.flag_abrosexual_inst.pix_y[7] ;
 wire \flag.flag_abrosexual_inst.pix_y[8] ;
 wire hsync;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_buf_1 _4603_ (.A(_0002_),
    .X(_4583_));
 sg13g2_buf_1 _4604_ (.A(net316),
    .X(_0051_));
 sg13g2_buf_1 _4605_ (.A(\flag.flag_abrosexual_inst.pix_y[5] ),
    .X(_0062_));
 sg13g2_buf_1 _4606_ (.A(net315),
    .X(_0073_));
 sg13g2_buf_1 _4607_ (.A(_0073_),
    .X(_0084_));
 sg13g2_buf_1 _4608_ (.A(net261),
    .X(_0095_));
 sg13g2_buf_8 _4609_ (.A(\flag.flag_abrosexual_inst.pix_y[1] ),
    .X(_0106_));
 sg13g2_buf_8 _4610_ (.A(_0106_),
    .X(_0117_));
 sg13g2_buf_1 _4611_ (.A(net295),
    .X(_0128_));
 sg13g2_buf_8 _4612_ (.A(\flag.flag_abrosexual_inst.pix_y[0] ),
    .X(_0139_));
 sg13g2_buf_1 _4613_ (.A(_0139_),
    .X(_0150_));
 sg13g2_buf_1 _4614_ (.A(net294),
    .X(_0161_));
 sg13g2_buf_1 _4615_ (.A(net259),
    .X(_0172_));
 sg13g2_buf_1 _4616_ (.A(net223),
    .X(_0183_));
 sg13g2_buf_1 _4617_ (.A(net190),
    .X(_0194_));
 sg13g2_nand2_2 _4618_ (.Y(_0205_),
    .A(net260),
    .B(net170));
 sg13g2_buf_1 _4619_ (.A(\flag.flag_abrosexual_inst.pix_y[2] ),
    .X(_0216_));
 sg13g2_buf_1 _4620_ (.A(_0216_),
    .X(_0227_));
 sg13g2_buf_8 _4621_ (.A(\flag.flag_abrosexual_inst.pix_y[3] ),
    .X(_0238_));
 sg13g2_nor2b_1 _4622_ (.A(net293),
    .B_N(_0238_),
    .Y(_0249_));
 sg13g2_buf_1 _4623_ (.A(_0249_),
    .X(_0260_));
 sg13g2_nand3_1 _4624_ (.B(_0205_),
    .C(_0260_),
    .A(net224),
    .Y(_0271_));
 sg13g2_nand2b_1 _4625_ (.Y(_0282_),
    .B(_0271_),
    .A_N(net297));
 sg13g2_buf_8 _4626_ (.A(\flag.flag_abrosexual_inst.pix_y[7] ),
    .X(_0293_));
 sg13g2_buf_1 _4627_ (.A(_0293_),
    .X(_0304_));
 sg13g2_buf_1 _4628_ (.A(_0304_),
    .X(_0315_));
 sg13g2_buf_8 _4629_ (.A(\flag.flag_abrosexual_inst.pix_y[6] ),
    .X(_0326_));
 sg13g2_buf_1 _4630_ (.A(_0326_),
    .X(_0337_));
 sg13g2_buf_1 _4631_ (.A(net291),
    .X(_0348_));
 sg13g2_buf_1 _4632_ (.A(net257),
    .X(_0359_));
 sg13g2_buf_1 _4633_ (.A(_0359_),
    .X(_0370_));
 sg13g2_buf_8 _4634_ (.A(\flag.flag_abrosexual_inst.pix_y[8] ),
    .X(_0381_));
 sg13g2_buf_1 _4635_ (.A(net313),
    .X(_0392_));
 sg13g2_buf_1 _4636_ (.A(net290),
    .X(_0403_));
 sg13g2_buf_1 _4637_ (.A(net256),
    .X(_0414_));
 sg13g2_inv_1 _4638_ (.Y(_0425_),
    .A(_0238_));
 sg13g2_buf_1 _4639_ (.A(_0425_),
    .X(_0436_));
 sg13g2_buf_1 _4640_ (.A(net293),
    .X(_0447_));
 sg13g2_buf_1 _4641_ (.A(net254),
    .X(_0458_));
 sg13g2_buf_8 _4642_ (.A(\flag.flag_abrosexual_inst.pix_y[4] ),
    .X(_0469_));
 sg13g2_buf_1 _4643_ (.A(_0469_),
    .X(_0480_));
 sg13g2_nand2b_1 _4644_ (.Y(_0491_),
    .B(net315),
    .A_N(_0480_));
 sg13g2_buf_1 _4645_ (.A(_0491_),
    .X(_0502_));
 sg13g2_nand2b_1 _4646_ (.Y(_0513_),
    .B(net295),
    .A_N(net294));
 sg13g2_buf_2 _4647_ (.A(_0513_),
    .X(_0524_));
 sg13g2_nor4_2 _4648_ (.A(_0436_),
    .B(net220),
    .C(_0502_),
    .Y(_0535_),
    .D(_0524_));
 sg13g2_nand4_1 _4649_ (.B(net189),
    .C(net221),
    .A(net258),
    .Y(_0546_),
    .D(_0535_));
 sg13g2_inv_2 _4650_ (.Y(_0557_),
    .A(_0293_));
 sg13g2_buf_1 _4651_ (.A(_0557_),
    .X(_0568_));
 sg13g2_inv_1 _4652_ (.Y(_0579_),
    .A(net313));
 sg13g2_buf_1 _4653_ (.A(_0579_),
    .X(_0590_));
 sg13g2_nor2_1 _4654_ (.A(net253),
    .B(net252),
    .Y(_0601_));
 sg13g2_buf_1 _4655_ (.A(_0601_),
    .X(_0612_));
 sg13g2_buf_1 _4656_ (.A(net188),
    .X(_0623_));
 sg13g2_and2_1 _4657_ (.A(net261),
    .B(net257),
    .X(_0634_));
 sg13g2_buf_1 _4658_ (.A(_0634_),
    .X(_0645_));
 sg13g2_buf_1 _4659_ (.A(_0238_),
    .X(_0656_));
 sg13g2_buf_1 _4660_ (.A(net288),
    .X(_0667_));
 sg13g2_nand2_1 _4661_ (.Y(_0678_),
    .A(_0667_),
    .B(_0227_));
 sg13g2_buf_1 _4662_ (.A(_0678_),
    .X(_0689_));
 sg13g2_buf_1 _4663_ (.A(net289),
    .X(_0700_));
 sg13g2_buf_1 _4664_ (.A(net250),
    .X(_0711_));
 sg13g2_buf_1 _4665_ (.A(net219),
    .X(_0722_));
 sg13g2_buf_1 _4666_ (.A(\hvsync_gen.vpos[9] ),
    .X(_0733_));
 sg13g2_nor2_1 _4667_ (.A(net186),
    .B(_0733_),
    .Y(_0744_));
 sg13g2_nand4_1 _4668_ (.B(_0645_),
    .C(_0689_),
    .A(net169),
    .Y(_0755_),
    .D(_0744_));
 sg13g2_a21oi_1 _4669_ (.A1(_0282_),
    .A2(_0546_),
    .Y(_0001_),
    .B1(_0755_));
 sg13g2_buf_1 _4670_ (.A(\flag.flag_abrosexual_inst.pix_x[9] ),
    .X(_0776_));
 sg13g2_inv_1 _4671_ (.Y(_0787_),
    .A(net312));
 sg13g2_buf_1 _4672_ (.A(_0787_),
    .X(_0798_));
 sg13g2_buf_8 _4673_ (.A(net249),
    .X(_0809_));
 sg13g2_buf_1 _4674_ (.A(_0004_),
    .X(_0820_));
 sg13g2_buf_1 _4675_ (.A(_0820_),
    .X(_0831_));
 sg13g2_buf_8 _4676_ (.A(\flag.flag_abrosexual_inst.pix_x[8] ),
    .X(_0842_));
 sg13g2_buf_1 _4677_ (.A(net311),
    .X(_0853_));
 sg13g2_buf_1 _4678_ (.A(net286),
    .X(_0864_));
 sg13g2_buf_1 _4679_ (.A(\flag.flag_abrosexual_inst.pix_x[7] ),
    .X(_0875_));
 sg13g2_buf_1 _4680_ (.A(net310),
    .X(_0886_));
 sg13g2_buf_8 _4681_ (.A(\flag.flag_abrosexual_inst.pix_x[6] ),
    .X(_0897_));
 sg13g2_buf_1 _4682_ (.A(_0897_),
    .X(_0908_));
 sg13g2_buf_1 _4683_ (.A(net284),
    .X(_0919_));
 sg13g2_buf_1 _4684_ (.A(net247),
    .X(_0930_));
 sg13g2_nand2_2 _4685_ (.Y(_0941_),
    .A(net285),
    .B(net217));
 sg13g2_buf_8 _4686_ (.A(\flag.flag_abrosexual_inst.pix_x[4] ),
    .X(_0952_));
 sg13g2_buf_1 _4687_ (.A(net309),
    .X(_0963_));
 sg13g2_buf_8 _4688_ (.A(\flag.flag_abrosexual_inst.pix_x[5] ),
    .X(_0974_));
 sg13g2_buf_1 _4689_ (.A(net308),
    .X(_0985_));
 sg13g2_nand2_2 _4690_ (.Y(_0996_),
    .A(net283),
    .B(net282));
 sg13g2_nor2_1 _4691_ (.A(_0941_),
    .B(_0996_),
    .Y(_1007_));
 sg13g2_nor2_1 _4692_ (.A(net248),
    .B(_1007_),
    .Y(_1018_));
 sg13g2_nor2_1 _4693_ (.A(net287),
    .B(_1018_),
    .Y(_1029_));
 sg13g2_buf_1 _4694_ (.A(net285),
    .X(_1040_));
 sg13g2_buf_1 _4695_ (.A(_1040_),
    .X(_1051_));
 sg13g2_inv_1 _4696_ (.Y(_1062_),
    .A(_0897_));
 sg13g2_buf_1 _4697_ (.A(_1062_),
    .X(_1073_));
 sg13g2_buf_1 _4698_ (.A(_0963_),
    .X(_1084_));
 sg13g2_buf_1 _4699_ (.A(net282),
    .X(_1095_));
 sg13g2_nor2_2 _4700_ (.A(net244),
    .B(net243),
    .Y(_1106_));
 sg13g2_nand2_1 _4701_ (.Y(_1117_),
    .A(net245),
    .B(_1106_));
 sg13g2_a21oi_1 _4702_ (.A1(net216),
    .A2(_1117_),
    .Y(_1128_),
    .B1(net248));
 sg13g2_nor3_1 _4703_ (.A(net218),
    .B(_1029_),
    .C(_1128_),
    .Y(_0000_));
 sg13g2_buf_1 _4704_ (.A(net312),
    .X(_1149_));
 sg13g2_nor2_1 _4705_ (.A(net285),
    .B(net217),
    .Y(_1160_));
 sg13g2_nand3_1 _4706_ (.B(net281),
    .C(_1160_),
    .A(net286),
    .Y(_1171_));
 sg13g2_inv_1 _4707_ (.Y(_1182_),
    .A(net308));
 sg13g2_buf_1 _4708_ (.A(net280),
    .X(_1193_));
 sg13g2_buf_1 _4709_ (.A(net244),
    .X(_1204_));
 sg13g2_buf_8 _4710_ (.A(\flag.flag_abrosexual_inst.pix_x[3] ),
    .X(_1215_));
 sg13g2_buf_1 _4711_ (.A(_1215_),
    .X(_1226_));
 sg13g2_inv_1 _4712_ (.Y(_1237_),
    .A(net279));
 sg13g2_buf_1 _4713_ (.A(_1237_),
    .X(_1248_));
 sg13g2_buf_8 _4714_ (.A(\flag.flag_abrosexual_inst.pix_x[2] ),
    .X(_1259_));
 sg13g2_buf_1 _4715_ (.A(_1259_),
    .X(_1270_));
 sg13g2_inv_2 _4716_ (.Y(_1281_),
    .A(net278));
 sg13g2_buf_1 _4717_ (.A(_1281_),
    .X(_1292_));
 sg13g2_nor2_1 _4718_ (.A(net214),
    .B(net213),
    .Y(_1303_));
 sg13g2_buf_2 _4719_ (.A(_1303_),
    .X(_1314_));
 sg13g2_nand2_2 _4720_ (.Y(_1325_),
    .A(net215),
    .B(_1314_));
 sg13g2_buf_2 _4721_ (.A(\flag.flag_abrosexual_inst.pix_x[1] ),
    .X(_1336_));
 sg13g2_buf_8 _4722_ (.A(_1336_),
    .X(_1347_));
 sg13g2_buf_1 _4723_ (.A(net277),
    .X(_1358_));
 sg13g2_buf_1 _4724_ (.A(\flag.flag_abrosexual_inst.pix_x[0] ),
    .X(_1369_));
 sg13g2_buf_1 _4725_ (.A(net307),
    .X(_1380_));
 sg13g2_buf_1 _4726_ (.A(net276),
    .X(_1391_));
 sg13g2_nand2_2 _4727_ (.Y(_1402_),
    .A(net241),
    .B(net240));
 sg13g2_nor2_2 _4728_ (.A(_1325_),
    .B(_1402_),
    .Y(_1413_));
 sg13g2_nand3b_1 _4729_ (.B(net242),
    .C(_1413_),
    .Y(_1424_),
    .A_N(_1171_));
 sg13g2_buf_1 _4730_ (.A(_1424_),
    .X(_1435_));
 sg13g2_buf_1 _4731_ (.A(_0022_),
    .X(_1446_));
 sg13g2_buf_1 _4732_ (.A(net306),
    .X(_1457_));
 sg13g2_buf_1 _4733_ (.A(net275),
    .X(_1468_));
 sg13g2_buf_1 _4734_ (.A(net239),
    .X(_1479_));
 sg13g2_buf_2 _4735_ (.A(rst_n),
    .X(_1490_));
 sg13g2_nor2_1 _4736_ (.A(net295),
    .B(_0139_),
    .Y(_1501_));
 sg13g2_buf_1 _4737_ (.A(_1501_),
    .X(_1512_));
 sg13g2_nor2b_1 _4738_ (.A(net187),
    .B_N(net211),
    .Y(_1523_));
 sg13g2_nor4_1 _4739_ (.A(net261),
    .B(_0722_),
    .C(net292),
    .D(net189),
    .Y(_1534_));
 sg13g2_nand4_1 _4740_ (.B(_0733_),
    .C(_1523_),
    .A(net252),
    .Y(_1545_),
    .D(_1534_));
 sg13g2_nand2_2 _4741_ (.Y(_1556_),
    .A(_1490_),
    .B(_1545_));
 sg13g2_inv_1 _4742_ (.Y(_1567_),
    .A(_1556_));
 sg13g2_nand2_1 _4743_ (.Y(_1578_),
    .A(net212),
    .B(_1567_));
 sg13g2_nand3_1 _4744_ (.B(net170),
    .C(_1435_),
    .A(_1490_),
    .Y(_1589_));
 sg13g2_o21ai_1 _4745_ (.B1(_1589_),
    .Y(_0041_),
    .A1(_1435_),
    .A2(_1578_));
 sg13g2_nand2_1 _4746_ (.Y(_1610_),
    .A(_1490_),
    .B(_1435_));
 sg13g2_nand2_1 _4747_ (.Y(_1621_),
    .A(_1567_),
    .B(_1610_));
 sg13g2_nand2b_1 _4748_ (.Y(_1632_),
    .B(net294),
    .A_N(net295));
 sg13g2_buf_1 _4749_ (.A(_1610_),
    .X(_1643_));
 sg13g2_o21ai_1 _4750_ (.B1(net40),
    .Y(_1654_),
    .A1(net170),
    .A2(_1556_));
 sg13g2_nand2_1 _4751_ (.Y(_1665_),
    .A(net260),
    .B(_1654_));
 sg13g2_o21ai_1 _4752_ (.B1(_1665_),
    .Y(_0042_),
    .A1(_1621_),
    .A2(_1632_));
 sg13g2_inv_2 _4753_ (.Y(_1686_),
    .A(net293));
 sg13g2_buf_1 _4754_ (.A(_1686_),
    .X(_1697_));
 sg13g2_inv_1 _4755_ (.Y(_1708_),
    .A(net260));
 sg13g2_inv_1 _4756_ (.Y(_1719_),
    .A(net294));
 sg13g2_buf_1 _4757_ (.A(_1719_),
    .X(_1730_));
 sg13g2_buf_1 _4758_ (.A(net208),
    .X(_1741_));
 sg13g2_nor2_1 _4759_ (.A(net209),
    .B(net185),
    .Y(_1752_));
 sg13g2_nand2_1 _4760_ (.Y(_1763_),
    .A(net210),
    .B(_1752_));
 sg13g2_o21ai_1 _4761_ (.B1(_1610_),
    .Y(_1774_),
    .A1(_1752_),
    .A2(_1556_));
 sg13g2_nand2_1 _4762_ (.Y(_1785_),
    .A(net220),
    .B(_1774_));
 sg13g2_o21ai_1 _4763_ (.B1(_1785_),
    .Y(_0043_),
    .A1(_1621_),
    .A2(_1763_));
 sg13g2_buf_1 _4764_ (.A(_0667_),
    .X(_1806_));
 sg13g2_nor2_1 _4765_ (.A(net210),
    .B(_0205_),
    .Y(_1817_));
 sg13g2_o21ai_1 _4766_ (.B1(net40),
    .Y(_1828_),
    .A1(_1556_),
    .A2(_1817_));
 sg13g2_nor4_1 _4767_ (.A(net207),
    .B(net210),
    .C(_0205_),
    .D(_1621_),
    .Y(_1839_));
 sg13g2_a21o_1 _4768_ (.A2(_1828_),
    .A1(net207),
    .B1(_1839_),
    .X(_0044_));
 sg13g2_nor2_1 _4769_ (.A(net187),
    .B(_0205_),
    .Y(_1860_));
 sg13g2_o21ai_1 _4770_ (.B1(net40),
    .Y(_1871_),
    .A1(_1556_),
    .A2(_1860_));
 sg13g2_nor4_1 _4771_ (.A(net186),
    .B(net187),
    .C(_0205_),
    .D(_1621_),
    .Y(_1882_));
 sg13g2_a21o_1 _4772_ (.A2(_1871_),
    .A1(net186),
    .B1(_1882_),
    .X(_0045_));
 sg13g2_a21oi_2 _4773_ (.B1(_1567_),
    .Y(_1903_),
    .A2(_1435_),
    .A1(_1490_));
 sg13g2_inv_2 _4774_ (.Y(_1914_),
    .A(net296));
 sg13g2_buf_1 _4775_ (.A(_1914_),
    .X(_1925_));
 sg13g2_nand2_1 _4776_ (.Y(_1936_),
    .A(net186),
    .B(_1860_));
 sg13g2_nand2b_1 _4777_ (.Y(_1947_),
    .B(_1610_),
    .A_N(_1936_));
 sg13g2_buf_1 _4778_ (.A(_1947_),
    .X(_1958_));
 sg13g2_xnor2_1 _4779_ (.Y(_1969_),
    .A(_1925_),
    .B(_1958_));
 sg13g2_nor2_1 _4780_ (.A(_1903_),
    .B(_1969_),
    .Y(_0046_));
 sg13g2_nor2_1 _4781_ (.A(net206),
    .B(_1958_),
    .Y(_1990_));
 sg13g2_xnor2_1 _4782_ (.Y(_2001_),
    .A(net189),
    .B(_1990_));
 sg13g2_nor2_1 _4783_ (.A(_1903_),
    .B(_2001_),
    .Y(_0047_));
 sg13g2_nand2_1 _4784_ (.Y(_2022_),
    .A(net296),
    .B(net257));
 sg13g2_buf_1 _4785_ (.A(_2022_),
    .X(_2033_));
 sg13g2_nor2_1 _4786_ (.A(net184),
    .B(_1958_),
    .Y(_2044_));
 sg13g2_xnor2_1 _4787_ (.Y(_2055_),
    .A(_0315_),
    .B(_2044_));
 sg13g2_nor2_1 _4788_ (.A(_1903_),
    .B(_2055_),
    .Y(_0048_));
 sg13g2_nand3_1 _4789_ (.B(net314),
    .C(_0326_),
    .A(net315),
    .Y(_2076_));
 sg13g2_buf_1 _4790_ (.A(_2076_),
    .X(_2087_));
 sg13g2_nor2_1 _4791_ (.A(_1958_),
    .B(_2087_),
    .Y(_2098_));
 sg13g2_xnor2_1 _4792_ (.Y(_2109_),
    .A(net221),
    .B(_2098_));
 sg13g2_nor2_1 _4793_ (.A(_1903_),
    .B(_2109_),
    .Y(_0049_));
 sg13g2_nand2_1 _4794_ (.Y(_2130_),
    .A(net258),
    .B(net256));
 sg13g2_buf_1 _4795_ (.A(_2130_),
    .X(_2141_));
 sg13g2_nor3_1 _4796_ (.A(net183),
    .B(_2033_),
    .C(_1958_),
    .Y(_2152_));
 sg13g2_xnor2_1 _4797_ (.Y(_2163_),
    .A(_0733_),
    .B(_2152_));
 sg13g2_nor2_1 _4798_ (.A(_1903_),
    .B(_2163_),
    .Y(_0050_));
 sg13g2_buf_1 _4799_ (.A(\counter[0] ),
    .X(_2184_));
 sg13g2_inv_1 _4800_ (.Y(_2195_),
    .A(_2184_));
 sg13g2_buf_2 _4801_ (.A(ui_in[6]),
    .X(_2206_));
 sg13g2_inv_1 _4802_ (.Y(_2217_),
    .A(_2206_));
 sg13g2_buf_2 _4803_ (.A(\counter[5] ),
    .X(_2228_));
 sg13g2_buf_1 _4804_ (.A(\counter[1] ),
    .X(_2239_));
 sg13g2_buf_1 _4805_ (.A(_2239_),
    .X(_2250_));
 sg13g2_buf_2 _4806_ (.A(\counter[2] ),
    .X(_2261_));
 sg13g2_buf_1 _4807_ (.A(\counter[3] ),
    .X(_2272_));
 sg13g2_nor4_1 _4808_ (.A(net205),
    .B(net182),
    .C(_2261_),
    .D(_2272_),
    .Y(_2283_));
 sg13g2_buf_1 _4809_ (.A(\counter[4] ),
    .X(_2294_));
 sg13g2_nor2b_1 _4810_ (.A(_2283_),
    .B_N(_2294_),
    .Y(_2305_));
 sg13g2_buf_2 _4811_ (.A(\counter[6] ),
    .X(_2316_));
 sg13g2_o21ai_1 _4812_ (.B1(_2316_),
    .Y(_2327_),
    .A1(_2228_),
    .A2(_2305_));
 sg13g2_buf_2 _4813_ (.A(ui_in[4]),
    .X(_2338_));
 sg13g2_buf_2 _4814_ (.A(ui_in[5]),
    .X(_2349_));
 sg13g2_nor2_1 _4815_ (.A(_2349_),
    .B(_2206_),
    .Y(_2360_));
 sg13g2_buf_2 _4816_ (.A(_2360_),
    .X(_2371_));
 sg13g2_nand2b_1 _4817_ (.Y(_2382_),
    .B(_2371_),
    .A_N(_2338_));
 sg13g2_buf_1 _4818_ (.A(_2382_),
    .X(_2393_));
 sg13g2_o21ai_1 _4819_ (.B1(_2393_),
    .Y(_2404_),
    .A1(_2217_),
    .A2(_2327_));
 sg13g2_buf_1 _4820_ (.A(uio_in[0]),
    .X(_2415_));
 sg13g2_nor2b_1 _4821_ (.A(_2415_),
    .B_N(_2338_),
    .Y(_2426_));
 sg13g2_buf_2 _4822_ (.A(ui_in[7]),
    .X(_2437_));
 sg13g2_a21oi_1 _4823_ (.A1(_2371_),
    .A2(_2426_),
    .Y(_2448_),
    .B1(_2437_));
 sg13g2_o21ai_1 _4824_ (.B1(_2448_),
    .Y(_2459_),
    .A1(_2195_),
    .A2(_2371_));
 sg13g2_a21oi_1 _4825_ (.A1(_2195_),
    .A2(_2404_),
    .Y(_0024_),
    .B1(_2459_));
 sg13g2_buf_1 _4826_ (.A(uio_in[1]),
    .X(_2480_));
 sg13g2_nand2b_1 _4827_ (.Y(_2491_),
    .B(_2338_),
    .A_N(_2480_));
 sg13g2_inv_1 _4828_ (.Y(_2502_),
    .A(_2327_));
 sg13g2_nor2_1 _4829_ (.A(_2217_),
    .B(_2502_),
    .Y(_2513_));
 sg13g2_buf_2 _4830_ (.A(_2513_),
    .X(_2524_));
 sg13g2_nand2b_1 _4831_ (.Y(_2535_),
    .B(_2239_),
    .A_N(\counter[0] ));
 sg13g2_nand2b_1 _4832_ (.Y(_2546_),
    .B(net205),
    .A_N(_2239_));
 sg13g2_nand2_1 _4833_ (.Y(_2557_),
    .A(_2535_),
    .B(_2546_));
 sg13g2_a22oi_1 _4834_ (.Y(_2568_),
    .B1(_2524_),
    .B2(_2557_),
    .A2(_2491_),
    .A1(_2371_));
 sg13g2_nor3_2 _4835_ (.A(_2349_),
    .B(_2338_),
    .C(_2206_),
    .Y(_2579_));
 sg13g2_a21oi_1 _4836_ (.A1(net205),
    .A2(_2568_),
    .Y(_2590_),
    .B1(_2579_));
 sg13g2_nor2_1 _4837_ (.A(net182),
    .B(_2590_),
    .Y(_2601_));
 sg13g2_inv_1 _4838_ (.Y(_2612_),
    .A(_2349_));
 sg13g2_nand2b_1 _4839_ (.Y(_2623_),
    .B(_2283_),
    .A_N(_2294_));
 sg13g2_buf_1 _4840_ (.A(_2623_),
    .X(_2634_));
 sg13g2_nor3_1 _4841_ (.A(_2228_),
    .B(_2316_),
    .C(_2634_),
    .Y(_2644_));
 sg13g2_nor3_1 _4842_ (.A(_2612_),
    .B(_2206_),
    .C(_2644_),
    .Y(_2655_));
 sg13g2_buf_1 _4843_ (.A(_2655_),
    .X(_2666_));
 sg13g2_inv_1 _4844_ (.Y(_2677_),
    .A(_2568_));
 sg13g2_a21oi_1 _4845_ (.A1(_2535_),
    .A2(net66),
    .Y(_2688_),
    .B1(_2677_));
 sg13g2_nor3_1 _4846_ (.A(_2437_),
    .B(_2601_),
    .C(_2688_),
    .Y(_0025_));
 sg13g2_inv_1 _4847_ (.Y(_2709_),
    .A(_0019_));
 sg13g2_nand2_1 _4848_ (.Y(_2720_),
    .A(_2206_),
    .B(_2327_));
 sg13g2_buf_1 _4849_ (.A(_2720_),
    .X(_2731_));
 sg13g2_nand2_1 _4850_ (.Y(_2742_),
    .A(net182),
    .B(net66));
 sg13g2_o21ai_1 _4851_ (.B1(_2742_),
    .Y(_2753_),
    .A1(net182),
    .A2(_2731_));
 sg13g2_nand2b_1 _4852_ (.Y(_2764_),
    .B(_2338_),
    .A_N(net1));
 sg13g2_nor2b_1 _4853_ (.A(_2250_),
    .B_N(net66),
    .Y(_2775_));
 sg13g2_and2_1 _4854_ (.A(_2250_),
    .B(_2524_),
    .X(_2786_));
 sg13g2_mux4_1 _4855_ (.S0(net205),
    .A0(_2524_),
    .A1(net66),
    .A2(_2775_),
    .A3(_2786_),
    .S1(_0019_),
    .X(_2797_));
 sg13g2_a221oi_1 _4856_ (.B2(_2371_),
    .C1(_2797_),
    .B1(_2764_),
    .A1(_2709_),
    .Y(_2808_),
    .A2(_2753_));
 sg13g2_nor2_1 _4857_ (.A(_2261_),
    .B(_2393_),
    .Y(_2819_));
 sg13g2_nor3_1 _4858_ (.A(_2437_),
    .B(_2808_),
    .C(_2819_),
    .Y(_0026_));
 sg13g2_inv_1 _4859_ (.Y(_2840_),
    .A(_2272_));
 sg13g2_buf_1 _4860_ (.A(_0020_),
    .X(_2851_));
 sg13g2_nor2_1 _4861_ (.A(net182),
    .B(_2261_),
    .Y(_2862_));
 sg13g2_nand3_1 _4862_ (.B(_2862_),
    .C(net66),
    .A(_2851_),
    .Y(_2873_));
 sg13g2_o21ai_1 _4863_ (.B1(_2873_),
    .Y(_2884_),
    .A1(_2851_),
    .A2(_2731_));
 sg13g2_nand2b_1 _4864_ (.Y(_2895_),
    .B(net66),
    .A_N(_2851_));
 sg13g2_nand4_1 _4865_ (.B(_2261_),
    .C(_2851_),
    .A(net182),
    .Y(_2906_),
    .D(_2524_));
 sg13g2_nand3_1 _4866_ (.B(_2895_),
    .C(_2906_),
    .A(net205),
    .Y(_2917_));
 sg13g2_o21ai_1 _4867_ (.B1(_2917_),
    .Y(_2928_),
    .A1(net205),
    .A2(_2884_));
 sg13g2_a21oi_1 _4868_ (.A1(_2862_),
    .A2(_2731_),
    .Y(_2939_),
    .B1(_2851_));
 sg13g2_a21oi_1 _4869_ (.A1(net182),
    .A2(_2261_),
    .Y(_2950_),
    .B1(_2731_));
 sg13g2_or2_1 _4870_ (.X(_2961_),
    .B(_2950_),
    .A(net66));
 sg13g2_inv_1 _4871_ (.Y(_2972_),
    .A(net2));
 sg13g2_nand2_1 _4872_ (.Y(_2983_),
    .A(_2338_),
    .B(_2972_));
 sg13g2_a22oi_1 _4873_ (.Y(_2994_),
    .B1(_2983_),
    .B2(_2371_),
    .A2(_2961_),
    .A1(_2939_));
 sg13g2_a221oi_1 _4874_ (.B2(_2994_),
    .C1(_2437_),
    .B1(_2928_),
    .A1(_2840_),
    .Y(_0027_),
    .A2(_2579_));
 sg13g2_nand3b_1 _4875_ (.B(_2634_),
    .C(_2349_),
    .Y(_3015_),
    .A_N(_2305_));
 sg13g2_o21ai_1 _4876_ (.B1(_3015_),
    .Y(_3026_),
    .A1(_2349_),
    .A2(net3));
 sg13g2_and4_1 _4877_ (.A(_2184_),
    .B(net182),
    .C(_2261_),
    .D(_2272_),
    .X(_3037_));
 sg13g2_buf_1 _4878_ (.A(_3037_),
    .X(_3048_));
 sg13g2_nand3b_1 _4879_ (.B(_2524_),
    .C(_3048_),
    .Y(_3059_),
    .A_N(_2294_));
 sg13g2_o21ai_1 _4880_ (.B1(_3059_),
    .Y(_3070_),
    .A1(_2206_),
    .A2(_3026_));
 sg13g2_o21ai_1 _4881_ (.B1(_2393_),
    .Y(_3081_),
    .A1(_2731_),
    .A2(_3048_));
 sg13g2_a22oi_1 _4882_ (.Y(_3092_),
    .B1(_3081_),
    .B2(_2294_),
    .A2(_3070_),
    .A1(_2393_));
 sg13g2_nor2_1 _4883_ (.A(_2437_),
    .B(_3092_),
    .Y(_0028_));
 sg13g2_nand2b_1 _4884_ (.Y(_3113_),
    .B(_2338_),
    .A_N(net4));
 sg13g2_inv_1 _4885_ (.Y(_3124_),
    .A(_2634_));
 sg13g2_and2_1 _4886_ (.A(_2294_),
    .B(_3048_),
    .X(_3135_));
 sg13g2_buf_1 _4887_ (.A(_3135_),
    .X(_3146_));
 sg13g2_a22oi_1 _4888_ (.Y(_3157_),
    .B1(_3146_),
    .B2(_2524_),
    .A2(net66),
    .A1(_3124_));
 sg13g2_inv_1 _4889_ (.Y(_3168_),
    .A(_3146_));
 sg13g2_a221oi_1 _4890_ (.B2(_2524_),
    .C1(_0021_),
    .B1(_3168_),
    .A1(_2634_),
    .Y(_3179_),
    .A2(_2666_));
 sg13g2_a21oi_1 _4891_ (.A1(_0021_),
    .A2(_3157_),
    .Y(_3190_),
    .B1(_3179_));
 sg13g2_a21oi_1 _4892_ (.A1(_2371_),
    .A2(_3113_),
    .Y(_3201_),
    .B1(_3190_));
 sg13g2_nor2_1 _4893_ (.A(_2228_),
    .B(_2393_),
    .Y(_3212_));
 sg13g2_nor3_1 _4894_ (.A(_2437_),
    .B(_3201_),
    .C(_3212_),
    .Y(_0029_));
 sg13g2_inv_1 _4895_ (.Y(_3233_),
    .A(_2316_));
 sg13g2_nand4_1 _4896_ (.B(_2228_),
    .C(_3233_),
    .A(_2206_),
    .Y(_3244_),
    .D(_3146_));
 sg13g2_and2_1 _4897_ (.A(_2228_),
    .B(_3146_),
    .X(_3255_));
 sg13g2_o21ai_1 _4898_ (.B1(_2393_),
    .Y(_3266_),
    .A1(_2731_),
    .A2(_3255_));
 sg13g2_o21ai_1 _4899_ (.B1(_2316_),
    .Y(_3277_),
    .A1(_2228_),
    .A2(_2634_));
 sg13g2_nor2b_1 _4900_ (.A(_2644_),
    .B_N(_3277_),
    .Y(_3288_));
 sg13g2_a21oi_1 _4901_ (.A1(_2338_),
    .A2(net5),
    .Y(_3299_),
    .B1(_2349_));
 sg13g2_a21oi_1 _4902_ (.A1(_2349_),
    .A2(_3288_),
    .Y(_3310_),
    .B1(_3299_));
 sg13g2_a22oi_1 _4903_ (.Y(_3321_),
    .B1(_3310_),
    .B2(_2217_),
    .A2(_3266_),
    .A1(_2316_));
 sg13g2_a21oi_1 _4904_ (.A1(_3244_),
    .A2(_3321_),
    .Y(_0030_),
    .B1(_2437_));
 sg13g2_buf_2 _4905_ (.A(_0023_),
    .X(_3342_));
 sg13g2_inv_1 _4906_ (.Y(_3353_),
    .A(_3342_));
 sg13g2_buf_1 _4907_ (.A(net274),
    .X(_3364_));
 sg13g2_nor2_1 _4908_ (.A(net238),
    .B(net40),
    .Y(_0031_));
 sg13g2_inv_1 _4909_ (.Y(_3384_),
    .A(_1490_));
 sg13g2_nor2b_1 _4910_ (.A(net277),
    .B_N(_1369_),
    .Y(_3395_));
 sg13g2_nor2b_1 _4911_ (.A(net307),
    .B_N(net277),
    .Y(_3406_));
 sg13g2_nor2_1 _4912_ (.A(_3395_),
    .B(_3406_),
    .Y(_3417_));
 sg13g2_nor2_1 _4913_ (.A(_3384_),
    .B(_3417_),
    .Y(_0032_));
 sg13g2_buf_1 _4914_ (.A(net278),
    .X(_3438_));
 sg13g2_buf_1 _4915_ (.A(net237),
    .X(_3449_));
 sg13g2_buf_1 _4916_ (.A(net204),
    .X(_3460_));
 sg13g2_buf_1 _4917_ (.A(net181),
    .X(_3471_));
 sg13g2_buf_1 _4918_ (.A(net168),
    .X(_3482_));
 sg13g2_nand2_1 _4919_ (.Y(_3492_),
    .A(net160),
    .B(_1402_));
 sg13g2_buf_1 _4920_ (.A(net240),
    .X(_3503_));
 sg13g2_buf_1 _4921_ (.A(net241),
    .X(_3514_));
 sg13g2_nand3b_1 _4922_ (.B(net203),
    .C(_3514_),
    .Y(_3525_),
    .A_N(net204));
 sg13g2_a21oi_1 _4923_ (.A1(_3492_),
    .A2(_3525_),
    .Y(_0033_),
    .B1(net40));
 sg13g2_buf_1 _4924_ (.A(_1226_),
    .X(_3546_));
 sg13g2_buf_1 _4925_ (.A(_3546_),
    .X(_3557_));
 sg13g2_buf_1 _4926_ (.A(net201),
    .X(_3568_));
 sg13g2_buf_1 _4927_ (.A(_3342_),
    .X(_3579_));
 sg13g2_buf_1 _4928_ (.A(_3579_),
    .X(_3590_));
 sg13g2_nand2_1 _4929_ (.Y(_3601_),
    .A(net241),
    .B(net278));
 sg13g2_nor2_1 _4930_ (.A(net235),
    .B(_3601_),
    .Y(_3612_));
 sg13g2_xnor2_1 _4931_ (.Y(_3623_),
    .A(_3568_),
    .B(_3612_));
 sg13g2_nor2_1 _4932_ (.A(net40),
    .B(_3623_),
    .Y(_0034_));
 sg13g2_inv_1 _4933_ (.Y(_3644_),
    .A(net283));
 sg13g2_nand2_2 _4934_ (.Y(_3655_),
    .A(net279),
    .B(net237));
 sg13g2_and2_1 _4935_ (.A(net241),
    .B(net276),
    .X(_3666_));
 sg13g2_buf_1 _4936_ (.A(_3666_),
    .X(_3677_));
 sg13g2_nand2b_1 _4937_ (.Y(_3688_),
    .B(_3677_),
    .A_N(_3655_));
 sg13g2_and2_1 _4938_ (.A(_3644_),
    .B(_3688_),
    .X(_3699_));
 sg13g2_nor3_1 _4939_ (.A(_3384_),
    .B(_1413_),
    .C(_3699_),
    .Y(_0035_));
 sg13g2_buf_1 _4940_ (.A(net243),
    .X(_3720_));
 sg13g2_buf_1 _4941_ (.A(net200),
    .X(_3731_));
 sg13g2_xnor2_1 _4942_ (.Y(_3742_),
    .A(net179),
    .B(_1413_));
 sg13g2_nor2_1 _4943_ (.A(net40),
    .B(_3742_),
    .Y(_0036_));
 sg13g2_nand2_1 _4944_ (.Y(_3763_),
    .A(net179),
    .B(_1413_));
 sg13g2_xnor2_1 _4945_ (.Y(_3774_),
    .A(net245),
    .B(_3763_));
 sg13g2_nor2_1 _4946_ (.A(_3384_),
    .B(_3774_),
    .Y(_0037_));
 sg13g2_inv_1 _4947_ (.Y(_3794_),
    .A(net277));
 sg13g2_buf_1 _4948_ (.A(_3794_),
    .X(_3805_));
 sg13g2_buf_1 _4949_ (.A(net199),
    .X(_3816_));
 sg13g2_nand2_1 _4950_ (.Y(_3827_),
    .A(net282),
    .B(net284));
 sg13g2_nor4_1 _4951_ (.A(net178),
    .B(net235),
    .C(_1325_),
    .D(_3827_),
    .Y(_3838_));
 sg13g2_xnor2_1 _4952_ (.Y(_3849_),
    .A(_1051_),
    .B(_3838_));
 sg13g2_nor2_1 _4953_ (.A(_1643_),
    .B(_3849_),
    .Y(_0038_));
 sg13g2_inv_2 _4954_ (.Y(_3870_),
    .A(_0842_));
 sg13g2_buf_1 _4955_ (.A(_3870_),
    .X(_3881_));
 sg13g2_or2_1 _4956_ (.X(_3892_),
    .B(_3763_),
    .A(_0941_));
 sg13g2_xnor2_1 _4957_ (.Y(_3903_),
    .A(net234),
    .B(_3892_));
 sg13g2_nor2_1 _4958_ (.A(_1643_),
    .B(_3903_),
    .Y(_0039_));
 sg13g2_or2_1 _4959_ (.X(_3924_),
    .B(_3892_),
    .A(net234));
 sg13g2_xnor2_1 _4960_ (.Y(_3935_),
    .A(net218),
    .B(_3924_));
 sg13g2_nor2_1 _4961_ (.A(net40),
    .B(_3935_),
    .Y(_0040_));
 sg13g2_nand2b_2 _4962_ (.Y(counter_clk),
    .B(_2579_),
    .A_N(_2437_));
 sg13g2_buf_1 _4963_ (.A(_0009_),
    .X(_3965_));
 sg13g2_inv_2 _4964_ (.Y(_3976_),
    .A(_3965_));
 sg13g2_and3_1 _4965_ (.X(_3987_),
    .A(net315),
    .B(net314),
    .C(_0326_));
 sg13g2_buf_1 _4966_ (.A(_3987_),
    .X(_3998_));
 sg13g2_a21oi_1 _4967_ (.A1(_3976_),
    .A2(_3998_),
    .Y(_4009_),
    .B1(net313));
 sg13g2_inv_1 _4968_ (.Y(_4020_),
    .A(_0469_));
 sg13g2_or2_1 _4969_ (.X(_4031_),
    .B(_0216_),
    .A(_0106_));
 sg13g2_buf_2 _4970_ (.A(_4031_),
    .X(_4042_));
 sg13g2_nand2b_1 _4971_ (.Y(_4053_),
    .B(_1446_),
    .A_N(_0238_));
 sg13g2_nor4_1 _4972_ (.A(_4020_),
    .B(net313),
    .C(_4042_),
    .D(_4053_),
    .Y(_4061_));
 sg13g2_and2_1 _4973_ (.A(net315),
    .B(_0469_),
    .X(_4062_));
 sg13g2_buf_1 _4974_ (.A(_4062_),
    .X(_4063_));
 sg13g2_nor4_1 _4975_ (.A(_0106_),
    .B(_0139_),
    .C(_0238_),
    .D(_0216_),
    .Y(_4064_));
 sg13g2_buf_2 _4976_ (.A(_4064_),
    .X(_4065_));
 sg13g2_buf_1 _4977_ (.A(_0005_),
    .X(_4066_));
 sg13g2_and3_1 _4978_ (.X(_4067_),
    .A(net314),
    .B(_0326_),
    .C(_4066_));
 sg13g2_buf_1 _4979_ (.A(_4067_),
    .X(_4068_));
 sg13g2_nand3_1 _4980_ (.B(_4065_),
    .C(_4068_),
    .A(_4063_),
    .Y(_4069_));
 sg13g2_o21ai_1 _4981_ (.B1(_4069_),
    .Y(_4070_),
    .A1(_4009_),
    .A2(_4061_));
 sg13g2_buf_8 _4982_ (.A(_4070_),
    .X(_4071_));
 sg13g2_buf_1 _4983_ (.A(net167),
    .X(_4072_));
 sg13g2_buf_1 _4984_ (.A(_0010_),
    .X(_4073_));
 sg13g2_inv_1 _4985_ (.Y(_4074_),
    .A(_4073_));
 sg13g2_nand3_1 _4986_ (.B(_0469_),
    .C(net291),
    .A(net315),
    .Y(_4075_));
 sg13g2_xnor2_1 _4987_ (.Y(_4076_),
    .A(_4074_),
    .B(_4075_));
 sg13g2_buf_1 _4988_ (.A(_4076_),
    .X(_4077_));
 sg13g2_buf_1 _4989_ (.A(_3965_),
    .X(_4078_));
 sg13g2_o21ai_1 _4990_ (.B1(_0579_),
    .Y(_4079_),
    .A1(net272),
    .A2(_2087_));
 sg13g2_buf_8 _4991_ (.A(_4079_),
    .X(_4080_));
 sg13g2_nor2_1 _4992_ (.A(_0106_),
    .B(_0216_),
    .Y(_4081_));
 sg13g2_buf_2 _4993_ (.A(_4081_),
    .X(_4082_));
 sg13g2_nor2b_1 _4994_ (.A(_0238_),
    .B_N(net306),
    .Y(_4083_));
 sg13g2_nor2b_1 _4995_ (.A(net313),
    .B_N(_0469_),
    .Y(_4084_));
 sg13g2_nand3_1 _4996_ (.B(_4083_),
    .C(_4084_),
    .A(_4082_),
    .Y(_4085_));
 sg13g2_buf_2 _4997_ (.A(_4085_),
    .X(_4086_));
 sg13g2_buf_8 _4998_ (.A(_4063_),
    .X(_4087_));
 sg13g2_or4_1 _4999_ (.A(_0106_),
    .B(_0139_),
    .C(_0238_),
    .D(_0216_),
    .X(_4088_));
 sg13g2_buf_2 _5000_ (.A(_4088_),
    .X(_4089_));
 sg13g2_nand3_1 _5001_ (.B(_0326_),
    .C(_4066_),
    .A(net314),
    .Y(_4090_));
 sg13g2_buf_1 _5002_ (.A(_4090_),
    .X(_4091_));
 sg13g2_nor2_1 _5003_ (.A(_4089_),
    .B(_4091_),
    .Y(_4092_));
 sg13g2_buf_8 _5004_ (.A(_4092_),
    .X(_4093_));
 sg13g2_a22oi_1 _5005_ (.Y(_4094_),
    .B1(net198),
    .B2(_4093_),
    .A2(_4086_),
    .A1(_4080_));
 sg13g2_buf_2 _5006_ (.A(_4094_),
    .X(_4095_));
 sg13g2_buf_8 _5007_ (.A(_4095_),
    .X(_4096_));
 sg13g2_buf_1 _5008_ (.A(net148),
    .X(_4097_));
 sg13g2_nor2_2 _5009_ (.A(_4042_),
    .B(_4053_),
    .Y(_4098_));
 sg13g2_nor2_1 _5010_ (.A(_4020_),
    .B(_0557_),
    .Y(_4099_));
 sg13g2_nand3b_1 _5011_ (.B(_0337_),
    .C(net315),
    .Y(_4100_),
    .A_N(net272));
 sg13g2_nor2_1 _5012_ (.A(net314),
    .B(_4100_),
    .Y(_4101_));
 sg13g2_nand3_1 _5013_ (.B(_4082_),
    .C(_4083_),
    .A(_0480_),
    .Y(_4102_));
 sg13g2_and2_1 _5014_ (.A(net314),
    .B(_4100_),
    .X(_4103_));
 sg13g2_a221oi_1 _5015_ (.B2(_4102_),
    .C1(_4103_),
    .B1(_4101_),
    .A1(_4098_),
    .Y(_4104_),
    .A2(_4099_));
 sg13g2_buf_2 _5016_ (.A(_4104_),
    .X(_4105_));
 sg13g2_and2_1 _5017_ (.A(net130),
    .B(_4105_),
    .X(_4106_));
 sg13g2_a21oi_1 _5018_ (.A1(net159),
    .A2(_4077_),
    .Y(_4107_),
    .B1(_4106_));
 sg13g2_buf_2 _5019_ (.A(_4107_),
    .X(_4108_));
 sg13g2_nor2_1 _5020_ (.A(_1336_),
    .B(net307),
    .Y(_4109_));
 sg13g2_buf_2 _5021_ (.A(_4109_),
    .X(_4110_));
 sg13g2_nor4_2 _5022_ (.A(_1215_),
    .B(_1259_),
    .C(net309),
    .Y(_4111_),
    .D(net308));
 sg13g2_nand2_1 _5023_ (.Y(_4112_),
    .A(_4110_),
    .B(_4111_));
 sg13g2_buf_2 _5024_ (.A(_4112_),
    .X(_4113_));
 sg13g2_buf_1 _5025_ (.A(_0011_),
    .X(_4114_));
 sg13g2_nor4_1 _5026_ (.A(_1062_),
    .B(net311),
    .C(net312),
    .D(net304),
    .Y(_4115_));
 sg13g2_inv_1 _5027_ (.Y(_4116_),
    .A(net304));
 sg13g2_or2_1 _5028_ (.X(_4117_),
    .B(net312),
    .A(net311));
 sg13g2_buf_1 _5029_ (.A(_4117_),
    .X(_4118_));
 sg13g2_or2_1 _5030_ (.X(_4119_),
    .B(net307),
    .A(_1336_));
 sg13g2_buf_1 _5031_ (.A(_4119_),
    .X(_4120_));
 sg13g2_or4_1 _5032_ (.A(_1215_),
    .B(_1259_),
    .C(net309),
    .D(net308),
    .X(_4121_));
 sg13g2_nor4_1 _5033_ (.A(_4116_),
    .B(_4118_),
    .C(_4120_),
    .D(_4121_),
    .Y(_4122_));
 sg13g2_a21oi_1 _5034_ (.A1(_4113_),
    .A2(_4115_),
    .Y(_4123_),
    .B1(_4122_));
 sg13g2_buf_2 _5035_ (.A(_4123_),
    .X(_4124_));
 sg13g2_nor2_1 _5036_ (.A(_0897_),
    .B(_0776_),
    .Y(_4125_));
 sg13g2_xor2_1 _5037_ (.B(_0897_),
    .A(net310),
    .X(_4126_));
 sg13g2_and2_1 _5038_ (.A(_4118_),
    .B(_4126_),
    .X(_4127_));
 sg13g2_a21oi_1 _5039_ (.A1(net304),
    .A2(_4125_),
    .Y(_4128_),
    .B1(_4127_));
 sg13g2_buf_2 _5040_ (.A(_4128_),
    .X(_4129_));
 sg13g2_nand2_1 _5041_ (.Y(_4130_),
    .A(_4124_),
    .B(_4129_));
 sg13g2_buf_2 _5042_ (.A(_4130_),
    .X(_4131_));
 sg13g2_o21ai_1 _5043_ (.B1(\flag.flag_abrosexual_inst.pix_x[8] ),
    .Y(_4132_),
    .A1(net310),
    .A2(_0897_));
 sg13g2_buf_1 _5044_ (.A(_4132_),
    .X(_4133_));
 sg13g2_buf_8 _5045_ (.A(_4133_),
    .X(_4134_));
 sg13g2_nand2_2 _5046_ (.Y(_4135_),
    .A(net249),
    .B(net197));
 sg13g2_buf_1 _5047_ (.A(_4135_),
    .X(_4136_));
 sg13g2_or4_1 _5048_ (.A(_1336_),
    .B(_1215_),
    .C(_1259_),
    .D(_0952_),
    .X(_4137_));
 sg13g2_buf_1 _5049_ (.A(_4137_),
    .X(_4138_));
 sg13g2_nor2_1 _5050_ (.A(net274),
    .B(_4138_),
    .Y(_4139_));
 sg13g2_nor2_1 _5051_ (.A(net166),
    .B(_4139_),
    .Y(_4140_));
 sg13g2_xnor2_1 _5052_ (.Y(_4141_),
    .A(_0985_),
    .B(_4140_));
 sg13g2_buf_1 _5053_ (.A(_4141_),
    .X(_4142_));
 sg13g2_nor2_1 _5054_ (.A(_4131_),
    .B(net129),
    .Y(_4143_));
 sg13g2_mux2_1 _5055_ (.A0(_4105_),
    .A1(_4077_),
    .S(_4071_),
    .X(_4144_));
 sg13g2_buf_1 _5056_ (.A(_4144_),
    .X(_4145_));
 sg13g2_buf_8 _5057_ (.A(net147),
    .X(_4146_));
 sg13g2_nand2_1 _5058_ (.Y(_4147_),
    .A(_3976_),
    .B(_3998_));
 sg13g2_nor2_1 _5059_ (.A(net313),
    .B(_4065_),
    .Y(_4148_));
 sg13g2_o21ai_1 _5060_ (.B1(_4148_),
    .Y(_4149_),
    .A1(_4147_),
    .A2(_4098_));
 sg13g2_nor2_1 _5061_ (.A(net272),
    .B(_2087_),
    .Y(_4150_));
 sg13g2_nor4_1 _5062_ (.A(net289),
    .B(net313),
    .C(_4150_),
    .D(_4065_),
    .Y(_4151_));
 sg13g2_a21oi_1 _5063_ (.A1(net289),
    .A2(_4149_),
    .Y(_4152_),
    .B1(_4151_));
 sg13g2_buf_1 _5064_ (.A(_4152_),
    .X(_4153_));
 sg13g2_buf_1 _5065_ (.A(net158),
    .X(_4154_));
 sg13g2_nand2_1 _5066_ (.Y(_4155_),
    .A(net128),
    .B(net146));
 sg13g2_nand2_1 _5067_ (.Y(_4156_),
    .A(net315),
    .B(_0469_));
 sg13g2_buf_2 _5068_ (.A(_4156_),
    .X(_4157_));
 sg13g2_o21ai_1 _5069_ (.B1(net291),
    .Y(_4158_),
    .A1(_4157_),
    .A2(_4065_));
 sg13g2_nand3b_1 _5070_ (.B(_4087_),
    .C(_4089_),
    .Y(_4159_),
    .A_N(net291));
 sg13g2_a22oi_1 _5071_ (.Y(_4160_),
    .B1(_4158_),
    .B2(_4159_),
    .A2(_4086_),
    .A1(_4080_));
 sg13g2_nand2b_1 _5072_ (.Y(_4161_),
    .B(_4157_),
    .A_N(net291));
 sg13g2_buf_1 _5073_ (.A(_4009_),
    .X(_4162_));
 sg13g2_a221oi_1 _5074_ (.B2(_4161_),
    .C1(net177),
    .B1(_4075_),
    .A1(_4098_),
    .Y(_4163_),
    .A2(_4084_));
 sg13g2_or2_1 _5075_ (.X(_4164_),
    .B(_4163_),
    .A(_4160_));
 sg13g2_buf_2 _5076_ (.A(_4164_),
    .X(_4165_));
 sg13g2_o21ai_1 _5077_ (.B1(net296),
    .Y(_4166_),
    .A1(net289),
    .A2(_4009_));
 sg13g2_nor2_1 _5078_ (.A(_0062_),
    .B(_0469_),
    .Y(_4167_));
 sg13g2_buf_2 _5079_ (.A(_4167_),
    .X(_4168_));
 sg13g2_a21oi_1 _5080_ (.A1(_4082_),
    .A2(_4083_),
    .Y(_4169_),
    .B1(_4020_));
 sg13g2_a22oi_1 _5081_ (.Y(_4170_),
    .B1(net177),
    .B2(_4169_),
    .A2(_4168_),
    .A1(_0381_));
 sg13g2_nor4_1 _5082_ (.A(_4080_),
    .B(_4098_),
    .C(_4157_),
    .D(_4093_),
    .Y(_4171_));
 sg13g2_a21o_1 _5083_ (.A2(_4170_),
    .A1(_4166_),
    .B1(_4171_),
    .X(_4172_));
 sg13g2_buf_2 _5084_ (.A(_4172_),
    .X(_4173_));
 sg13g2_buf_1 _5085_ (.A(_4173_),
    .X(_4174_));
 sg13g2_buf_1 _5086_ (.A(net127),
    .X(_4175_));
 sg13g2_nor2_2 _5087_ (.A(_4165_),
    .B(net104),
    .Y(_4176_));
 sg13g2_xor2_1 _5088_ (.B(_4176_),
    .A(_4155_),
    .X(_4177_));
 sg13g2_xnor2_1 _5089_ (.Y(_4178_),
    .A(_4143_),
    .B(_4177_));
 sg13g2_inv_1 _5090_ (.Y(_4179_),
    .A(_4178_));
 sg13g2_a21o_1 _5091_ (.A2(_4115_),
    .A1(_4113_),
    .B1(_4122_),
    .X(_4180_));
 sg13g2_buf_2 _5092_ (.A(_4180_),
    .X(_4181_));
 sg13g2_a21o_1 _5093_ (.A2(_4125_),
    .A1(net304),
    .B1(_4127_),
    .X(_4182_));
 sg13g2_buf_2 _5094_ (.A(_4182_),
    .X(_4183_));
 sg13g2_nor2_1 _5095_ (.A(_4181_),
    .B(_4183_),
    .Y(_4184_));
 sg13g2_buf_2 _5096_ (.A(_4184_),
    .X(_4185_));
 sg13g2_buf_1 _5097_ (.A(_0014_),
    .X(_4186_));
 sg13g2_inv_1 _5098_ (.Y(_4187_),
    .A(_4186_));
 sg13g2_or4_1 _5099_ (.A(net277),
    .B(net307),
    .C(_1215_),
    .D(net278),
    .X(_4188_));
 sg13g2_nand3_1 _5100_ (.B(net197),
    .C(_4188_),
    .A(net249),
    .Y(_4189_));
 sg13g2_xnor2_1 _5101_ (.Y(_4190_),
    .A(_4187_),
    .B(_4189_));
 sg13g2_buf_1 _5102_ (.A(_4190_),
    .X(_4191_));
 sg13g2_buf_1 _5103_ (.A(net157),
    .X(_4192_));
 sg13g2_nand2_1 _5104_ (.Y(_4193_),
    .A(_4185_),
    .B(net145));
 sg13g2_nand2_1 _5105_ (.Y(_4194_),
    .A(_4082_),
    .B(_4083_));
 sg13g2_buf_2 _5106_ (.A(_4194_),
    .X(_4195_));
 sg13g2_inv_1 _5107_ (.Y(_4196_),
    .A(net306));
 sg13g2_o21ai_1 _5108_ (.B1(_0238_),
    .Y(_4197_),
    .A1(_4196_),
    .A2(_4042_));
 sg13g2_buf_2 _5109_ (.A(_4197_),
    .X(_4198_));
 sg13g2_nand2_1 _5110_ (.Y(_4199_),
    .A(_4195_),
    .B(_4198_));
 sg13g2_mux2_1 _5111_ (.A0(net316),
    .A1(_4199_),
    .S(net148),
    .X(_4200_));
 sg13g2_buf_2 _5112_ (.A(_4200_),
    .X(_4201_));
 sg13g2_nor2_2 _5113_ (.A(_4165_),
    .B(_4201_),
    .Y(_4202_));
 sg13g2_nand2b_1 _5114_ (.Y(_4203_),
    .B(_4202_),
    .A_N(_4155_));
 sg13g2_buf_2 _5115_ (.A(_4203_),
    .X(_4204_));
 sg13g2_xnor2_1 _5116_ (.Y(_4205_),
    .A(_4193_),
    .B(_4204_));
 sg13g2_buf_1 _5117_ (.A(net146),
    .X(_4206_));
 sg13g2_nor2_1 _5118_ (.A(_4160_),
    .B(_4163_),
    .Y(_4207_));
 sg13g2_buf_1 _5119_ (.A(_4207_),
    .X(_4208_));
 sg13g2_nand2_1 _5120_ (.Y(_4209_),
    .A(net126),
    .B(net144));
 sg13g2_nand4_1 _5121_ (.B(_4195_),
    .C(_4069_),
    .A(net177),
    .Y(_4210_),
    .D(_4198_));
 sg13g2_o21ai_1 _5122_ (.B1(_4210_),
    .Y(_4211_),
    .A1(net316),
    .A2(_4095_));
 sg13g2_buf_2 _5123_ (.A(_4211_),
    .X(_4212_));
 sg13g2_buf_1 _5124_ (.A(_4212_),
    .X(_4213_));
 sg13g2_buf_1 _5125_ (.A(net103),
    .X(_4214_));
 sg13g2_a21o_1 _5126_ (.A2(_4149_),
    .A1(net289),
    .B1(_4151_),
    .X(_4215_));
 sg13g2_buf_2 _5127_ (.A(_4215_),
    .X(_4216_));
 sg13g2_buf_1 _5128_ (.A(_4216_),
    .X(_4217_));
 sg13g2_a21oi_1 _5129_ (.A1(_4166_),
    .A2(_4170_),
    .Y(_4218_),
    .B1(_4171_));
 sg13g2_buf_1 _5130_ (.A(_4218_),
    .X(_4219_));
 sg13g2_buf_1 _5131_ (.A(_0008_),
    .X(_4220_));
 sg13g2_buf_1 _5132_ (.A(_4220_),
    .X(_4221_));
 sg13g2_xnor2_1 _5133_ (.Y(_4222_),
    .A(_1686_),
    .B(net211));
 sg13g2_mux2_1 _5134_ (.A0(net271),
    .A1(_4222_),
    .S(net148),
    .X(_4223_));
 sg13g2_buf_8 _5135_ (.A(_4223_),
    .X(_4224_));
 sg13g2_nor3_1 _5136_ (.A(net143),
    .B(net142),
    .C(_4224_),
    .Y(_4225_));
 sg13g2_o21ai_1 _5137_ (.B1(net128),
    .Y(_4226_),
    .A1(_4214_),
    .A2(_4225_));
 sg13g2_xnor2_1 _5138_ (.Y(_4227_),
    .A(net293),
    .B(_1501_));
 sg13g2_buf_1 _5139_ (.A(_4227_),
    .X(_4228_));
 sg13g2_inv_2 _5140_ (.Y(_4229_),
    .A(_4220_));
 sg13g2_and3_1 _5141_ (.X(_4230_),
    .A(_4229_),
    .B(_4071_),
    .C(_4077_));
 sg13g2_buf_1 _5142_ (.A(_4230_),
    .X(_4231_));
 sg13g2_a221oi_1 _5143_ (.B2(_4106_),
    .C1(_4231_),
    .B1(net176),
    .A1(net146),
    .Y(_4232_),
    .A2(net103));
 sg13g2_mux2_1 _5144_ (.A0(_4229_),
    .A1(net176),
    .S(_4095_),
    .X(_4233_));
 sg13g2_buf_1 _5145_ (.A(_4233_),
    .X(_4234_));
 sg13g2_buf_8 _5146_ (.A(_4234_),
    .X(_4235_));
 sg13g2_nand3_1 _5147_ (.B(net103),
    .C(net102),
    .A(net126),
    .Y(_4236_));
 sg13g2_o21ai_1 _5148_ (.B1(_4236_),
    .Y(_4237_),
    .A1(_4165_),
    .A2(_4232_));
 sg13g2_a22oi_1 _5149_ (.Y(_4238_),
    .B1(_4237_),
    .B2(net104),
    .A2(_4226_),
    .A1(_4209_));
 sg13g2_nor2b_1 _5150_ (.A(_4205_),
    .B_N(_4238_),
    .Y(_4239_));
 sg13g2_and3_1 _5151_ (.X(_4240_),
    .A(net148),
    .B(_4105_),
    .C(net176));
 sg13g2_buf_1 _5152_ (.A(_4240_),
    .X(_4241_));
 sg13g2_nor2_1 _5153_ (.A(_4241_),
    .B(_4231_),
    .Y(_4242_));
 sg13g2_nand2b_1 _5154_ (.Y(_4243_),
    .B(_4202_),
    .A_N(_4242_));
 sg13g2_buf_1 _5155_ (.A(_4201_),
    .X(_4244_));
 sg13g2_a21oi_1 _5156_ (.A1(_4165_),
    .A2(_4244_),
    .Y(_4245_),
    .B1(_4242_));
 sg13g2_buf_1 _5157_ (.A(net126),
    .X(_4246_));
 sg13g2_o21ai_1 _5158_ (.B1(net101),
    .Y(_4247_),
    .A1(_4202_),
    .A2(_4245_));
 sg13g2_buf_1 _5159_ (.A(net142),
    .X(_4248_));
 sg13g2_a21oi_1 _5160_ (.A1(_4243_),
    .A2(_4247_),
    .Y(_4249_),
    .B1(net125));
 sg13g2_nor2_1 _5161_ (.A(_4239_),
    .B(_4249_),
    .Y(_4250_));
 sg13g2_nor2_1 _5162_ (.A(_4179_),
    .B(_4250_),
    .Y(_4251_));
 sg13g2_buf_2 _5163_ (.A(_0012_),
    .X(_4252_));
 sg13g2_o21ai_1 _5164_ (.B1(_4252_),
    .Y(_4253_),
    .A1(_4120_),
    .A2(_4121_));
 sg13g2_or2_1 _5165_ (.X(_4254_),
    .B(_0897_),
    .A(net310));
 sg13g2_buf_1 _5166_ (.A(_4254_),
    .X(_4255_));
 sg13g2_nor3_1 _5167_ (.A(_1347_),
    .B(_1369_),
    .C(_4252_),
    .Y(_4256_));
 sg13g2_a221oi_1 _5168_ (.B2(_4256_),
    .C1(net312),
    .B1(_4111_),
    .A1(net311),
    .Y(_4257_),
    .A2(_4255_));
 sg13g2_a21oi_1 _5169_ (.A1(_0798_),
    .A2(_4134_),
    .Y(_4258_),
    .B1(_0897_));
 sg13g2_a21o_1 _5170_ (.A2(_4257_),
    .A1(_4253_),
    .B1(_4258_),
    .X(_4259_));
 sg13g2_buf_2 _5171_ (.A(_4259_),
    .X(_4260_));
 sg13g2_buf_1 _5172_ (.A(_4260_),
    .X(_4261_));
 sg13g2_xnor2_1 _5173_ (.Y(_4262_),
    .A(_4186_),
    .B(_4189_));
 sg13g2_buf_2 _5174_ (.A(_4262_),
    .X(_4263_));
 sg13g2_buf_1 _5175_ (.A(_4263_),
    .X(_4264_));
 sg13g2_nor2_1 _5176_ (.A(net140),
    .B(_4204_),
    .Y(_4265_));
 sg13g2_xnor2_1 _5177_ (.Y(_4266_),
    .A(net129),
    .B(_4265_));
 sg13g2_nand2_2 _5178_ (.Y(_4267_),
    .A(_4185_),
    .B(_4260_));
 sg13g2_nor2_1 _5179_ (.A(net140),
    .B(_4267_),
    .Y(_4268_));
 sg13g2_nand2_1 _5180_ (.Y(_4269_),
    .A(net141),
    .B(net129));
 sg13g2_a22oi_1 _5181_ (.Y(_4270_),
    .B1(_4269_),
    .B2(_4131_),
    .A2(_4268_),
    .A1(_4204_));
 sg13g2_o21ai_1 _5182_ (.B1(_4270_),
    .Y(_4271_),
    .A1(net141),
    .A2(_4266_));
 sg13g2_a21oi_1 _5183_ (.A1(_4179_),
    .A2(_4250_),
    .Y(_4272_),
    .B1(_4271_));
 sg13g2_nor2_2 _5184_ (.A(_4251_),
    .B(_4272_),
    .Y(_4273_));
 sg13g2_a21oi_1 _5185_ (.A1(_4253_),
    .A2(_4257_),
    .Y(_4274_),
    .B1(_4258_));
 sg13g2_buf_2 _5186_ (.A(_4274_),
    .X(_4275_));
 sg13g2_o21ai_1 _5187_ (.B1(_4275_),
    .Y(_4276_),
    .A1(_4142_),
    .A2(_4204_));
 sg13g2_nand2b_1 _5188_ (.Y(_4277_),
    .B(_4276_),
    .A_N(_4193_));
 sg13g2_buf_1 _5189_ (.A(_4277_),
    .X(_4278_));
 sg13g2_nor3_2 _5190_ (.A(_4181_),
    .B(_4183_),
    .C(_4275_),
    .Y(_4279_));
 sg13g2_buf_1 _5191_ (.A(net144),
    .X(_4280_));
 sg13g2_xnor2_1 _5192_ (.Y(_4281_),
    .A(_1182_),
    .B(_4140_));
 sg13g2_nand2_1 _5193_ (.Y(_4282_),
    .A(_4185_),
    .B(_4281_));
 sg13g2_nor2_2 _5194_ (.A(net146),
    .B(net142),
    .Y(_4283_));
 sg13g2_nand2_1 _5195_ (.Y(_4284_),
    .A(_4108_),
    .B(net104));
 sg13g2_o21ai_1 _5196_ (.B1(_4284_),
    .Y(_4285_),
    .A1(_4282_),
    .A2(_4283_));
 sg13g2_nor2_1 _5197_ (.A(net143),
    .B(net127),
    .Y(_4286_));
 sg13g2_o21ai_1 _5198_ (.B1(_4286_),
    .Y(_4287_),
    .A1(net124),
    .A2(_4143_));
 sg13g2_nor2_1 _5199_ (.A(net144),
    .B(net125),
    .Y(_4288_));
 sg13g2_o21ai_1 _5200_ (.B1(_4288_),
    .Y(_4289_),
    .A1(net143),
    .A2(_4282_));
 sg13g2_nand2_1 _5201_ (.Y(_4290_),
    .A(_4287_),
    .B(_4289_));
 sg13g2_a22oi_1 _5202_ (.Y(_4291_),
    .B1(_4290_),
    .B2(net128),
    .A2(_4285_),
    .A1(net124));
 sg13g2_xnor2_1 _5203_ (.Y(_4292_),
    .A(_4279_),
    .B(_4291_));
 sg13g2_nor4_2 _5204_ (.A(net277),
    .B(_1215_),
    .C(_1270_),
    .Y(_4293_),
    .D(_0952_));
 sg13g2_a21oi_1 _5205_ (.A1(_3342_),
    .A2(_4293_),
    .Y(_4294_),
    .B1(net280));
 sg13g2_nor3_1 _5206_ (.A(net308),
    .B(net274),
    .C(_4138_),
    .Y(_4295_));
 sg13g2_and2_1 _5207_ (.A(_0787_),
    .B(_4133_),
    .X(_4296_));
 sg13g2_buf_2 _5208_ (.A(_4296_),
    .X(_4297_));
 sg13g2_o21ai_1 _5209_ (.B1(_4297_),
    .Y(_4298_),
    .A1(_4294_),
    .A2(_4295_));
 sg13g2_buf_2 _5210_ (.A(_4298_),
    .X(_4299_));
 sg13g2_buf_1 _5211_ (.A(_0013_),
    .X(_4300_));
 sg13g2_nand2_2 _5212_ (.Y(_4301_),
    .A(_4300_),
    .B(_4135_));
 sg13g2_nand2_2 _5213_ (.Y(_4302_),
    .A(_4299_),
    .B(_4301_));
 sg13g2_nand2_2 _5214_ (.Y(_4303_),
    .A(net129),
    .B(_4302_));
 sg13g2_and2_1 _5215_ (.A(_4299_),
    .B(_4301_),
    .X(_4304_));
 sg13g2_buf_2 _5216_ (.A(_4304_),
    .X(_4305_));
 sg13g2_nand2_1 _5217_ (.Y(_4306_),
    .A(_4131_),
    .B(_4305_));
 sg13g2_o21ai_1 _5218_ (.B1(_4306_),
    .Y(_4307_),
    .A1(_4131_),
    .A2(_4303_));
 sg13g2_nand2_1 _5219_ (.Y(_4308_),
    .A(net141),
    .B(_4307_));
 sg13g2_inv_1 _5220_ (.Y(_4309_),
    .A(_4308_));
 sg13g2_xnor2_1 _5221_ (.Y(_4310_),
    .A(_4292_),
    .B(_4309_));
 sg13g2_and2_1 _5222_ (.A(_4278_),
    .B(_4310_),
    .X(_4311_));
 sg13g2_o21ai_1 _5223_ (.B1(_4273_),
    .Y(_4312_),
    .A1(_4278_),
    .A2(_4310_));
 sg13g2_nand2b_1 _5224_ (.Y(_4313_),
    .B(_4312_),
    .A_N(_4311_));
 sg13g2_buf_1 _5225_ (.A(_0016_),
    .X(_4314_));
 sg13g2_buf_1 _5226_ (.A(_4314_),
    .X(_4315_));
 sg13g2_or3_1 _5227_ (.A(_1336_),
    .B(\flag.flag_abrosexual_inst.pix_x[0] ),
    .C(_1259_),
    .X(_4316_));
 sg13g2_buf_2 _5228_ (.A(_4316_),
    .X(_4317_));
 sg13g2_nand3_1 _5229_ (.B(net197),
    .C(_4317_),
    .A(net249),
    .Y(_4318_));
 sg13g2_buf_1 _5230_ (.A(_4318_),
    .X(_4319_));
 sg13g2_xnor2_1 _5231_ (.Y(_4320_),
    .A(net270),
    .B(_4319_));
 sg13g2_buf_2 _5232_ (.A(_4320_),
    .X(_4321_));
 sg13g2_nor3_1 _5233_ (.A(_4181_),
    .B(_4183_),
    .C(_4321_),
    .Y(_4322_));
 sg13g2_buf_2 _5234_ (.A(_4322_),
    .X(_4323_));
 sg13g2_nand4_1 _5235_ (.B(_4208_),
    .C(net103),
    .A(net146),
    .Y(_4324_),
    .D(net127));
 sg13g2_a22oi_1 _5236_ (.Y(_4325_),
    .B1(net127),
    .B2(net146),
    .A2(_4213_),
    .A1(_4208_));
 sg13g2_a21oi_1 _5237_ (.A1(_4242_),
    .A2(_4324_),
    .Y(_4326_),
    .B1(_4325_));
 sg13g2_and2_1 _5238_ (.A(_4323_),
    .B(_4326_),
    .X(_4327_));
 sg13g2_buf_1 _5239_ (.A(_4327_),
    .X(_4328_));
 sg13g2_a21oi_2 _5240_ (.B1(_4260_),
    .Y(_4329_),
    .A2(_4129_),
    .A1(_4124_));
 sg13g2_nor2_1 _5241_ (.A(_4305_),
    .B(_4328_),
    .Y(_4330_));
 sg13g2_nor3_1 _5242_ (.A(_4279_),
    .B(_4329_),
    .C(_4330_),
    .Y(_4331_));
 sg13g2_a21o_1 _5243_ (.A2(_4328_),
    .A1(_4305_),
    .B1(_4331_),
    .X(_4332_));
 sg13g2_nor2_2 _5244_ (.A(_4191_),
    .B(net129),
    .Y(_4333_));
 sg13g2_a22oi_1 _5245_ (.Y(_4334_),
    .B1(_4333_),
    .B2(_4328_),
    .A2(_4332_),
    .A1(net145));
 sg13g2_xnor2_1 _5246_ (.Y(_4335_),
    .A(_4179_),
    .B(_4250_));
 sg13g2_xnor2_1 _5247_ (.Y(_4336_),
    .A(_4271_),
    .B(_4335_));
 sg13g2_nor2_1 _5248_ (.A(_4334_),
    .B(_4336_),
    .Y(_4337_));
 sg13g2_xnor2_1 _5249_ (.Y(_4338_),
    .A(_4238_),
    .B(_4205_));
 sg13g2_buf_1 _5250_ (.A(_4338_),
    .X(_4339_));
 sg13g2_inv_1 _5251_ (.Y(_4340_),
    .A(_4339_));
 sg13g2_xnor2_1 _5252_ (.Y(_4341_),
    .A(net129),
    .B(_4326_));
 sg13g2_and2_1 _5253_ (.A(net140),
    .B(_4323_),
    .X(_4342_));
 sg13g2_o21ai_1 _5254_ (.B1(_4302_),
    .Y(_4343_),
    .A1(_4279_),
    .A2(_4329_));
 sg13g2_or3_1 _5255_ (.A(_4279_),
    .B(_4329_),
    .C(_4302_),
    .X(_4344_));
 sg13g2_a21oi_1 _5256_ (.A1(_4343_),
    .A2(_4344_),
    .Y(_4345_),
    .B1(net140));
 sg13g2_nand3_1 _5257_ (.B(_4343_),
    .C(_4344_),
    .A(_4192_),
    .Y(_4346_));
 sg13g2_a21oi_1 _5258_ (.A1(_4323_),
    .A2(_4326_),
    .Y(_4347_),
    .B1(_4346_));
 sg13g2_a221oi_1 _5259_ (.B2(_4328_),
    .C1(_4347_),
    .B1(_4345_),
    .A1(_4341_),
    .Y(_4348_),
    .A2(_4342_));
 sg13g2_buf_2 _5260_ (.A(_4348_),
    .X(_4349_));
 sg13g2_buf_1 _5261_ (.A(net104),
    .X(_4350_));
 sg13g2_nand2b_1 _5262_ (.Y(_4351_),
    .B(_4072_),
    .A_N(_4583_));
 sg13g2_nand3_1 _5263_ (.B(_4105_),
    .C(net176),
    .A(net130),
    .Y(_4352_));
 sg13g2_nand3_1 _5264_ (.B(net159),
    .C(_4077_),
    .A(_4229_),
    .Y(_4353_));
 sg13g2_a221oi_1 _5265_ (.B2(_4353_),
    .C1(_4165_),
    .B1(_4352_),
    .A1(_4210_),
    .Y(_4354_),
    .A2(_4351_));
 sg13g2_xnor2_1 _5266_ (.Y(_4355_),
    .A(_4202_),
    .B(_4242_));
 sg13g2_mux2_1 _5267_ (.A0(_4354_),
    .A1(_4355_),
    .S(net101),
    .X(_4356_));
 sg13g2_o21ai_1 _5268_ (.B1(_4323_),
    .Y(_4357_),
    .A1(_4241_),
    .A2(_4231_));
 sg13g2_nor3_1 _5269_ (.A(_4241_),
    .B(_4231_),
    .C(_4323_),
    .Y(_4358_));
 sg13g2_a22oi_1 _5270_ (.Y(_4359_),
    .B1(_4358_),
    .B2(_4217_),
    .A2(_4357_),
    .A1(_4219_));
 sg13g2_a22oi_1 _5271_ (.Y(_4360_),
    .B1(_4358_),
    .B2(net125),
    .A2(_4323_),
    .A1(_4354_));
 sg13g2_o21ai_1 _5272_ (.B1(_4360_),
    .Y(_4361_),
    .A1(_4202_),
    .A2(_4359_));
 sg13g2_a21oi_1 _5273_ (.A1(net63),
    .A2(_4356_),
    .Y(_4362_),
    .B1(_4361_));
 sg13g2_buf_2 _5274_ (.A(_4362_),
    .X(_4363_));
 sg13g2_nand2b_1 _5275_ (.Y(_4364_),
    .B(_4363_),
    .A_N(_4349_));
 sg13g2_nor2b_1 _5276_ (.A(_4363_),
    .B_N(_4349_),
    .Y(_4365_));
 sg13g2_a21oi_1 _5277_ (.A1(_4340_),
    .A2(_4364_),
    .Y(_4366_),
    .B1(_4365_));
 sg13g2_nand2_1 _5278_ (.Y(_4367_),
    .A(_4334_),
    .B(_4336_));
 sg13g2_o21ai_1 _5279_ (.B1(_4367_),
    .Y(_4368_),
    .A1(_4337_),
    .A2(_4366_));
 sg13g2_nor4_1 _5280_ (.A(_4278_),
    .B(_4273_),
    .C(_4310_),
    .D(_4368_),
    .Y(_4369_));
 sg13g2_a221oi_1 _5281_ (.B2(_4368_),
    .C1(_4369_),
    .B1(_4313_),
    .A1(_4273_),
    .Y(_4370_),
    .A2(_4311_));
 sg13g2_nor2_1 _5282_ (.A(_4282_),
    .B(_4267_),
    .Y(_4371_));
 sg13g2_nor2_1 _5283_ (.A(_4282_),
    .B(_4288_),
    .Y(_4372_));
 sg13g2_o21ai_1 _5284_ (.B1(_4279_),
    .Y(_4373_),
    .A1(_4176_),
    .A2(_4372_));
 sg13g2_nand3_1 _5285_ (.B(_4267_),
    .C(_4288_),
    .A(_4143_),
    .Y(_4374_));
 sg13g2_a21oi_1 _5286_ (.A1(_4373_),
    .A2(_4374_),
    .Y(_4375_),
    .B1(_4155_));
 sg13g2_a221oi_1 _5287_ (.B2(_4176_),
    .C1(_4375_),
    .B1(_4371_),
    .A1(_4292_),
    .Y(_4376_),
    .A2(_4309_));
 sg13g2_a21oi_1 _5288_ (.A1(net141),
    .A2(_4288_),
    .Y(_4377_),
    .B1(_4176_));
 sg13g2_nand3_1 _5289_ (.B(_4350_),
    .C(_4303_),
    .A(net141),
    .Y(_4378_));
 sg13g2_o21ai_1 _5290_ (.B1(_4378_),
    .Y(_4379_),
    .A1(net141),
    .A2(_4350_));
 sg13g2_o21ai_1 _5291_ (.B1(net141),
    .Y(_4380_),
    .A1(net124),
    .A2(_4303_));
 sg13g2_a22oi_1 _5292_ (.Y(_4381_),
    .B1(_4380_),
    .B2(_4108_),
    .A2(_4379_),
    .A1(net124));
 sg13g2_o21ai_1 _5293_ (.B1(_4381_),
    .Y(_4382_),
    .A1(_4303_),
    .A2(_4377_));
 sg13g2_nand4_1 _5294_ (.B(_4165_),
    .C(net125),
    .A(_4261_),
    .Y(_4383_),
    .D(_4303_));
 sg13g2_o21ai_1 _5295_ (.B1(_4383_),
    .Y(_4384_),
    .A1(_4185_),
    .A2(_4176_));
 sg13g2_a22oi_1 _5296_ (.Y(_4385_),
    .B1(_4384_),
    .B2(net128),
    .A2(_4382_),
    .A1(_4185_));
 sg13g2_xnor2_1 _5297_ (.Y(_4386_),
    .A(_4376_),
    .B(_4385_));
 sg13g2_xnor2_1 _5298_ (.Y(_4387_),
    .A(_4370_),
    .B(_4386_));
 sg13g2_buf_1 _5299_ (.A(_0015_),
    .X(_4388_));
 sg13g2_inv_1 _5300_ (.Y(_4389_),
    .A(net303));
 sg13g2_and2_1 _5301_ (.A(net269),
    .B(_4077_),
    .X(_4390_));
 sg13g2_nor2b_1 _5302_ (.A(_0139_),
    .B_N(net295),
    .Y(_4391_));
 sg13g2_buf_2 _5303_ (.A(_4391_),
    .X(_4392_));
 sg13g2_nor2b_2 _5304_ (.A(_0117_),
    .B_N(_0139_),
    .Y(_4393_));
 sg13g2_nor2_2 _5305_ (.A(_4392_),
    .B(_4393_),
    .Y(_4394_));
 sg13g2_a221oi_1 _5306_ (.B2(_4093_),
    .C1(_4394_),
    .B1(net198),
    .A1(_4080_),
    .Y(_4395_),
    .A2(_4086_));
 sg13g2_buf_1 _5307_ (.A(_4395_),
    .X(_4396_));
 sg13g2_a22oi_1 _5308_ (.Y(_4397_),
    .B1(_4396_),
    .B2(_4105_),
    .A2(_4390_),
    .A1(net167));
 sg13g2_buf_2 _5309_ (.A(_4397_),
    .X(_4398_));
 sg13g2_buf_8 _5310_ (.A(_4398_),
    .X(_4399_));
 sg13g2_nand2_1 _5311_ (.Y(_4400_),
    .A(_4216_),
    .B(net100));
 sg13g2_xnor2_1 _5312_ (.Y(_4401_),
    .A(net291),
    .B(net198));
 sg13g2_buf_1 _5313_ (.A(_4401_),
    .X(_4402_));
 sg13g2_nand2_1 _5314_ (.Y(_4403_),
    .A(_0524_),
    .B(_1632_));
 sg13g2_and2_1 _5315_ (.A(net165),
    .B(_4403_),
    .X(_4404_));
 sg13g2_nor2_1 _5316_ (.A(net303),
    .B(net165),
    .Y(_4405_));
 sg13g2_mux2_1 _5317_ (.A0(_4404_),
    .A1(_4405_),
    .S(net167),
    .X(_4406_));
 sg13g2_buf_2 _5318_ (.A(_4406_),
    .X(_4407_));
 sg13g2_a21oi_2 _5319_ (.B1(_4407_),
    .Y(_4408_),
    .A2(net128),
    .A1(net223));
 sg13g2_and2_1 _5320_ (.A(net167),
    .B(_4390_),
    .X(_4409_));
 sg13g2_buf_1 _5321_ (.A(_4409_),
    .X(_4410_));
 sg13g2_nor2_1 _5322_ (.A(_1719_),
    .B(net165),
    .Y(_4411_));
 sg13g2_and4_1 _5323_ (.A(net294),
    .B(_4105_),
    .C(net165),
    .D(_4396_),
    .X(_4412_));
 sg13g2_buf_1 _5324_ (.A(_4412_),
    .X(_4413_));
 sg13g2_a221oi_1 _5325_ (.B2(_4411_),
    .C1(_4413_),
    .B1(_4410_),
    .A1(_4173_),
    .Y(_4414_),
    .A2(_4234_));
 sg13g2_xnor2_1 _5326_ (.Y(_4415_),
    .A(net158),
    .B(net100));
 sg13g2_o21ai_1 _5327_ (.B1(_4415_),
    .Y(_4416_),
    .A1(_4408_),
    .A2(_4414_));
 sg13g2_buf_1 _5328_ (.A(_4416_),
    .X(_4417_));
 sg13g2_nand2_1 _5329_ (.Y(_4418_),
    .A(_4080_),
    .B(_4086_));
 sg13g2_and2_1 _5330_ (.A(net176),
    .B(_4402_),
    .X(_4419_));
 sg13g2_nor4_1 _5331_ (.A(net271),
    .B(net177),
    .C(_4061_),
    .D(net165),
    .Y(_4420_));
 sg13g2_a21oi_1 _5332_ (.A1(_4418_),
    .A2(_4419_),
    .Y(_4421_),
    .B1(_4420_));
 sg13g2_o21ai_1 _5333_ (.B1(_4421_),
    .Y(_4422_),
    .A1(_4201_),
    .A2(_4219_));
 sg13g2_buf_1 _5334_ (.A(_0018_),
    .X(_4423_));
 sg13g2_mux2_1 _5335_ (.A0(net302),
    .A1(_3417_),
    .S(_4297_),
    .X(_4424_));
 sg13g2_buf_2 _5336_ (.A(_4424_),
    .X(_4425_));
 sg13g2_buf_1 _5337_ (.A(_0017_),
    .X(_4426_));
 sg13g2_a21oi_1 _5338_ (.A1(_0798_),
    .A2(_4134_),
    .Y(_4427_),
    .B1(_4426_));
 sg13g2_o21ai_1 _5339_ (.B1(_1259_),
    .Y(_4428_),
    .A1(_1336_),
    .A2(net307));
 sg13g2_nand4_1 _5340_ (.B(net197),
    .C(_4317_),
    .A(net218),
    .Y(_4429_),
    .D(_4428_));
 sg13g2_nand2b_1 _5341_ (.Y(_4430_),
    .B(_4429_),
    .A_N(_4427_));
 sg13g2_buf_1 _5342_ (.A(_4430_),
    .X(_4431_));
 sg13g2_buf_1 _5343_ (.A(_4431_),
    .X(_4432_));
 sg13g2_o21ai_1 _5344_ (.B1(net139),
    .Y(_4433_),
    .A1(net100),
    .A2(_4425_));
 sg13g2_and4_1 _5345_ (.A(net249),
    .B(_4133_),
    .C(_4317_),
    .D(_4428_),
    .X(_4434_));
 sg13g2_buf_1 _5346_ (.A(_4434_),
    .X(_4435_));
 sg13g2_nor2_1 _5347_ (.A(_4427_),
    .B(_4435_),
    .Y(_4436_));
 sg13g2_buf_2 _5348_ (.A(_4436_),
    .X(_4437_));
 sg13g2_inv_2 _5349_ (.Y(_4438_),
    .A(net302));
 sg13g2_xor2_1 _5350_ (.B(net307),
    .A(_1336_),
    .X(_4439_));
 sg13g2_buf_2 _5351_ (.A(_4439_),
    .X(_4440_));
 sg13g2_mux2_1 _5352_ (.A0(_4438_),
    .A1(_4440_),
    .S(_4297_),
    .X(_4441_));
 sg13g2_buf_2 _5353_ (.A(_4441_),
    .X(_4442_));
 sg13g2_nand3b_1 _5354_ (.B(_4437_),
    .C(_4442_),
    .Y(_4443_),
    .A_N(net100));
 sg13g2_a21oi_2 _5355_ (.B1(_4131_),
    .Y(_4444_),
    .A2(_4443_),
    .A1(_4433_));
 sg13g2_a21o_1 _5356_ (.A2(_4419_),
    .A1(_4418_),
    .B1(_4420_),
    .X(_4445_));
 sg13g2_buf_1 _5357_ (.A(_4445_),
    .X(_4446_));
 sg13g2_a22oi_1 _5358_ (.Y(_4447_),
    .B1(_4446_),
    .B2(net158),
    .A2(net127),
    .A1(_4212_));
 sg13g2_buf_2 _5359_ (.A(_4447_),
    .X(_4448_));
 sg13g2_nor2_1 _5360_ (.A(net158),
    .B(_4446_),
    .Y(_4449_));
 sg13g2_or2_1 _5361_ (.X(_4450_),
    .B(_4449_),
    .A(_4448_));
 sg13g2_xnor2_1 _5362_ (.Y(_4451_),
    .A(_4444_),
    .B(_4450_));
 sg13g2_a22oi_1 _5363_ (.Y(_4452_),
    .B1(_4422_),
    .B2(_4451_),
    .A2(_4417_),
    .A1(_4400_));
 sg13g2_nand3_1 _5364_ (.B(_4174_),
    .C(_4446_),
    .A(_4212_),
    .Y(_4453_));
 sg13g2_buf_1 _5365_ (.A(_4453_),
    .X(_4454_));
 sg13g2_nand3b_1 _5366_ (.B(_4454_),
    .C(net100),
    .Y(_4455_),
    .A_N(_4417_));
 sg13g2_nand3b_1 _5367_ (.B(_4448_),
    .C(net126),
    .Y(_4456_),
    .A_N(_4444_));
 sg13g2_nand4_1 _5368_ (.B(_4454_),
    .C(_4444_),
    .A(_4206_),
    .Y(_4457_),
    .D(_4422_));
 sg13g2_nand2_1 _5369_ (.Y(_4458_),
    .A(_4213_),
    .B(net127));
 sg13g2_nand3b_1 _5370_ (.B(_4421_),
    .C(_4458_),
    .Y(_4459_),
    .A_N(_4444_));
 sg13g2_nand4_1 _5371_ (.B(_4456_),
    .C(_4457_),
    .A(_4455_),
    .Y(_4460_),
    .D(_4459_));
 sg13g2_nor3_1 _5372_ (.A(_4181_),
    .B(_4183_),
    .C(_4437_),
    .Y(_4461_));
 sg13g2_buf_2 _5373_ (.A(_4461_),
    .X(_4462_));
 sg13g2_nor3_1 _5374_ (.A(_4181_),
    .B(_4183_),
    .C(_4425_),
    .Y(_4463_));
 sg13g2_buf_2 _5375_ (.A(_4463_),
    .X(_4464_));
 sg13g2_nand3b_1 _5376_ (.B(_4462_),
    .C(_4464_),
    .Y(_4465_),
    .A_N(net100));
 sg13g2_o21ai_1 _5377_ (.B1(_4465_),
    .Y(_4466_),
    .A1(_4448_),
    .A2(_4449_));
 sg13g2_buf_1 _5378_ (.A(_4466_),
    .X(_4467_));
 sg13g2_nand3_1 _5379_ (.B(_4129_),
    .C(_4431_),
    .A(_4124_),
    .Y(_4468_));
 sg13g2_nand2b_1 _5380_ (.Y(_4469_),
    .B(_4464_),
    .A_N(net100));
 sg13g2_nand2_1 _5381_ (.Y(_4470_),
    .A(_4468_),
    .B(_4469_));
 sg13g2_inv_2 _5382_ (.Y(_4471_),
    .A(_4314_));
 sg13g2_xnor2_1 _5383_ (.Y(_4472_),
    .A(_4471_),
    .B(_4319_));
 sg13g2_buf_8 _5384_ (.A(_4472_),
    .X(_4473_));
 sg13g2_nand2_1 _5385_ (.Y(_4474_),
    .A(_4260_),
    .B(net138));
 sg13g2_a21oi_2 _5386_ (.B1(_4474_),
    .Y(_4475_),
    .A2(_4462_),
    .A1(_4302_));
 sg13g2_nand3_1 _5387_ (.B(_4281_),
    .C(_4475_),
    .A(_4264_),
    .Y(_4476_));
 sg13g2_nand4_1 _5388_ (.B(_4299_),
    .C(_4301_),
    .A(_4190_),
    .Y(_4477_),
    .D(_4472_));
 sg13g2_buf_1 _5389_ (.A(_4477_),
    .X(_4478_));
 sg13g2_nand2_1 _5390_ (.Y(_4479_),
    .A(_4191_),
    .B(_4260_));
 sg13g2_a21oi_1 _5391_ (.A1(_4478_),
    .A2(_4479_),
    .Y(_4480_),
    .B1(_4468_));
 sg13g2_or3_1 _5392_ (.A(_4333_),
    .B(_4475_),
    .C(_4480_),
    .X(_4481_));
 sg13g2_buf_1 _5393_ (.A(_4481_),
    .X(_4482_));
 sg13g2_a22oi_1 _5394_ (.Y(_4483_),
    .B1(_4476_),
    .B2(_4482_),
    .A2(_4470_),
    .A1(_4467_));
 sg13g2_and4_1 _5395_ (.A(_4467_),
    .B(_4470_),
    .C(_4476_),
    .D(_4482_),
    .X(_4484_));
 sg13g2_xnor2_1 _5396_ (.Y(_4485_),
    .A(_4283_),
    .B(_4355_));
 sg13g2_nor3_2 _5397_ (.A(_4483_),
    .B(_4484_),
    .C(_4485_),
    .Y(_4486_));
 sg13g2_nor3_1 _5398_ (.A(_4448_),
    .B(_4449_),
    .C(_4469_),
    .Y(_4487_));
 sg13g2_o21ai_1 _5399_ (.B1(_4462_),
    .Y(_4488_),
    .A1(_4154_),
    .A2(_4446_));
 sg13g2_o21ai_1 _5400_ (.B1(_4465_),
    .Y(_4489_),
    .A1(_4448_),
    .A2(_4488_));
 sg13g2_and3_1 _5401_ (.X(_4490_),
    .A(net140),
    .B(_4281_),
    .C(_4475_));
 sg13g2_nor3_1 _5402_ (.A(_4333_),
    .B(_4475_),
    .C(_4480_),
    .Y(_4491_));
 sg13g2_nor4_1 _5403_ (.A(_4487_),
    .B(_4489_),
    .C(_4490_),
    .D(_4491_),
    .Y(_4492_));
 sg13g2_and2_1 _5404_ (.A(_4468_),
    .B(_4469_),
    .X(_4493_));
 sg13g2_a221oi_1 _5405_ (.B2(_4482_),
    .C1(_4493_),
    .B1(_4476_),
    .A1(_4450_),
    .Y(_4494_),
    .A2(_4465_));
 sg13g2_xor2_1 _5406_ (.B(_4355_),
    .A(_4283_),
    .X(_4495_));
 sg13g2_nor3_2 _5407_ (.A(_4492_),
    .B(_4494_),
    .C(_4495_),
    .Y(_4496_));
 sg13g2_nor4_2 _5408_ (.A(_4452_),
    .B(_4460_),
    .C(_4486_),
    .Y(_4497_),
    .D(_4496_));
 sg13g2_mux2_1 _5409_ (.A0(_4486_),
    .A1(_4496_),
    .S(_4323_),
    .X(_4498_));
 sg13g2_buf_1 _5410_ (.A(_4498_),
    .X(_4499_));
 sg13g2_nor2_1 _5411_ (.A(_4497_),
    .B(_4499_),
    .Y(_4500_));
 sg13g2_xor2_1 _5412_ (.B(_4349_),
    .A(_4339_),
    .X(_4501_));
 sg13g2_or2_1 _5413_ (.X(_4502_),
    .B(_4480_),
    .A(_4475_));
 sg13g2_nand3_1 _5414_ (.B(_4470_),
    .C(_4502_),
    .A(_4467_),
    .Y(_4503_));
 sg13g2_xnor2_1 _5415_ (.Y(_4504_),
    .A(_4323_),
    .B(_4333_));
 sg13g2_a21oi_1 _5416_ (.A1(_4467_),
    .A2(_4470_),
    .Y(_4505_),
    .B1(_4502_));
 sg13g2_a21oi_2 _5417_ (.B1(_4505_),
    .Y(_4506_),
    .A2(_4504_),
    .A1(_4503_));
 sg13g2_xor2_1 _5418_ (.B(_4506_),
    .A(_4363_),
    .X(_4507_));
 sg13g2_xnor2_1 _5419_ (.Y(_4508_),
    .A(_4501_),
    .B(_4507_));
 sg13g2_xnor2_1 _5420_ (.Y(_4509_),
    .A(_4500_),
    .B(_4508_));
 sg13g2_nand3_1 _5421_ (.B(_4129_),
    .C(_4442_),
    .A(_4124_),
    .Y(_4510_));
 sg13g2_buf_2 _5422_ (.A(_4510_),
    .X(_4511_));
 sg13g2_buf_1 _5423_ (.A(_4297_),
    .X(_4512_));
 sg13g2_inv_2 _5424_ (.Y(_4513_),
    .A(_4252_));
 sg13g2_o21ai_1 _5425_ (.B1(net308),
    .Y(_4514_),
    .A1(net274),
    .A2(_4138_));
 sg13g2_nand3_1 _5426_ (.B(_3342_),
    .C(_4293_),
    .A(net280),
    .Y(_4515_));
 sg13g2_nand3_1 _5427_ (.B(_4514_),
    .C(_4515_),
    .A(_4315_),
    .Y(_4516_));
 sg13g2_a21o_1 _5428_ (.A2(_4515_),
    .A1(_4514_),
    .B1(_4317_),
    .X(_4517_));
 sg13g2_nand4_1 _5429_ (.B(_4428_),
    .C(_4516_),
    .A(_4513_),
    .Y(_4518_),
    .D(_4517_));
 sg13g2_o21ai_1 _5430_ (.B1(_4252_),
    .Y(_4519_),
    .A1(_1347_),
    .A2(net276));
 sg13g2_o21ai_1 _5431_ (.B1(_4519_),
    .Y(_4520_),
    .A1(_1281_),
    .A2(_4256_));
 sg13g2_nor2_1 _5432_ (.A(_1270_),
    .B(net270),
    .Y(_4521_));
 sg13g2_a22oi_1 _5433_ (.Y(_4522_),
    .B1(_4521_),
    .B2(_4110_),
    .A2(_4520_),
    .A1(_4315_));
 sg13g2_or3_1 _5434_ (.A(_4294_),
    .B(_4295_),
    .C(_4522_),
    .X(_4523_));
 sg13g2_nand3_1 _5435_ (.B(_4518_),
    .C(_4523_),
    .A(net164),
    .Y(_4524_));
 sg13g2_buf_1 _5436_ (.A(_4426_),
    .X(_4525_));
 sg13g2_nor2_1 _5437_ (.A(net284),
    .B(net268),
    .Y(_4526_));
 sg13g2_buf_1 _5438_ (.A(_4300_),
    .X(_4527_));
 sg13g2_nor2_1 _5439_ (.A(net267),
    .B(net270),
    .Y(_4528_));
 sg13g2_xnor2_1 _5440_ (.Y(_4529_),
    .A(_4526_),
    .B(_4528_));
 sg13g2_nand2_1 _5441_ (.Y(_4530_),
    .A(net166),
    .B(_4529_));
 sg13g2_nand3_1 _5442_ (.B(_4524_),
    .C(_4530_),
    .A(_4511_),
    .Y(_4531_));
 sg13g2_a22oi_1 _5443_ (.Y(_4532_),
    .B1(_4526_),
    .B2(_4136_),
    .A2(_4435_),
    .A1(_4513_));
 sg13g2_nor2_1 _5444_ (.A(_4511_),
    .B(_4532_),
    .Y(_4533_));
 sg13g2_a21oi_1 _5445_ (.A1(_4305_),
    .A2(_4533_),
    .Y(_4534_),
    .B1(net157));
 sg13g2_nor2_1 _5446_ (.A(net140),
    .B(_4464_),
    .Y(_4535_));
 sg13g2_nor2_1 _5447_ (.A(_4263_),
    .B(_4321_),
    .Y(_4536_));
 sg13g2_nor2_1 _5448_ (.A(_4275_),
    .B(_4425_),
    .Y(_4537_));
 sg13g2_a22oi_1 _5449_ (.Y(_4538_),
    .B1(_4536_),
    .B2(_4537_),
    .A2(_4431_),
    .A1(_4305_));
 sg13g2_or2_1 _5450_ (.X(_4539_),
    .B(_4537_),
    .A(_4536_));
 sg13g2_nand2b_1 _5451_ (.Y(_4540_),
    .B(_4539_),
    .A_N(_4538_));
 sg13g2_buf_2 _5452_ (.A(_4540_),
    .X(_4541_));
 sg13g2_and4_1 _5453_ (.A(net157),
    .B(_4464_),
    .C(_4524_),
    .D(_4530_),
    .X(_4542_));
 sg13g2_a221oi_1 _5454_ (.B2(_4541_),
    .C1(_4542_),
    .B1(_4535_),
    .A1(_4531_),
    .Y(_4543_),
    .A2(_4534_));
 sg13g2_nor2_1 _5455_ (.A(_4462_),
    .B(_4478_),
    .Y(_4544_));
 sg13g2_inv_1 _5456_ (.Y(_4545_),
    .A(net268));
 sg13g2_nand2_1 _5457_ (.Y(_4546_),
    .A(_4545_),
    .B(net166));
 sg13g2_nor2_1 _5458_ (.A(_4300_),
    .B(_4297_),
    .Y(_4547_));
 sg13g2_nor3_1 _5459_ (.A(_4135_),
    .B(_4294_),
    .C(_4295_),
    .Y(_4548_));
 sg13g2_o21ai_1 _5460_ (.B1(net138),
    .Y(_4549_),
    .A1(_4547_),
    .A2(_4548_));
 sg13g2_o21ai_1 _5461_ (.B1(_4260_),
    .Y(_4550_),
    .A1(_4181_),
    .A2(_4183_));
 sg13g2_a221oi_1 _5462_ (.B2(_4263_),
    .C1(_4550_),
    .B1(_4549_),
    .A1(_4546_),
    .Y(_4551_),
    .A2(_4429_));
 sg13g2_nor2_1 _5463_ (.A(_4544_),
    .B(_4551_),
    .Y(_4552_));
 sg13g2_nand4_1 _5464_ (.B(_4299_),
    .C(_4301_),
    .A(_4260_),
    .Y(_4553_),
    .D(_4472_));
 sg13g2_nand4_1 _5465_ (.B(_4478_),
    .C(_4479_),
    .A(_4462_),
    .Y(_4554_),
    .D(_4553_));
 sg13g2_inv_1 _5466_ (.Y(_4555_),
    .A(net276));
 sg13g2_nor3_1 _5467_ (.A(_4555_),
    .B(_4181_),
    .C(_4183_),
    .Y(_4556_));
 sg13g2_buf_1 _5468_ (.A(_4556_),
    .X(_4557_));
 sg13g2_nand3_1 _5469_ (.B(_4145_),
    .C(net123),
    .A(_0150_),
    .Y(_4558_));
 sg13g2_a221oi_1 _5470_ (.B2(_4407_),
    .C1(_4413_),
    .B1(net123),
    .A1(_4410_),
    .Y(_4559_),
    .A2(_4411_));
 sg13g2_xnor2_1 _5471_ (.Y(_4560_),
    .A(_4398_),
    .B(_4511_));
 sg13g2_a21o_1 _5472_ (.A2(_4559_),
    .A1(_4558_),
    .B1(_4560_),
    .X(_4561_));
 sg13g2_nand2_1 _5473_ (.Y(_4562_),
    .A(_4152_),
    .B(_4212_));
 sg13g2_buf_1 _5474_ (.A(_4562_),
    .X(_4563_));
 sg13g2_and3_1 _5475_ (.X(_4564_),
    .A(_4560_),
    .B(_4558_),
    .C(_4559_));
 sg13g2_a221oi_1 _5476_ (.B2(_4563_),
    .C1(_4564_),
    .B1(_4561_),
    .A1(_4552_),
    .Y(_4565_),
    .A2(_4554_));
 sg13g2_and4_1 _5477_ (.A(_4462_),
    .B(_4478_),
    .C(_4479_),
    .D(_4553_),
    .X(_4566_));
 sg13g2_nor3_1 _5478_ (.A(_4544_),
    .B(_4551_),
    .C(_4566_),
    .Y(_4567_));
 sg13g2_a21o_1 _5479_ (.A2(_4559_),
    .A1(_4558_),
    .B1(_4563_),
    .X(_4568_));
 sg13g2_or2_1 _5480_ (.X(_4569_),
    .B(_4560_),
    .A(_4563_));
 sg13g2_and4_1 _5481_ (.A(_4567_),
    .B(_4561_),
    .C(_4568_),
    .D(_4569_),
    .X(_4570_));
 sg13g2_buf_1 _5482_ (.A(_4570_),
    .X(_4571_));
 sg13g2_or3_1 _5483_ (.A(_4543_),
    .B(_4565_),
    .C(_4571_),
    .X(_4572_));
 sg13g2_buf_1 _5484_ (.A(_4572_),
    .X(_4573_));
 sg13g2_o21ai_1 _5485_ (.B1(_4543_),
    .Y(_4574_),
    .A1(_4565_),
    .A2(_4571_));
 sg13g2_and2_1 _5486_ (.A(_4573_),
    .B(_4574_),
    .X(_4575_));
 sg13g2_and2_1 _5487_ (.A(net223),
    .B(net128),
    .X(_4576_));
 sg13g2_a22oi_1 _5488_ (.Y(_4577_),
    .B1(_4405_),
    .B2(net167),
    .A2(_4396_),
    .A1(net165));
 sg13g2_buf_2 _5489_ (.A(_4577_),
    .X(_4578_));
 sg13g2_mux2_1 _5490_ (.A0(net275),
    .A1(_4224_),
    .S(_4578_),
    .X(_4579_));
 sg13g2_nand4_1 _5491_ (.B(net128),
    .C(net102),
    .A(net223),
    .Y(_4580_),
    .D(_4407_));
 sg13g2_o21ai_1 _5492_ (.B1(_4580_),
    .Y(_4581_),
    .A1(_4576_),
    .A2(_4579_));
 sg13g2_and2_1 _5493_ (.A(net104),
    .B(_4581_),
    .X(_4582_));
 sg13g2_xnor2_1 _5494_ (.Y(_4584_),
    .A(_4216_),
    .B(net100));
 sg13g2_o21ai_1 _5495_ (.B1(_4584_),
    .Y(_4585_),
    .A1(_4408_),
    .A2(_4414_));
 sg13g2_or3_1 _5496_ (.A(_4584_),
    .B(_4408_),
    .C(_4414_),
    .X(_4586_));
 sg13g2_buf_1 _5497_ (.A(_4586_),
    .X(_4587_));
 sg13g2_and2_1 _5498_ (.A(_4585_),
    .B(_4587_),
    .X(_4588_));
 sg13g2_or2_1 _5499_ (.X(_4589_),
    .B(_4588_),
    .A(_4582_));
 sg13g2_nand2_1 _5500_ (.Y(_4590_),
    .A(_4563_),
    .B(_4464_));
 sg13g2_nand3_1 _5501_ (.B(_4212_),
    .C(_4511_),
    .A(_4153_),
    .Y(_4591_));
 sg13g2_o21ai_1 _5502_ (.B1(net294),
    .Y(_4592_),
    .A1(net144),
    .A2(net123));
 sg13g2_a21oi_1 _5503_ (.A1(net144),
    .A2(net123),
    .Y(_4593_),
    .B1(_4398_));
 sg13g2_nand2_1 _5504_ (.Y(_0052_),
    .A(net165),
    .B(_4396_));
 sg13g2_or4_1 _5505_ (.A(_4074_),
    .B(_4388_),
    .C(_4096_),
    .D(net165),
    .X(_0053_));
 sg13g2_o21ai_1 _5506_ (.B1(_0053_),
    .Y(_0054_),
    .A1(_4105_),
    .A2(_0052_));
 sg13g2_nand3_1 _5507_ (.B(_4096_),
    .C(_4105_),
    .A(net295),
    .Y(_0055_));
 sg13g2_nand3_1 _5508_ (.B(net167),
    .C(_4077_),
    .A(net303),
    .Y(_0056_));
 sg13g2_nand4_1 _5509_ (.B(_1380_),
    .C(_4124_),
    .A(net294),
    .Y(_0057_),
    .D(_4129_));
 sg13g2_a21oi_1 _5510_ (.A1(_0055_),
    .A2(_0056_),
    .Y(_0058_),
    .B1(_0057_));
 sg13g2_a221oi_1 _5511_ (.B2(net123),
    .C1(_0058_),
    .B1(_0054_),
    .A1(_4592_),
    .Y(_0059_),
    .A2(_4593_));
 sg13g2_buf_1 _5512_ (.A(_0059_),
    .X(_0060_));
 sg13g2_a21o_1 _5513_ (.A2(_4591_),
    .A1(_4590_),
    .B1(_0060_),
    .X(_0061_));
 sg13g2_buf_1 _5514_ (.A(_0061_),
    .X(_0063_));
 sg13g2_a21oi_1 _5515_ (.A1(_4153_),
    .A2(_4212_),
    .Y(_0064_),
    .B1(_4464_));
 sg13g2_nor2_1 _5516_ (.A(_4563_),
    .B(_4511_),
    .Y(_0065_));
 sg13g2_o21ai_1 _5517_ (.B1(_0060_),
    .Y(_0066_),
    .A1(_0064_),
    .A2(_0065_));
 sg13g2_buf_1 _5518_ (.A(_0066_),
    .X(_0067_));
 sg13g2_and4_1 _5519_ (.A(_4175_),
    .B(_4581_),
    .C(_4585_),
    .D(_4587_),
    .X(_0068_));
 sg13g2_a21o_1 _5520_ (.A2(_0067_),
    .A1(_0063_),
    .B1(_0068_),
    .X(_0069_));
 sg13g2_a21oi_1 _5521_ (.A1(_4212_),
    .A2(_4174_),
    .Y(_0070_),
    .B1(_4446_));
 sg13g2_a21oi_1 _5522_ (.A1(_4454_),
    .A2(_4399_),
    .Y(_0071_),
    .B1(_0070_));
 sg13g2_or3_1 _5523_ (.A(_4154_),
    .B(_4399_),
    .C(_0070_),
    .X(_0072_));
 sg13g2_mux2_1 _5524_ (.A0(_0071_),
    .A1(_0072_),
    .S(_4417_),
    .X(_0074_));
 sg13g2_nor2_1 _5525_ (.A(_4217_),
    .B(_4454_),
    .Y(_0075_));
 sg13g2_nor2_1 _5526_ (.A(_4400_),
    .B(_4422_),
    .Y(_0076_));
 sg13g2_a21oi_1 _5527_ (.A1(_4417_),
    .A2(_0075_),
    .Y(_0077_),
    .B1(_0076_));
 sg13g2_a21o_1 _5528_ (.A2(_0077_),
    .A1(_0074_),
    .B1(_4451_),
    .X(_0078_));
 sg13g2_nand3_1 _5529_ (.B(_0074_),
    .C(_0077_),
    .A(_4451_),
    .Y(_0079_));
 sg13g2_a22oi_1 _5530_ (.Y(_0080_),
    .B1(_0078_),
    .B2(_0079_),
    .A2(_0069_),
    .A1(_4589_));
 sg13g2_nor2_1 _5531_ (.A(_4575_),
    .B(_0080_),
    .Y(_0081_));
 sg13g2_nand4_1 _5532_ (.B(_0069_),
    .C(_0078_),
    .A(_4589_),
    .Y(_0082_),
    .D(_0079_));
 sg13g2_nor2b_1 _5533_ (.A(_0081_),
    .B_N(_0082_),
    .Y(_0083_));
 sg13g2_or2_1 _5534_ (.X(_0085_),
    .B(_4460_),
    .A(_4452_));
 sg13g2_nor2_1 _5535_ (.A(_4486_),
    .B(_4496_),
    .Y(_0086_));
 sg13g2_xnor2_1 _5536_ (.Y(_0087_),
    .A(_0085_),
    .B(_0086_));
 sg13g2_buf_2 _5537_ (.A(_0087_),
    .X(_0088_));
 sg13g2_nor2_1 _5538_ (.A(_4314_),
    .B(_4426_),
    .Y(_0089_));
 sg13g2_a22oi_1 _5539_ (.Y(_0090_),
    .B1(_0089_),
    .B2(_4135_),
    .A2(_4435_),
    .A1(net270));
 sg13g2_buf_2 _5540_ (.A(_0090_),
    .X(_0091_));
 sg13g2_nor2_1 _5541_ (.A(_4267_),
    .B(_0091_),
    .Y(_0092_));
 sg13g2_nor2_1 _5542_ (.A(_4543_),
    .B(_4565_),
    .Y(_0093_));
 sg13g2_or2_1 _5543_ (.X(_0094_),
    .B(_0093_),
    .A(_4571_));
 sg13g2_buf_1 _5544_ (.A(_0094_),
    .X(_0096_));
 sg13g2_nand2b_1 _5545_ (.Y(_0097_),
    .B(_0096_),
    .A_N(_0092_));
 sg13g2_nor2b_1 _5546_ (.A(_0096_),
    .B_N(_0092_),
    .Y(_0098_));
 sg13g2_a21oi_1 _5547_ (.A1(_0088_),
    .A2(_0097_),
    .Y(_0099_),
    .B1(_0098_));
 sg13g2_o21ai_1 _5548_ (.B1(_0082_),
    .Y(_0100_),
    .A1(_4575_),
    .A2(_0080_));
 sg13g2_and2_1 _5549_ (.A(_0100_),
    .B(_0088_),
    .X(_0101_));
 sg13g2_nor2_1 _5550_ (.A(_0088_),
    .B(_0097_),
    .Y(_0102_));
 sg13g2_a221oi_1 _5551_ (.B2(_0098_),
    .C1(_0102_),
    .B1(_0101_),
    .A1(_0083_),
    .Y(_0103_),
    .A2(_0099_));
 sg13g2_xnor2_1 _5552_ (.Y(_0104_),
    .A(_4509_),
    .B(_0103_));
 sg13g2_buf_1 _5553_ (.A(_0104_),
    .X(_0105_));
 sg13g2_xor2_1 _5554_ (.B(_0092_),
    .A(_0096_),
    .X(_0107_));
 sg13g2_xnor2_1 _5555_ (.Y(_0108_),
    .A(_0088_),
    .B(_0107_));
 sg13g2_xnor2_1 _5556_ (.Y(_0109_),
    .A(_0083_),
    .B(_0108_));
 sg13g2_nand2_1 _5557_ (.Y(_0110_),
    .A(_4582_),
    .B(_4588_));
 sg13g2_a22oi_1 _5558_ (.Y(_0111_),
    .B1(_4585_),
    .B2(_4587_),
    .A2(_4581_),
    .A1(_4175_));
 sg13g2_nand3b_1 _5559_ (.B(_0067_),
    .C(_0063_),
    .Y(_0112_),
    .A_N(_0111_));
 sg13g2_a22oi_1 _5560_ (.Y(_0113_),
    .B1(_4573_),
    .B2(_4574_),
    .A2(_0112_),
    .A1(_0110_));
 sg13g2_and4_1 _5561_ (.A(_0110_),
    .B(_0112_),
    .C(_4573_),
    .D(_4574_),
    .X(_0114_));
 sg13g2_and2_1 _5562_ (.A(_0078_),
    .B(_0079_),
    .X(_0115_));
 sg13g2_o21ai_1 _5563_ (.B1(_0115_),
    .Y(_0116_),
    .A1(_0113_),
    .A2(_0114_));
 sg13g2_or3_1 _5564_ (.A(_0115_),
    .B(_0113_),
    .C(_0114_),
    .X(_0118_));
 sg13g2_and2_1 _5565_ (.A(_0116_),
    .B(_0118_),
    .X(_0119_));
 sg13g2_buf_8 _5566_ (.A(_0119_),
    .X(_0120_));
 sg13g2_nand3_1 _5567_ (.B(_4124_),
    .C(_4129_),
    .A(_1380_),
    .Y(_0121_));
 sg13g2_buf_1 _5568_ (.A(_0121_),
    .X(_0122_));
 sg13g2_nand3_1 _5569_ (.B(net147),
    .C(_0122_),
    .A(net259),
    .Y(_0123_));
 sg13g2_buf_1 _5570_ (.A(_0123_),
    .X(_0124_));
 sg13g2_a21o_1 _5571_ (.A2(net147),
    .A1(_0150_),
    .B1(_0122_),
    .X(_0125_));
 sg13g2_buf_1 _5572_ (.A(_0125_),
    .X(_0126_));
 sg13g2_nand2_1 _5573_ (.Y(_0127_),
    .A(_4229_),
    .B(net167));
 sg13g2_nand2_1 _5574_ (.Y(_0129_),
    .A(net148),
    .B(net176));
 sg13g2_nand2_1 _5575_ (.Y(_0130_),
    .A(net296),
    .B(_0579_));
 sg13g2_a21oi_1 _5576_ (.A1(_4150_),
    .A2(_4195_),
    .Y(_0131_),
    .B1(_0130_));
 sg13g2_o21ai_1 _5577_ (.B1(net289),
    .Y(_0132_),
    .A1(net296),
    .A2(net252));
 sg13g2_nor2_1 _5578_ (.A(net313),
    .B(_0502_),
    .Y(_0133_));
 sg13g2_nand2_1 _5579_ (.Y(_0134_),
    .A(net314),
    .B(_0337_));
 sg13g2_nand2b_1 _5580_ (.Y(_0135_),
    .B(_3976_),
    .A_N(_0134_));
 sg13g2_a21o_1 _5581_ (.A2(_4168_),
    .A1(_0381_),
    .B1(net306),
    .X(_0136_));
 sg13g2_a221oi_1 _5582_ (.B2(_0135_),
    .C1(_0136_),
    .B1(_0133_),
    .A1(net198),
    .Y(_0137_),
    .A2(_4093_));
 sg13g2_o21ai_1 _5583_ (.B1(_0137_),
    .Y(_0138_),
    .A1(_0131_),
    .A2(_0132_));
 sg13g2_buf_1 _5584_ (.A(_0138_),
    .X(_0140_));
 sg13g2_buf_1 _5585_ (.A(_0140_),
    .X(_0141_));
 sg13g2_a221oi_1 _5586_ (.B2(_0141_),
    .C1(_4216_),
    .B1(_4407_),
    .A1(_0127_),
    .Y(_0142_),
    .A2(_0129_));
 sg13g2_a21oi_2 _5587_ (.B1(_0142_),
    .Y(_0143_),
    .A2(_0126_),
    .A1(_0124_));
 sg13g2_a21o_1 _5588_ (.A2(_4195_),
    .A1(_4150_),
    .B1(_0130_),
    .X(_0144_));
 sg13g2_buf_1 _5589_ (.A(_4020_),
    .X(_0145_));
 sg13g2_a21oi_1 _5590_ (.A1(_1914_),
    .A2(net290),
    .Y(_0146_),
    .B1(net233));
 sg13g2_a21o_1 _5591_ (.A2(_0135_),
    .A1(_0133_),
    .B1(_0136_),
    .X(_0147_));
 sg13g2_a221oi_1 _5592_ (.B2(_0146_),
    .C1(_0147_),
    .B1(_0144_),
    .A1(net198),
    .Y(_0148_),
    .A2(_4093_));
 sg13g2_buf_2 _5593_ (.A(_0148_),
    .X(_0149_));
 sg13g2_a21oi_1 _5594_ (.A1(net158),
    .A2(net102),
    .Y(_0151_),
    .B1(_0149_));
 sg13g2_a221oi_1 _5595_ (.B2(net259),
    .C1(_4407_),
    .B1(net147),
    .A1(_1391_),
    .Y(_0152_),
    .A2(_4185_));
 sg13g2_and4_1 _5596_ (.A(net259),
    .B(net147),
    .C(_4578_),
    .D(_4557_),
    .X(_0153_));
 sg13g2_or3_1 _5597_ (.A(_0151_),
    .B(_0152_),
    .C(_0153_),
    .X(_0154_));
 sg13g2_buf_1 _5598_ (.A(_0154_),
    .X(_0155_));
 sg13g2_o21ai_1 _5599_ (.B1(net139),
    .Y(_0156_),
    .A1(_4547_),
    .A2(_4548_));
 sg13g2_xnor2_1 _5600_ (.Y(_0157_),
    .A(_0156_),
    .B(_4537_));
 sg13g2_xnor2_1 _5601_ (.Y(_0158_),
    .A(_4536_),
    .B(_0157_));
 sg13g2_o21ai_1 _5602_ (.B1(_0158_),
    .Y(_0159_),
    .A1(_0143_),
    .A2(_0155_));
 sg13g2_xnor2_1 _5603_ (.Y(_0160_),
    .A(net145),
    .B(_4464_));
 sg13g2_xor2_1 _5604_ (.B(_0160_),
    .A(_4541_),
    .X(_0162_));
 sg13g2_nor3_1 _5605_ (.A(_0143_),
    .B(_0155_),
    .C(_0158_),
    .Y(_0163_));
 sg13g2_a21oi_2 _5606_ (.B1(_0163_),
    .Y(_0164_),
    .A2(_0162_),
    .A1(_0159_));
 sg13g2_nand2_1 _5607_ (.Y(_0165_),
    .A(_0124_),
    .B(_0126_));
 sg13g2_nand2_1 _5608_ (.Y(_0166_),
    .A(net158),
    .B(net102));
 sg13g2_nor2_1 _5609_ (.A(_4578_),
    .B(_0149_),
    .Y(_0167_));
 sg13g2_xnor2_1 _5610_ (.Y(_0168_),
    .A(_0166_),
    .B(_0167_));
 sg13g2_xor2_1 _5611_ (.B(_0168_),
    .A(_0165_),
    .X(_0169_));
 sg13g2_mux2_1 _5612_ (.A0(net303),
    .A1(_4394_),
    .S(_4095_),
    .X(_0170_));
 sg13g2_buf_1 _5613_ (.A(_0170_),
    .X(_0171_));
 sg13g2_buf_1 _5614_ (.A(_0171_),
    .X(_0173_));
 sg13g2_nand2_1 _5615_ (.Y(_0174_),
    .A(net306),
    .B(_4082_));
 sg13g2_buf_2 _5616_ (.A(_0174_),
    .X(_0175_));
 sg13g2_and4_1 _5617_ (.A(_0425_),
    .B(net177),
    .C(_0175_),
    .D(_4069_),
    .X(_0176_));
 sg13g2_buf_1 _5618_ (.A(_0176_),
    .X(_0177_));
 sg13g2_a21oi_2 _5619_ (.B1(net255),
    .Y(_0178_),
    .A2(_0175_),
    .A1(net177));
 sg13g2_nor2_1 _5620_ (.A(net291),
    .B(net306),
    .Y(_0179_));
 sg13g2_o21ai_1 _5621_ (.B1(_0179_),
    .Y(_0180_),
    .A1(_4157_),
    .A2(_4065_));
 sg13g2_nor2b_1 _5622_ (.A(net306),
    .B_N(net291),
    .Y(_0181_));
 sg13g2_nand3_1 _5623_ (.B(_4089_),
    .C(_0181_),
    .A(net198),
    .Y(_0182_));
 sg13g2_a22oi_1 _5624_ (.Y(_0184_),
    .B1(_0180_),
    .B2(_0182_),
    .A2(_4086_),
    .A1(_4080_));
 sg13g2_nand2_1 _5625_ (.Y(_0185_),
    .A(_4157_),
    .B(_0181_));
 sg13g2_nand2_1 _5626_ (.Y(_0186_),
    .A(net198),
    .B(_0179_));
 sg13g2_a221oi_1 _5627_ (.B2(_0186_),
    .C1(net177),
    .B1(_0185_),
    .A1(_4098_),
    .Y(_0187_),
    .A2(_4084_));
 sg13g2_buf_1 _5628_ (.A(_0187_),
    .X(_0188_));
 sg13g2_nor4_1 _5629_ (.A(_0177_),
    .B(_0178_),
    .C(_0184_),
    .D(_0188_),
    .Y(_0189_));
 sg13g2_nor3_1 _5630_ (.A(net142),
    .B(_0173_),
    .C(_0189_),
    .Y(_0190_));
 sg13g2_nor2_2 _5631_ (.A(_0177_),
    .B(_0178_),
    .Y(_0191_));
 sg13g2_nor2_1 _5632_ (.A(_0184_),
    .B(_0188_),
    .Y(_0192_));
 sg13g2_nor2_1 _5633_ (.A(_0191_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_or2_1 _5634_ (.X(_0195_),
    .B(_0193_),
    .A(_0190_));
 sg13g2_a21o_1 _5635_ (.A2(_4411_),
    .A1(_4410_),
    .B1(_4413_),
    .X(_0196_));
 sg13g2_nor2_1 _5636_ (.A(_4408_),
    .B(_0196_),
    .Y(_0197_));
 sg13g2_a21o_1 _5637_ (.A2(_0195_),
    .A1(_0169_),
    .B1(_0197_),
    .X(_0198_));
 sg13g2_buf_2 _5638_ (.A(_0198_),
    .X(_0199_));
 sg13g2_xnor2_1 _5639_ (.Y(_0200_),
    .A(_0165_),
    .B(_0168_));
 sg13g2_mux2_1 _5640_ (.A0(net269),
    .A1(_4403_),
    .S(_4095_),
    .X(_0201_));
 sg13g2_buf_2 _5641_ (.A(_0201_),
    .X(_0202_));
 sg13g2_or2_1 _5642_ (.X(_0203_),
    .B(_0188_),
    .A(_0184_));
 sg13g2_buf_1 _5643_ (.A(_0203_),
    .X(_0204_));
 sg13g2_a21oi_1 _5644_ (.A1(_4173_),
    .A2(_0202_),
    .Y(_0206_),
    .B1(_0204_));
 sg13g2_or2_1 _5645_ (.X(_0207_),
    .B(_0206_),
    .A(_0191_));
 sg13g2_xnor2_1 _5646_ (.Y(_0208_),
    .A(_0196_),
    .B(_0141_));
 sg13g2_nor2_1 _5647_ (.A(_4578_),
    .B(_4576_),
    .Y(_0209_));
 sg13g2_a22oi_1 _5648_ (.Y(_0210_),
    .B1(_0208_),
    .B2(_0209_),
    .A2(_0207_),
    .A1(_0200_));
 sg13g2_buf_1 _5649_ (.A(_0210_),
    .X(_0211_));
 sg13g2_a21o_1 _5650_ (.A2(_0126_),
    .A1(_0124_),
    .B1(_0142_),
    .X(_0212_));
 sg13g2_nor3_1 _5651_ (.A(_0151_),
    .B(_0152_),
    .C(_0153_),
    .Y(_0213_));
 sg13g2_a21oi_1 _5652_ (.A1(_0212_),
    .A2(_0213_),
    .Y(_0214_),
    .B1(_0158_));
 sg13g2_nand2_1 _5653_ (.Y(_0215_),
    .A(net157),
    .B(net138));
 sg13g2_xnor2_1 _5654_ (.Y(_0217_),
    .A(_0215_),
    .B(_0157_));
 sg13g2_nor3_1 _5655_ (.A(_0143_),
    .B(_0155_),
    .C(_0217_),
    .Y(_0218_));
 sg13g2_o21ai_1 _5656_ (.B1(_0162_),
    .Y(_0219_),
    .A1(_0214_),
    .A2(_0218_));
 sg13g2_xnor2_1 _5657_ (.Y(_0220_),
    .A(_4541_),
    .B(_0160_));
 sg13g2_o21ai_1 _5658_ (.B1(_0217_),
    .Y(_0221_),
    .A1(_0143_),
    .A2(_0155_));
 sg13g2_nand3_1 _5659_ (.B(_0213_),
    .C(_0158_),
    .A(_0212_),
    .Y(_0222_));
 sg13g2_nand3_1 _5660_ (.B(_0221_),
    .C(_0222_),
    .A(_0220_),
    .Y(_0223_));
 sg13g2_nand4_1 _5661_ (.B(_0211_),
    .C(_0219_),
    .A(_0199_),
    .Y(_0224_),
    .D(_0223_));
 sg13g2_a21oi_1 _5662_ (.A1(net259),
    .A2(net147),
    .Y(_0225_),
    .B1(_0149_));
 sg13g2_nand2_1 _5663_ (.Y(_0226_),
    .A(_4224_),
    .B(_4407_));
 sg13g2_nand4_1 _5664_ (.B(net147),
    .C(net142),
    .A(_0161_),
    .Y(_0228_),
    .D(_4407_));
 sg13g2_o21ai_1 _5665_ (.B1(_0228_),
    .Y(_0229_),
    .A1(_0225_),
    .A2(_0226_));
 sg13g2_buf_1 _5666_ (.A(_4196_),
    .X(_0230_));
 sg13g2_a21o_1 _5667_ (.A2(net147),
    .A1(_0161_),
    .B1(net232),
    .X(_0231_));
 sg13g2_nand2_2 _5668_ (.Y(_0232_),
    .A(net127),
    .B(_4235_));
 sg13g2_a21oi_1 _5669_ (.A1(_4407_),
    .A2(_0231_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_o21ai_1 _5670_ (.B1(_4415_),
    .Y(_0234_),
    .A1(_0229_),
    .A2(_0233_));
 sg13g2_or3_1 _5671_ (.A(_4415_),
    .B(_0229_),
    .C(_0233_),
    .X(_0235_));
 sg13g2_buf_1 _5672_ (.A(_0235_),
    .X(_0236_));
 sg13g2_and4_1 _5673_ (.A(_0063_),
    .B(_0067_),
    .C(_0234_),
    .D(_0236_),
    .X(_0237_));
 sg13g2_buf_1 _5674_ (.A(_0237_),
    .X(_0239_));
 sg13g2_a22oi_1 _5675_ (.Y(_0240_),
    .B1(_0234_),
    .B2(_0236_),
    .A2(_0067_),
    .A1(_0063_));
 sg13g2_a21oi_1 _5676_ (.A1(_0221_),
    .A2(_0222_),
    .Y(_0241_),
    .B1(_0220_));
 sg13g2_nor3_1 _5677_ (.A(_0162_),
    .B(_0214_),
    .C(_0218_),
    .Y(_0242_));
 sg13g2_or4_1 _5678_ (.A(_0239_),
    .B(_0240_),
    .C(_0241_),
    .D(_0242_),
    .X(_0243_));
 sg13g2_buf_1 _5679_ (.A(_0243_),
    .X(_0244_));
 sg13g2_a21oi_1 _5680_ (.A1(_0169_),
    .A2(_0195_),
    .Y(_0245_),
    .B1(_0197_));
 sg13g2_nor2_1 _5681_ (.A(_0191_),
    .B(_0206_),
    .Y(_0246_));
 sg13g2_nand2_1 _5682_ (.Y(_0247_),
    .A(_0208_),
    .B(_0209_));
 sg13g2_o21ai_1 _5683_ (.B1(_0247_),
    .Y(_0248_),
    .A1(_0169_),
    .A2(_0246_));
 sg13g2_or4_1 _5684_ (.A(_0245_),
    .B(_0248_),
    .C(_0239_),
    .D(_0240_),
    .X(_0250_));
 sg13g2_buf_1 _5685_ (.A(_0250_),
    .X(_0251_));
 sg13g2_nand4_1 _5686_ (.B(_0224_),
    .C(_0244_),
    .A(_0164_),
    .Y(_0252_),
    .D(_0251_));
 sg13g2_a21oi_1 _5687_ (.A1(_4511_),
    .A2(_4532_),
    .Y(_0253_),
    .B1(_4549_));
 sg13g2_nor2_2 _5688_ (.A(_4533_),
    .B(_0253_),
    .Y(_0254_));
 sg13g2_inv_1 _5689_ (.Y(_0255_),
    .A(_0254_));
 sg13g2_a22oi_1 _5690_ (.Y(_0256_),
    .B1(_0219_),
    .B2(_0223_),
    .A2(_0211_),
    .A1(_0199_));
 sg13g2_or3_1 _5691_ (.A(_0239_),
    .B(_0240_),
    .C(_0164_),
    .X(_0257_));
 sg13g2_and2_1 _5692_ (.A(_0162_),
    .B(_0163_),
    .X(_0258_));
 sg13g2_nand3_1 _5693_ (.B(_0211_),
    .C(_0258_),
    .A(_0199_),
    .Y(_0259_));
 sg13g2_o21ai_1 _5694_ (.B1(_0259_),
    .Y(_0261_),
    .A1(_0256_),
    .A2(_0257_));
 sg13g2_a21oi_1 _5695_ (.A1(_0252_),
    .A2(_0255_),
    .Y(_0262_),
    .B1(_0261_));
 sg13g2_a21oi_1 _5696_ (.A1(_0116_),
    .A2(_0118_),
    .Y(_0263_),
    .B1(_0254_));
 sg13g2_nor2_1 _5697_ (.A(_0252_),
    .B(_0255_),
    .Y(_0264_));
 sg13g2_a221oi_1 _5698_ (.B2(_0261_),
    .C1(_0264_),
    .B1(_0263_),
    .A1(_0120_),
    .Y(_0265_),
    .A2(_0262_));
 sg13g2_xor2_1 _5699_ (.B(_0265_),
    .A(_0109_),
    .X(_0266_));
 sg13g2_or2_1 _5700_ (.X(_0267_),
    .B(_3342_),
    .A(net312));
 sg13g2_a221oi_1 _5701_ (.B2(_4256_),
    .C1(_0267_),
    .B1(_4111_),
    .A1(net311),
    .Y(_0268_),
    .A2(_4255_));
 sg13g2_a22oi_1 _5702_ (.Y(_0269_),
    .B1(_0268_),
    .B2(_4253_),
    .A2(_4258_),
    .A1(net274));
 sg13g2_buf_2 _5703_ (.A(_0269_),
    .X(_0270_));
 sg13g2_and4_1 _5704_ (.A(net280),
    .B(net249),
    .C(_4440_),
    .D(net197),
    .X(_0272_));
 sg13g2_or2_1 _5705_ (.X(_0273_),
    .B(net302),
    .A(_4300_));
 sg13g2_a21oi_1 _5706_ (.A1(net249),
    .A2(net197),
    .Y(_0274_),
    .B1(_0273_));
 sg13g2_o21ai_1 _5707_ (.B1(_3353_),
    .Y(_0275_),
    .A1(_0272_),
    .A2(_0274_));
 sg13g2_buf_1 _5708_ (.A(_0275_),
    .X(_0276_));
 sg13g2_nor2_1 _5709_ (.A(_0270_),
    .B(_0276_),
    .Y(_0277_));
 sg13g2_and3_1 _5710_ (.X(_0278_),
    .A(net249),
    .B(_4440_),
    .C(net197));
 sg13g2_buf_1 _5711_ (.A(_0278_),
    .X(_0279_));
 sg13g2_a21oi_1 _5712_ (.A1(_3342_),
    .A2(_4293_),
    .Y(_0280_),
    .B1(net308));
 sg13g2_a21oi_1 _5713_ (.A1(net218),
    .A2(net197),
    .Y(_0281_),
    .B1(net302));
 sg13g2_a22oi_1 _5714_ (.Y(_0283_),
    .B1(_0281_),
    .B2(_0974_),
    .A2(_0280_),
    .A1(_0279_));
 sg13g2_nand3_1 _5715_ (.B(_4139_),
    .C(_0279_),
    .A(_0974_),
    .Y(_0284_));
 sg13g2_nand3_1 _5716_ (.B(_0283_),
    .C(_0284_),
    .A(_4437_),
    .Y(_0285_));
 sg13g2_nand3_1 _5717_ (.B(_0277_),
    .C(_0285_),
    .A(_4321_),
    .Y(_0286_));
 sg13g2_nor2_1 _5718_ (.A(_0091_),
    .B(_0276_),
    .Y(_0287_));
 sg13g2_nor2_1 _5719_ (.A(_0091_),
    .B(_0270_),
    .Y(_0288_));
 sg13g2_nand2_1 _5720_ (.Y(_0289_),
    .A(_0283_),
    .B(_0284_));
 sg13g2_o21ai_1 _5721_ (.B1(_0289_),
    .Y(_0290_),
    .A1(_0287_),
    .A2(_0288_));
 sg13g2_a21o_1 _5722_ (.A2(_0290_),
    .A1(_0286_),
    .B1(_4263_),
    .X(_0291_));
 sg13g2_buf_1 _5723_ (.A(_0291_),
    .X(_0292_));
 sg13g2_nor2_1 _5724_ (.A(_4218_),
    .B(_0171_),
    .Y(_0294_));
 sg13g2_buf_1 _5725_ (.A(_0294_),
    .X(_0295_));
 sg13g2_nor2_1 _5726_ (.A(net316),
    .B(net271),
    .Y(_0296_));
 sg13g2_and3_1 _5727_ (.X(_0297_),
    .A(_4195_),
    .B(_4198_),
    .C(net176));
 sg13g2_buf_1 _5728_ (.A(_0297_),
    .X(_0298_));
 sg13g2_mux2_1 _5729_ (.A0(_0296_),
    .A1(_0298_),
    .S(_4095_),
    .X(_0299_));
 sg13g2_buf_2 _5730_ (.A(_0299_),
    .X(_0300_));
 sg13g2_nand3_1 _5731_ (.B(_0295_),
    .C(_0300_),
    .A(_0192_),
    .Y(_0301_));
 sg13g2_nor2_1 _5732_ (.A(_4165_),
    .B(_0300_),
    .Y(_0302_));
 sg13g2_a21oi_1 _5733_ (.A1(_4173_),
    .A2(_0202_),
    .Y(_0303_),
    .B1(net144));
 sg13g2_nor3_1 _5734_ (.A(net158),
    .B(net142),
    .C(_0171_),
    .Y(_0305_));
 sg13g2_or4_1 _5735_ (.A(net275),
    .B(_0302_),
    .C(_0303_),
    .D(_0305_),
    .X(_0306_));
 sg13g2_and2_1 _5736_ (.A(_0301_),
    .B(_0306_),
    .X(_0307_));
 sg13g2_buf_1 _5737_ (.A(_0307_),
    .X(_0308_));
 sg13g2_a21o_1 _5738_ (.A2(_0289_),
    .A1(net139),
    .B1(_0277_),
    .X(_0309_));
 sg13g2_or2_1 _5739_ (.X(_0310_),
    .B(_0276_),
    .A(_4263_));
 sg13g2_and2_1 _5740_ (.A(_4472_),
    .B(_0270_),
    .X(_0311_));
 sg13g2_and2_1 _5741_ (.A(_0283_),
    .B(_0284_),
    .X(_0312_));
 sg13g2_a21oi_1 _5742_ (.A1(net157),
    .A2(_4431_),
    .Y(_0313_),
    .B1(net138));
 sg13g2_a22oi_1 _5743_ (.Y(_0314_),
    .B1(_0312_),
    .B2(_0313_),
    .A2(_0311_),
    .A1(_0310_));
 sg13g2_a21oi_2 _5744_ (.B1(_0314_),
    .Y(_0316_),
    .A2(_0309_),
    .A1(net157));
 sg13g2_a21oi_2 _5745_ (.B1(_0316_),
    .Y(_0317_),
    .A2(_0308_),
    .A1(_0292_));
 sg13g2_a21o_1 _5746_ (.A2(_0309_),
    .A1(net157),
    .B1(_0314_),
    .X(_0318_));
 sg13g2_nor3_1 _5747_ (.A(_0302_),
    .B(_0303_),
    .C(_0305_),
    .Y(_0319_));
 sg13g2_nand2_2 _5748_ (.Y(_0320_),
    .A(_4173_),
    .B(_0202_));
 sg13g2_nand2_1 _5749_ (.Y(_0321_),
    .A(_4212_),
    .B(_4234_));
 sg13g2_nor3_1 _5750_ (.A(_0204_),
    .B(_0320_),
    .C(_0321_),
    .Y(_0322_));
 sg13g2_a221oi_1 _5751_ (.B2(_0230_),
    .C1(_0322_),
    .B1(_0319_),
    .A1(_0318_),
    .Y(_0323_),
    .A2(_0292_));
 sg13g2_nand2_1 _5752_ (.Y(_0324_),
    .A(_0286_),
    .B(_0290_));
 sg13g2_a221oi_1 _5753_ (.B2(_0306_),
    .C1(_0316_),
    .B1(_0301_),
    .A1(net157),
    .Y(_0325_),
    .A2(_0324_));
 sg13g2_nor2_1 _5754_ (.A(_0191_),
    .B(_0321_),
    .Y(_0327_));
 sg13g2_xnor2_1 _5755_ (.Y(_0328_),
    .A(net144),
    .B(_0300_));
 sg13g2_or2_1 _5756_ (.X(_0329_),
    .B(_0178_),
    .A(_0177_));
 sg13g2_nand3_1 _5757_ (.B(_0329_),
    .C(_0300_),
    .A(net144),
    .Y(_0330_));
 sg13g2_o21ai_1 _5758_ (.B1(_0330_),
    .Y(_0331_),
    .A1(_4216_),
    .A2(_0328_));
 sg13g2_nor2_1 _5759_ (.A(net275),
    .B(_0320_),
    .Y(_0332_));
 sg13g2_nor3_1 _5760_ (.A(net142),
    .B(_0192_),
    .C(_0173_),
    .Y(_0333_));
 sg13g2_nor4_1 _5761_ (.A(_0329_),
    .B(_0206_),
    .C(_0333_),
    .D(_0300_),
    .Y(_0334_));
 sg13g2_a221oi_1 _5762_ (.B2(_0332_),
    .C1(_0334_),
    .B1(_0331_),
    .A1(_0206_),
    .Y(_0335_),
    .A2(_0327_));
 sg13g2_o21ai_1 _5763_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0323_),
    .A2(_0325_));
 sg13g2_buf_1 _5764_ (.A(_0336_),
    .X(_0338_));
 sg13g2_or3_1 _5765_ (.A(_0335_),
    .B(_0323_),
    .C(_0325_),
    .X(_0339_));
 sg13g2_buf_1 _5766_ (.A(_0339_),
    .X(_0340_));
 sg13g2_nand2_1 _5767_ (.Y(_0341_),
    .A(_0204_),
    .B(net62));
 sg13g2_nor2_2 _5768_ (.A(_4216_),
    .B(_4224_),
    .Y(_0342_));
 sg13g2_o21ai_1 _5769_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0190_),
    .A2(_0193_));
 sg13g2_or3_1 _5770_ (.A(_0342_),
    .B(_0190_),
    .C(_0193_),
    .X(_0344_));
 sg13g2_nand3_1 _5771_ (.B(_0343_),
    .C(_0344_),
    .A(_0341_),
    .Y(_0345_));
 sg13g2_nand3_1 _5772_ (.B(_0204_),
    .C(net62),
    .A(_0342_),
    .Y(_0346_));
 sg13g2_nand3_1 _5773_ (.B(_0345_),
    .C(_0346_),
    .A(net123),
    .Y(_0347_));
 sg13g2_and3_1 _5774_ (.X(_0349_),
    .A(_0341_),
    .B(_0343_),
    .C(_0344_));
 sg13g2_nor3_1 _5775_ (.A(_0166_),
    .B(_0192_),
    .C(_0320_),
    .Y(_0350_));
 sg13g2_o21ai_1 _5776_ (.B1(_0122_),
    .Y(_0351_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_nand3_1 _5777_ (.B(_0347_),
    .C(_0351_),
    .A(_0340_),
    .Y(_0352_));
 sg13g2_and2_1 _5778_ (.A(_0338_),
    .B(_0352_),
    .X(_0353_));
 sg13g2_buf_1 _5779_ (.A(_0353_),
    .X(_0354_));
 sg13g2_nand2_1 _5780_ (.Y(_0355_),
    .A(_0317_),
    .B(_0354_));
 sg13g2_nand3_1 _5781_ (.B(_0244_),
    .C(_0251_),
    .A(_0224_),
    .Y(_0356_));
 sg13g2_xnor2_1 _5782_ (.Y(_0357_),
    .A(_0164_),
    .B(_0254_));
 sg13g2_xnor2_1 _5783_ (.Y(_0358_),
    .A(_0356_),
    .B(_0357_));
 sg13g2_xor2_1 _5784_ (.B(_0358_),
    .A(_0120_),
    .X(_0360_));
 sg13g2_xnor2_1 _5785_ (.Y(_0361_),
    .A(_4563_),
    .B(_0060_));
 sg13g2_xnor2_1 _5786_ (.Y(_0362_),
    .A(net145),
    .B(_0361_));
 sg13g2_nand3_1 _5787_ (.B(_0211_),
    .C(_0362_),
    .A(_0199_),
    .Y(_0363_));
 sg13g2_xnor2_1 _5788_ (.Y(_0364_),
    .A(net140),
    .B(_0361_));
 sg13g2_o21ai_1 _5789_ (.B1(_0364_),
    .Y(_0365_),
    .A1(_0245_),
    .A2(_0248_));
 sg13g2_and2_1 _5790_ (.A(_0234_),
    .B(_0236_),
    .X(_0366_));
 sg13g2_nor2_1 _5791_ (.A(_0214_),
    .B(_0218_),
    .Y(_0367_));
 sg13g2_xnor2_1 _5792_ (.Y(_0368_),
    .A(_0366_),
    .B(_0367_));
 sg13g2_a21oi_2 _5793_ (.B1(_0368_),
    .Y(_0369_),
    .A2(_0365_),
    .A1(_0363_));
 sg13g2_o21ai_1 _5794_ (.B1(_0362_),
    .Y(_0371_),
    .A1(_0245_),
    .A2(_0248_));
 sg13g2_nand3_1 _5795_ (.B(_0211_),
    .C(_0364_),
    .A(_0199_),
    .Y(_0372_));
 sg13g2_xor2_1 _5796_ (.B(_0367_),
    .A(_0366_),
    .X(_0373_));
 sg13g2_a21oi_2 _5797_ (.B1(_0373_),
    .Y(_0374_),
    .A2(_0372_),
    .A1(_0371_));
 sg13g2_nor2_1 _5798_ (.A(_0369_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_or2_1 _5799_ (.X(_0376_),
    .B(_0375_),
    .A(_4541_));
 sg13g2_a21o_1 _5800_ (.A2(_0360_),
    .A1(_0355_),
    .B1(_0376_),
    .X(_0377_));
 sg13g2_o21ai_1 _5801_ (.B1(_0375_),
    .Y(_0378_),
    .A1(_0317_),
    .A2(_0354_));
 sg13g2_a21o_1 _5802_ (.A2(_0378_),
    .A1(_0355_),
    .B1(_0360_),
    .X(_0379_));
 sg13g2_nand2_1 _5803_ (.Y(_0380_),
    .A(_0377_),
    .B(_0379_));
 sg13g2_nand2_1 _5804_ (.Y(_0382_),
    .A(_0091_),
    .B(_0270_));
 sg13g2_nand2b_1 _5805_ (.Y(_0383_),
    .B(_0117_),
    .A_N(net290));
 sg13g2_a21oi_2 _5806_ (.B1(_0383_),
    .Y(_0384_),
    .A2(_3998_),
    .A1(_3976_));
 sg13g2_nor2_1 _5807_ (.A(net208),
    .B(_0384_),
    .Y(_0385_));
 sg13g2_nor3_1 _5808_ (.A(net316),
    .B(net271),
    .C(net303),
    .Y(_0386_));
 sg13g2_mux2_1 _5809_ (.A0(_0298_),
    .A1(_0386_),
    .S(net167),
    .X(_0387_));
 sg13g2_mux2_1 _5810_ (.A0(net282),
    .A1(_4300_),
    .S(net166),
    .X(_0388_));
 sg13g2_nor2_2 _5811_ (.A(_3342_),
    .B(_0388_),
    .Y(_0389_));
 sg13g2_a21o_1 _5812_ (.A2(_0387_),
    .A1(_0385_),
    .B1(_0389_),
    .X(_0390_));
 sg13g2_nand2b_1 _5813_ (.Y(_0391_),
    .B(net307),
    .A_N(_4186_));
 sg13g2_nor2_1 _5814_ (.A(net268),
    .B(_0391_),
    .Y(_0393_));
 sg13g2_buf_1 _5815_ (.A(_4186_),
    .X(_0394_));
 sg13g2_nor2b_1 _5816_ (.A(net237),
    .B_N(net276),
    .Y(_0395_));
 sg13g2_and2_1 _5817_ (.A(net266),
    .B(_0395_),
    .X(_0396_));
 sg13g2_mux2_1 _5818_ (.A0(_0393_),
    .A1(_0396_),
    .S(net164),
    .X(_0397_));
 sg13g2_and3_1 _5819_ (.X(_0398_),
    .A(_0389_),
    .B(_0385_),
    .C(_0387_));
 sg13g2_a21o_1 _5820_ (.A2(_0397_),
    .A1(_0390_),
    .B1(_0398_),
    .X(_0399_));
 sg13g2_a21oi_2 _5821_ (.B1(_0288_),
    .Y(_0400_),
    .A2(_0399_),
    .A1(_0382_));
 sg13g2_inv_1 _5822_ (.Y(_0401_),
    .A(_0400_));
 sg13g2_nand2_1 _5823_ (.Y(_0402_),
    .A(_0345_),
    .B(_0346_));
 sg13g2_a21o_1 _5824_ (.A2(_0338_),
    .A1(_0340_),
    .B1(_0402_),
    .X(_0404_));
 sg13g2_buf_1 _5825_ (.A(_0404_),
    .X(_0405_));
 sg13g2_nand3_1 _5826_ (.B(_0402_),
    .C(_0338_),
    .A(_0340_),
    .Y(_0406_));
 sg13g2_buf_2 _5827_ (.A(_0406_),
    .X(_0407_));
 sg13g2_nand2_1 _5828_ (.Y(_0408_),
    .A(_0405_),
    .B(_0407_));
 sg13g2_xnor2_1 _5829_ (.Y(_0409_),
    .A(_0191_),
    .B(_0300_));
 sg13g2_o21ai_1 _5830_ (.B1(_0149_),
    .Y(_0410_),
    .A1(_4216_),
    .A2(_0171_));
 sg13g2_buf_1 _5831_ (.A(_0410_),
    .X(_0411_));
 sg13g2_nand3_1 _5832_ (.B(_0140_),
    .C(_0202_),
    .A(_4152_),
    .Y(_0412_));
 sg13g2_buf_1 _5833_ (.A(_0412_),
    .X(_0413_));
 sg13g2_nand2_1 _5834_ (.Y(_0415_),
    .A(_0411_),
    .B(_0413_));
 sg13g2_nand2_1 _5835_ (.Y(_0416_),
    .A(net208),
    .B(net275));
 sg13g2_or2_1 _5836_ (.X(_0417_),
    .B(net303),
    .A(net316));
 sg13g2_nand4_1 _5837_ (.B(_4195_),
    .C(_4198_),
    .A(net177),
    .Y(_0418_),
    .D(_4403_));
 sg13g2_o21ai_1 _5838_ (.B1(_0418_),
    .Y(_0419_),
    .A1(net148),
    .A2(_0417_));
 sg13g2_buf_1 _5839_ (.A(_0419_),
    .X(_0420_));
 sg13g2_and2_1 _5840_ (.A(net158),
    .B(_0420_),
    .X(_0421_));
 sg13g2_o21ai_1 _5841_ (.B1(net252),
    .Y(_0422_),
    .A1(_4147_),
    .A2(_4098_));
 sg13g2_o21ai_1 _5842_ (.B1(net294),
    .Y(_0423_),
    .A1(net250),
    .A2(_4080_));
 sg13g2_a21oi_2 _5843_ (.B1(_0423_),
    .Y(_0424_),
    .A2(_0422_),
    .A1(net250));
 sg13g2_o21ai_1 _5844_ (.B1(net102),
    .Y(_0426_),
    .A1(net98),
    .A2(_0424_));
 sg13g2_a21o_1 _5845_ (.A2(_0421_),
    .A1(_0416_),
    .B1(_0426_),
    .X(_0427_));
 sg13g2_nand3_1 _5846_ (.B(_0415_),
    .C(_0427_),
    .A(_0409_),
    .Y(_0428_));
 sg13g2_a21oi_1 _5847_ (.A1(_0415_),
    .A2(_0427_),
    .Y(_0429_),
    .B1(_0409_));
 sg13g2_nor2_1 _5848_ (.A(net289),
    .B(_4150_),
    .Y(_0430_));
 sg13g2_a221oi_1 _5849_ (.B2(_4148_),
    .C1(net306),
    .B1(_0430_),
    .A1(net289),
    .Y(_0431_),
    .A2(_4149_));
 sg13g2_buf_2 _5850_ (.A(_0431_),
    .X(_0432_));
 sg13g2_and2_1 _5851_ (.A(net98),
    .B(_0432_),
    .X(_0433_));
 sg13g2_buf_2 _5852_ (.A(_0433_),
    .X(_0434_));
 sg13g2_xnor2_1 _5853_ (.Y(_0435_),
    .A(_0420_),
    .B(_0424_));
 sg13g2_a221oi_1 _5854_ (.B2(_0413_),
    .C1(_0435_),
    .B1(_0411_),
    .A1(_0127_),
    .Y(_0437_),
    .A2(_0129_));
 sg13g2_buf_1 _5855_ (.A(_0437_),
    .X(_0438_));
 sg13g2_nor2_1 _5856_ (.A(_4440_),
    .B(net166),
    .Y(_0439_));
 sg13g2_o21ai_1 _5857_ (.B1(_4319_),
    .Y(_0440_),
    .A1(net302),
    .A2(net164));
 sg13g2_buf_1 _5858_ (.A(_4187_),
    .X(_0441_));
 sg13g2_a22oi_1 _5859_ (.Y(_0442_),
    .B1(_0440_),
    .B2(net231),
    .A2(_0439_),
    .A1(_4317_));
 sg13g2_xnor2_1 _5860_ (.Y(_0443_),
    .A(_4471_),
    .B(_0442_));
 sg13g2_xnor2_1 _5861_ (.Y(_0444_),
    .A(_0270_),
    .B(_0443_));
 sg13g2_o21ai_1 _5862_ (.B1(_0444_),
    .Y(_0445_),
    .A1(_0434_),
    .A2(_0438_));
 sg13g2_or3_1 _5863_ (.A(_0434_),
    .B(_0438_),
    .C(_0444_),
    .X(_0446_));
 sg13g2_nand3b_1 _5864_ (.B(_0445_),
    .C(_0446_),
    .Y(_0448_),
    .A_N(_0429_));
 sg13g2_nand2_1 _5865_ (.Y(_0449_),
    .A(_0428_),
    .B(_0448_));
 sg13g2_a22oi_1 _5866_ (.Y(_0450_),
    .B1(_0289_),
    .B2(net138),
    .A2(net139),
    .A1(net145));
 sg13g2_a21o_1 _5867_ (.A2(_0312_),
    .A1(_4321_),
    .B1(_0450_),
    .X(_0451_));
 sg13g2_xnor2_1 _5868_ (.Y(_0452_),
    .A(net138),
    .B(_0270_));
 sg13g2_nor2_1 _5869_ (.A(net266),
    .B(net302),
    .Y(_0453_));
 sg13g2_a22oi_1 _5870_ (.Y(_0454_),
    .B1(_0453_),
    .B2(net166),
    .A2(_0279_),
    .A1(net266));
 sg13g2_nor2_1 _5871_ (.A(_0452_),
    .B(_0454_),
    .Y(_0455_));
 sg13g2_o21ai_1 _5872_ (.B1(_0455_),
    .Y(_0456_),
    .A1(_0434_),
    .A2(_0438_));
 sg13g2_nand2b_1 _5873_ (.Y(_0457_),
    .B(_0454_),
    .A_N(_0434_));
 sg13g2_and2_1 _5874_ (.A(_0310_),
    .B(_0452_),
    .X(_0459_));
 sg13g2_o21ai_1 _5875_ (.B1(_0459_),
    .Y(_0460_),
    .A1(_0438_),
    .A2(_0457_));
 sg13g2_nand3_1 _5876_ (.B(_0456_),
    .C(_0460_),
    .A(_0451_),
    .Y(_0461_));
 sg13g2_buf_1 _5877_ (.A(_0461_),
    .X(_0462_));
 sg13g2_a21o_1 _5878_ (.A2(_0460_),
    .A1(_0456_),
    .B1(_0451_),
    .X(_0463_));
 sg13g2_buf_1 _5879_ (.A(_0463_),
    .X(_0464_));
 sg13g2_and2_1 _5880_ (.A(_0462_),
    .B(_0464_),
    .X(_0465_));
 sg13g2_xnor2_1 _5881_ (.Y(_0466_),
    .A(_0449_),
    .B(_0465_));
 sg13g2_xnor2_1 _5882_ (.Y(_0467_),
    .A(_0408_),
    .B(_0466_));
 sg13g2_xor2_1 _5883_ (.B(_0443_),
    .A(_0434_),
    .X(_0468_));
 sg13g2_xnor2_1 _5884_ (.Y(_0470_),
    .A(_0415_),
    .B(_0468_));
 sg13g2_xnor2_1 _5885_ (.Y(_0471_),
    .A(_0409_),
    .B(_0470_));
 sg13g2_xor2_1 _5886_ (.B(_0399_),
    .A(_0091_),
    .X(_0472_));
 sg13g2_nand3_1 _5887_ (.B(_0298_),
    .C(_0385_),
    .A(net148),
    .Y(_0473_));
 sg13g2_nand2_1 _5888_ (.Y(_0474_),
    .A(net166),
    .B(_0393_));
 sg13g2_nand2_1 _5889_ (.Y(_0475_),
    .A(net164),
    .B(_0396_));
 sg13g2_inv_1 _5890_ (.Y(_0476_),
    .A(_0386_));
 sg13g2_nor3_1 _5891_ (.A(net208),
    .B(_0384_),
    .C(_0476_),
    .Y(_0477_));
 sg13g2_a22oi_1 _5892_ (.Y(_0478_),
    .B1(_0477_),
    .B2(net159),
    .A2(_0475_),
    .A1(_0474_));
 sg13g2_nand2b_1 _5893_ (.Y(_0479_),
    .B(net259),
    .A_N(_0384_));
 sg13g2_nor2_1 _5894_ (.A(_0479_),
    .B(_0397_),
    .Y(_0481_));
 sg13g2_a22oi_1 _5895_ (.Y(_0482_),
    .B1(_0481_),
    .B2(_0387_),
    .A2(_0478_),
    .A1(_0473_));
 sg13g2_buf_1 _5896_ (.A(_0482_),
    .X(_0483_));
 sg13g2_xnor2_1 _5897_ (.Y(_0484_),
    .A(_0389_),
    .B(_0483_));
 sg13g2_o21ai_1 _5898_ (.B1(net208),
    .Y(_0485_),
    .A1(net275),
    .A2(_4224_));
 sg13g2_nor2_1 _5899_ (.A(net98),
    .B(_0424_),
    .Y(_0486_));
 sg13g2_a21oi_2 _5900_ (.B1(_0486_),
    .Y(_0487_),
    .A2(_0485_),
    .A1(_0421_));
 sg13g2_nand2_2 _5901_ (.Y(_0488_),
    .A(_0484_),
    .B(_0487_));
 sg13g2_xnor2_1 _5902_ (.Y(_0489_),
    .A(_0472_),
    .B(_0488_));
 sg13g2_xnor2_1 _5903_ (.Y(_0490_),
    .A(_0471_),
    .B(_0489_));
 sg13g2_nand2_2 _5904_ (.Y(_0492_),
    .A(net138),
    .B(_4442_));
 sg13g2_nand3_1 _5905_ (.B(_4229_),
    .C(net269),
    .A(net259),
    .Y(_0493_));
 sg13g2_nand2_1 _5906_ (.Y(_0494_),
    .A(net259),
    .B(_4082_));
 sg13g2_mux2_1 _5907_ (.A0(_0493_),
    .A1(_0494_),
    .S(net148),
    .X(_0495_));
 sg13g2_and2_1 _5908_ (.A(net268),
    .B(_0391_),
    .X(_0496_));
 sg13g2_or3_1 _5909_ (.A(net164),
    .B(_0393_),
    .C(_0496_),
    .X(_0497_));
 sg13g2_buf_1 _5910_ (.A(_0497_),
    .X(_0498_));
 sg13g2_nand2_1 _5911_ (.Y(_0499_),
    .A(net276),
    .B(_4186_));
 sg13g2_a21oi_1 _5912_ (.A1(_4120_),
    .A2(_0499_),
    .Y(_0500_),
    .B1(_1281_));
 sg13g2_and3_1 _5913_ (.X(_0501_),
    .A(_1281_),
    .B(_4120_),
    .C(_0499_));
 sg13g2_o21ai_1 _5914_ (.B1(net164),
    .Y(_0503_),
    .A1(_0500_),
    .A2(_0501_));
 sg13g2_and2_1 _5915_ (.A(_0498_),
    .B(_0503_),
    .X(_0504_));
 sg13g2_buf_1 _5916_ (.A(_0504_),
    .X(_0505_));
 sg13g2_or3_1 _5917_ (.A(net103),
    .B(_0495_),
    .C(_0505_),
    .X(_0506_));
 sg13g2_buf_2 _5918_ (.A(_0506_),
    .X(_0507_));
 sg13g2_xor2_1 _5919_ (.B(_0507_),
    .A(_0492_),
    .X(_0508_));
 sg13g2_nand2_1 _5920_ (.Y(_0509_),
    .A(net269),
    .B(net159));
 sg13g2_nand3_1 _5921_ (.B(_0498_),
    .C(_0503_),
    .A(net316),
    .Y(_0510_));
 sg13g2_a21oi_1 _5922_ (.A1(_4195_),
    .A2(_4198_),
    .Y(_0511_),
    .B1(_1632_));
 sg13g2_nand4_1 _5923_ (.B(_0498_),
    .C(_0503_),
    .A(_4097_),
    .Y(_0512_),
    .D(_0511_));
 sg13g2_o21ai_1 _5924_ (.B1(_0512_),
    .Y(_0514_),
    .A1(_0509_),
    .A2(_0510_));
 sg13g2_nand2_1 _5925_ (.Y(_0515_),
    .A(_4392_),
    .B(net130));
 sg13g2_o21ai_1 _5926_ (.B1(_0515_),
    .Y(_0516_),
    .A1(_0172_),
    .A2(_0509_));
 sg13g2_o21ai_1 _5927_ (.B1(_4235_),
    .Y(_0517_),
    .A1(_0514_),
    .A2(_0516_));
 sg13g2_nor2_1 _5928_ (.A(_1730_),
    .B(_4201_),
    .Y(_0518_));
 sg13g2_nor2_1 _5929_ (.A(net303),
    .B(_0479_),
    .Y(_0519_));
 sg13g2_nand3_1 _5930_ (.B(_4228_),
    .C(_0479_),
    .A(_4097_),
    .Y(_0520_));
 sg13g2_o21ai_1 _5931_ (.B1(_0520_),
    .Y(_0521_),
    .A1(_0127_),
    .A2(_0519_));
 sg13g2_nor2_1 _5932_ (.A(net288),
    .B(net293),
    .Y(_0522_));
 sg13g2_nand2_1 _5933_ (.Y(_0523_),
    .A(net295),
    .B(_0522_));
 sg13g2_nand2_1 _5934_ (.Y(_0525_),
    .A(net303),
    .B(_0296_));
 sg13g2_mux2_1 _5935_ (.A0(_0523_),
    .A1(_0525_),
    .S(net159),
    .X(_0526_));
 sg13g2_o21ai_1 _5936_ (.B1(_0505_),
    .Y(_0527_),
    .A1(_1730_),
    .A2(_0526_));
 sg13g2_o21ai_1 _5937_ (.B1(_0527_),
    .Y(_0528_),
    .A1(_0518_),
    .A2(_0521_));
 sg13g2_nand2_1 _5938_ (.Y(_0529_),
    .A(_0517_),
    .B(_0528_));
 sg13g2_xor2_1 _5939_ (.B(_0487_),
    .A(_0483_),
    .X(_0530_));
 sg13g2_nor3_1 _5940_ (.A(_0508_),
    .B(_0529_),
    .C(_0530_),
    .Y(_0531_));
 sg13g2_xnor2_1 _5941_ (.Y(_0532_),
    .A(_0492_),
    .B(_0507_));
 sg13g2_xnor2_1 _5942_ (.Y(_0533_),
    .A(_0483_),
    .B(_0487_));
 sg13g2_buf_2 _5943_ (.A(_0533_),
    .X(_0534_));
 sg13g2_nor3_1 _5944_ (.A(_0532_),
    .B(_0529_),
    .C(_0534_),
    .Y(_0536_));
 sg13g2_nor4_1 _5945_ (.A(_3579_),
    .B(_0388_),
    .C(_0532_),
    .D(_0530_),
    .Y(_0537_));
 sg13g2_nor3_1 _5946_ (.A(_0389_),
    .B(_0508_),
    .C(_0534_),
    .Y(_0538_));
 sg13g2_nor4_1 _5947_ (.A(_0531_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0539_));
 sg13g2_nor2_1 _5948_ (.A(_0492_),
    .B(_0507_),
    .Y(_0540_));
 sg13g2_nor2_1 _5949_ (.A(_0389_),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_and2_1 _5950_ (.A(_0492_),
    .B(_0507_),
    .X(_0542_));
 sg13g2_buf_1 _5951_ (.A(_0542_),
    .X(_0543_));
 sg13g2_nor2_1 _5952_ (.A(_0541_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_a21o_1 _5953_ (.A2(_0539_),
    .A1(_0490_),
    .B1(_0544_),
    .X(_0545_));
 sg13g2_o21ai_1 _5954_ (.B1(_0545_),
    .Y(_0547_),
    .A1(_0490_),
    .A2(_0539_));
 sg13g2_buf_1 _5955_ (.A(_0547_),
    .X(_0548_));
 sg13g2_nand2_1 _5956_ (.Y(_0549_),
    .A(_0467_),
    .B(_0548_));
 sg13g2_a21o_1 _5957_ (.A2(_0308_),
    .A1(_0292_),
    .B1(_0316_),
    .X(_0550_));
 sg13g2_nand4_1 _5958_ (.B(_0340_),
    .C(_0347_),
    .A(_0550_),
    .Y(_0551_),
    .D(_0351_));
 sg13g2_or2_1 _5959_ (.X(_0552_),
    .B(_0340_),
    .A(_0550_));
 sg13g2_nand3_1 _5960_ (.B(_0308_),
    .C(_0335_),
    .A(_0316_),
    .Y(_0553_));
 sg13g2_o21ai_1 _5961_ (.B1(net123),
    .Y(_0554_),
    .A1(_0349_),
    .A2(_0350_));
 sg13g2_nand3_1 _5962_ (.B(_0345_),
    .C(_0346_),
    .A(_0122_),
    .Y(_0555_));
 sg13g2_nand4_1 _5963_ (.B(_0554_),
    .C(_0555_),
    .A(_0317_),
    .Y(_0556_),
    .D(_0338_));
 sg13g2_nand4_1 _5964_ (.B(_0552_),
    .C(_0553_),
    .A(_0551_),
    .Y(_0558_),
    .D(_0556_));
 sg13g2_nor3_1 _5965_ (.A(_0369_),
    .B(_0374_),
    .C(_0558_),
    .Y(_0559_));
 sg13g2_a21o_1 _5966_ (.A2(_0365_),
    .A1(_0363_),
    .B1(_0368_),
    .X(_0560_));
 sg13g2_buf_1 _5967_ (.A(_0560_),
    .X(_0561_));
 sg13g2_a21o_1 _5968_ (.A2(_0372_),
    .A1(_0371_),
    .B1(_0373_),
    .X(_0562_));
 sg13g2_buf_1 _5969_ (.A(_0562_),
    .X(_0563_));
 sg13g2_and4_1 _5970_ (.A(_0551_),
    .B(_0552_),
    .C(_0553_),
    .D(_0556_),
    .X(_0564_));
 sg13g2_a21oi_1 _5971_ (.A1(_0561_),
    .A2(_0563_),
    .Y(_0565_),
    .B1(_0564_));
 sg13g2_nand2_1 _5972_ (.Y(_0566_),
    .A(net123),
    .B(_0462_));
 sg13g2_nand2_1 _5973_ (.Y(_0567_),
    .A(_0464_),
    .B(_0566_));
 sg13g2_inv_1 _5974_ (.Y(_0569_),
    .A(_0567_));
 sg13g2_o21ai_1 _5975_ (.B1(_0569_),
    .Y(_0570_),
    .A1(_0559_),
    .A2(_0565_));
 sg13g2_nand3_1 _5976_ (.B(_0563_),
    .C(_0564_),
    .A(_0561_),
    .Y(_0571_));
 sg13g2_o21ai_1 _5977_ (.B1(_0558_),
    .Y(_0572_),
    .A1(_0369_),
    .A2(_0374_));
 sg13g2_nand3_1 _5978_ (.B(_0572_),
    .C(_0567_),
    .A(_0571_),
    .Y(_0573_));
 sg13g2_nand2_1 _5979_ (.Y(_0574_),
    .A(_0462_),
    .B(_0464_));
 sg13g2_and4_1 _5980_ (.A(_0405_),
    .B(_0407_),
    .C(_0449_),
    .D(_0574_),
    .X(_0575_));
 sg13g2_a221oi_1 _5981_ (.B2(_0448_),
    .C1(_0574_),
    .B1(_0428_),
    .A1(_0405_),
    .Y(_0576_),
    .A2(_0407_));
 sg13g2_a221oi_1 _5982_ (.B2(_0464_),
    .C1(_0122_),
    .B1(_0462_),
    .A1(_0405_),
    .Y(_0577_),
    .A2(_0407_));
 sg13g2_and4_1 _5983_ (.A(_0122_),
    .B(_0405_),
    .C(_0407_),
    .D(_0465_),
    .X(_0578_));
 sg13g2_or4_1 _5984_ (.A(_0575_),
    .B(_0576_),
    .C(_0577_),
    .D(_0578_),
    .X(_0580_));
 sg13g2_buf_1 _5985_ (.A(_0580_),
    .X(_0581_));
 sg13g2_a221oi_1 _5986_ (.B2(_0573_),
    .C1(_0581_),
    .B1(_0570_),
    .A1(_0401_),
    .Y(_0582_),
    .A2(_0549_));
 sg13g2_a21oi_1 _5987_ (.A1(_0467_),
    .A2(_0548_),
    .Y(_0583_),
    .B1(_0400_));
 sg13g2_a21oi_1 _5988_ (.A1(_0571_),
    .A2(_0572_),
    .Y(_0584_),
    .B1(_0567_));
 sg13g2_nor3_1 _5989_ (.A(_0559_),
    .B(_0565_),
    .C(_0569_),
    .Y(_0585_));
 sg13g2_inv_1 _5990_ (.Y(_0586_),
    .A(_0581_));
 sg13g2_nor4_1 _5991_ (.A(_0583_),
    .B(_0584_),
    .C(_0585_),
    .D(_0586_),
    .Y(_0587_));
 sg13g2_nor2_1 _5992_ (.A(_3438_),
    .B(net166),
    .Y(_0588_));
 sg13g2_o21ai_1 _5993_ (.B1(net203),
    .Y(_0589_),
    .A1(_4427_),
    .A2(_0588_));
 sg13g2_nor2_1 _5994_ (.A(_0492_),
    .B(_0589_),
    .Y(_0591_));
 sg13g2_buf_1 _5995_ (.A(net270),
    .X(_0592_));
 sg13g2_nor2_1 _5996_ (.A(_4555_),
    .B(net230),
    .Y(_0593_));
 sg13g2_nor2_1 _5997_ (.A(_4555_),
    .B(_4471_),
    .Y(_0594_));
 sg13g2_nor2_1 _5998_ (.A(net268),
    .B(_4423_),
    .Y(_0595_));
 sg13g2_nand2_1 _5999_ (.Y(_0596_),
    .A(_1281_),
    .B(_1402_));
 sg13g2_mux2_1 _6000_ (.A0(_0595_),
    .A1(_0596_),
    .S(net164),
    .X(_0597_));
 sg13g2_mux2_1 _6001_ (.A0(_0593_),
    .A1(_0594_),
    .S(_0597_),
    .X(_0598_));
 sg13g2_nor2_2 _6002_ (.A(_4437_),
    .B(_4425_),
    .Y(_0599_));
 sg13g2_o21ai_1 _6003_ (.B1(_0524_),
    .Y(_0600_),
    .A1(net139),
    .A2(_4442_));
 sg13g2_nand2b_1 _6004_ (.Y(_0602_),
    .B(_0600_),
    .A_N(_0599_));
 sg13g2_a21o_1 _6005_ (.A2(_0602_),
    .A1(net203),
    .B1(_0598_),
    .X(_0603_));
 sg13g2_nor2_2 _6006_ (.A(net273),
    .B(_4321_),
    .Y(_0604_));
 sg13g2_xnor2_1 _6007_ (.Y(_0605_),
    .A(net295),
    .B(net293));
 sg13g2_nand2_1 _6008_ (.Y(_0606_),
    .A(net130),
    .B(_0605_));
 sg13g2_nor2_1 _6009_ (.A(net271),
    .B(_4389_),
    .Y(_0607_));
 sg13g2_buf_1 _6010_ (.A(_4388_),
    .X(_0608_));
 sg13g2_nor2_1 _6011_ (.A(_4229_),
    .B(net265),
    .Y(_0609_));
 sg13g2_or3_1 _6012_ (.A(net130),
    .B(_0607_),
    .C(_0609_),
    .X(_0610_));
 sg13g2_nand3_1 _6013_ (.B(_0606_),
    .C(_0610_),
    .A(_0172_),
    .Y(_0611_));
 sg13g2_xnor2_1 _6014_ (.Y(_0613_),
    .A(_0604_),
    .B(_0611_));
 sg13g2_nand2_1 _6015_ (.Y(_0614_),
    .A(_4392_),
    .B(_0598_));
 sg13g2_nand2_1 _6016_ (.Y(_0615_),
    .A(_4392_),
    .B(_0604_));
 sg13g2_xnor2_1 _6017_ (.Y(_0616_),
    .A(_4425_),
    .B(_0589_));
 sg13g2_a21oi_1 _6018_ (.A1(_0614_),
    .A2(_0615_),
    .Y(_0617_),
    .B1(_0616_));
 sg13g2_a221oi_1 _6019_ (.B2(_0613_),
    .C1(_0617_),
    .B1(_0603_),
    .A1(_0598_),
    .Y(_0618_),
    .A2(_0602_));
 sg13g2_nand2b_1 _6020_ (.Y(_0619_),
    .B(_0618_),
    .A_N(_0591_));
 sg13g2_nor3_1 _6021_ (.A(net159),
    .B(_4222_),
    .C(_4403_),
    .Y(_0620_));
 sg13g2_a21oi_1 _6022_ (.A1(net159),
    .A2(_0607_),
    .Y(_0621_),
    .B1(_0620_));
 sg13g2_xor2_1 _6023_ (.B(_0621_),
    .A(_0505_),
    .X(_0622_));
 sg13g2_xnor2_1 _6024_ (.Y(_0624_),
    .A(_0518_),
    .B(_0622_));
 sg13g2_nand2_1 _6025_ (.Y(_0625_),
    .A(net223),
    .B(net102));
 sg13g2_nor2_1 _6026_ (.A(_0202_),
    .B(_0604_),
    .Y(_0626_));
 sg13g2_nand2_1 _6027_ (.Y(_0627_),
    .A(_0608_),
    .B(net159));
 sg13g2_nand4_1 _6028_ (.B(_0627_),
    .C(_0385_),
    .A(_4224_),
    .Y(_0628_),
    .D(_0604_));
 sg13g2_buf_1 _6029_ (.A(_0628_),
    .X(_0629_));
 sg13g2_o21ai_1 _6030_ (.B1(_0629_),
    .Y(_0630_),
    .A1(_0625_),
    .A2(_0626_));
 sg13g2_mux2_1 _6031_ (.A0(_0391_),
    .A1(_0499_),
    .S(net164),
    .X(_0631_));
 sg13g2_xor2_1 _6032_ (.B(_0631_),
    .A(_0599_),
    .X(_0632_));
 sg13g2_xnor2_1 _6033_ (.Y(_0633_),
    .A(_0630_),
    .B(_0632_));
 sg13g2_xnor2_1 _6034_ (.Y(_0635_),
    .A(_0624_),
    .B(_0633_));
 sg13g2_nor2b_1 _6035_ (.A(_0618_),
    .B_N(_0591_),
    .Y(_0636_));
 sg13g2_a21oi_1 _6036_ (.A1(_0619_),
    .A2(_0635_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_nor2b_1 _6037_ (.A(_0599_),
    .B_N(_0631_),
    .Y(_0638_));
 sg13g2_nand2b_1 _6038_ (.Y(_0639_),
    .B(_0599_),
    .A_N(_0631_));
 sg13g2_o21ai_1 _6039_ (.B1(_0639_),
    .Y(_0640_),
    .A1(_0629_),
    .A2(_0638_));
 sg13g2_buf_1 _6040_ (.A(_0640_),
    .X(_0641_));
 sg13g2_nor2_1 _6041_ (.A(_0530_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nor2_1 _6042_ (.A(_0534_),
    .B(_0641_),
    .Y(_0643_));
 sg13g2_and2_1 _6043_ (.A(_0517_),
    .B(_0528_),
    .X(_0644_));
 sg13g2_buf_1 _6044_ (.A(_0644_),
    .X(_0646_));
 sg13g2_xnor2_1 _6045_ (.Y(_0647_),
    .A(_0532_),
    .B(_0646_));
 sg13g2_mux2_1 _6046_ (.A0(_0642_),
    .A1(_0643_),
    .S(_0647_),
    .X(_0648_));
 sg13g2_nor2_1 _6047_ (.A(_0625_),
    .B(_0626_),
    .Y(_0649_));
 sg13g2_xor2_1 _6048_ (.B(_0632_),
    .A(_0629_),
    .X(_0650_));
 sg13g2_nand2_1 _6049_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nand2_1 _6050_ (.Y(_0652_),
    .A(_0624_),
    .B(_0651_));
 sg13g2_o21ai_1 _6051_ (.B1(_0652_),
    .Y(_0653_),
    .A1(_0649_),
    .A2(_0650_));
 sg13g2_a21oi_1 _6052_ (.A1(_0637_),
    .A2(_0648_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_nor2_1 _6053_ (.A(_0637_),
    .B(_0648_),
    .Y(_0655_));
 sg13g2_nand2b_1 _6054_ (.Y(_0657_),
    .B(_0543_),
    .A_N(_0389_));
 sg13g2_nor2_1 _6055_ (.A(_4321_),
    .B(_0276_),
    .Y(_0658_));
 sg13g2_nand3_1 _6056_ (.B(_0517_),
    .C(_0528_),
    .A(_0507_),
    .Y(_0659_));
 sg13g2_a221oi_1 _6057_ (.B2(_0659_),
    .C1(_0534_),
    .B1(_0658_),
    .A1(_0541_),
    .Y(_0660_),
    .A2(_0646_));
 sg13g2_nand2_1 _6058_ (.Y(_0661_),
    .A(_0543_),
    .B(_0646_));
 sg13g2_a22oi_1 _6059_ (.Y(_0662_),
    .B1(_0661_),
    .B2(_0534_),
    .A2(_0660_),
    .A1(_0657_));
 sg13g2_xnor2_1 _6060_ (.Y(_0663_),
    .A(_0490_),
    .B(_0662_));
 sg13g2_o21ai_1 _6061_ (.B1(_0663_),
    .Y(_0664_),
    .A1(_0654_),
    .A2(_0655_));
 sg13g2_nor2_1 _6062_ (.A(_0637_),
    .B(_0653_),
    .Y(_0665_));
 sg13g2_nand2_1 _6063_ (.Y(_0666_),
    .A(_0530_),
    .B(_0641_));
 sg13g2_nand3_1 _6064_ (.B(_0641_),
    .C(_0647_),
    .A(_0534_),
    .Y(_0668_));
 sg13g2_o21ai_1 _6065_ (.B1(_0668_),
    .Y(_0669_),
    .A1(_0647_),
    .A2(_0666_));
 sg13g2_o21ai_1 _6066_ (.B1(_0669_),
    .Y(_0670_),
    .A1(_0663_),
    .A2(_0665_));
 sg13g2_nand2_1 _6067_ (.Y(_0671_),
    .A(_0664_),
    .B(_0670_));
 sg13g2_a21oi_1 _6068_ (.A1(_0400_),
    .A2(_0467_),
    .Y(_0672_),
    .B1(_0548_));
 sg13g2_nor2_1 _6069_ (.A(net235),
    .B(_4275_),
    .Y(_0673_));
 sg13g2_nand2b_1 _6070_ (.Y(_0674_),
    .B(_0472_),
    .A_N(_0488_));
 sg13g2_nor2b_1 _6071_ (.A(_0472_),
    .B_N(_0488_),
    .Y(_0675_));
 sg13g2_a21oi_1 _6072_ (.A1(_0471_),
    .A2(_0674_),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_nor2_1 _6073_ (.A(_0472_),
    .B(_0488_),
    .Y(_0677_));
 sg13g2_nor2_1 _6074_ (.A(_0471_),
    .B(_0677_),
    .Y(_0679_));
 sg13g2_a221oi_1 _6075_ (.B2(_0488_),
    .C1(_0679_),
    .B1(_0472_),
    .A1(net238),
    .Y(_0680_),
    .A2(_4261_));
 sg13g2_a21oi_1 _6076_ (.A1(_0673_),
    .A2(_0676_),
    .Y(_0681_),
    .B1(_0680_));
 sg13g2_o21ai_1 _6077_ (.B1(_0681_),
    .Y(_0682_),
    .A1(_0400_),
    .A2(_0467_));
 sg13g2_nor3_1 _6078_ (.A(_0671_),
    .B(_0672_),
    .C(_0682_),
    .Y(_0683_));
 sg13g2_a21oi_1 _6079_ (.A1(_0664_),
    .A2(_0670_),
    .Y(_0684_),
    .B1(_0681_));
 sg13g2_nor3_1 _6080_ (.A(_0401_),
    .B(_0549_),
    .C(_0684_),
    .Y(_0685_));
 sg13g2_nor4_2 _6081_ (.A(_0582_),
    .B(_0587_),
    .C(_0683_),
    .Y(_0686_),
    .D(_0685_));
 sg13g2_a21o_1 _6082_ (.A2(_0676_),
    .A1(_0673_),
    .B1(_0680_),
    .X(_0687_));
 sg13g2_a221oi_1 _6083_ (.B2(_0687_),
    .C1(_0581_),
    .B1(_0671_),
    .A1(_0570_),
    .Y(_0688_),
    .A2(_0573_));
 sg13g2_nor4_1 _6084_ (.A(_0584_),
    .B(_0585_),
    .C(_0586_),
    .D(_0684_),
    .Y(_0690_));
 sg13g2_nor2_1 _6085_ (.A(_0467_),
    .B(_0548_),
    .Y(_0691_));
 sg13g2_o21ai_1 _6086_ (.B1(_0691_),
    .Y(_0692_),
    .A1(_0671_),
    .A2(_0687_));
 sg13g2_o21ai_1 _6087_ (.B1(_0692_),
    .Y(_0693_),
    .A1(_0688_),
    .A2(_0690_));
 sg13g2_a22oi_1 _6088_ (.Y(_0694_),
    .B1(_0567_),
    .B2(_0581_),
    .A2(_0572_),
    .A1(_0571_));
 sg13g2_a21o_1 _6089_ (.A2(_0586_),
    .A1(_0569_),
    .B1(_0694_),
    .X(_0695_));
 sg13g2_buf_1 _6090_ (.A(_0695_),
    .X(_0696_));
 sg13g2_inv_1 _6091_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_a221oi_1 _6092_ (.B2(_0693_),
    .C1(_0697_),
    .B1(_0686_),
    .A1(_0266_),
    .Y(_0698_),
    .A2(_0380_));
 sg13g2_nor3_1 _6093_ (.A(_0550_),
    .B(_0369_),
    .C(_0374_),
    .Y(_0699_));
 sg13g2_a221oi_1 _6094_ (.B2(_0563_),
    .C1(_4541_),
    .B1(_0561_),
    .A1(_0317_),
    .Y(_0701_),
    .A2(_0354_));
 sg13g2_and3_1 _6095_ (.X(_0702_),
    .A(_0354_),
    .B(_0561_),
    .C(_0563_));
 sg13g2_and3_1 _6096_ (.X(_0703_),
    .A(_4541_),
    .B(_0317_),
    .C(_0354_));
 sg13g2_nor4_1 _6097_ (.A(_0699_),
    .B(_0701_),
    .C(_0702_),
    .D(_0703_),
    .Y(_0704_));
 sg13g2_xnor2_1 _6098_ (.Y(_0705_),
    .A(_0360_),
    .B(_0704_));
 sg13g2_inv_1 _6099_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_a221oi_1 _6100_ (.B2(_0693_),
    .C1(_0706_),
    .B1(_0686_),
    .A1(_0266_),
    .Y(_0707_),
    .A2(_0380_));
 sg13g2_xnor2_1 _6101_ (.Y(_0708_),
    .A(_0109_),
    .B(_0265_));
 sg13g2_a21oi_1 _6102_ (.A1(_0377_),
    .A2(_0379_),
    .Y(_0709_),
    .B1(_0708_));
 sg13g2_nand2_1 _6103_ (.Y(_0710_),
    .A(_0696_),
    .B(_0705_));
 sg13g2_nand3_1 _6104_ (.B(_0377_),
    .C(_0379_),
    .A(_0708_),
    .Y(_0712_));
 sg13g2_o21ai_1 _6105_ (.B1(_0712_),
    .Y(_0713_),
    .A1(_0709_),
    .A2(_0710_));
 sg13g2_or4_1 _6106_ (.A(_0105_),
    .B(_0698_),
    .C(_0707_),
    .D(_0713_),
    .X(_0714_));
 sg13g2_buf_1 _6107_ (.A(_0714_),
    .X(_0715_));
 sg13g2_and4_1 _6108_ (.A(_0164_),
    .B(_0224_),
    .C(_0244_),
    .D(_0251_),
    .X(_0716_));
 sg13g2_a21oi_1 _6109_ (.A1(_0120_),
    .A2(_0716_),
    .Y(_0717_),
    .B1(_0254_));
 sg13g2_nor2_1 _6110_ (.A(_0120_),
    .B(_0716_),
    .Y(_0718_));
 sg13g2_o21ai_1 _6111_ (.B1(_0109_),
    .Y(_0719_),
    .A1(_0717_),
    .A2(_0718_));
 sg13g2_o21ai_1 _6112_ (.B1(_0261_),
    .Y(_0720_),
    .A1(_0109_),
    .A2(_0263_));
 sg13g2_nand2_2 _6113_ (.Y(_0721_),
    .A(_0719_),
    .B(_0720_));
 sg13g2_inv_1 _6114_ (.Y(_0723_),
    .A(_0721_));
 sg13g2_xor2_1 _6115_ (.B(_4310_),
    .A(_4278_),
    .X(_0724_));
 sg13g2_xnor2_1 _6116_ (.Y(_0725_),
    .A(_4273_),
    .B(_0724_));
 sg13g2_xnor2_1 _6117_ (.Y(_0726_),
    .A(_4368_),
    .B(_0725_));
 sg13g2_buf_2 _6118_ (.A(_0726_),
    .X(_0727_));
 sg13g2_a21o_1 _6119_ (.A2(_0097_),
    .A1(_0088_),
    .B1(_0098_),
    .X(_0728_));
 sg13g2_o21ai_1 _6120_ (.B1(_0088_),
    .Y(_0729_),
    .A1(_4509_),
    .A2(_0098_));
 sg13g2_nand2_1 _6121_ (.Y(_0730_),
    .A(_4509_),
    .B(_0097_));
 sg13g2_nand2_1 _6122_ (.Y(_0731_),
    .A(_0729_),
    .B(_0730_));
 sg13g2_a22oi_1 _6123_ (.Y(_0732_),
    .B1(_0731_),
    .B2(_0100_),
    .A2(_0728_),
    .A1(_4509_));
 sg13g2_buf_1 _6124_ (.A(_0732_),
    .X(_0734_));
 sg13g2_inv_1 _6125_ (.Y(_0735_),
    .A(net14));
 sg13g2_nand2_1 _6126_ (.Y(_0736_),
    .A(_0727_),
    .B(_0735_));
 sg13g2_xor2_1 _6127_ (.B(_4336_),
    .A(_4334_),
    .X(_0737_));
 sg13g2_nor2_1 _6128_ (.A(_4340_),
    .B(_4349_),
    .Y(_0738_));
 sg13g2_and2_1 _6129_ (.A(_4340_),
    .B(_4365_),
    .X(_0739_));
 sg13g2_o21ai_1 _6130_ (.B1(_4506_),
    .Y(_0740_),
    .A1(_4497_),
    .A2(_4499_));
 sg13g2_mux2_1 _6131_ (.A0(_0738_),
    .A1(_0739_),
    .S(_0740_),
    .X(_0741_));
 sg13g2_nand2_1 _6132_ (.Y(_0742_),
    .A(_4339_),
    .B(_4363_));
 sg13g2_a21oi_1 _6133_ (.A1(_4364_),
    .A2(_0742_),
    .Y(_0743_),
    .B1(_0740_));
 sg13g2_nor2_1 _6134_ (.A(_0741_),
    .B(_0743_),
    .Y(_0745_));
 sg13g2_nor3_1 _6135_ (.A(_4497_),
    .B(_4499_),
    .C(_4506_),
    .Y(_0746_));
 sg13g2_nand3_1 _6136_ (.B(_4349_),
    .C(_0746_),
    .A(_4340_),
    .Y(_0747_));
 sg13g2_nand2b_1 _6137_ (.Y(_0748_),
    .B(_4500_),
    .A_N(_4506_));
 sg13g2_or2_1 _6138_ (.X(_0749_),
    .B(_4364_),
    .A(_4340_));
 sg13g2_inv_1 _6139_ (.Y(_0750_),
    .A(_0749_));
 sg13g2_nand2_1 _6140_ (.Y(_0751_),
    .A(_0748_),
    .B(_0750_));
 sg13g2_nor2_1 _6141_ (.A(_4339_),
    .B(_4363_),
    .Y(_0752_));
 sg13g2_o21ai_1 _6142_ (.B1(_0746_),
    .Y(_0753_),
    .A1(_4365_),
    .A2(_0752_));
 sg13g2_nand4_1 _6143_ (.B(_0747_),
    .C(_0751_),
    .A(_0745_),
    .Y(_0754_),
    .D(_0753_));
 sg13g2_xnor2_1 _6144_ (.Y(_0756_),
    .A(_0737_),
    .B(_0754_));
 sg13g2_buf_1 _6145_ (.A(_0756_),
    .X(_0757_));
 sg13g2_nand2_1 _6146_ (.Y(_0758_),
    .A(_0727_),
    .B(_0757_));
 sg13g2_nand3_1 _6147_ (.B(_0696_),
    .C(_0705_),
    .A(_0105_),
    .Y(_0759_));
 sg13g2_nand3_1 _6148_ (.B(_0693_),
    .C(_0759_),
    .A(_0686_),
    .Y(_0760_));
 sg13g2_o21ai_1 _6149_ (.B1(_0105_),
    .Y(_0761_),
    .A1(_0696_),
    .A2(_0705_));
 sg13g2_nor2_1 _6150_ (.A(_0709_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_nor2b_1 _6151_ (.A(_0712_),
    .B_N(_0105_),
    .Y(_0763_));
 sg13g2_a21o_1 _6152_ (.A2(_0762_),
    .A1(_0760_),
    .B1(_0763_),
    .X(_0764_));
 sg13g2_buf_2 _6153_ (.A(_0764_),
    .X(_0765_));
 sg13g2_a221oi_1 _6154_ (.B2(_0758_),
    .C1(_0765_),
    .B1(_0736_),
    .A1(_0715_),
    .Y(_0766_),
    .A2(_0723_));
 sg13g2_nor4_1 _6155_ (.A(_0105_),
    .B(_0698_),
    .C(_0707_),
    .D(_0713_),
    .Y(_0767_));
 sg13g2_buf_2 _6156_ (.A(_0767_),
    .X(_0768_));
 sg13g2_nor2_1 _6157_ (.A(_0266_),
    .B(_0380_),
    .Y(_0769_));
 sg13g2_a221oi_1 _6158_ (.B2(_0762_),
    .C1(_0723_),
    .B1(_0760_),
    .A1(_0105_),
    .Y(_0770_),
    .A2(_0769_));
 sg13g2_nor2b_1 _6159_ (.A(_4500_),
    .B_N(_4506_),
    .Y(_0771_));
 sg13g2_mux2_1 _6160_ (.A0(_4366_),
    .A1(_4365_),
    .S(_0737_),
    .X(_0772_));
 sg13g2_xnor2_1 _6161_ (.Y(_0773_),
    .A(_4339_),
    .B(_4363_));
 sg13g2_nor2_1 _6162_ (.A(_4349_),
    .B(_0752_),
    .Y(_0774_));
 sg13g2_a21oi_1 _6163_ (.A1(_4349_),
    .A2(_0773_),
    .Y(_0775_),
    .B1(_0774_));
 sg13g2_mux2_1 _6164_ (.A0(_0750_),
    .A1(_0775_),
    .S(_0737_),
    .X(_0777_));
 sg13g2_a22oi_1 _6165_ (.Y(_0778_),
    .B1(_0777_),
    .B2(_0748_),
    .A2(_0772_),
    .A1(_0771_));
 sg13g2_buf_1 _6166_ (.A(_0778_),
    .X(_0779_));
 sg13g2_nor2_1 _6167_ (.A(net14),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_o21ai_1 _6168_ (.B1(_0780_),
    .Y(_0781_),
    .A1(_0768_),
    .A2(_0770_));
 sg13g2_inv_1 _6169_ (.Y(_0782_),
    .A(_0779_));
 sg13g2_nor2b_1 _6170_ (.A(net14),
    .B_N(_0757_),
    .Y(_0783_));
 sg13g2_buf_1 _6171_ (.A(_0783_),
    .X(_0784_));
 sg13g2_o21ai_1 _6172_ (.B1(_0727_),
    .Y(_0785_),
    .A1(_0782_),
    .A2(_0784_));
 sg13g2_nand3b_1 _6173_ (.B(_0781_),
    .C(_0785_),
    .Y(_0786_),
    .A_N(_0766_));
 sg13g2_xnor2_1 _6174_ (.Y(_0788_),
    .A(_4387_),
    .B(_0786_));
 sg13g2_xnor2_1 _6175_ (.Y(_0789_),
    .A(_0727_),
    .B(_0779_));
 sg13g2_nor2_1 _6176_ (.A(_0721_),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_a22oi_1 _6177_ (.Y(_0791_),
    .B1(_0790_),
    .B2(_0765_),
    .A2(_0789_),
    .A1(_0768_));
 sg13g2_nor2_1 _6178_ (.A(net14),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_nand3_1 _6179_ (.B(net14),
    .C(_0757_),
    .A(_0721_),
    .Y(_0793_));
 sg13g2_inv_1 _6180_ (.Y(_0794_),
    .A(_0793_));
 sg13g2_nor2_1 _6181_ (.A(_0782_),
    .B(_0784_),
    .Y(_0795_));
 sg13g2_xnor2_1 _6182_ (.Y(_0796_),
    .A(_0727_),
    .B(_0795_));
 sg13g2_a21oi_1 _6183_ (.A1(_0768_),
    .A2(_0794_),
    .Y(_0797_),
    .B1(_0796_));
 sg13g2_nand2_1 _6184_ (.Y(_0799_),
    .A(_0735_),
    .B(_0789_));
 sg13g2_a21oi_1 _6185_ (.A1(_0758_),
    .A2(_0799_),
    .Y(_0800_),
    .B1(_0723_));
 sg13g2_inv_1 _6186_ (.Y(_0801_),
    .A(_0757_));
 sg13g2_nand2_1 _6187_ (.Y(_0802_),
    .A(_0734_),
    .B(_0801_));
 sg13g2_nor2_1 _6188_ (.A(_0721_),
    .B(_0802_),
    .Y(_0803_));
 sg13g2_mux2_1 _6189_ (.A0(_0800_),
    .A1(_0803_),
    .S(_0765_),
    .X(_0804_));
 sg13g2_nor2_1 _6190_ (.A(_0715_),
    .B(_0758_),
    .Y(_0805_));
 sg13g2_or4_1 _6191_ (.A(_0792_),
    .B(_0797_),
    .C(_0804_),
    .D(_0805_),
    .X(_0806_));
 sg13g2_buf_1 _6192_ (.A(_0806_),
    .X(_0807_));
 sg13g2_buf_1 _6193_ (.A(net281),
    .X(_0808_));
 sg13g2_xnor2_1 _6194_ (.Y(_0810_),
    .A(net234),
    .B(_0941_));
 sg13g2_nor2_1 _6195_ (.A(net229),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_and4_1 _6196_ (.A(_4108_),
    .B(_0788_),
    .C(_0807_),
    .D(_0811_),
    .X(_0812_));
 sg13g2_and2_1 _6197_ (.A(_0723_),
    .B(_0784_),
    .X(_0813_));
 sg13g2_a22oi_1 _6198_ (.Y(_0814_),
    .B1(_0813_),
    .B2(_0715_),
    .A2(_0784_),
    .A1(_0765_));
 sg13g2_nor2_1 _6199_ (.A(net14),
    .B(_0757_),
    .Y(_0815_));
 sg13g2_and2_1 _6200_ (.A(_0721_),
    .B(_0815_),
    .X(_0816_));
 sg13g2_a21oi_1 _6201_ (.A1(_0760_),
    .A2(_0762_),
    .Y(_0817_),
    .B1(_0763_));
 sg13g2_a22oi_1 _6202_ (.Y(_0818_),
    .B1(_0816_),
    .B2(_0817_),
    .A2(_0815_),
    .A1(_0768_));
 sg13g2_nand3_1 _6203_ (.B(net14),
    .C(_0757_),
    .A(_0768_),
    .Y(_0819_));
 sg13g2_nand2_1 _6204_ (.Y(_0821_),
    .A(_0817_),
    .B(_0794_));
 sg13g2_nand4_1 _6205_ (.B(_0818_),
    .C(_0819_),
    .A(_0814_),
    .Y(_0822_),
    .D(_0821_));
 sg13g2_nor2_1 _6206_ (.A(_0789_),
    .B(_0802_),
    .Y(_0823_));
 sg13g2_nor2_2 _6207_ (.A(_0768_),
    .B(_0770_),
    .Y(_0824_));
 sg13g2_a22oi_1 _6208_ (.Y(_0825_),
    .B1(_0823_),
    .B2(_0824_),
    .A2(_0822_),
    .A1(_0789_));
 sg13g2_buf_1 _6209_ (.A(_0825_),
    .X(_0826_));
 sg13g2_nand2_1 _6210_ (.Y(_0827_),
    .A(_0812_),
    .B(_0826_));
 sg13g2_nor2_1 _6211_ (.A(net261),
    .B(net222),
    .Y(_0828_));
 sg13g2_nand2_2 _6212_ (.Y(_0829_),
    .A(net253),
    .B(net290));
 sg13g2_nor2_1 _6213_ (.A(_0828_),
    .B(_0829_),
    .Y(_0830_));
 sg13g2_buf_2 _6214_ (.A(_0830_),
    .X(_0832_));
 sg13g2_nor2_1 _6215_ (.A(net188),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_buf_2 _6216_ (.A(_0833_),
    .X(_0834_));
 sg13g2_nand4_1 _6217_ (.B(_0788_),
    .C(_0807_),
    .A(_4108_),
    .Y(_0835_),
    .D(_0811_));
 sg13g2_buf_1 _6218_ (.A(_0835_),
    .X(_0836_));
 sg13g2_or2_1 _6219_ (.X(_0837_),
    .B(net257),
    .A(_0073_));
 sg13g2_buf_2 _6220_ (.A(_0837_),
    .X(_0838_));
 sg13g2_nor2_1 _6221_ (.A(_0838_),
    .B(_0829_),
    .Y(_0839_));
 sg13g2_nor2_2 _6222_ (.A(net288),
    .B(net250),
    .Y(_0840_));
 sg13g2_nand2_1 _6223_ (.Y(_0841_),
    .A(net271),
    .B(_0840_));
 sg13g2_nor3_2 _6224_ (.A(_0700_),
    .B(_4042_),
    .C(_4053_),
    .Y(_0843_));
 sg13g2_nor2_1 _6225_ (.A(net184),
    .B(_0843_),
    .Y(_0844_));
 sg13g2_nor2_2 _6226_ (.A(_0502_),
    .B(_4089_),
    .Y(_0845_));
 sg13g2_nor2b_1 _6227_ (.A(net292),
    .B_N(_4066_),
    .Y(_0846_));
 sg13g2_and2_1 _6228_ (.A(net222),
    .B(_0846_),
    .X(_0847_));
 sg13g2_nand2_1 _6229_ (.Y(_0848_),
    .A(_0557_),
    .B(net252));
 sg13g2_buf_1 _6230_ (.A(_0848_),
    .X(_0849_));
 sg13g2_a21oi_1 _6231_ (.A1(_0845_),
    .A2(_0847_),
    .Y(_0850_),
    .B1(net175));
 sg13g2_nor2b_1 _6232_ (.A(_0844_),
    .B_N(_0850_),
    .Y(_0851_));
 sg13g2_buf_1 _6233_ (.A(_0851_),
    .X(_0852_));
 sg13g2_buf_1 _6234_ (.A(_0852_),
    .X(_0854_));
 sg13g2_a21oi_1 _6235_ (.A1(_0839_),
    .A2(_0841_),
    .Y(_0855_),
    .B1(net121));
 sg13g2_and2_1 _6236_ (.A(_0836_),
    .B(_0855_),
    .X(_0856_));
 sg13g2_buf_1 _6237_ (.A(net203),
    .X(_0857_));
 sg13g2_buf_1 _6238_ (.A(net174),
    .X(_0858_));
 sg13g2_buf_1 _6239_ (.A(_0858_),
    .X(_0859_));
 sg13g2_xnor2_1 _6240_ (.Y(_0860_),
    .A(net170),
    .B(net156));
 sg13g2_buf_1 _6241_ (.A(_0860_),
    .X(_0861_));
 sg13g2_buf_1 _6242_ (.A(net120),
    .X(_0862_));
 sg13g2_buf_1 _6243_ (.A(net97),
    .X(_0863_));
 sg13g2_buf_1 _6244_ (.A(net61),
    .X(_0865_));
 sg13g2_nand2_1 _6245_ (.Y(_0866_),
    .A(_1914_),
    .B(net219));
 sg13g2_nor2_1 _6246_ (.A(_4091_),
    .B(_0866_),
    .Y(_0867_));
 sg13g2_buf_2 _6247_ (.A(_0006_),
    .X(_0868_));
 sg13g2_o21ai_1 _6248_ (.B1(net252),
    .Y(_0869_),
    .A1(net253),
    .A2(_0868_));
 sg13g2_nand2_2 _6249_ (.Y(_0870_),
    .A(net288),
    .B(net250));
 sg13g2_nand2_1 _6250_ (.Y(_0871_),
    .A(_0447_),
    .B(_1479_));
 sg13g2_o21ai_1 _6251_ (.B1(_4229_),
    .Y(_0872_),
    .A1(net260),
    .A2(_0871_));
 sg13g2_buf_1 _6252_ (.A(_0872_),
    .X(_0873_));
 sg13g2_nor3_2 _6253_ (.A(_0084_),
    .B(net290),
    .C(_0134_),
    .Y(_0874_));
 sg13g2_o21ai_1 _6254_ (.B1(_0874_),
    .Y(_0876_),
    .A1(_0870_),
    .A2(_0873_));
 sg13g2_a22oi_1 _6255_ (.Y(_0877_),
    .B1(_0869_),
    .B2(_0876_),
    .A2(_0867_),
    .A1(_1523_));
 sg13g2_nand2_1 _6256_ (.Y(_0878_),
    .A(net39),
    .B(_0877_));
 sg13g2_nand3_1 _6257_ (.B(_0856_),
    .C(_0878_),
    .A(_0834_),
    .Y(_0879_));
 sg13g2_buf_1 _6258_ (.A(ui_in[0]),
    .X(_0880_));
 sg13g2_buf_1 _6259_ (.A(_0880_),
    .X(_0881_));
 sg13g2_nand2b_1 _6260_ (.Y(_0882_),
    .B(_0881_),
    .A_N(net1));
 sg13g2_buf_1 _6261_ (.A(_0880_),
    .X(_0883_));
 sg13g2_nor2_1 _6262_ (.A(net300),
    .B(_2261_),
    .Y(_0884_));
 sg13g2_nand2_1 _6263_ (.Y(_0885_),
    .A(_2840_),
    .B(_0884_));
 sg13g2_o21ai_1 _6264_ (.B1(_0885_),
    .Y(_0887_),
    .A1(net2),
    .A2(_0882_));
 sg13g2_buf_2 _6265_ (.A(_0887_),
    .X(_0888_));
 sg13g2_nand3b_1 _6266_ (.B(net301),
    .C(_2415_),
    .Y(_0889_),
    .A_N(_2480_));
 sg13g2_o21ai_1 _6267_ (.B1(_0889_),
    .Y(_0890_),
    .A1(net301),
    .A2(_2546_));
 sg13g2_buf_2 _6268_ (.A(_0890_),
    .X(_0891_));
 sg13g2_nand2_1 _6269_ (.Y(_0892_),
    .A(_0888_),
    .B(_0891_));
 sg13g2_buf_1 _6270_ (.A(_0892_),
    .X(_0893_));
 sg13g2_mux2_1 _6271_ (.A0(_2294_),
    .A1(net3),
    .S(net300),
    .X(_0894_));
 sg13g2_buf_1 _6272_ (.A(_0894_),
    .X(_0895_));
 sg13g2_buf_1 _6273_ (.A(_0895_),
    .X(_0896_));
 sg13g2_inv_1 _6274_ (.Y(_0898_),
    .A(net5));
 sg13g2_nand2b_1 _6275_ (.Y(_0899_),
    .B(_0883_),
    .A_N(net4));
 sg13g2_nor2_1 _6276_ (.A(net300),
    .B(_2228_),
    .Y(_0900_));
 sg13g2_nand2_1 _6277_ (.Y(_0901_),
    .A(_2316_),
    .B(_0900_));
 sg13g2_o21ai_1 _6278_ (.B1(_0901_),
    .Y(_0902_),
    .A1(_0898_),
    .A2(_0899_));
 sg13g2_nand2_1 _6279_ (.Y(_0903_),
    .A(net155),
    .B(_0902_));
 sg13g2_or2_1 _6280_ (.X(_0904_),
    .B(_0903_),
    .A(_0893_));
 sg13g2_buf_1 _6281_ (.A(_0904_),
    .X(_0905_));
 sg13g2_a21o_1 _6282_ (.A2(_0879_),
    .A1(_0827_),
    .B1(_0905_),
    .X(_0906_));
 sg13g2_nand2_1 _6283_ (.Y(_0907_),
    .A(net202),
    .B(_3644_));
 sg13g2_o21ai_1 _6284_ (.B1(_0394_),
    .Y(_0909_),
    .A1(_3655_),
    .A2(_0907_));
 sg13g2_nor3_1 _6285_ (.A(net310),
    .B(net311),
    .C(net312),
    .Y(_0910_));
 sg13g2_buf_1 _6286_ (.A(_0910_),
    .X(_0911_));
 sg13g2_buf_1 _6287_ (.A(net228),
    .X(_0912_));
 sg13g2_and3_1 _6288_ (.X(_0913_),
    .A(net241),
    .B(net279),
    .C(net237));
 sg13g2_and2_1 _6289_ (.A(net282),
    .B(net284),
    .X(_0914_));
 sg13g2_o21ai_1 _6290_ (.B1(_0914_),
    .Y(_0915_),
    .A1(net309),
    .A2(_0913_));
 sg13g2_nand2_1 _6291_ (.Y(_0916_),
    .A(net196),
    .B(_0915_));
 sg13g2_buf_2 _6292_ (.A(_0916_),
    .X(_0917_));
 sg13g2_mux2_1 _6293_ (.A0(_3699_),
    .A1(_0909_),
    .S(_0917_),
    .X(_0918_));
 sg13g2_xnor2_1 _6294_ (.Y(_0920_),
    .A(net280),
    .B(_0918_));
 sg13g2_buf_2 _6295_ (.A(_0920_),
    .X(_0921_));
 sg13g2_buf_1 _6296_ (.A(net266),
    .X(_0922_));
 sg13g2_a221oi_1 _6297_ (.B2(net227),
    .C1(net283),
    .B1(net196),
    .A1(net202),
    .Y(_0923_),
    .A2(_1314_));
 sg13g2_xnor2_1 _6298_ (.Y(_0924_),
    .A(_0394_),
    .B(_3688_));
 sg13g2_nand2_1 _6299_ (.Y(_0925_),
    .A(net283),
    .B(_0913_));
 sg13g2_nand2_1 _6300_ (.Y(_0926_),
    .A(_3827_),
    .B(_0911_));
 sg13g2_mux2_1 _6301_ (.A0(_0924_),
    .A1(_0925_),
    .S(_0926_),
    .X(_0927_));
 sg13g2_nor2b_1 _6302_ (.A(_0923_),
    .B_N(_0927_),
    .Y(_0928_));
 sg13g2_buf_2 _6303_ (.A(_0928_),
    .X(_0929_));
 sg13g2_and2_1 _6304_ (.A(net196),
    .B(_0915_),
    .X(_0931_));
 sg13g2_buf_1 _6305_ (.A(_0931_),
    .X(_0932_));
 sg13g2_and3_1 _6306_ (.X(_0933_),
    .A(net241),
    .B(net276),
    .C(net278));
 sg13g2_buf_1 _6307_ (.A(_0933_),
    .X(_0934_));
 sg13g2_xnor2_1 _6308_ (.Y(_0935_),
    .A(net214),
    .B(_0934_));
 sg13g2_and2_1 _6309_ (.A(net277),
    .B(net278),
    .X(_0936_));
 sg13g2_buf_1 _6310_ (.A(_0936_),
    .X(_0937_));
 sg13g2_xnor2_1 _6311_ (.Y(_0938_),
    .A(net230),
    .B(_0937_));
 sg13g2_nor2_1 _6312_ (.A(net154),
    .B(_0938_),
    .Y(_0939_));
 sg13g2_a21o_1 _6313_ (.A2(_0935_),
    .A1(net154),
    .B1(_0939_),
    .X(_0940_));
 sg13g2_buf_1 _6314_ (.A(_0940_),
    .X(_0942_));
 sg13g2_buf_1 _6315_ (.A(_0942_),
    .X(_0943_));
 sg13g2_xnor2_1 _6316_ (.Y(_0944_),
    .A(net282),
    .B(_0918_));
 sg13g2_nor2_1 _6317_ (.A(net273),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_or2_1 _6318_ (.X(_0946_),
    .B(_0924_),
    .A(_0917_));
 sg13g2_nor2_1 _6319_ (.A(net283),
    .B(net154),
    .Y(_0947_));
 sg13g2_nor3_1 _6320_ (.A(net203),
    .B(net227),
    .C(_0917_),
    .Y(_0948_));
 sg13g2_o21ai_1 _6321_ (.B1(net178),
    .Y(_0949_),
    .A1(_0947_),
    .A2(_0948_));
 sg13g2_o21ai_1 _6322_ (.B1(_0949_),
    .Y(_0950_),
    .A1(_1402_),
    .A2(_0946_));
 sg13g2_nor2_1 _6323_ (.A(_0945_),
    .B(_0950_),
    .Y(_0951_));
 sg13g2_a21oi_2 _6324_ (.B1(_0939_),
    .Y(_0953_),
    .A2(_0935_),
    .A1(net154));
 sg13g2_and3_1 _6325_ (.X(_0954_),
    .A(net240),
    .B(net228),
    .C(_0915_));
 sg13g2_buf_1 _6326_ (.A(_0954_),
    .X(_0955_));
 sg13g2_mux2_1 _6327_ (.A0(_0917_),
    .A1(_0955_),
    .S(net202),
    .X(_0956_));
 sg13g2_xnor2_1 _6328_ (.Y(_0957_),
    .A(net213),
    .B(_0956_));
 sg13g2_buf_1 _6329_ (.A(_0957_),
    .X(_0958_));
 sg13g2_nand2_2 _6330_ (.Y(_0959_),
    .A(_0953_),
    .B(net96));
 sg13g2_a22oi_1 _6331_ (.Y(_0960_),
    .B1(_0945_),
    .B2(_0950_),
    .A2(_0958_),
    .A1(_0953_));
 sg13g2_or2_1 _6332_ (.X(_0961_),
    .B(_0960_),
    .A(_0951_));
 sg13g2_or2_1 _6333_ (.X(_0962_),
    .B(net236),
    .A(net203));
 sg13g2_buf_1 _6334_ (.A(_0962_),
    .X(_0964_));
 sg13g2_nor3_1 _6335_ (.A(net181),
    .B(_0917_),
    .C(_0964_),
    .Y(_0965_));
 sg13g2_nor3_1 _6336_ (.A(net213),
    .B(net230),
    .C(_0932_),
    .Y(_0966_));
 sg13g2_o21ai_1 _6337_ (.B1(net178),
    .Y(_0967_),
    .A1(_0965_),
    .A2(_0966_));
 sg13g2_o21ai_1 _6338_ (.B1(_0967_),
    .Y(_0968_),
    .A1(_3688_),
    .A2(_0917_));
 sg13g2_buf_1 _6339_ (.A(_0968_),
    .X(_0969_));
 sg13g2_nand2b_1 _6340_ (.Y(_0970_),
    .B(_0927_),
    .A_N(_0923_));
 sg13g2_buf_1 _6341_ (.A(_0970_),
    .X(_0971_));
 sg13g2_xnor2_1 _6342_ (.Y(_0972_),
    .A(net199),
    .B(_0955_));
 sg13g2_nand2_1 _6343_ (.Y(_0973_),
    .A(net96),
    .B(_0972_));
 sg13g2_o21ai_1 _6344_ (.B1(_0942_),
    .Y(_0975_),
    .A1(net96),
    .A2(_0972_));
 sg13g2_nand4_1 _6345_ (.B(_0971_),
    .C(_0973_),
    .A(net174),
    .Y(_0976_),
    .D(_0975_));
 sg13g2_nor2b_1 _6346_ (.A(_0969_),
    .B_N(_0976_),
    .Y(_0977_));
 sg13g2_a22oi_1 _6347_ (.Y(_0978_),
    .B1(_0961_),
    .B2(_0977_),
    .A2(_0959_),
    .A1(_0951_));
 sg13g2_buf_2 _6348_ (.A(_0978_),
    .X(_0979_));
 sg13g2_xnor2_1 _6349_ (.Y(_0980_),
    .A(net181),
    .B(_0956_));
 sg13g2_buf_2 _6350_ (.A(_0980_),
    .X(_0981_));
 sg13g2_a21oi_1 _6351_ (.A1(net60),
    .A2(_0979_),
    .Y(_0982_),
    .B1(_0981_));
 sg13g2_nor2_1 _6352_ (.A(net95),
    .B(net60),
    .Y(_0983_));
 sg13g2_o21ai_1 _6353_ (.B1(_0983_),
    .Y(_0984_),
    .A1(net96),
    .A2(_0972_));
 sg13g2_o21ai_1 _6354_ (.B1(_0984_),
    .Y(_0986_),
    .A1(_0929_),
    .A2(_0982_));
 sg13g2_a22oi_1 _6355_ (.Y(_0987_),
    .B1(_0981_),
    .B2(_0979_),
    .A2(_0953_),
    .A1(_0944_));
 sg13g2_nor2_1 _6356_ (.A(_0929_),
    .B(_0987_),
    .Y(_0988_));
 sg13g2_a21oi_1 _6357_ (.A1(_0921_),
    .A2(_0986_),
    .Y(_0989_),
    .B1(_0988_));
 sg13g2_nor4_2 _6358_ (.A(_1914_),
    .B(_0557_),
    .C(net257),
    .Y(_0990_),
    .D(_0392_));
 sg13g2_a21oi_2 _6359_ (.B1(net290),
    .Y(_0991_),
    .A2(_0838_),
    .A1(net292));
 sg13g2_a21o_1 _6360_ (.A2(_0990_),
    .A1(_0843_),
    .B1(_0991_),
    .X(_0992_));
 sg13g2_buf_2 _6361_ (.A(_0992_),
    .X(_0993_));
 sg13g2_nor2b_1 _6362_ (.A(net257),
    .B_N(net314),
    .Y(_0994_));
 sg13g2_and2_1 _6363_ (.A(_4066_),
    .B(_0994_),
    .X(_0995_));
 sg13g2_nand2_2 _6364_ (.Y(_0997_),
    .A(_0845_),
    .B(_0995_));
 sg13g2_nand2_1 _6365_ (.Y(_0998_),
    .A(_0260_),
    .B(net211));
 sg13g2_nor2_1 _6366_ (.A(_4091_),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_nor4_2 _6367_ (.A(net296),
    .B(net250),
    .C(net290),
    .Y(_1000_),
    .D(_0134_));
 sg13g2_inv_2 _6368_ (.Y(_1001_),
    .A(_0868_));
 sg13g2_a21oi_2 _6369_ (.B1(net290),
    .Y(_1002_),
    .A2(_1001_),
    .A1(net292));
 sg13g2_a21oi_1 _6370_ (.A1(_4198_),
    .A2(_1000_),
    .Y(_1003_),
    .B1(_1002_));
 sg13g2_a221oi_1 _6371_ (.B2(_4168_),
    .C1(_1003_),
    .B1(_0999_),
    .A1(_0993_),
    .Y(_1004_),
    .A2(_0997_));
 sg13g2_buf_1 _6372_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nand2_1 _6373_ (.Y(_1006_),
    .A(_0348_),
    .B(_0846_));
 sg13g2_nor3_1 _6374_ (.A(_4157_),
    .B(_1006_),
    .C(_0998_),
    .Y(_1008_));
 sg13g2_nor2_1 _6375_ (.A(net184),
    .B(_0870_),
    .Y(_1009_));
 sg13g2_a21oi_1 _6376_ (.A1(_0175_),
    .A2(_1009_),
    .Y(_1010_),
    .B1(net175));
 sg13g2_nor2b_1 _6377_ (.A(_1008_),
    .B_N(_1010_),
    .Y(_1011_));
 sg13g2_buf_2 _6378_ (.A(_1011_),
    .X(_1012_));
 sg13g2_or3_1 _6379_ (.A(net271),
    .B(_1005_),
    .C(_1012_),
    .X(_1013_));
 sg13g2_buf_1 _6380_ (.A(_1013_),
    .X(_1014_));
 sg13g2_buf_1 _6381_ (.A(_1014_),
    .X(_1015_));
 sg13g2_buf_1 _6382_ (.A(_1005_),
    .X(_1016_));
 sg13g2_o21ai_1 _6383_ (.B1(net176),
    .Y(_1017_),
    .A1(net59),
    .A2(_1012_));
 sg13g2_buf_1 _6384_ (.A(_1017_),
    .X(_1019_));
 sg13g2_buf_8 _6385_ (.A(_1019_),
    .X(_1020_));
 sg13g2_or3_1 _6386_ (.A(net288),
    .B(net59),
    .C(_1012_),
    .X(_1021_));
 sg13g2_buf_1 _6387_ (.A(_1021_),
    .X(_1022_));
 sg13g2_xor2_1 _6388_ (.B(_0175_),
    .A(net297),
    .X(_1023_));
 sg13g2_o21ai_1 _6389_ (.B1(_1023_),
    .Y(_1024_),
    .A1(net59),
    .A2(_1012_));
 sg13g2_a22oi_1 _6390_ (.Y(_1025_),
    .B1(_1022_),
    .B2(_1024_),
    .A2(net22),
    .A1(net25));
 sg13g2_nand2b_1 _6391_ (.Y(_1026_),
    .B(_1010_),
    .A_N(_1008_));
 sg13g2_buf_1 _6392_ (.A(_1026_),
    .X(_1027_));
 sg13g2_nand3b_1 _6393_ (.B(_1027_),
    .C(net265),
    .Y(_1028_),
    .A_N(net59));
 sg13g2_buf_2 _6394_ (.A(_1028_),
    .X(_1030_));
 sg13g2_o21ai_1 _6395_ (.B1(_4394_),
    .Y(_1031_),
    .A1(net59),
    .A2(_1012_));
 sg13g2_buf_2 _6396_ (.A(_1031_),
    .X(_1032_));
 sg13g2_and2_1 _6397_ (.A(_1030_),
    .B(_1032_),
    .X(_1033_));
 sg13g2_buf_2 _6398_ (.A(_1033_),
    .X(_1034_));
 sg13g2_nand2_1 _6399_ (.Y(_1035_),
    .A(_1025_),
    .B(_1034_));
 sg13g2_a21oi_1 _6400_ (.A1(_0260_),
    .A2(net211),
    .Y(_1036_),
    .B1(net316));
 sg13g2_xnor2_1 _6401_ (.Y(_1037_),
    .A(_3976_),
    .B(_1036_));
 sg13g2_nand2_1 _6402_ (.Y(_1038_),
    .A(_1016_),
    .B(_1037_));
 sg13g2_a21oi_1 _6403_ (.A1(_1457_),
    .A2(_4082_),
    .Y(_1039_),
    .B1(_4075_));
 sg13g2_o21ai_1 _6404_ (.B1(net288),
    .Y(_1041_),
    .A1(net175),
    .A2(_1039_));
 sg13g2_or2_1 _6405_ (.X(_1042_),
    .B(_1036_),
    .A(net175));
 sg13g2_and4_1 _6406_ (.A(_0993_),
    .B(_0997_),
    .C(_1041_),
    .D(_1042_),
    .X(_1043_));
 sg13g2_a21o_1 _6407_ (.A2(_1000_),
    .A1(_4198_),
    .B1(_1002_),
    .X(_1044_));
 sg13g2_buf_1 _6408_ (.A(_1044_),
    .X(_1045_));
 sg13g2_nand4_1 _6409_ (.B(_1512_),
    .C(_4168_),
    .A(_0260_),
    .Y(_1046_),
    .D(_4068_));
 sg13g2_buf_1 _6410_ (.A(_1046_),
    .X(_1047_));
 sg13g2_a221oi_1 _6411_ (.B2(_1047_),
    .C1(_0436_),
    .B1(_1045_),
    .A1(_0993_),
    .Y(_1048_),
    .A2(_0997_));
 sg13g2_o21ai_1 _6412_ (.B1(net233),
    .Y(_1049_),
    .A1(_1043_),
    .A2(_1048_));
 sg13g2_a21oi_1 _6413_ (.A1(_0843_),
    .A2(_0990_),
    .Y(_1050_),
    .B1(_0991_));
 sg13g2_a221oi_1 _6414_ (.B2(_1042_),
    .C1(_1050_),
    .B1(_1041_),
    .A1(_0845_),
    .Y(_1052_),
    .A2(_0995_));
 sg13g2_a221oi_1 _6415_ (.B2(_1047_),
    .C1(_0656_),
    .B1(_1045_),
    .A1(_0993_),
    .Y(_1053_),
    .A2(_0997_));
 sg13g2_o21ai_1 _6416_ (.B1(_0700_),
    .Y(_1054_),
    .A1(_1052_),
    .A2(_1053_));
 sg13g2_nand4_1 _6417_ (.B(_1038_),
    .C(_1049_),
    .A(net190),
    .Y(_1055_),
    .D(_1054_));
 sg13g2_buf_1 _6418_ (.A(_1055_),
    .X(_1056_));
 sg13g2_nor2_1 _6419_ (.A(_1035_),
    .B(_1056_),
    .Y(_1057_));
 sg13g2_nand4_1 _6420_ (.B(net22),
    .C(_1022_),
    .A(net25),
    .Y(_1058_),
    .D(_1024_));
 sg13g2_a21oi_1 _6421_ (.A1(net190),
    .A2(_1058_),
    .Y(_1059_),
    .B1(_1025_));
 sg13g2_nand3_1 _6422_ (.B(_1049_),
    .C(_1054_),
    .A(_1038_),
    .Y(_1060_));
 sg13g2_buf_1 _6423_ (.A(_1060_),
    .X(_1061_));
 sg13g2_nand2_1 _6424_ (.Y(_1063_),
    .A(_1030_),
    .B(_1032_));
 sg13g2_buf_1 _6425_ (.A(_1063_),
    .X(_1064_));
 sg13g2_nor2_1 _6426_ (.A(net21),
    .B(net19),
    .Y(_1065_));
 sg13g2_nor2b_1 _6427_ (.A(_1059_),
    .B_N(_1065_),
    .Y(_1066_));
 sg13g2_nand3b_1 _6428_ (.B(_1027_),
    .C(net288),
    .Y(_1067_),
    .A_N(net59));
 sg13g2_buf_1 _6429_ (.A(_1067_),
    .X(_1068_));
 sg13g2_xnor2_1 _6430_ (.Y(_1069_),
    .A(net297),
    .B(_0175_));
 sg13g2_o21ai_1 _6431_ (.B1(_1069_),
    .Y(_1070_),
    .A1(_1016_),
    .A2(_1012_));
 sg13g2_buf_1 _6432_ (.A(_1070_),
    .X(_1071_));
 sg13g2_nand4_1 _6433_ (.B(net22),
    .C(_1068_),
    .A(net25),
    .Y(_1072_),
    .D(_1071_));
 sg13g2_buf_2 _6434_ (.A(_1072_),
    .X(_1074_));
 sg13g2_and2_1 _6435_ (.A(_0993_),
    .B(_0997_),
    .X(_1075_));
 sg13g2_buf_1 _6436_ (.A(_1075_),
    .X(_1076_));
 sg13g2_nand2_1 _6437_ (.Y(_1077_),
    .A(_0840_),
    .B(_1003_));
 sg13g2_nand2_1 _6438_ (.Y(_1078_),
    .A(net233),
    .B(_4198_));
 sg13g2_nand3_1 _6439_ (.B(_1047_),
    .C(_1078_),
    .A(_1045_),
    .Y(_1079_));
 sg13g2_buf_1 _6440_ (.A(_0003_),
    .X(_1080_));
 sg13g2_inv_1 _6441_ (.Y(_1081_),
    .A(net299));
 sg13g2_a21oi_1 _6442_ (.A1(_1077_),
    .A2(_1079_),
    .Y(_1082_),
    .B1(_1081_));
 sg13g2_and3_1 _6443_ (.X(_1083_),
    .A(_1081_),
    .B(_1077_),
    .C(_1079_));
 sg13g2_or3_1 _6444_ (.A(_1076_),
    .B(_1082_),
    .C(_1083_),
    .X(_1085_));
 sg13g2_buf_1 _6445_ (.A(_1085_),
    .X(_1086_));
 sg13g2_nor2_2 _6446_ (.A(net255),
    .B(net233),
    .Y(_1087_));
 sg13g2_nand3_1 _6447_ (.B(_1087_),
    .C(_0175_),
    .A(net184),
    .Y(_1088_));
 sg13g2_nand2_1 _6448_ (.Y(_1089_),
    .A(_0870_),
    .B(net175));
 sg13g2_o21ai_1 _6449_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net175),
    .A2(_1088_));
 sg13g2_xnor2_1 _6450_ (.Y(_1091_),
    .A(_1914_),
    .B(_1090_));
 sg13g2_nand2_1 _6451_ (.Y(_1092_),
    .A(_1076_),
    .B(_1091_));
 sg13g2_buf_2 _6452_ (.A(_1092_),
    .X(_1093_));
 sg13g2_nand3_1 _6453_ (.B(_1086_),
    .C(_1093_),
    .A(net232),
    .Y(_1094_));
 sg13g2_xnor2_1 _6454_ (.Y(_1096_),
    .A(_1074_),
    .B(_1094_));
 sg13g2_and2_1 _6455_ (.A(_1014_),
    .B(_1019_),
    .X(_1097_));
 sg13g2_buf_2 _6456_ (.A(_1097_),
    .X(_1098_));
 sg13g2_nand2_1 _6457_ (.Y(_1099_),
    .A(_1068_),
    .B(_1071_));
 sg13g2_buf_1 _6458_ (.A(_1099_),
    .X(_1100_));
 sg13g2_and3_1 _6459_ (.X(_1101_),
    .A(_1038_),
    .B(_1049_),
    .C(_1054_));
 sg13g2_buf_1 _6460_ (.A(_1101_),
    .X(_1102_));
 sg13g2_buf_1 _6461_ (.A(_1102_),
    .X(_1103_));
 sg13g2_mux2_1 _6462_ (.A0(net17),
    .A1(_1056_),
    .S(net19),
    .X(_1104_));
 sg13g2_nor4_1 _6463_ (.A(_1098_),
    .B(net18),
    .C(_1094_),
    .D(_1104_),
    .Y(_1105_));
 sg13g2_a221oi_1 _6464_ (.B2(_1096_),
    .C1(_1105_),
    .B1(_1066_),
    .A1(net232),
    .Y(_1107_),
    .A2(_1057_));
 sg13g2_buf_1 _6465_ (.A(_1107_),
    .X(_1108_));
 sg13g2_nand2_1 _6466_ (.Y(_1109_),
    .A(_1022_),
    .B(_1024_));
 sg13g2_buf_1 _6467_ (.A(_1109_),
    .X(_1110_));
 sg13g2_nand2_1 _6468_ (.Y(_1111_),
    .A(net17),
    .B(_1110_));
 sg13g2_and3_1 _6469_ (.X(_1112_),
    .A(_1086_),
    .B(_1093_),
    .C(_1034_));
 sg13g2_buf_1 _6470_ (.A(_1112_),
    .X(_1113_));
 sg13g2_nand4_1 _6471_ (.B(_1098_),
    .C(_1111_),
    .A(net212),
    .Y(_1114_),
    .D(_1113_));
 sg13g2_nor2_1 _6472_ (.A(net17),
    .B(_1110_),
    .Y(_1115_));
 sg13g2_a21oi_1 _6473_ (.A1(_1086_),
    .A2(_1093_),
    .Y(_1116_),
    .B1(net21));
 sg13g2_nor2_1 _6474_ (.A(net19),
    .B(_1074_),
    .Y(_1118_));
 sg13g2_a22oi_1 _6475_ (.Y(_1119_),
    .B1(_1116_),
    .B2(_1118_),
    .A2(_1115_),
    .A1(_1113_));
 sg13g2_nand2_2 _6476_ (.Y(_1120_),
    .A(net25),
    .B(net22));
 sg13g2_nor2_1 _6477_ (.A(net21),
    .B(_1099_),
    .Y(_1121_));
 sg13g2_nand4_1 _6478_ (.B(_1120_),
    .C(_1121_),
    .A(net239),
    .Y(_1122_),
    .D(_1113_));
 sg13g2_nand3_1 _6479_ (.B(_1093_),
    .C(_1034_),
    .A(_1086_),
    .Y(_1123_));
 sg13g2_buf_1 _6480_ (.A(_1123_),
    .X(_1124_));
 sg13g2_nand2_1 _6481_ (.Y(_1125_),
    .A(net21),
    .B(net18));
 sg13g2_nand4_1 _6482_ (.B(_1111_),
    .C(_1124_),
    .A(_1120_),
    .Y(_1126_),
    .D(_1125_));
 sg13g2_and4_1 _6483_ (.A(_1015_),
    .B(_1020_),
    .C(_1068_),
    .D(_1071_),
    .X(_1127_));
 sg13g2_nand4_1 _6484_ (.B(_1093_),
    .C(_1064_),
    .A(_1086_),
    .Y(_1129_),
    .D(_1127_));
 sg13g2_nand3_1 _6485_ (.B(_1120_),
    .C(_1100_),
    .A(_1103_),
    .Y(_1130_));
 sg13g2_a21o_1 _6486_ (.A2(_1130_),
    .A1(_1129_),
    .B1(net239),
    .X(_1131_));
 sg13g2_and3_1 _6487_ (.X(_1132_),
    .A(_1122_),
    .B(_1126_),
    .C(_1131_));
 sg13g2_nand3_1 _6488_ (.B(_1119_),
    .C(_1132_),
    .A(_1114_),
    .Y(_1133_));
 sg13g2_xnor2_1 _6489_ (.Y(_1134_),
    .A(_1108_),
    .B(_1133_));
 sg13g2_and3_1 _6490_ (.X(_1135_),
    .A(net239),
    .B(_1030_),
    .C(_1032_));
 sg13g2_a21o_1 _6491_ (.A2(net22),
    .A1(net25),
    .B1(net208),
    .X(_1136_));
 sg13g2_nor2_1 _6492_ (.A(_1135_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_nor4_1 _6493_ (.A(_1102_),
    .B(_1098_),
    .C(net18),
    .D(net19),
    .Y(_1138_));
 sg13g2_a221oi_1 _6494_ (.B2(_1137_),
    .C1(_1138_),
    .B1(_1121_),
    .A1(_1059_),
    .Y(_1139_),
    .A2(_1065_));
 sg13g2_xor2_1 _6495_ (.B(_1139_),
    .A(_1096_),
    .X(_1140_));
 sg13g2_xnor2_1 _6496_ (.Y(_1141_),
    .A(_0945_),
    .B(_0950_));
 sg13g2_xnor2_1 _6497_ (.Y(_1142_),
    .A(_0959_),
    .B(_1141_));
 sg13g2_nand2_1 _6498_ (.Y(_1143_),
    .A(net174),
    .B(_0970_));
 sg13g2_nand2b_1 _6499_ (.Y(_1144_),
    .B(_3449_),
    .A_N(_3503_));
 sg13g2_buf_1 _6500_ (.A(net202),
    .X(_1145_));
 sg13g2_a221oi_1 _6501_ (.B2(net173),
    .C1(_0395_),
    .B1(_1144_),
    .A1(net181),
    .Y(_1146_),
    .A2(_4110_));
 sg13g2_nor2_2 _6502_ (.A(net214),
    .B(net181),
    .Y(_1147_));
 sg13g2_nand2_1 _6503_ (.Y(_1148_),
    .A(_4110_),
    .B(_1147_));
 sg13g2_o21ai_1 _6504_ (.B1(_1148_),
    .Y(_1150_),
    .A1(net236),
    .A2(_1146_));
 sg13g2_nor2b_1 _6505_ (.A(_3514_),
    .B_N(net204),
    .Y(_1151_));
 sg13g2_a21oi_1 _6506_ (.A1(net230),
    .A2(_1151_),
    .Y(_1152_),
    .B1(_4521_));
 sg13g2_nor2_1 _6507_ (.A(net154),
    .B(_1152_),
    .Y(_1153_));
 sg13g2_a21oi_1 _6508_ (.A1(_0932_),
    .A2(_1150_),
    .Y(_1154_),
    .B1(_1153_));
 sg13g2_o21ai_1 _6509_ (.B1(_0969_),
    .Y(_1155_),
    .A1(net235),
    .A2(_1143_));
 sg13g2_o21ai_1 _6510_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_1143_),
    .A2(_1154_));
 sg13g2_xnor2_1 _6511_ (.Y(_1157_),
    .A(_1142_),
    .B(_1156_));
 sg13g2_a21oi_2 _6512_ (.B1(net239),
    .Y(_1158_),
    .A2(net22),
    .A1(net25));
 sg13g2_mux2_1 _6513_ (.A0(_1098_),
    .A1(_1158_),
    .S(net19),
    .X(_1159_));
 sg13g2_nand2_1 _6514_ (.Y(_1161_),
    .A(net190),
    .B(net239));
 sg13g2_a21oi_1 _6515_ (.A1(net25),
    .A2(net22),
    .Y(_1162_),
    .B1(_1161_));
 sg13g2_mux2_1 _6516_ (.A0(_1098_),
    .A1(_1162_),
    .S(_1102_),
    .X(_1163_));
 sg13g2_nor3_1 _6517_ (.A(net17),
    .B(_1135_),
    .C(_1136_),
    .Y(_1164_));
 sg13g2_a221oi_1 _6518_ (.B2(_1034_),
    .C1(_1164_),
    .B1(_1163_),
    .A1(net185),
    .Y(_1165_),
    .A2(_1159_));
 sg13g2_nor2_1 _6519_ (.A(_1034_),
    .B(_1056_),
    .Y(_1166_));
 sg13g2_nand2b_1 _6520_ (.Y(_1167_),
    .B(_1027_),
    .A_N(net59));
 sg13g2_buf_1 _6521_ (.A(_1012_),
    .X(_1168_));
 sg13g2_nor3_1 _6522_ (.A(net269),
    .B(net59),
    .C(net94),
    .Y(_1169_));
 sg13g2_a221oi_1 _6523_ (.B2(net22),
    .C1(_1169_),
    .B1(net25),
    .A1(_4394_),
    .Y(_1170_),
    .A2(_1167_));
 sg13g2_xnor2_1 _6524_ (.Y(_1172_),
    .A(_1170_),
    .B(_1056_));
 sg13g2_a22oi_1 _6525_ (.Y(_1173_),
    .B1(_1172_),
    .B2(net18),
    .A2(_1166_),
    .A1(_1098_));
 sg13g2_o21ai_1 _6526_ (.B1(_1173_),
    .Y(_1174_),
    .A1(net18),
    .A2(_1165_));
 sg13g2_buf_1 _6527_ (.A(_1174_),
    .X(_1175_));
 sg13g2_o21ai_1 _6528_ (.B1(net273),
    .Y(_1176_),
    .A1(_0929_),
    .A2(net60));
 sg13g2_xnor2_1 _6529_ (.Y(_1177_),
    .A(net178),
    .B(net154));
 sg13g2_a21oi_1 _6530_ (.A1(net238),
    .A2(net95),
    .Y(_1178_),
    .B1(_1177_));
 sg13g2_or2_1 _6531_ (.X(_1179_),
    .B(_0935_),
    .A(_0917_));
 sg13g2_nand3b_1 _6532_ (.B(_1179_),
    .C(net173),
    .Y(_1180_),
    .A_N(_0939_));
 sg13g2_o21ai_1 _6533_ (.B1(_1180_),
    .Y(_1181_),
    .A1(net173),
    .A2(_1179_));
 sg13g2_buf_1 _6534_ (.A(_4555_),
    .X(_1183_));
 sg13g2_a221oi_1 _6535_ (.B2(_0929_),
    .C1(net195),
    .B1(_1181_),
    .A1(_1176_),
    .Y(_1184_),
    .A2(_1178_));
 sg13g2_nor3_1 _6536_ (.A(net178),
    .B(net273),
    .C(net60),
    .Y(_1185_));
 sg13g2_nor2_1 _6537_ (.A(net173),
    .B(_0953_),
    .Y(_1186_));
 sg13g2_nor3_1 _6538_ (.A(net174),
    .B(_1185_),
    .C(_1186_),
    .Y(_1187_));
 sg13g2_nor2_1 _6539_ (.A(net173),
    .B(net154),
    .Y(_1188_));
 sg13g2_nand3_1 _6540_ (.B(net60),
    .C(_1188_),
    .A(_0929_),
    .Y(_1189_));
 sg13g2_o21ai_1 _6541_ (.B1(_1189_),
    .Y(_1190_),
    .A1(_1184_),
    .A2(_1187_));
 sg13g2_o21ai_1 _6542_ (.B1(_1143_),
    .Y(_1191_),
    .A1(_0972_),
    .A2(_0959_));
 sg13g2_a22oi_1 _6543_ (.Y(_1192_),
    .B1(_1191_),
    .B2(_0976_),
    .A2(_1190_),
    .A1(_0981_));
 sg13g2_buf_1 _6544_ (.A(_1192_),
    .X(_1194_));
 sg13g2_inv_1 _6545_ (.Y(_1195_),
    .A(_1194_));
 sg13g2_buf_1 _6546_ (.A(_4120_),
    .X(_1196_));
 sg13g2_nand2_1 _6547_ (.Y(_1197_),
    .A(net174),
    .B(net273));
 sg13g2_o21ai_1 _6548_ (.B1(_1197_),
    .Y(_1198_),
    .A1(net273),
    .A2(_1144_));
 sg13g2_nand2_1 _6549_ (.Y(_1199_),
    .A(net174),
    .B(net154));
 sg13g2_nand2_1 _6550_ (.Y(_1200_),
    .A(net213),
    .B(net238));
 sg13g2_o21ai_1 _6551_ (.B1(_1200_),
    .Y(_1201_),
    .A1(_3364_),
    .A2(_1199_));
 sg13g2_a21oi_1 _6552_ (.A1(net195),
    .A2(_0917_),
    .Y(_1202_),
    .B1(_1200_));
 sg13g2_a221oi_1 _6553_ (.B2(_1145_),
    .C1(_1202_),
    .B1(_1201_),
    .A1(_1188_),
    .Y(_1203_),
    .A2(_1198_));
 sg13g2_o21ai_1 _6554_ (.B1(_1203_),
    .Y(_1205_),
    .A1(net194),
    .A2(_1064_));
 sg13g2_nor3_1 _6555_ (.A(net194),
    .B(net19),
    .C(_1203_),
    .Y(_1206_));
 sg13g2_a21o_1 _6556_ (.A2(_1205_),
    .A1(_1158_),
    .B1(_1206_),
    .X(_1207_));
 sg13g2_nand2_1 _6557_ (.Y(_1208_),
    .A(net19),
    .B(_1158_));
 sg13g2_nand3b_1 _6558_ (.B(_1034_),
    .C(net190),
    .Y(_1209_),
    .A_N(_1158_));
 sg13g2_a21oi_1 _6559_ (.A1(_1208_),
    .A2(_1209_),
    .Y(_1210_),
    .B1(_1203_));
 sg13g2_a21oi_1 _6560_ (.A1(net185),
    .A2(_1207_),
    .Y(_1211_),
    .B1(_1210_));
 sg13g2_a22oi_1 _6561_ (.Y(_1212_),
    .B1(_1030_),
    .B2(_1032_),
    .A2(_1020_),
    .A1(_1015_));
 sg13g2_and4_1 _6562_ (.A(_1068_),
    .B(_1071_),
    .C(_1030_),
    .D(_1032_),
    .X(_1213_));
 sg13g2_mux2_1 _6563_ (.A0(_1212_),
    .A1(_1213_),
    .S(net232),
    .X(_1214_));
 sg13g2_o21ai_1 _6564_ (.B1(_1074_),
    .Y(_1216_),
    .A1(_1110_),
    .A2(_1136_));
 sg13g2_and2_1 _6565_ (.A(_1099_),
    .B(_1212_),
    .X(_1217_));
 sg13g2_a221oi_1 _6566_ (.B2(net232),
    .C1(_1217_),
    .B1(_1216_),
    .A1(net185),
    .Y(_1218_),
    .A2(_1214_));
 sg13g2_xnor2_1 _6567_ (.Y(_1219_),
    .A(net173),
    .B(_0955_));
 sg13g2_nor2_1 _6568_ (.A(net96),
    .B(_1219_),
    .Y(_1220_));
 sg13g2_nor3_1 _6569_ (.A(net273),
    .B(_0942_),
    .C(_0972_),
    .Y(_1221_));
 sg13g2_a21o_1 _6570_ (.A2(_1220_),
    .A1(net273),
    .B1(_1221_),
    .X(_1222_));
 sg13g2_nand3_1 _6571_ (.B(_0943_),
    .C(_0981_),
    .A(net174),
    .Y(_1223_));
 sg13g2_a21oi_1 _6572_ (.A1(_0959_),
    .A2(_1223_),
    .Y(_1224_),
    .B1(net235));
 sg13g2_a221oi_1 _6573_ (.B2(net195),
    .C1(_1224_),
    .B1(_1222_),
    .A1(net60),
    .Y(_1225_),
    .A2(_1220_));
 sg13g2_or2_1 _6574_ (.X(_1227_),
    .B(_1225_),
    .A(_1218_));
 sg13g2_and2_1 _6575_ (.A(_1218_),
    .B(_1225_),
    .X(_1228_));
 sg13g2_a21oi_1 _6576_ (.A1(_1211_),
    .A2(_1227_),
    .Y(_1229_),
    .B1(_1228_));
 sg13g2_buf_2 _6577_ (.A(_1229_),
    .X(_1230_));
 sg13g2_a221oi_1 _6578_ (.B2(_1195_),
    .C1(_1230_),
    .B1(net15),
    .A1(_1140_),
    .Y(_1231_),
    .A2(_1157_));
 sg13g2_a21o_1 _6579_ (.A2(_1157_),
    .A1(_1140_),
    .B1(net15),
    .X(_1232_));
 sg13g2_xnor2_1 _6580_ (.Y(_1233_),
    .A(_1096_),
    .B(_1139_));
 sg13g2_xor2_1 _6581_ (.B(_1156_),
    .A(_1142_),
    .X(_1234_));
 sg13g2_nand2_1 _6582_ (.Y(_1235_),
    .A(_1233_),
    .B(_1234_));
 sg13g2_o21ai_1 _6583_ (.B1(_1235_),
    .Y(_1236_),
    .A1(_1195_),
    .A2(_1232_));
 sg13g2_nand4_1 _6584_ (.B(net238),
    .C(net95),
    .A(net163),
    .Y(_1238_),
    .D(_0969_));
 sg13g2_o21ai_1 _6585_ (.B1(_1238_),
    .Y(_1239_),
    .A1(_0977_),
    .A2(_1142_));
 sg13g2_nand2_1 _6586_ (.Y(_1240_),
    .A(_0921_),
    .B(_1219_));
 sg13g2_inv_1 _6587_ (.Y(_1241_),
    .A(_0983_));
 sg13g2_nand2_1 _6588_ (.Y(_1242_),
    .A(net95),
    .B(_0943_));
 sg13g2_a21oi_1 _6589_ (.A1(_1241_),
    .A2(_1242_),
    .Y(_1243_),
    .B1(net96));
 sg13g2_xnor2_1 _6590_ (.Y(_1244_),
    .A(_1240_),
    .B(_1243_));
 sg13g2_xnor2_1 _6591_ (.Y(_1245_),
    .A(_0961_),
    .B(_1244_));
 sg13g2_xnor2_1 _6592_ (.Y(_1246_),
    .A(_1239_),
    .B(_1245_));
 sg13g2_nor3_1 _6593_ (.A(_1231_),
    .B(_1236_),
    .C(_1246_),
    .Y(_1247_));
 sg13g2_o21ai_1 _6594_ (.B1(_1246_),
    .Y(_1249_),
    .A1(_1231_),
    .A2(_1236_));
 sg13g2_o21ai_1 _6595_ (.B1(_1249_),
    .Y(_1250_),
    .A1(_1134_),
    .A2(_1247_));
 sg13g2_nor2_1 _6596_ (.A(net21),
    .B(_1074_),
    .Y(_1251_));
 sg13g2_o21ai_1 _6597_ (.B1(_1098_),
    .Y(_1252_),
    .A1(net17),
    .A2(_1110_));
 sg13g2_a21oi_1 _6598_ (.A1(_1111_),
    .A2(_1252_),
    .Y(_1253_),
    .B1(net212));
 sg13g2_o21ai_1 _6599_ (.B1(_1113_),
    .Y(_1254_),
    .A1(_1251_),
    .A2(_1253_));
 sg13g2_nand2_1 _6600_ (.Y(_1255_),
    .A(_1103_),
    .B(_1127_));
 sg13g2_a221oi_1 _6601_ (.B2(_1111_),
    .C1(_1124_),
    .B1(_1252_),
    .A1(net239),
    .Y(_1256_),
    .A2(_1255_));
 sg13g2_nor4_1 _6602_ (.A(net232),
    .B(_1120_),
    .C(_1121_),
    .D(_1124_),
    .Y(_1257_));
 sg13g2_nor2_1 _6603_ (.A(_1124_),
    .B(_1125_),
    .Y(_1258_));
 sg13g2_and2_1 _6604_ (.A(_1116_),
    .B(_1118_),
    .X(_1260_));
 sg13g2_nor4_1 _6605_ (.A(_1256_),
    .B(_1257_),
    .C(_1258_),
    .D(_1260_),
    .Y(_1261_));
 sg13g2_a221oi_1 _6606_ (.B2(_1261_),
    .C1(_1110_),
    .B1(_1132_),
    .A1(_1254_),
    .Y(_1262_),
    .A2(_1108_));
 sg13g2_nand2_1 _6607_ (.Y(_1263_),
    .A(net212),
    .B(_1061_));
 sg13g2_a21oi_1 _6608_ (.A1(_1113_),
    .A2(_1263_),
    .Y(_1264_),
    .B1(_1074_));
 sg13g2_and2_1 _6609_ (.A(_1086_),
    .B(_1093_),
    .X(_1265_));
 sg13g2_buf_1 _6610_ (.A(_1265_),
    .X(_1266_));
 sg13g2_a21oi_1 _6611_ (.A1(_1266_),
    .A2(_1058_),
    .Y(_1267_),
    .B1(net17));
 sg13g2_nor3_1 _6612_ (.A(_1262_),
    .B(_1264_),
    .C(_1267_),
    .Y(_1268_));
 sg13g2_nor2_1 _6613_ (.A(net18),
    .B(_1256_),
    .Y(_1269_));
 sg13g2_and4_1 _6614_ (.A(_1114_),
    .B(_1119_),
    .C(_1122_),
    .D(_1126_),
    .X(_1271_));
 sg13g2_a21oi_1 _6615_ (.A1(_1129_),
    .A2(_1130_),
    .Y(_1272_),
    .B1(net212));
 sg13g2_nor3_1 _6616_ (.A(_1100_),
    .B(_1256_),
    .C(_1272_),
    .Y(_1273_));
 sg13g2_a221oi_1 _6617_ (.B2(_1273_),
    .C1(_1217_),
    .B1(_1271_),
    .A1(_1108_),
    .Y(_1274_),
    .A2(_1269_));
 sg13g2_nand2_1 _6618_ (.Y(_1275_),
    .A(_1086_),
    .B(_1093_));
 sg13g2_a21oi_1 _6619_ (.A1(net21),
    .A2(net19),
    .Y(_1276_),
    .B1(_1275_));
 sg13g2_nand2b_1 _6620_ (.Y(_1277_),
    .B(_1276_),
    .A_N(_1274_));
 sg13g2_nand2_1 _6621_ (.Y(_1278_),
    .A(_1268_),
    .B(_1277_));
 sg13g2_a21o_1 _6622_ (.A2(_0979_),
    .A1(_0981_),
    .B1(_0929_),
    .X(_1279_));
 sg13g2_o21ai_1 _6623_ (.B1(_0959_),
    .Y(_1280_),
    .A1(net95),
    .A2(_0979_));
 sg13g2_a21o_1 _6624_ (.A2(_1279_),
    .A1(net60),
    .B1(_1280_),
    .X(_1282_));
 sg13g2_nand2_1 _6625_ (.Y(_1283_),
    .A(_1219_),
    .B(_0979_));
 sg13g2_nand3_1 _6626_ (.B(net95),
    .C(_0953_),
    .A(_0921_),
    .Y(_1284_));
 sg13g2_o21ai_1 _6627_ (.B1(_1284_),
    .Y(_1285_),
    .A1(net95),
    .A2(_0981_));
 sg13g2_nand4_1 _6628_ (.B(net60),
    .C(net96),
    .A(net95),
    .Y(_1286_),
    .D(_0979_));
 sg13g2_nand4_1 _6629_ (.B(_0981_),
    .C(_0983_),
    .A(_0921_),
    .Y(_1287_),
    .D(_0979_));
 sg13g2_nor4_1 _6630_ (.A(_0944_),
    .B(_0929_),
    .C(net96),
    .D(_1219_),
    .Y(_1288_));
 sg13g2_nand2b_1 _6631_ (.Y(_1289_),
    .B(_1288_),
    .A_N(_0979_));
 sg13g2_nand4_1 _6632_ (.B(_0981_),
    .C(_1219_),
    .A(_0921_),
    .Y(_1290_),
    .D(_0983_));
 sg13g2_nand4_1 _6633_ (.B(_1287_),
    .C(_1289_),
    .A(_1286_),
    .Y(_1291_),
    .D(_1290_));
 sg13g2_a221oi_1 _6634_ (.B2(_1285_),
    .C1(_1291_),
    .B1(_1283_),
    .A1(_0944_),
    .Y(_1293_),
    .A2(_1282_));
 sg13g2_buf_1 _6635_ (.A(_1293_),
    .X(_1294_));
 sg13g2_xnor2_1 _6636_ (.Y(_1295_),
    .A(_1278_),
    .B(_1294_));
 sg13g2_xnor2_1 _6637_ (.Y(_1296_),
    .A(_1250_),
    .B(_1295_));
 sg13g2_nand2_1 _6638_ (.Y(_1297_),
    .A(_1230_),
    .B(net15));
 sg13g2_o21ai_1 _6639_ (.B1(_1195_),
    .Y(_1298_),
    .A1(_1230_),
    .A2(net15));
 sg13g2_a21oi_1 _6640_ (.A1(_1297_),
    .A2(_1298_),
    .Y(_1299_),
    .B1(_1234_));
 sg13g2_o21ai_1 _6641_ (.B1(_1157_),
    .Y(_1300_),
    .A1(_1230_),
    .A2(net15));
 sg13g2_a21oi_1 _6642_ (.A1(_1230_),
    .A2(net15),
    .Y(_1301_),
    .B1(_1157_));
 sg13g2_a21o_1 _6643_ (.A2(_1300_),
    .A1(_1194_),
    .B1(_1301_),
    .X(_1302_));
 sg13g2_xor2_1 _6644_ (.B(_1246_),
    .A(_1134_),
    .X(_1304_));
 sg13g2_mux2_1 _6645_ (.A0(_1299_),
    .A1(_1302_),
    .S(_1304_),
    .X(_1305_));
 sg13g2_nand2_1 _6646_ (.Y(_1306_),
    .A(_1234_),
    .B(_1194_));
 sg13g2_nor3_1 _6647_ (.A(_1230_),
    .B(net15),
    .C(_1306_),
    .Y(_1307_));
 sg13g2_nor3_1 _6648_ (.A(_1157_),
    .B(_1230_),
    .C(net15),
    .Y(_1308_));
 sg13g2_a21oi_1 _6649_ (.A1(_1230_),
    .A2(_1175_),
    .Y(_1309_),
    .B1(_1306_));
 sg13g2_or2_1 _6650_ (.X(_1310_),
    .B(_1309_),
    .A(_1308_));
 sg13g2_nor3_1 _6651_ (.A(_1234_),
    .B(_1297_),
    .C(_1194_),
    .Y(_1311_));
 sg13g2_nor4_1 _6652_ (.A(_1233_),
    .B(_1304_),
    .C(_1310_),
    .D(_1311_),
    .Y(_1312_));
 sg13g2_a221oi_1 _6653_ (.B2(_1304_),
    .C1(_1312_),
    .B1(_1307_),
    .A1(_1233_),
    .Y(_1313_),
    .A2(_1305_));
 sg13g2_nand2_1 _6654_ (.Y(_1315_),
    .A(_1296_),
    .B(_1313_));
 sg13g2_nand2b_1 _6655_ (.Y(_1316_),
    .B(_1294_),
    .A_N(_1278_));
 sg13g2_a21oi_1 _6656_ (.A1(_1268_),
    .A2(_1277_),
    .Y(_1317_),
    .B1(_1294_));
 sg13g2_a21oi_2 _6657_ (.B1(_1317_),
    .Y(_1318_),
    .A2(_1250_),
    .A1(_1316_));
 sg13g2_a21oi_1 _6658_ (.A1(_1266_),
    .A2(_1120_),
    .Y(_1319_),
    .B1(_1262_));
 sg13g2_o21ai_1 _6659_ (.B1(_1319_),
    .Y(_1320_),
    .A1(_1266_),
    .A2(net18));
 sg13g2_nor4_1 _6660_ (.A(_1275_),
    .B(net17),
    .C(net18),
    .D(_1170_),
    .Y(_1321_));
 sg13g2_a21oi_1 _6661_ (.A1(net17),
    .A2(_1320_),
    .Y(_1322_),
    .B1(_1321_));
 sg13g2_inv_1 _6662_ (.Y(_1323_),
    .A(_1322_));
 sg13g2_nor2_1 _6663_ (.A(_1318_),
    .B(_1323_),
    .Y(_1324_));
 sg13g2_nand2_1 _6664_ (.Y(_1326_),
    .A(_1318_),
    .B(_1323_));
 sg13g2_o21ai_1 _6665_ (.B1(_1326_),
    .Y(_1327_),
    .A1(_1315_),
    .A2(_1324_));
 sg13g2_nand2b_1 _6666_ (.Y(_1328_),
    .B(_1327_),
    .A_N(_0989_));
 sg13g2_nor2_1 _6667_ (.A(_1326_),
    .B(_1315_),
    .Y(_1329_));
 sg13g2_nor2_1 _6668_ (.A(_0971_),
    .B(_0969_),
    .Y(_1330_));
 sg13g2_nor2_1 _6669_ (.A(_0944_),
    .B(_1330_),
    .Y(_1331_));
 sg13g2_nor2_1 _6670_ (.A(_1329_),
    .B(_1331_),
    .Y(_1332_));
 sg13g2_nand2_1 _6671_ (.Y(_1333_),
    .A(_0921_),
    .B(_1242_));
 sg13g2_a21oi_2 _6672_ (.B1(_1333_),
    .Y(_1334_),
    .A2(_0969_),
    .A1(_0929_));
 sg13g2_a21oi_1 _6673_ (.A1(net21),
    .A2(_1035_),
    .Y(_1335_),
    .B1(_1275_));
 sg13g2_and2_1 _6674_ (.A(_1335_),
    .B(_1331_),
    .X(_1337_));
 sg13g2_nand2_1 _6675_ (.Y(_1338_),
    .A(_0989_),
    .B(_1322_));
 sg13g2_nor4_1 _6676_ (.A(_1318_),
    .B(_1334_),
    .C(_1337_),
    .D(_1338_),
    .Y(_1339_));
 sg13g2_nand2_1 _6677_ (.Y(_1340_),
    .A(_1315_),
    .B(_1339_));
 sg13g2_buf_1 _6678_ (.A(_1076_),
    .X(_1341_));
 sg13g2_buf_1 _6679_ (.A(_1341_),
    .X(_1342_));
 sg13g2_nand2_1 _6680_ (.Y(_1343_),
    .A(net305),
    .B(net38));
 sg13g2_buf_1 _6681_ (.A(_1081_),
    .X(_1344_));
 sg13g2_nand3_1 _6682_ (.B(net226),
    .C(_1050_),
    .A(net189),
    .Y(_1345_));
 sg13g2_a21o_1 _6683_ (.A2(_1345_),
    .A1(_1343_),
    .B1(net253),
    .X(_1346_));
 sg13g2_o21ai_1 _6684_ (.B1(_1346_),
    .Y(_1348_),
    .A1(_0645_),
    .A2(_1343_));
 sg13g2_xnor2_1 _6685_ (.Y(_1349_),
    .A(_0590_),
    .B(_1348_));
 sg13g2_nand2_1 _6686_ (.Y(_1350_),
    .A(_0829_),
    .B(_1343_));
 sg13g2_xnor2_1 _6687_ (.Y(_1351_),
    .A(net184),
    .B(_1350_));
 sg13g2_buf_1 _6688_ (.A(_1351_),
    .X(_1352_));
 sg13g2_xnor2_1 _6689_ (.Y(_1353_),
    .A(net296),
    .B(net257));
 sg13g2_xnor2_1 _6690_ (.Y(_1354_),
    .A(_1342_),
    .B(_1353_));
 sg13g2_xnor2_1 _6691_ (.Y(_1355_),
    .A(net226),
    .B(_1341_));
 sg13g2_nor2_1 _6692_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sg13g2_buf_1 _6693_ (.A(net233),
    .X(_1357_));
 sg13g2_o21ai_1 _6694_ (.B1(net193),
    .Y(_1359_),
    .A1(net187),
    .A2(_0205_));
 sg13g2_nand3_1 _6695_ (.B(_4089_),
    .C(_0993_),
    .A(net186),
    .Y(_1360_));
 sg13g2_o21ai_1 _6696_ (.B1(_1360_),
    .Y(_1361_),
    .A1(net38),
    .A2(_1359_));
 sg13g2_nand3_1 _6697_ (.B(_1356_),
    .C(_1361_),
    .A(_1352_),
    .Y(_1362_));
 sg13g2_o21ai_1 _6698_ (.B1(net216),
    .Y(_1363_),
    .A1(net217),
    .A2(_4113_));
 sg13g2_nor2_1 _6699_ (.A(net286),
    .B(net281),
    .Y(_1364_));
 sg13g2_buf_1 _6700_ (.A(_1364_),
    .X(_1365_));
 sg13g2_a22oi_1 _6701_ (.Y(_1366_),
    .B1(_1363_),
    .B2(net192),
    .A2(_1362_),
    .A1(_1349_));
 sg13g2_inv_1 _6702_ (.Y(_1367_),
    .A(_1366_));
 sg13g2_nand3_1 _6703_ (.B(_1340_),
    .C(_1367_),
    .A(_0921_),
    .Y(_1368_));
 sg13g2_a21o_1 _6704_ (.A2(_1332_),
    .A1(_1328_),
    .B1(_1368_),
    .X(_1370_));
 sg13g2_nand3_1 _6705_ (.B(_1340_),
    .C(_1367_),
    .A(_1335_),
    .Y(_1371_));
 sg13g2_o21ai_1 _6706_ (.B1(_1266_),
    .Y(_1372_),
    .A1(net21),
    .A2(_1110_));
 sg13g2_nor3_1 _6707_ (.A(_1138_),
    .B(_1366_),
    .C(_1372_),
    .Y(_1373_));
 sg13g2_nor2_1 _6708_ (.A(_0989_),
    .B(_1322_),
    .Y(_1374_));
 sg13g2_o21ai_1 _6709_ (.B1(_1338_),
    .Y(_1375_),
    .A1(_1318_),
    .A2(_1374_));
 sg13g2_nand2b_1 _6710_ (.Y(_1376_),
    .B(_1375_),
    .A_N(_1334_));
 sg13g2_a21oi_1 _6711_ (.A1(_1334_),
    .A2(_1338_),
    .Y(_1377_),
    .B1(_1318_));
 sg13g2_nor2_1 _6712_ (.A(_1374_),
    .B(_1334_),
    .Y(_1378_));
 sg13g2_o21ai_1 _6713_ (.B1(_1315_),
    .Y(_1379_),
    .A1(_1377_),
    .A2(_1378_));
 sg13g2_nand3_1 _6714_ (.B(_1376_),
    .C(_1379_),
    .A(_1373_),
    .Y(_1381_));
 sg13g2_nand2_1 _6715_ (.Y(_1382_),
    .A(_0993_),
    .B(_0997_));
 sg13g2_buf_1 _6716_ (.A(_1382_),
    .X(_1383_));
 sg13g2_mux2_1 _6717_ (.A0(_4438_),
    .A1(net93),
    .S(_0183_),
    .X(_1384_));
 sg13g2_mux2_1 _6718_ (.A0(_4438_),
    .A1(net58),
    .S(net185),
    .X(_1385_));
 sg13g2_mux2_1 _6719_ (.A0(_1384_),
    .A1(_1385_),
    .S(net209),
    .X(_1386_));
 sg13g2_xnor2_1 _6720_ (.Y(_1387_),
    .A(net209),
    .B(net58));
 sg13g2_a22oi_1 _6721_ (.Y(_1388_),
    .B1(_1387_),
    .B2(_4438_),
    .A2(_1386_),
    .A1(net163));
 sg13g2_nor2_1 _6722_ (.A(net236),
    .B(net181),
    .Y(_1389_));
 sg13g2_buf_2 _6723_ (.A(_1389_),
    .X(_1390_));
 sg13g2_a22oi_1 _6724_ (.Y(_1392_),
    .B1(_1390_),
    .B2(net58),
    .A2(_1314_),
    .A1(_1686_));
 sg13g2_a221oi_1 _6725_ (.B2(net93),
    .C1(net251),
    .B1(_1390_),
    .A1(net254),
    .Y(_1393_),
    .A2(_1314_));
 sg13g2_a21oi_1 _6726_ (.A1(net251),
    .A2(_1392_),
    .Y(_1394_),
    .B1(_1393_));
 sg13g2_a21oi_1 _6727_ (.A1(_3471_),
    .A2(_1388_),
    .Y(_1395_),
    .B1(_1394_));
 sg13g2_xnor2_1 _6728_ (.Y(_1396_),
    .A(net254),
    .B(net58));
 sg13g2_o21ai_1 _6729_ (.B1(_1396_),
    .Y(_1397_),
    .A1(_3471_),
    .A2(_1388_));
 sg13g2_xnor2_1 _6730_ (.Y(_1398_),
    .A(net250),
    .B(net244));
 sg13g2_a21oi_1 _6731_ (.A1(net251),
    .A2(_3655_),
    .Y(_1399_),
    .B1(_1390_));
 sg13g2_nor2_1 _6732_ (.A(net93),
    .B(_1399_),
    .Y(_1400_));
 sg13g2_xnor2_1 _6733_ (.Y(_1401_),
    .A(net93),
    .B(_1398_));
 sg13g2_a21oi_1 _6734_ (.A1(net255),
    .A2(_3655_),
    .Y(_1403_),
    .B1(_1390_));
 sg13g2_nor3_1 _6735_ (.A(net58),
    .B(_1398_),
    .C(_1403_),
    .Y(_1404_));
 sg13g2_a221oi_1 _6736_ (.B2(_1314_),
    .C1(_1404_),
    .B1(_1401_),
    .A1(_1398_),
    .Y(_1405_),
    .A2(_1400_));
 sg13g2_a21oi_1 _6737_ (.A1(_1395_),
    .A2(_1397_),
    .Y(_1406_),
    .B1(_1405_));
 sg13g2_buf_1 _6738_ (.A(_3644_),
    .X(_1407_));
 sg13g2_nor2_1 _6739_ (.A(net191),
    .B(_3655_),
    .Y(_1408_));
 sg13g2_nor2_1 _6740_ (.A(net244),
    .B(_1314_),
    .Y(_1409_));
 sg13g2_xnor2_1 _6741_ (.Y(_1410_),
    .A(net250),
    .B(net58));
 sg13g2_o21ai_1 _6742_ (.B1(_1410_),
    .Y(_1411_),
    .A1(_1408_),
    .A2(_1409_));
 sg13g2_inv_1 _6743_ (.Y(_1412_),
    .A(_1411_));
 sg13g2_xnor2_1 _6744_ (.Y(_1414_),
    .A(net260),
    .B(net302));
 sg13g2_xnor2_1 _6745_ (.Y(_1415_),
    .A(_0183_),
    .B(net235));
 sg13g2_nand2_1 _6746_ (.Y(_1416_),
    .A(_1414_),
    .B(_1415_));
 sg13g2_nor2_1 _6747_ (.A(_1414_),
    .B(_1415_),
    .Y(_1417_));
 sg13g2_nand2_1 _6748_ (.Y(_1418_),
    .A(net58),
    .B(_1417_));
 sg13g2_o21ai_1 _6749_ (.B1(_1418_),
    .Y(_1419_),
    .A1(net58),
    .A2(_1416_));
 sg13g2_buf_1 _6750_ (.A(net214),
    .X(_1420_));
 sg13g2_nand2_1 _6751_ (.Y(_1421_),
    .A(_1420_),
    .B(net213));
 sg13g2_nor2_1 _6752_ (.A(_0656_),
    .B(_1686_),
    .Y(_1422_));
 sg13g2_nor2_1 _6753_ (.A(_0260_),
    .B(_1422_),
    .Y(_1423_));
 sg13g2_mux2_1 _6754_ (.A0(_3655_),
    .A1(_1421_),
    .S(_1423_),
    .X(_1425_));
 sg13g2_xnor2_1 _6755_ (.Y(_1426_),
    .A(net168),
    .B(_1396_));
 sg13g2_nor2_1 _6756_ (.A(_1405_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_nand3_1 _6757_ (.B(_1425_),
    .C(_1427_),
    .A(_1419_),
    .Y(_1428_));
 sg13g2_o21ai_1 _6758_ (.B1(_1428_),
    .Y(_1429_),
    .A1(_1406_),
    .A2(_1412_));
 sg13g2_nand2_1 _6759_ (.Y(_1430_),
    .A(_1355_),
    .B(_1429_));
 sg13g2_nand2_1 _6760_ (.Y(_1431_),
    .A(_3557_),
    .B(_1204_));
 sg13g2_nor2_1 _6761_ (.A(net268),
    .B(_1431_),
    .Y(_1432_));
 sg13g2_xnor2_1 _6762_ (.Y(_1433_),
    .A(net200),
    .B(_1432_));
 sg13g2_o21ai_1 _6763_ (.B1(_1433_),
    .Y(_1434_),
    .A1(_1355_),
    .A2(_1429_));
 sg13g2_nand2_1 _6764_ (.Y(_1436_),
    .A(_1430_),
    .B(_1434_));
 sg13g2_buf_1 _6765_ (.A(_4252_),
    .X(_1437_));
 sg13g2_inv_2 _6766_ (.Y(_1438_),
    .A(net267));
 sg13g2_nor2_1 _6767_ (.A(net200),
    .B(_1325_),
    .Y(_1439_));
 sg13g2_nor2_1 _6768_ (.A(_1438_),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_xnor2_1 _6769_ (.Y(_1441_),
    .A(net264),
    .B(_1440_));
 sg13g2_a21o_1 _6770_ (.A2(_1436_),
    .A1(_1354_),
    .B1(_1441_),
    .X(_1442_));
 sg13g2_o21ai_1 _6771_ (.B1(_1442_),
    .Y(_1443_),
    .A1(_1354_),
    .A2(_1436_));
 sg13g2_nor2_1 _6772_ (.A(_1352_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_nor2_1 _6773_ (.A(_3720_),
    .B(net217),
    .Y(_1445_));
 sg13g2_nand2_1 _6774_ (.Y(_1447_),
    .A(_1325_),
    .B(_1445_));
 sg13g2_xnor2_1 _6775_ (.Y(_1448_),
    .A(net246),
    .B(_1447_));
 sg13g2_a21oi_1 _6776_ (.A1(_1352_),
    .A2(_1443_),
    .Y(_1449_),
    .B1(_1448_));
 sg13g2_nor2_1 _6777_ (.A(_1444_),
    .B(_1449_),
    .Y(_1450_));
 sg13g2_buf_1 _6778_ (.A(net93),
    .X(_1451_));
 sg13g2_buf_1 _6779_ (.A(net57),
    .X(_1452_));
 sg13g2_nor2_1 _6780_ (.A(_4089_),
    .B(net37),
    .Y(_1453_));
 sg13g2_nand2_1 _6781_ (.Y(_1454_),
    .A(net245),
    .B(net267));
 sg13g2_o21ai_1 _6782_ (.B1(net246),
    .Y(_1455_),
    .A1(_1439_),
    .A2(_1454_));
 sg13g2_xnor2_1 _6783_ (.Y(_1456_),
    .A(net234),
    .B(_1455_));
 sg13g2_o21ai_1 _6784_ (.B1(_1456_),
    .Y(_1458_),
    .A1(_1936_),
    .A2(net38));
 sg13g2_a21oi_1 _6785_ (.A1(net193),
    .A2(_1453_),
    .Y(_1459_),
    .B1(_1458_));
 sg13g2_nand4_1 _6786_ (.B(_1356_),
    .C(_1450_),
    .A(_1352_),
    .Y(_1460_),
    .D(_1459_));
 sg13g2_inv_1 _6787_ (.Y(_1461_),
    .A(_1349_));
 sg13g2_o21ai_1 _6788_ (.B1(_1461_),
    .Y(_1462_),
    .A1(_1450_),
    .A2(_1456_));
 sg13g2_xor2_1 _6789_ (.B(_1331_),
    .A(_1335_),
    .X(_1463_));
 sg13g2_nand4_1 _6790_ (.B(net248),
    .C(net229),
    .A(net216),
    .Y(_1464_),
    .D(_1454_));
 sg13g2_nor4_2 _6791_ (.A(net310),
    .B(_0908_),
    .C(net311),
    .Y(_1465_),
    .D(net281));
 sg13g2_inv_1 _6792_ (.Y(_1466_),
    .A(net310));
 sg13g2_buf_1 _6793_ (.A(_1466_),
    .X(_1467_));
 sg13g2_nor4_1 _6794_ (.A(net225),
    .B(net234),
    .C(net218),
    .D(_1325_),
    .Y(_1469_));
 sg13g2_nand2_1 _6795_ (.Y(_1470_),
    .A(_3731_),
    .B(_1408_));
 sg13g2_o21ai_1 _6796_ (.B1(_1470_),
    .Y(_1471_),
    .A1(_1465_),
    .A2(_1469_));
 sg13g2_o21ai_1 _6797_ (.B1(_1445_),
    .Y(_1472_),
    .A1(net268),
    .A2(_1431_));
 sg13g2_nand3_1 _6798_ (.B(net248),
    .C(_1472_),
    .A(net216),
    .Y(_1473_));
 sg13g2_xnor2_1 _6799_ (.Y(_1474_),
    .A(net287),
    .B(_1473_));
 sg13g2_nand3_1 _6800_ (.B(_1471_),
    .C(_1474_),
    .A(_1464_),
    .Y(_1475_));
 sg13g2_a221oi_1 _6801_ (.B2(_1373_),
    .C1(_1475_),
    .B1(_1463_),
    .A1(_1460_),
    .Y(_1476_),
    .A2(_1462_));
 sg13g2_nand4_1 _6802_ (.B(_1371_),
    .C(_1381_),
    .A(_1370_),
    .Y(_1477_),
    .D(_1476_));
 sg13g2_a21oi_1 _6803_ (.A1(net253),
    .A2(_0868_),
    .Y(_1478_),
    .B1(net252));
 sg13g2_buf_1 _6804_ (.A(_1478_),
    .X(_1480_));
 sg13g2_buf_1 _6805_ (.A(_1480_),
    .X(_1481_));
 sg13g2_nor2_2 _6806_ (.A(net38),
    .B(net162),
    .Y(_1482_));
 sg13g2_buf_1 _6807_ (.A(_0007_),
    .X(_1483_));
 sg13g2_xnor2_1 _6808_ (.Y(_1484_),
    .A(net298),
    .B(_1349_));
 sg13g2_nand2_1 _6809_ (.Y(_1485_),
    .A(net287),
    .B(_1484_));
 sg13g2_xnor2_1 _6810_ (.Y(_1486_),
    .A(net304),
    .B(_1352_));
 sg13g2_xnor2_1 _6811_ (.Y(_1487_),
    .A(_4513_),
    .B(_1354_));
 sg13g2_nor3_1 _6812_ (.A(_1485_),
    .B(_1486_),
    .C(_1487_),
    .Y(_1488_));
 sg13g2_nor2_1 _6813_ (.A(net193),
    .B(net227),
    .Y(_1489_));
 sg13g2_nor2_1 _6814_ (.A(net219),
    .B(net231),
    .Y(_1491_));
 sg13g2_nor2_1 _6815_ (.A(_1489_),
    .B(_1491_),
    .Y(_1492_));
 sg13g2_xnor2_1 _6816_ (.Y(_1493_),
    .A(net220),
    .B(net268));
 sg13g2_xor2_1 _6817_ (.B(net299),
    .A(net243),
    .X(_1494_));
 sg13g2_buf_1 _6818_ (.A(_1494_),
    .X(_1495_));
 sg13g2_xnor2_1 _6819_ (.Y(_1496_),
    .A(net251),
    .B(net230));
 sg13g2_nand4_1 _6820_ (.B(_1493_),
    .C(_1495_),
    .A(_1492_),
    .Y(_1497_),
    .D(_1496_));
 sg13g2_nor4_1 _6821_ (.A(_1492_),
    .B(_1493_),
    .C(_1495_),
    .D(_1496_),
    .Y(_1498_));
 sg13g2_nand2_1 _6822_ (.Y(_1499_),
    .A(net38),
    .B(_1498_));
 sg13g2_o21ai_1 _6823_ (.B1(_1499_),
    .Y(_1500_),
    .A1(net38),
    .A2(_1497_));
 sg13g2_xor2_1 _6824_ (.B(net230),
    .A(net251),
    .X(_1502_));
 sg13g2_nand2_1 _6825_ (.Y(_1503_),
    .A(net254),
    .B(_1502_));
 sg13g2_nor2_1 _6826_ (.A(net220),
    .B(_1502_),
    .Y(_1504_));
 sg13g2_nand2_1 _6827_ (.Y(_1505_),
    .A(net93),
    .B(_1504_));
 sg13g2_o21ai_1 _6828_ (.B1(_1505_),
    .Y(_1506_),
    .A1(net93),
    .A2(_1503_));
 sg13g2_xnor2_1 _6829_ (.Y(_1507_),
    .A(net207),
    .B(net38));
 sg13g2_a22oi_1 _6830_ (.Y(_1508_),
    .B1(_1507_),
    .B2(net172),
    .A2(_1506_),
    .A1(_4525_));
 sg13g2_o21ai_1 _6831_ (.B1(net215),
    .Y(_1509_),
    .A1(net227),
    .A2(_1508_));
 sg13g2_nor3_1 _6832_ (.A(net231),
    .B(_1410_),
    .C(_1508_),
    .Y(_1510_));
 sg13g2_a21o_1 _6833_ (.A2(_1509_),
    .A1(_1410_),
    .B1(_1510_),
    .X(_1511_));
 sg13g2_nand2_1 _6834_ (.Y(_1513_),
    .A(net179),
    .B(_1355_));
 sg13g2_a22oi_1 _6835_ (.Y(_1514_),
    .B1(_1511_),
    .B2(_1513_),
    .A2(_1500_),
    .A1(_1388_));
 sg13g2_o21ai_1 _6836_ (.B1(_1514_),
    .Y(_1515_),
    .A1(net179),
    .A2(_1355_));
 sg13g2_nor3_1 _6837_ (.A(_4513_),
    .B(_1354_),
    .C(_1486_),
    .Y(_1516_));
 sg13g2_a21oi_1 _6838_ (.A1(net225),
    .A2(_1352_),
    .Y(_1517_),
    .B1(_1516_));
 sg13g2_nand2_1 _6839_ (.Y(_1518_),
    .A(net192),
    .B(_1461_));
 sg13g2_o21ai_1 _6840_ (.B1(_1518_),
    .Y(_1519_),
    .A1(_1485_),
    .A2(_1517_));
 sg13g2_a21oi_1 _6841_ (.A1(_1488_),
    .A2(_1515_),
    .Y(_1520_),
    .B1(_1519_));
 sg13g2_nand3_1 _6842_ (.B(_1488_),
    .C(_1500_),
    .A(_1419_),
    .Y(_1521_));
 sg13g2_nor2b_2 _6843_ (.A(_1520_),
    .B_N(_1521_),
    .Y(_1522_));
 sg13g2_nor2_1 _6844_ (.A(_1482_),
    .B(_1522_),
    .Y(_1524_));
 sg13g2_nor2b_1 _6845_ (.A(net155),
    .B_N(_0902_),
    .Y(_1525_));
 sg13g2_buf_1 _6846_ (.A(_1525_),
    .X(_1526_));
 sg13g2_buf_1 _6847_ (.A(_1526_),
    .X(_1527_));
 sg13g2_nand2_1 _6848_ (.Y(_1528_),
    .A(net205),
    .B(_2239_));
 sg13g2_nand3_1 _6849_ (.B(net301),
    .C(_2480_),
    .A(_2415_),
    .Y(_1529_));
 sg13g2_o21ai_1 _6850_ (.B1(_1529_),
    .Y(_1530_),
    .A1(net301),
    .A2(_1528_));
 sg13g2_buf_2 _6851_ (.A(_1530_),
    .X(_1531_));
 sg13g2_and2_1 _6852_ (.A(_1531_),
    .B(_0888_),
    .X(_1532_));
 sg13g2_buf_2 _6853_ (.A(_1532_),
    .X(_1533_));
 sg13g2_nand2_1 _6854_ (.Y(_1535_),
    .A(net92),
    .B(_1533_));
 sg13g2_a21oi_1 _6855_ (.A1(_1477_),
    .A2(_1524_),
    .Y(_1536_),
    .B1(_1535_));
 sg13g2_nand2b_1 _6856_ (.Y(_1537_),
    .B(_0902_),
    .A_N(net155));
 sg13g2_buf_2 _6857_ (.A(_1537_),
    .X(_1538_));
 sg13g2_buf_1 _6858_ (.A(_1538_),
    .X(_1539_));
 sg13g2_buf_1 _6859_ (.A(_1539_),
    .X(_1540_));
 sg13g2_nand2b_1 _6860_ (.Y(_1541_),
    .B(_2261_),
    .A_N(net300));
 sg13g2_nand3_1 _6861_ (.B(net1),
    .C(_2972_),
    .A(_0881_),
    .Y(_1542_));
 sg13g2_o21ai_1 _6862_ (.B1(_1542_),
    .Y(_1543_),
    .A1(_2272_),
    .A2(_1541_));
 sg13g2_buf_2 _6863_ (.A(_1543_),
    .X(_1544_));
 sg13g2_and2_1 _6864_ (.A(_1544_),
    .B(_0891_),
    .X(_1546_));
 sg13g2_buf_1 _6865_ (.A(_1546_),
    .X(_1547_));
 sg13g2_buf_1 _6866_ (.A(net38),
    .X(_1548_));
 sg13g2_nand2_1 _6867_ (.Y(_1549_),
    .A(net253),
    .B(_0868_));
 sg13g2_nand2_1 _6868_ (.Y(_1550_),
    .A(net256),
    .B(_1549_));
 sg13g2_buf_1 _6869_ (.A(_1550_),
    .X(_1551_));
 sg13g2_buf_1 _6870_ (.A(_1551_),
    .X(_1552_));
 sg13g2_nand3b_1 _6871_ (.B(net300),
    .C(_2480_),
    .Y(_1553_),
    .A_N(_2415_));
 sg13g2_o21ai_1 _6872_ (.B1(_1553_),
    .Y(_1554_),
    .A1(net301),
    .A2(_2535_));
 sg13g2_buf_1 _6873_ (.A(_1554_),
    .X(_1555_));
 sg13g2_nand2_1 _6874_ (.Y(_1557_),
    .A(net152),
    .B(_0888_));
 sg13g2_buf_1 _6875_ (.A(_1557_),
    .X(_1558_));
 sg13g2_buf_1 _6876_ (.A(_0893_),
    .X(_1559_));
 sg13g2_o21ai_1 _6877_ (.B1(net55),
    .Y(_1560_),
    .A1(net90),
    .A2(_1548_));
 sg13g2_nor2_1 _6878_ (.A(_2415_),
    .B(_2480_),
    .Y(_1561_));
 sg13g2_nor3_1 _6879_ (.A(net205),
    .B(net300),
    .C(_2239_),
    .Y(_1562_));
 sg13g2_a21o_1 _6880_ (.A2(_1561_),
    .A1(net301),
    .B1(_1562_),
    .X(_1563_));
 sg13g2_buf_2 _6881_ (.A(_1563_),
    .X(_1564_));
 sg13g2_and2_1 _6882_ (.A(_1564_),
    .B(_0888_),
    .X(_1565_));
 sg13g2_buf_2 _6883_ (.A(_1565_),
    .X(_1566_));
 sg13g2_a221oi_1 _6884_ (.B2(_1560_),
    .C1(_1566_),
    .B1(net153),
    .A1(_1547_),
    .Y(_1568_),
    .A2(net24));
 sg13g2_nor2_1 _6885_ (.A(net56),
    .B(_1568_),
    .Y(_1569_));
 sg13g2_and2_1 _6886_ (.A(_1544_),
    .B(_1531_),
    .X(_1570_));
 sg13g2_buf_2 _6887_ (.A(_1570_),
    .X(_1571_));
 sg13g2_nor2_1 _6888_ (.A(net188),
    .B(_0852_),
    .Y(_1572_));
 sg13g2_buf_2 _6889_ (.A(_1572_),
    .X(_1573_));
 sg13g2_nand2_1 _6890_ (.Y(_1574_),
    .A(_1571_),
    .B(_1573_));
 sg13g2_and2_1 _6891_ (.A(net152),
    .B(_0888_),
    .X(_1575_));
 sg13g2_buf_2 _6892_ (.A(_1575_),
    .X(_1576_));
 sg13g2_buf_1 _6893_ (.A(net130),
    .X(_1577_));
 sg13g2_buf_1 _6894_ (.A(net89),
    .X(_1579_));
 sg13g2_buf_1 _6895_ (.A(net54),
    .X(_1580_));
 sg13g2_nor2_1 _6896_ (.A(_1708_),
    .B(_1468_),
    .Y(_1581_));
 sg13g2_o21ai_1 _6897_ (.B1(net207),
    .Y(_1582_),
    .A1(net220),
    .A2(_1581_));
 sg13g2_nand2_1 _6898_ (.Y(_1583_),
    .A(_1357_),
    .B(_1582_));
 sg13g2_nand3_1 _6899_ (.B(_4392_),
    .C(_1534_),
    .A(_0260_),
    .Y(_1584_));
 sg13g2_nand2_1 _6900_ (.Y(_1585_),
    .A(_0839_),
    .B(_1584_));
 sg13g2_o21ai_1 _6901_ (.B1(net221),
    .Y(_1586_),
    .A1(_1583_),
    .A2(_1585_));
 sg13g2_buf_2 _6902_ (.A(_1586_),
    .X(_1587_));
 sg13g2_a22oi_1 _6903_ (.Y(_1588_),
    .B1(_1587_),
    .B2(_1533_),
    .A2(net36),
    .A1(_1576_));
 sg13g2_nand2_1 _6904_ (.Y(_1590_),
    .A(_3233_),
    .B(_0900_));
 sg13g2_o21ai_1 _6905_ (.B1(_1590_),
    .Y(_1591_),
    .A1(net5),
    .A2(_0899_));
 sg13g2_buf_1 _6906_ (.A(_1591_),
    .X(_1592_));
 sg13g2_nand2b_1 _6907_ (.Y(_1593_),
    .B(_1592_),
    .A_N(net155));
 sg13g2_buf_1 _6908_ (.A(_1593_),
    .X(_1594_));
 sg13g2_buf_1 _6909_ (.A(net88),
    .X(_1595_));
 sg13g2_a21oi_1 _6910_ (.A1(_1574_),
    .A2(_1588_),
    .Y(_1596_),
    .B1(net53));
 sg13g2_nor3_1 _6911_ (.A(_1536_),
    .B(_1569_),
    .C(_1596_),
    .Y(_1597_));
 sg13g2_nor2b_1 _6912_ (.A(net155),
    .B_N(_1592_),
    .Y(_1598_));
 sg13g2_buf_1 _6913_ (.A(_1598_),
    .X(_1599_));
 sg13g2_buf_1 _6914_ (.A(_1599_),
    .X(_1600_));
 sg13g2_nand2_1 _6915_ (.Y(_1601_),
    .A(_1544_),
    .B(_0891_));
 sg13g2_buf_1 _6916_ (.A(_1601_),
    .X(_1602_));
 sg13g2_buf_1 _6917_ (.A(_4072_),
    .X(_1603_));
 sg13g2_xnor2_1 _6918_ (.Y(_1604_),
    .A(_0557_),
    .B(_0645_));
 sg13g2_nand2_1 _6919_ (.Y(_1605_),
    .A(net137),
    .B(_1604_));
 sg13g2_o21ai_1 _6920_ (.B1(_1605_),
    .Y(_1606_),
    .A1(_4074_),
    .A2(net137));
 sg13g2_buf_2 _6921_ (.A(_1606_),
    .X(_1607_));
 sg13g2_buf_1 _6922_ (.A(_1607_),
    .X(_1608_));
 sg13g2_or3_1 _6923_ (.A(net279),
    .B(net309),
    .C(net308),
    .X(_1609_));
 sg13g2_buf_2 _6924_ (.A(_1609_),
    .X(_1611_));
 sg13g2_o21ai_1 _6925_ (.B1(net217),
    .Y(_1612_),
    .A1(_4545_),
    .A2(_1611_));
 sg13g2_xnor2_1 _6926_ (.Y(_1613_),
    .A(net225),
    .B(_1612_));
 sg13g2_inv_1 _6927_ (.Y(_1614_),
    .A(_1613_));
 sg13g2_nor2_1 _6928_ (.A(net35),
    .B(_1614_),
    .Y(_1615_));
 sg13g2_or2_1 _6929_ (.X(_1616_),
    .B(net309),
    .A(_1226_));
 sg13g2_buf_1 _6930_ (.A(_1616_),
    .X(_1617_));
 sg13g2_nor2_1 _6931_ (.A(_3482_),
    .B(_1617_),
    .Y(_1618_));
 sg13g2_xnor2_1 _6932_ (.Y(_1619_),
    .A(_1438_),
    .B(_1618_));
 sg13g2_xnor2_1 _6933_ (.Y(_1620_),
    .A(net267),
    .B(net299));
 sg13g2_nand2_1 _6934_ (.Y(_1622_),
    .A(_1421_),
    .B(_1620_));
 sg13g2_xnor2_1 _6935_ (.Y(_1623_),
    .A(net244),
    .B(_1620_));
 sg13g2_nand3_1 _6936_ (.B(_1390_),
    .C(_1623_),
    .A(net231),
    .Y(_1624_));
 sg13g2_o21ai_1 _6937_ (.B1(_1624_),
    .Y(_1625_),
    .A1(net231),
    .A2(_1622_));
 sg13g2_nand2_1 _6938_ (.Y(_1626_),
    .A(net233),
    .B(_4080_));
 sg13g2_a21oi_1 _6939_ (.A1(net296),
    .A2(_4093_),
    .Y(_1627_),
    .B1(net233));
 sg13g2_nand2_1 _6940_ (.Y(_1628_),
    .A(_4418_),
    .B(_1627_));
 sg13g2_nand2_1 _6941_ (.Y(_1629_),
    .A(_1626_),
    .B(_1628_));
 sg13g2_buf_1 _6942_ (.A(_1629_),
    .X(_1630_));
 sg13g2_buf_1 _6943_ (.A(net118),
    .X(_1631_));
 sg13g2_a22oi_1 _6944_ (.Y(_1633_),
    .B1(_1625_),
    .B2(net87),
    .A2(_1619_),
    .A1(net224));
 sg13g2_xnor2_1 _6945_ (.Y(_1634_),
    .A(net288),
    .B(net89));
 sg13g2_buf_1 _6946_ (.A(_1634_),
    .X(_1635_));
 sg13g2_xnor2_1 _6947_ (.Y(_1636_),
    .A(net293),
    .B(net89));
 sg13g2_buf_1 _6948_ (.A(_1636_),
    .X(_1637_));
 sg13g2_a21oi_1 _6949_ (.A1(net209),
    .A2(net137),
    .Y(_1638_),
    .B1(_0384_));
 sg13g2_nor2_1 _6950_ (.A(_3805_),
    .B(net302),
    .Y(_1639_));
 sg13g2_nand2_1 _6951_ (.Y(_1640_),
    .A(net208),
    .B(_1639_));
 sg13g2_o21ai_1 _6952_ (.B1(_1640_),
    .Y(_1641_),
    .A1(net208),
    .A2(net130));
 sg13g2_mux2_1 _6953_ (.A0(net130),
    .A1(_1639_),
    .S(net190),
    .X(_1642_));
 sg13g2_mux2_1 _6954_ (.A0(_1641_),
    .A1(_1642_),
    .S(net209),
    .X(_1644_));
 sg13g2_nor3_1 _6955_ (.A(net178),
    .B(_4438_),
    .C(_1638_),
    .Y(_1645_));
 sg13g2_a221oi_1 _6956_ (.B2(_3364_),
    .C1(_1645_),
    .B1(_1644_),
    .A1(_4438_),
    .Y(_1646_),
    .A2(_1638_));
 sg13g2_buf_1 _6957_ (.A(_1646_),
    .X(_1647_));
 sg13g2_or2_1 _6958_ (.X(_1648_),
    .B(_1647_),
    .A(net33));
 sg13g2_nand2_1 _6959_ (.Y(_1649_),
    .A(net34),
    .B(_1648_));
 sg13g2_nand2_1 _6960_ (.Y(_1650_),
    .A(net33),
    .B(_1647_));
 sg13g2_xnor2_1 _6961_ (.Y(_1651_),
    .A(net255),
    .B(net89));
 sg13g2_buf_2 _6962_ (.A(_1651_),
    .X(_1652_));
 sg13g2_a22oi_1 _6963_ (.Y(_1653_),
    .B1(_1650_),
    .B2(_1652_),
    .A2(_1649_),
    .A1(net160));
 sg13g2_nand2_1 _6964_ (.Y(_1655_),
    .A(_1421_),
    .B(_1648_));
 sg13g2_nand2_1 _6965_ (.Y(_1656_),
    .A(_1390_),
    .B(_1623_));
 sg13g2_and2_1 _6966_ (.A(_1626_),
    .B(_1628_),
    .X(_1657_));
 sg13g2_buf_1 _6967_ (.A(_1657_),
    .X(_1658_));
 sg13g2_xnor2_1 _6968_ (.Y(_1659_),
    .A(net231),
    .B(net117));
 sg13g2_mux2_1 _6969_ (.A0(_1622_),
    .A1(_1656_),
    .S(_1659_),
    .X(_1660_));
 sg13g2_a221oi_1 _6970_ (.B2(_1652_),
    .C1(_1660_),
    .B1(_1655_),
    .A1(_1390_),
    .Y(_1661_),
    .A2(_1650_));
 sg13g2_o21ai_1 _6971_ (.B1(_1661_),
    .Y(_1662_),
    .A1(net172),
    .A2(_1653_));
 sg13g2_xnor2_1 _6972_ (.Y(_1663_),
    .A(net201),
    .B(net34));
 sg13g2_nand3b_1 _6973_ (.B(_1663_),
    .C(net160),
    .Y(_1664_),
    .A_N(net33));
 sg13g2_nand2_1 _6974_ (.Y(_1666_),
    .A(net213),
    .B(net33));
 sg13g2_or2_1 _6975_ (.X(_1667_),
    .B(_1663_),
    .A(_1666_));
 sg13g2_a21oi_1 _6976_ (.A1(_1664_),
    .A2(_1667_),
    .Y(_1668_),
    .B1(_1660_));
 sg13g2_nand2_1 _6977_ (.Y(_1669_),
    .A(net54),
    .B(_1417_));
 sg13g2_o21ai_1 _6978_ (.B1(_1669_),
    .Y(_1670_),
    .A1(net54),
    .A2(_1416_));
 sg13g2_buf_1 _6979_ (.A(_1670_),
    .X(_1671_));
 sg13g2_a22oi_1 _6980_ (.Y(_1672_),
    .B1(_1668_),
    .B2(_1671_),
    .A2(_1662_),
    .A1(_1633_));
 sg13g2_xnor2_1 _6981_ (.Y(_1673_),
    .A(_1073_),
    .B(_4111_));
 sg13g2_nand2_1 _6982_ (.Y(_1674_),
    .A(_1672_),
    .B(_1673_));
 sg13g2_nand2_1 _6983_ (.Y(_1675_),
    .A(_1001_),
    .B(_1577_));
 sg13g2_nand2_1 _6984_ (.Y(_1676_),
    .A(net137),
    .B(_1353_));
 sg13g2_nand2_1 _6985_ (.Y(_1677_),
    .A(_1675_),
    .B(_1676_));
 sg13g2_buf_1 _6986_ (.A(_1677_),
    .X(_1678_));
 sg13g2_o21ai_1 _6987_ (.B1(net23),
    .Y(_1679_),
    .A1(_1672_),
    .A2(_1673_));
 sg13g2_nand2_1 _6988_ (.Y(_1680_),
    .A(_1674_),
    .B(_1679_));
 sg13g2_nor2_1 _6989_ (.A(net286),
    .B(net298),
    .Y(_1681_));
 sg13g2_nor2_1 _6990_ (.A(_0941_),
    .B(_4111_),
    .Y(_1682_));
 sg13g2_mux2_1 _6991_ (.A0(net298),
    .A1(_1681_),
    .S(_1682_),
    .X(_1683_));
 sg13g2_nand2_1 _6992_ (.Y(_1684_),
    .A(net286),
    .B(net218));
 sg13g2_nor3_1 _6993_ (.A(net287),
    .B(net298),
    .C(_1684_),
    .Y(_1685_));
 sg13g2_a22oi_1 _6994_ (.Y(_1687_),
    .B1(_1685_),
    .B2(_1682_),
    .A2(_1683_),
    .A1(net287));
 sg13g2_a21oi_1 _6995_ (.A1(net35),
    .A2(_1614_),
    .Y(_1688_),
    .B1(_1687_));
 sg13g2_o21ai_1 _6996_ (.B1(_1688_),
    .Y(_1689_),
    .A1(_1615_),
    .A2(_1680_));
 sg13g2_buf_1 _6997_ (.A(_1689_),
    .X(_1690_));
 sg13g2_xnor2_1 _6998_ (.Y(_1691_),
    .A(net181),
    .B(net33));
 sg13g2_and2_1 _6999_ (.A(_4525_),
    .B(net33),
    .X(_1692_));
 sg13g2_a21o_1 _7000_ (.A2(_1691_),
    .A1(_1647_),
    .B1(_1692_),
    .X(_1693_));
 sg13g2_nand2b_1 _7001_ (.Y(_1694_),
    .B(_1652_),
    .A_N(_1693_));
 sg13g2_nor3_1 _7002_ (.A(net242),
    .B(_1617_),
    .C(_1620_),
    .Y(_1695_));
 sg13g2_a21oi_1 _7003_ (.A1(_1617_),
    .A2(_1620_),
    .Y(_1696_),
    .B1(_1695_));
 sg13g2_and2_1 _7004_ (.A(_1675_),
    .B(_1676_),
    .X(_1698_));
 sg13g2_buf_1 _7005_ (.A(_1698_),
    .X(_1699_));
 sg13g2_xnor2_1 _7006_ (.Y(_1700_),
    .A(_4252_),
    .B(_1699_));
 sg13g2_nor2b_1 _7007_ (.A(_1696_),
    .B_N(_1700_),
    .Y(_1701_));
 sg13g2_nor4_1 _7008_ (.A(net200),
    .B(_1700_),
    .C(_1617_),
    .D(_1620_),
    .Y(_1702_));
 sg13g2_or2_1 _7009_ (.X(_1703_),
    .B(_1702_),
    .A(_1701_));
 sg13g2_o21ai_1 _7010_ (.B1(_1703_),
    .Y(_1704_),
    .A1(net87),
    .A2(_1694_));
 sg13g2_a21oi_1 _7011_ (.A1(net87),
    .A2(_1694_),
    .Y(_1705_),
    .B1(_1431_));
 sg13g2_and2_1 _7012_ (.A(net34),
    .B(_1693_),
    .X(_1706_));
 sg13g2_buf_1 _7013_ (.A(_1706_),
    .X(_1707_));
 sg13g2_a21oi_1 _7014_ (.A1(net215),
    .A2(net118),
    .Y(_1709_),
    .B1(_1707_));
 sg13g2_a21oi_1 _7015_ (.A1(net191),
    .A2(net117),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_nor2_1 _7016_ (.A(net180),
    .B(_1710_),
    .Y(_1711_));
 sg13g2_nor3_1 _7017_ (.A(_1704_),
    .B(_1705_),
    .C(_1711_),
    .Y(_1712_));
 sg13g2_nor2_1 _7018_ (.A(net267),
    .B(net299),
    .Y(_1713_));
 sg13g2_nor2_1 _7019_ (.A(net23),
    .B(_1713_),
    .Y(_1714_));
 sg13g2_nor3_1 _7020_ (.A(net179),
    .B(net264),
    .C(_1714_),
    .Y(_1715_));
 sg13g2_a21oi_1 _7021_ (.A1(net23),
    .A2(_1713_),
    .Y(_1716_),
    .B1(_1715_));
 sg13g2_buf_1 _7022_ (.A(net299),
    .X(_1717_));
 sg13g2_nor2_2 _7023_ (.A(net279),
    .B(net309),
    .Y(_1718_));
 sg13g2_nor3_1 _7024_ (.A(_1438_),
    .B(net263),
    .C(_1718_),
    .Y(_1720_));
 sg13g2_a21oi_1 _7025_ (.A1(net267),
    .A2(net226),
    .Y(_1721_),
    .B1(net23));
 sg13g2_and2_1 _7026_ (.A(_1718_),
    .B(_1713_),
    .X(_1722_));
 sg13g2_o21ai_1 _7027_ (.B1(_3720_),
    .Y(_1723_),
    .A1(net23),
    .A2(_1722_));
 sg13g2_o21ai_1 _7028_ (.B1(_1723_),
    .Y(_1724_),
    .A1(_1718_),
    .A2(_1721_));
 sg13g2_a22oi_1 _7029_ (.Y(_1725_),
    .B1(_1724_),
    .B2(net264),
    .A2(_1720_),
    .A1(net23));
 sg13g2_o21ai_1 _7030_ (.B1(_1725_),
    .Y(_1726_),
    .A1(_1617_),
    .A2(_1716_));
 sg13g2_nand2_1 _7031_ (.Y(_1727_),
    .A(net172),
    .B(_1635_));
 sg13g2_xnor2_1 _7032_ (.Y(_1728_),
    .A(_1407_),
    .B(net117));
 sg13g2_nand3_1 _7033_ (.B(_1652_),
    .C(_1728_),
    .A(net180),
    .Y(_1729_));
 sg13g2_o21ai_1 _7034_ (.B1(_1729_),
    .Y(_1731_),
    .A1(_1727_),
    .A2(_1728_));
 sg13g2_nand4_1 _7035_ (.B(_1671_),
    .C(_1703_),
    .A(_1691_),
    .Y(_1732_),
    .D(_1731_));
 sg13g2_o21ai_1 _7036_ (.B1(_1732_),
    .Y(_1733_),
    .A1(_1712_),
    .A2(_1726_));
 sg13g2_a21o_1 _7037_ (.A2(_1718_),
    .A1(_1445_),
    .B1(net225),
    .X(_1734_));
 sg13g2_buf_1 _7038_ (.A(_1734_),
    .X(_1735_));
 sg13g2_nand3_1 _7039_ (.B(_1445_),
    .C(_1718_),
    .A(net225),
    .Y(_1736_));
 sg13g2_a22oi_1 _7040_ (.Y(_1737_),
    .B1(_1735_),
    .B2(_1736_),
    .A2(_1733_),
    .A1(net35));
 sg13g2_nor2_1 _7041_ (.A(net35),
    .B(_1733_),
    .Y(_1738_));
 sg13g2_mux2_1 _7042_ (.A0(_1681_),
    .A1(net298),
    .S(_1735_),
    .X(_1739_));
 sg13g2_nor4_1 _7043_ (.A(net287),
    .B(net298),
    .C(_1684_),
    .D(_1735_),
    .Y(_1740_));
 sg13g2_a21o_1 _7044_ (.A2(_1739_),
    .A1(net287),
    .B1(_1740_),
    .X(_1742_));
 sg13g2_o21ai_1 _7045_ (.B1(_1742_),
    .Y(_1743_),
    .A1(_1737_),
    .A2(_1738_));
 sg13g2_and2_1 _7046_ (.A(_1690_),
    .B(_1743_),
    .X(_1744_));
 sg13g2_buf_1 _7047_ (.A(_1744_),
    .X(_1745_));
 sg13g2_nor2_1 _7048_ (.A(net261),
    .B(net118),
    .Y(_1746_));
 sg13g2_nand2_1 _7049_ (.Y(_1747_),
    .A(_1686_),
    .B(net89));
 sg13g2_nand3_1 _7050_ (.B(net254),
    .C(net137),
    .A(net251),
    .Y(_1748_));
 sg13g2_o21ai_1 _7051_ (.B1(_1748_),
    .Y(_1749_),
    .A1(net251),
    .A2(_1747_));
 sg13g2_and2_1 _7052_ (.A(_1746_),
    .B(_1749_),
    .X(_1750_));
 sg13g2_xnor2_1 _7053_ (.Y(_1751_),
    .A(net23),
    .B(_1750_));
 sg13g2_nor2_1 _7054_ (.A(net264),
    .B(_1751_),
    .Y(_1753_));
 sg13g2_xnor2_1 _7055_ (.Y(_1754_),
    .A(_4116_),
    .B(_1607_));
 sg13g2_buf_2 _7056_ (.A(_1754_),
    .X(_1755_));
 sg13g2_buf_1 _7057_ (.A(_1699_),
    .X(_1756_));
 sg13g2_nand2_1 _7058_ (.Y(_1757_),
    .A(net117),
    .B(_1652_));
 sg13g2_buf_1 _7059_ (.A(_1757_),
    .X(_1758_));
 sg13g2_o21ai_1 _7060_ (.B1(net299),
    .Y(_1759_),
    .A1(net33),
    .A2(_1758_));
 sg13g2_o21ai_1 _7061_ (.B1(net184),
    .Y(_1760_),
    .A1(_1756_),
    .A2(_1759_));
 sg13g2_xor2_1 _7062_ (.B(_1760_),
    .A(_1755_),
    .X(_1761_));
 sg13g2_inv_1 _7063_ (.Y(_1762_),
    .A(_0820_));
 sg13g2_nor3_1 _7064_ (.A(_1607_),
    .B(net20),
    .C(_1750_),
    .Y(_1764_));
 sg13g2_xnor2_1 _7065_ (.Y(_1765_),
    .A(net298),
    .B(_1764_));
 sg13g2_nor2_1 _7066_ (.A(_1762_),
    .B(_1765_),
    .Y(_1766_));
 sg13g2_nand2_1 _7067_ (.Y(_1767_),
    .A(net137),
    .B(_1494_));
 sg13g2_o21ai_1 _7068_ (.B1(_1767_),
    .Y(_1768_),
    .A1(net171),
    .A2(_1747_));
 sg13g2_nand2_1 _7069_ (.Y(_1769_),
    .A(net255),
    .B(_1768_));
 sg13g2_o21ai_1 _7070_ (.B1(_1769_),
    .Y(_1770_),
    .A1(net220),
    .A2(_1767_));
 sg13g2_and2_1 _7071_ (.A(net89),
    .B(net171),
    .X(_1771_));
 sg13g2_nor3_1 _7072_ (.A(net210),
    .B(net89),
    .C(net171),
    .Y(_1772_));
 sg13g2_o21ai_1 _7073_ (.B1(net207),
    .Y(_1773_),
    .A1(_1771_),
    .A2(_1772_));
 sg13g2_nand2_1 _7074_ (.Y(_1775_),
    .A(_0447_),
    .B(_1771_));
 sg13g2_nand3_1 _7075_ (.B(_1773_),
    .C(_1775_),
    .A(net186),
    .Y(_1776_));
 sg13g2_o21ai_1 _7076_ (.B1(_1776_),
    .Y(_1777_),
    .A1(net186),
    .A2(_1770_));
 sg13g2_o21ai_1 _7077_ (.B1(net187),
    .Y(_1778_),
    .A1(_0522_),
    .A2(net137));
 sg13g2_xnor2_1 _7078_ (.Y(_1779_),
    .A(net193),
    .B(_1778_));
 sg13g2_nand3_1 _7079_ (.B(net171),
    .C(_1779_),
    .A(net227),
    .Y(_1780_));
 sg13g2_o21ai_1 _7080_ (.B1(_1780_),
    .Y(_1781_),
    .A1(net227),
    .A2(_1777_));
 sg13g2_nand2_1 _7081_ (.Y(_1782_),
    .A(_1437_),
    .B(_1751_));
 sg13g2_xnor2_1 _7082_ (.Y(_1783_),
    .A(net160),
    .B(net54));
 sg13g2_nand2_1 _7083_ (.Y(_1784_),
    .A(_1504_),
    .B(_1783_));
 sg13g2_o21ai_1 _7084_ (.B1(_1784_),
    .Y(_1786_),
    .A1(_1503_),
    .A2(_1783_));
 sg13g2_nand4_1 _7085_ (.B(_1781_),
    .C(_1782_),
    .A(_1766_),
    .Y(_1787_),
    .D(_1786_));
 sg13g2_nor3_1 _7086_ (.A(_1753_),
    .B(_1761_),
    .C(_1787_),
    .Y(_1788_));
 sg13g2_nor2_1 _7087_ (.A(net286),
    .B(_1762_),
    .Y(_1789_));
 sg13g2_nor2_1 _7088_ (.A(_1753_),
    .B(_1761_),
    .Y(_1790_));
 sg13g2_nor2_1 _7089_ (.A(net54),
    .B(_1503_),
    .Y(_1791_));
 sg13g2_a21oi_1 _7090_ (.A1(net54),
    .A2(_1504_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_nand2_1 _7091_ (.Y(_1793_),
    .A(net172),
    .B(_1423_));
 sg13g2_o21ai_1 _7092_ (.B1(_1793_),
    .Y(_1794_),
    .A1(net160),
    .A2(_1792_));
 sg13g2_nand2_1 _7093_ (.Y(_1795_),
    .A(_1781_),
    .B(_1794_));
 sg13g2_nor2_1 _7094_ (.A(net33),
    .B(_1758_),
    .Y(_1796_));
 sg13g2_nor2_1 _7095_ (.A(_0145_),
    .B(_0522_),
    .Y(_1797_));
 sg13g2_and2_1 _7096_ (.A(net187),
    .B(_1603_),
    .X(_1798_));
 sg13g2_a22oi_1 _7097_ (.Y(_1799_),
    .B1(_1798_),
    .B2(_1357_),
    .A2(_1797_),
    .A1(_1577_));
 sg13g2_a22oi_1 _7098_ (.Y(_1800_),
    .B1(_1799_),
    .B2(net179),
    .A2(_1796_),
    .A1(net215));
 sg13g2_nor2_1 _7099_ (.A(net200),
    .B(_1799_),
    .Y(_1801_));
 sg13g2_nor2_1 _7100_ (.A(_1759_),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_a21oi_1 _7101_ (.A1(net242),
    .A2(_1759_),
    .Y(_1803_),
    .B1(net191));
 sg13g2_nor2_1 _7102_ (.A(_1802_),
    .B(_1803_),
    .Y(_1804_));
 sg13g2_o21ai_1 _7103_ (.B1(_1804_),
    .Y(_1805_),
    .A1(net263),
    .A2(_1800_));
 sg13g2_nand3_1 _7104_ (.B(_1782_),
    .C(_1805_),
    .A(_1795_),
    .Y(_1807_));
 sg13g2_xnor2_1 _7105_ (.Y(_1808_),
    .A(_1608_),
    .B(_1760_));
 sg13g2_a22oi_1 _7106_ (.Y(_1809_),
    .B1(_1808_),
    .B2(net225),
    .A2(_1807_),
    .A1(_1790_));
 sg13g2_nor2b_1 _7107_ (.A(_1809_),
    .B_N(_1766_),
    .Y(_1810_));
 sg13g2_a221oi_1 _7108_ (.B2(_1764_),
    .C1(_1810_),
    .B1(_1789_),
    .A1(_1647_),
    .Y(_1811_),
    .A2(_1788_));
 sg13g2_a21oi_2 _7109_ (.B1(_1811_),
    .Y(_1812_),
    .A2(_1788_),
    .A1(_1671_));
 sg13g2_buf_1 _7110_ (.A(_1603_),
    .X(_1813_));
 sg13g2_buf_1 _7111_ (.A(net116),
    .X(_1814_));
 sg13g2_o21ai_1 _7112_ (.B1(net188),
    .Y(_1815_),
    .A1(_3976_),
    .A2(_0838_));
 sg13g2_buf_1 _7113_ (.A(_1815_),
    .X(_1816_));
 sg13g2_nor2_1 _7114_ (.A(net118),
    .B(net34),
    .Y(_1818_));
 sg13g2_nor2_2 _7115_ (.A(net261),
    .B(_1677_),
    .Y(_1819_));
 sg13g2_and2_1 _7116_ (.A(_1818_),
    .B(_1819_),
    .X(_1820_));
 sg13g2_nor2_1 _7117_ (.A(net35),
    .B(_1820_),
    .Y(_1821_));
 sg13g2_nand2_1 _7118_ (.Y(_1822_),
    .A(net299),
    .B(_1758_));
 sg13g2_nand2_1 _7119_ (.Y(_1823_),
    .A(_1819_),
    .B(_1822_));
 sg13g2_xor2_1 _7120_ (.B(_1823_),
    .A(net35),
    .X(_1824_));
 sg13g2_a21oi_1 _7121_ (.A1(net206),
    .A2(_1818_),
    .Y(_1825_),
    .B1(net20));
 sg13g2_o21ai_1 _7122_ (.B1(net264),
    .Y(_1826_),
    .A1(_1820_),
    .A2(_1825_));
 sg13g2_o21ai_1 _7123_ (.B1(_1106_),
    .Y(_1827_),
    .A1(_1087_),
    .A2(_0840_));
 sg13g2_o21ai_1 _7124_ (.B1(_1628_),
    .Y(_1829_),
    .A1(net219),
    .A2(_1095_));
 sg13g2_a21oi_1 _7125_ (.A1(net219),
    .A2(net200),
    .Y(_1830_),
    .B1(net207));
 sg13g2_nand2_1 _7126_ (.Y(_1831_),
    .A(net193),
    .B(_4162_));
 sg13g2_a221oi_1 _7127_ (.B2(_1831_),
    .C1(net299),
    .B1(_1830_),
    .A1(net207),
    .Y(_1832_),
    .A2(_1829_));
 sg13g2_a21oi_1 _7128_ (.A1(net263),
    .A2(_1758_),
    .Y(_1833_),
    .B1(_1832_));
 sg13g2_nand2_1 _7129_ (.Y(_1834_),
    .A(_0996_),
    .B(_1833_));
 sg13g2_nand3_1 _7130_ (.B(_1827_),
    .C(_1834_),
    .A(_1826_),
    .Y(_1835_));
 sg13g2_a21oi_1 _7131_ (.A1(net54),
    .A2(_1489_),
    .Y(_1836_),
    .B1(_1491_));
 sg13g2_nor3_1 _7132_ (.A(net219),
    .B(net227),
    .C(_4162_),
    .Y(_1837_));
 sg13g2_nor2_1 _7133_ (.A(net193),
    .B(net231),
    .Y(_1838_));
 sg13g2_nor3_1 _7134_ (.A(_1806_),
    .B(_1837_),
    .C(_1838_),
    .Y(_1840_));
 sg13g2_a21oi_1 _7135_ (.A1(_1806_),
    .A2(_1836_),
    .Y(_1841_),
    .B1(_1840_));
 sg13g2_nor2_1 _7136_ (.A(net227),
    .B(net171),
    .Y(_1842_));
 sg13g2_a22oi_1 _7137_ (.Y(_1843_),
    .B1(_1842_),
    .B2(_1818_),
    .A2(_1841_),
    .A1(net171));
 sg13g2_a21o_1 _7138_ (.A2(_1693_),
    .A1(net180),
    .B1(_0592_),
    .X(_1844_));
 sg13g2_a22oi_1 _7139_ (.Y(_1845_),
    .B1(_1844_),
    .B2(_1652_),
    .A2(_1707_),
    .A1(_1420_));
 sg13g2_nor2_1 _7140_ (.A(_1843_),
    .B(_1845_),
    .Y(_1846_));
 sg13g2_nand2_1 _7141_ (.Y(_1847_),
    .A(net20),
    .B(_1822_));
 sg13g2_a21oi_1 _7142_ (.A1(_4513_),
    .A2(net20),
    .Y(_1848_),
    .B1(net206));
 sg13g2_a221oi_1 _7143_ (.B2(net264),
    .C1(_1848_),
    .B1(_1847_),
    .A1(net23),
    .Y(_1849_),
    .A2(_1758_));
 sg13g2_o21ai_1 _7144_ (.B1(_1758_),
    .Y(_1850_),
    .A1(_4513_),
    .A2(net263));
 sg13g2_a21oi_1 _7145_ (.A1(_1819_),
    .A2(_1850_),
    .Y(_1851_),
    .B1(_1755_));
 sg13g2_a21oi_1 _7146_ (.A1(_1755_),
    .A2(_1849_),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_o21ai_1 _7147_ (.B1(_1852_),
    .Y(_1853_),
    .A1(_1835_),
    .A2(_1846_));
 sg13g2_o21ai_1 _7148_ (.B1(_1853_),
    .Y(_1854_),
    .A1(net246),
    .A2(_1824_));
 sg13g2_xor2_1 _7149_ (.B(_1821_),
    .A(net298),
    .X(_1855_));
 sg13g2_a22oi_1 _7150_ (.Y(_1856_),
    .B1(_1854_),
    .B2(_1855_),
    .A2(_1821_),
    .A1(_3881_));
 sg13g2_nand2_1 _7151_ (.Y(_1857_),
    .A(_1691_),
    .B(_1671_));
 sg13g2_nor3_1 _7152_ (.A(_1857_),
    .B(_1663_),
    .C(_1843_),
    .Y(_1858_));
 sg13g2_and4_1 _7153_ (.A(_1852_),
    .B(_1826_),
    .C(_1855_),
    .D(_1858_),
    .X(_1859_));
 sg13g2_nor3_1 _7154_ (.A(_1762_),
    .B(_1856_),
    .C(_1859_),
    .Y(_1861_));
 sg13g2_buf_1 _7155_ (.A(_1861_),
    .X(_1862_));
 sg13g2_a21oi_1 _7156_ (.A1(_1814_),
    .A2(_1816_),
    .Y(_1863_),
    .B1(_1862_));
 sg13g2_nand2_1 _7157_ (.Y(_1864_),
    .A(net206),
    .B(net179));
 sg13g2_a22oi_1 _7158_ (.Y(_1865_),
    .B1(_1694_),
    .B2(_0592_),
    .A2(_1707_),
    .A1(_3557_));
 sg13g2_nand2_1 _7159_ (.Y(_1866_),
    .A(net191),
    .B(net118));
 sg13g2_o21ai_1 _7160_ (.B1(_1866_),
    .Y(_1867_),
    .A1(_1865_),
    .A2(_1659_));
 sg13g2_nor2_1 _7161_ (.A(net206),
    .B(net179),
    .Y(_1868_));
 sg13g2_a21oi_1 _7162_ (.A1(_1864_),
    .A2(_1867_),
    .Y(_1869_),
    .B1(_1868_));
 sg13g2_inv_1 _7163_ (.Y(_1870_),
    .A(_1869_));
 sg13g2_a21oi_1 _7164_ (.A1(_4513_),
    .A2(_1869_),
    .Y(_1872_),
    .B1(net20));
 sg13g2_a21oi_1 _7165_ (.A1(net264),
    .A2(_1870_),
    .Y(_1873_),
    .B1(_1872_));
 sg13g2_nand2b_1 _7166_ (.Y(_1874_),
    .B(_1467_),
    .A_N(_1608_));
 sg13g2_o21ai_1 _7167_ (.B1(_1874_),
    .Y(_1875_),
    .A1(_1755_),
    .A2(_1873_));
 sg13g2_nand2_1 _7168_ (.Y(_1876_),
    .A(net180),
    .B(net34));
 sg13g2_o21ai_1 _7169_ (.B1(_1876_),
    .Y(_1877_),
    .A1(_4471_),
    .A2(net34));
 sg13g2_nand2b_1 _7170_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1857_));
 sg13g2_nand2_1 _7171_ (.Y(_1879_),
    .A(net224),
    .B(net242));
 sg13g2_nand3_1 _7172_ (.B(_1879_),
    .C(_1700_),
    .A(_1864_),
    .Y(_1880_));
 sg13g2_or4_1 _7173_ (.A(_1755_),
    .B(_1659_),
    .C(_1878_),
    .D(_1880_),
    .X(_1881_));
 sg13g2_nand3_1 _7174_ (.B(_1875_),
    .C(_1881_),
    .A(net192),
    .Y(_1883_));
 sg13g2_buf_1 _7175_ (.A(_1883_),
    .X(_1884_));
 sg13g2_o21ai_1 _7176_ (.B1(_1884_),
    .Y(_1885_),
    .A1(_1812_),
    .A2(_1863_));
 sg13g2_and2_1 _7177_ (.A(_1745_),
    .B(_1885_),
    .X(_1886_));
 sg13g2_inv_1 _7178_ (.Y(_1887_),
    .A(_1812_));
 sg13g2_nand3_1 _7179_ (.B(_1690_),
    .C(_1887_),
    .A(_1884_),
    .Y(_1888_));
 sg13g2_and2_1 _7180_ (.A(net34),
    .B(_1637_),
    .X(_1889_));
 sg13g2_buf_1 _7181_ (.A(_1889_),
    .X(_1890_));
 sg13g2_nor3_2 _7182_ (.A(net261),
    .B(net118),
    .C(_1890_),
    .Y(_1891_));
 sg13g2_xnor2_1 _7183_ (.Y(_1892_),
    .A(_1678_),
    .B(_1891_));
 sg13g2_nand2_1 _7184_ (.Y(_1893_),
    .A(net264),
    .B(_1892_));
 sg13g2_o21ai_1 _7185_ (.B1(net246),
    .Y(_1894_),
    .A1(net304),
    .A2(_1893_));
 sg13g2_nor2_2 _7186_ (.A(net118),
    .B(_1890_),
    .Y(_1895_));
 sg13g2_nand2_1 _7187_ (.Y(_1896_),
    .A(_1080_),
    .B(_1677_));
 sg13g2_o21ai_1 _7188_ (.B1(net184),
    .Y(_1897_),
    .A1(_1895_),
    .A2(_1896_));
 sg13g2_xnor2_1 _7189_ (.Y(_1898_),
    .A(_1607_),
    .B(_1897_));
 sg13g2_o21ai_1 _7190_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_4116_),
    .A2(_1893_));
 sg13g2_o21ai_1 _7191_ (.B1(_1899_),
    .Y(_1900_),
    .A1(_1894_),
    .A2(_1898_));
 sg13g2_o21ai_1 _7192_ (.B1(_1607_),
    .Y(_1901_),
    .A1(_1756_),
    .A2(_1891_));
 sg13g2_xor2_1 _7193_ (.B(_1901_),
    .A(_1483_),
    .X(_1902_));
 sg13g2_nand2_1 _7194_ (.Y(_1904_),
    .A(_0820_),
    .B(_1902_));
 sg13g2_nand2_1 _7195_ (.Y(_1905_),
    .A(_1364_),
    .B(_1901_));
 sg13g2_o21ai_1 _7196_ (.B1(_1905_),
    .Y(_1906_),
    .A1(_1900_),
    .A2(_1904_));
 sg13g2_nand2_1 _7197_ (.Y(_1907_),
    .A(_1630_),
    .B(_1890_));
 sg13g2_a21o_1 _7198_ (.A2(_1907_),
    .A1(net263),
    .B1(net215),
    .X(_1908_));
 sg13g2_o21ai_1 _7199_ (.B1(_1908_),
    .Y(_1909_),
    .A1(net263),
    .A2(_1895_));
 sg13g2_nand2b_1 _7200_ (.Y(_1910_),
    .B(_1907_),
    .A_N(_1895_));
 sg13g2_nand3_1 _7201_ (.B(_1630_),
    .C(_1890_),
    .A(_0441_),
    .Y(_1911_));
 sg13g2_o21ai_1 _7202_ (.B1(_1911_),
    .Y(_1912_),
    .A1(_0441_),
    .A2(_1910_));
 sg13g2_a22oi_1 _7203_ (.Y(_1913_),
    .B1(_1912_),
    .B2(net171),
    .A2(_1895_),
    .A1(_1842_));
 sg13g2_nor2_1 _7204_ (.A(net220),
    .B(_1496_),
    .Y(_1915_));
 sg13g2_nor2_1 _7205_ (.A(_1502_),
    .B(_1783_),
    .Y(_1916_));
 sg13g2_a22oi_1 _7206_ (.Y(_1917_),
    .B1(_1916_),
    .B2(_0458_),
    .A2(_1915_),
    .A1(_1783_));
 sg13g2_nor2_1 _7207_ (.A(_1913_),
    .B(_1917_),
    .Y(_1918_));
 sg13g2_nand2_1 _7208_ (.Y(_1919_),
    .A(net54),
    .B(_1915_));
 sg13g2_nand3_1 _7209_ (.B(net116),
    .C(_1496_),
    .A(_0458_),
    .Y(_1920_));
 sg13g2_a21oi_1 _7210_ (.A1(_1919_),
    .A2(_1920_),
    .Y(_1921_),
    .B1(_3482_));
 sg13g2_nor2_1 _7211_ (.A(net180),
    .B(_1423_),
    .Y(_1922_));
 sg13g2_nor2_1 _7212_ (.A(_0922_),
    .B(net118),
    .Y(_1923_));
 sg13g2_xnor2_1 _7213_ (.Y(_1924_),
    .A(net226),
    .B(_1923_));
 sg13g2_xnor2_1 _7214_ (.Y(_1926_),
    .A(_0922_),
    .B(_1910_));
 sg13g2_a21oi_1 _7215_ (.A1(_3731_),
    .A2(_1924_),
    .Y(_1927_),
    .B1(_1926_));
 sg13g2_o21ai_1 _7216_ (.B1(_1927_),
    .Y(_1928_),
    .A1(_1921_),
    .A2(_1922_));
 sg13g2_nand3_1 _7217_ (.B(_0996_),
    .C(_1895_),
    .A(net263),
    .Y(_1929_));
 sg13g2_nand4_1 _7218_ (.B(net226),
    .C(_1631_),
    .A(_1407_),
    .Y(_1930_),
    .D(_1890_));
 sg13g2_nand3_1 _7219_ (.B(_1929_),
    .C(_1930_),
    .A(_1928_),
    .Y(_1931_));
 sg13g2_a221oi_1 _7220_ (.B2(_1647_),
    .C1(_1931_),
    .B1(_1918_),
    .A1(net242),
    .Y(_1932_),
    .A2(_1909_));
 sg13g2_xor2_1 _7221_ (.B(_1891_),
    .A(_1700_),
    .X(_1933_));
 sg13g2_xnor2_1 _7222_ (.Y(_1934_),
    .A(_1755_),
    .B(_1897_));
 sg13g2_nor3_1 _7223_ (.A(_1904_),
    .B(_1933_),
    .C(_1934_),
    .Y(_1935_));
 sg13g2_nor2b_1 _7224_ (.A(_1932_),
    .B_N(_1935_),
    .Y(_1937_));
 sg13g2_nand3_1 _7225_ (.B(_1935_),
    .C(_1918_),
    .A(_1671_),
    .Y(_1938_));
 sg13g2_o21ai_1 _7226_ (.B1(_1938_),
    .Y(_1939_),
    .A1(_1906_),
    .A2(_1937_));
 sg13g2_nand2_1 _7227_ (.Y(_1940_),
    .A(net116),
    .B(_1816_));
 sg13g2_o21ai_1 _7228_ (.B1(net20),
    .Y(_1941_),
    .A1(net226),
    .A2(net117));
 sg13g2_a221oi_1 _7229_ (.B2(_1437_),
    .C1(_1848_),
    .B1(_1941_),
    .A1(_1678_),
    .Y(_1942_),
    .A2(net87));
 sg13g2_o21ai_1 _7230_ (.B1(_1631_),
    .Y(_1943_),
    .A1(_4513_),
    .A2(net263));
 sg13g2_nand3_1 _7231_ (.B(_1819_),
    .C(_1943_),
    .A(_1755_),
    .Y(_1944_));
 sg13g2_o21ai_1 _7232_ (.B1(_1944_),
    .Y(_1945_),
    .A1(_1755_),
    .A2(_1942_));
 sg13g2_nand3_1 _7233_ (.B(net117),
    .C(_1819_),
    .A(_1607_),
    .Y(_1946_));
 sg13g2_xor2_1 _7234_ (.B(_1946_),
    .A(_1483_),
    .X(_1948_));
 sg13g2_nand2_1 _7235_ (.Y(_1949_),
    .A(net287),
    .B(_1948_));
 sg13g2_nand2_1 _7236_ (.Y(_1950_),
    .A(_4252_),
    .B(_1677_));
 sg13g2_nand2_1 _7237_ (.Y(_1951_),
    .A(_1438_),
    .B(net87));
 sg13g2_nand3_1 _7238_ (.B(net267),
    .C(_1658_),
    .A(net215),
    .Y(_1952_));
 sg13g2_o21ai_1 _7239_ (.B1(_1952_),
    .Y(_1953_),
    .A1(net215),
    .A2(_1951_));
 sg13g2_nor3_1 _7240_ (.A(net224),
    .B(_1438_),
    .C(_1866_),
    .Y(_1954_));
 sg13g2_a21o_1 _7241_ (.A2(_1953_),
    .A1(net224),
    .B1(_1954_),
    .X(_1955_));
 sg13g2_nor4_1 _7242_ (.A(net224),
    .B(net191),
    .C(_4527_),
    .D(net87),
    .Y(_1956_));
 sg13g2_nand2_1 _7243_ (.Y(_1957_),
    .A(_4252_),
    .B(net20));
 sg13g2_a22oi_1 _7244_ (.Y(_1959_),
    .B1(_1956_),
    .B2(_1957_),
    .A2(_1955_),
    .A1(_1950_));
 sg13g2_nor3_1 _7245_ (.A(_1878_),
    .B(_1949_),
    .C(_1959_),
    .Y(_1960_));
 sg13g2_inv_1 _7246_ (.Y(_1961_),
    .A(_1949_));
 sg13g2_o21ai_1 _7247_ (.B1(_1819_),
    .Y(_1962_),
    .A1(net226),
    .A2(net117));
 sg13g2_xnor2_1 _7248_ (.Y(_1963_),
    .A(net35),
    .B(_1962_));
 sg13g2_o21ai_1 _7249_ (.B1(_1950_),
    .Y(_1964_),
    .A1(net200),
    .A2(net117));
 sg13g2_nand2_1 _7250_ (.Y(_1965_),
    .A(net200),
    .B(_1957_));
 sg13g2_a22oi_1 _7251_ (.Y(_1966_),
    .B1(_1965_),
    .B2(_1746_),
    .A2(_1964_),
    .A1(net224));
 sg13g2_o21ai_1 _7252_ (.B1(_1966_),
    .Y(_1967_),
    .A1(_1658_),
    .A2(_1950_));
 sg13g2_xnor2_1 _7253_ (.Y(_1968_),
    .A(net261),
    .B(_4527_));
 sg13g2_a21oi_1 _7254_ (.A1(_1204_),
    .A2(_1865_),
    .Y(_1970_),
    .B1(net87));
 sg13g2_nor3_1 _7255_ (.A(_1865_),
    .B(_1866_),
    .C(_1968_),
    .Y(_1971_));
 sg13g2_a21o_1 _7256_ (.A2(_1970_),
    .A1(_1968_),
    .B1(_1971_),
    .X(_1972_));
 sg13g2_o21ai_1 _7257_ (.B1(_1945_),
    .Y(_1973_),
    .A1(_1967_),
    .A2(_1972_));
 sg13g2_o21ai_1 _7258_ (.B1(_1973_),
    .Y(_1974_),
    .A1(net246),
    .A2(_1963_));
 sg13g2_a22oi_1 _7259_ (.Y(_1975_),
    .B1(_1961_),
    .B2(_1974_),
    .A2(_1946_),
    .A1(_1789_));
 sg13g2_a21o_1 _7260_ (.A2(_1960_),
    .A1(_1945_),
    .B1(_1975_),
    .X(_1976_));
 sg13g2_nand2_1 _7261_ (.Y(_1977_),
    .A(_1940_),
    .B(_1976_));
 sg13g2_a21oi_1 _7262_ (.A1(_1939_),
    .A2(_1977_),
    .Y(_1978_),
    .B1(_1862_));
 sg13g2_and2_1 _7263_ (.A(_1544_),
    .B(net152),
    .X(_1979_));
 sg13g2_buf_2 _7264_ (.A(_1979_),
    .X(_1980_));
 sg13g2_o21ai_1 _7265_ (.B1(_1980_),
    .Y(_1981_),
    .A1(_1888_),
    .A2(_1978_));
 sg13g2_o21ai_1 _7266_ (.B1(_1981_),
    .Y(_1982_),
    .A1(net119),
    .A2(_1886_));
 sg13g2_nand2_1 _7267_ (.Y(_1983_),
    .A(_1045_),
    .B(_1047_));
 sg13g2_nand3_1 _7268_ (.B(net256),
    .C(_0838_),
    .A(net253),
    .Y(_1984_));
 sg13g2_buf_1 _7269_ (.A(_1984_),
    .X(_1985_));
 sg13g2_buf_1 _7270_ (.A(_1985_),
    .X(_1986_));
 sg13g2_nand2_1 _7271_ (.Y(_1987_),
    .A(net183),
    .B(net136));
 sg13g2_a21oi_1 _7272_ (.A1(_1087_),
    .A2(_0839_),
    .Y(_1988_),
    .B1(_1987_));
 sg13g2_nand2_1 _7273_ (.Y(_1989_),
    .A(_1564_),
    .B(_0888_));
 sg13g2_buf_1 _7274_ (.A(_1989_),
    .X(_1991_));
 sg13g2_nand2b_1 _7275_ (.Y(_1992_),
    .B(_2228_),
    .A_N(net300));
 sg13g2_nand3_1 _7276_ (.B(net4),
    .C(_0898_),
    .A(_0883_),
    .Y(_1993_));
 sg13g2_o21ai_1 _7277_ (.B1(_1993_),
    .Y(_1994_),
    .A1(_2316_),
    .A2(_1992_));
 sg13g2_buf_1 _7278_ (.A(_1994_),
    .X(_1995_));
 sg13g2_nor2b_1 _7279_ (.A(net155),
    .B_N(_1995_),
    .Y(_1996_));
 sg13g2_buf_1 _7280_ (.A(_1996_),
    .X(_1997_));
 sg13g2_nand2_1 _7281_ (.Y(_1998_),
    .A(net115),
    .B(_1884_));
 sg13g2_a21o_1 _7282_ (.A2(net55),
    .A1(net85),
    .B1(_1998_),
    .X(_1999_));
 sg13g2_a21oi_1 _7283_ (.A1(_1983_),
    .A2(_1988_),
    .Y(_2000_),
    .B1(_1999_));
 sg13g2_nand2_1 _7284_ (.Y(_2002_),
    .A(_0896_),
    .B(_1592_));
 sg13g2_buf_1 _7285_ (.A(_2002_),
    .X(_2003_));
 sg13g2_buf_1 _7286_ (.A(net84),
    .X(_2004_));
 sg13g2_and2_1 _7287_ (.A(_0888_),
    .B(_0891_),
    .X(_2005_));
 sg13g2_buf_1 _7288_ (.A(_2005_),
    .X(_2006_));
 sg13g2_nor2_1 _7289_ (.A(net184),
    .B(_0840_),
    .Y(_2007_));
 sg13g2_nor2_1 _7290_ (.A(net258),
    .B(_2007_),
    .Y(_2008_));
 sg13g2_nor2_1 _7291_ (.A(net252),
    .B(_2008_),
    .Y(_2009_));
 sg13g2_buf_2 _7292_ (.A(_2009_),
    .X(_2010_));
 sg13g2_nor2_1 _7293_ (.A(net94),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_buf_2 _7294_ (.A(_2011_),
    .X(_2012_));
 sg13g2_nand2_1 _7295_ (.Y(_2013_),
    .A(_1544_),
    .B(_1564_));
 sg13g2_buf_1 _7296_ (.A(_2013_),
    .X(_2014_));
 sg13g2_a21oi_1 _7297_ (.A1(net260),
    .A2(_0227_),
    .Y(_2015_),
    .B1(net251));
 sg13g2_nand2b_1 _7298_ (.Y(_2016_),
    .B(_0711_),
    .A_N(_2015_));
 sg13g2_nand2_1 _7299_ (.Y(_2017_),
    .A(_1914_),
    .B(_2016_));
 sg13g2_a21oi_2 _7300_ (.B1(_0304_),
    .Y(_2018_),
    .A2(_2017_),
    .A1(_0359_));
 sg13g2_nor2_1 _7301_ (.A(_0590_),
    .B(_2018_),
    .Y(_2019_));
 sg13g2_buf_2 _7302_ (.A(_2019_),
    .X(_2020_));
 sg13g2_nand3_1 _7303_ (.B(_4136_),
    .C(net86),
    .A(_1533_),
    .Y(_2021_));
 sg13g2_o21ai_1 _7304_ (.B1(_2021_),
    .Y(_2023_),
    .A1(net114),
    .A2(_2020_));
 sg13g2_a221oi_1 _7305_ (.B2(_1576_),
    .C1(_2023_),
    .B1(_2012_),
    .A1(_2006_),
    .Y(_2024_),
    .A2(_1573_));
 sg13g2_a21oi_1 _7306_ (.A1(_0843_),
    .A2(_0874_),
    .Y(_2025_),
    .B1(_1002_));
 sg13g2_a21o_1 _7307_ (.A2(_4093_),
    .A1(_4168_),
    .B1(_2025_),
    .X(_2026_));
 sg13g2_buf_1 _7308_ (.A(_2026_),
    .X(_2027_));
 sg13g2_nand2_1 _7309_ (.Y(_2028_),
    .A(_0834_),
    .B(net151));
 sg13g2_buf_2 _7310_ (.A(_2028_),
    .X(_2029_));
 sg13g2_nand3_1 _7311_ (.B(net1),
    .C(net2),
    .A(net300),
    .Y(_2030_));
 sg13g2_o21ai_1 _7312_ (.B1(_2030_),
    .Y(_2031_),
    .A1(_2840_),
    .A2(_1541_));
 sg13g2_buf_1 _7313_ (.A(_2031_),
    .X(_2032_));
 sg13g2_nand2_1 _7314_ (.Y(_2034_),
    .A(net152),
    .B(net150));
 sg13g2_buf_2 _7315_ (.A(_2034_),
    .X(_2035_));
 sg13g2_nor2_2 _7316_ (.A(_1538_),
    .B(_2035_),
    .Y(_2036_));
 sg13g2_nand2_1 _7317_ (.Y(_2037_),
    .A(_2029_),
    .B(_2036_));
 sg13g2_o21ai_1 _7318_ (.B1(_2037_),
    .Y(_2038_),
    .A1(_2004_),
    .A2(_2024_));
 sg13g2_nor2_1 _7319_ (.A(net145),
    .B(_4305_),
    .Y(_2039_));
 sg13g2_inv_1 _7320_ (.Y(_2040_),
    .A(_2039_));
 sg13g2_nor3_1 _7321_ (.A(net238),
    .B(net139),
    .C(_4442_),
    .Y(_2041_));
 sg13g2_nor2_1 _7322_ (.A(_4321_),
    .B(_2041_),
    .Y(_2042_));
 sg13g2_o21ai_1 _7323_ (.B1(net141),
    .Y(_2043_),
    .A1(_2040_),
    .A2(_2042_));
 sg13g2_buf_1 _7324_ (.A(net143),
    .X(_2045_));
 sg13g2_nand2_1 _7325_ (.Y(_2046_),
    .A(_2045_),
    .B(net125));
 sg13g2_buf_1 _7326_ (.A(_4224_),
    .X(_2047_));
 sg13g2_buf_1 _7327_ (.A(net64),
    .X(_2048_));
 sg13g2_a21oi_1 _7328_ (.A1(net211),
    .A2(net50),
    .Y(_2049_),
    .B1(net32));
 sg13g2_nor2_1 _7329_ (.A(_2046_),
    .B(_2049_),
    .Y(_2050_));
 sg13g2_xnor2_1 _7330_ (.Y(_2051_),
    .A(net124),
    .B(_2050_));
 sg13g2_nor2_1 _7331_ (.A(net145),
    .B(_2051_),
    .Y(_2052_));
 sg13g2_nand3_1 _7332_ (.B(_4222_),
    .C(_4394_),
    .A(net89),
    .Y(_2053_));
 sg13g2_nand3_1 _7333_ (.B(_0608_),
    .C(net137),
    .A(net271),
    .Y(_2054_));
 sg13g2_nand2_1 _7334_ (.Y(_2056_),
    .A(_2053_),
    .B(_2054_));
 sg13g2_a21oi_1 _7335_ (.A1(_1468_),
    .A2(_2056_),
    .Y(_2057_),
    .B1(net32));
 sg13g2_nor2_1 _7336_ (.A(net101),
    .B(_2057_),
    .Y(_2058_));
 sg13g2_xnor2_1 _7337_ (.Y(_2059_),
    .A(_4248_),
    .B(_2058_));
 sg13g2_buf_1 _7338_ (.A(net102),
    .X(_2060_));
 sg13g2_o21ai_1 _7339_ (.B1(net211),
    .Y(_2061_),
    .A1(net235),
    .A2(_2060_));
 sg13g2_nand3_1 _7340_ (.B(net211),
    .C(_2060_),
    .A(net235),
    .Y(_2062_));
 sg13g2_o21ai_1 _7341_ (.B1(_2062_),
    .Y(_2063_),
    .A1(net211),
    .A2(net49));
 sg13g2_a21o_1 _7342_ (.A2(_2061_),
    .A1(net195),
    .B1(_2063_),
    .X(_2064_));
 sg13g2_nor2_1 _7343_ (.A(_4425_),
    .B(_2064_),
    .Y(_2065_));
 sg13g2_nand3_1 _7344_ (.B(net32),
    .C(_2056_),
    .A(_1479_),
    .Y(_2066_));
 sg13g2_nand2b_1 _7345_ (.Y(_2067_),
    .B(_2066_),
    .A_N(_2057_));
 sg13g2_a21oi_1 _7346_ (.A1(_4425_),
    .A2(_2064_),
    .Y(_2068_),
    .B1(_2067_));
 sg13g2_o21ai_1 _7347_ (.B1(net139),
    .Y(_2069_),
    .A1(_2065_),
    .A2(_2068_));
 sg13g2_xnor2_1 _7348_ (.Y(_2070_),
    .A(_2045_),
    .B(_2049_));
 sg13g2_nor3_1 _7349_ (.A(_4432_),
    .B(_2065_),
    .C(_2068_),
    .Y(_2071_));
 sg13g2_a21oi_1 _7350_ (.A1(_2069_),
    .A2(_2070_),
    .Y(_2072_),
    .B1(_2071_));
 sg13g2_a21o_1 _7351_ (.A2(_2072_),
    .A1(_2059_),
    .B1(_4473_),
    .X(_2073_));
 sg13g2_o21ai_1 _7352_ (.B1(_2073_),
    .Y(_2074_),
    .A1(_2059_),
    .A2(_2072_));
 sg13g2_nand2_1 _7353_ (.Y(_2075_),
    .A(net145),
    .B(_2051_));
 sg13g2_o21ai_1 _7354_ (.B1(_2075_),
    .Y(_2077_),
    .A1(_2052_),
    .A2(_2074_));
 sg13g2_o21ai_1 _7355_ (.B1(net124),
    .Y(_2078_),
    .A1(_2046_),
    .A2(_2057_));
 sg13g2_xnor2_1 _7356_ (.Y(_2079_),
    .A(_4108_),
    .B(_2078_));
 sg13g2_nor2_1 _7357_ (.A(net129),
    .B(_2079_),
    .Y(_2080_));
 sg13g2_nand2_1 _7358_ (.Y(_2081_),
    .A(net129),
    .B(_2079_));
 sg13g2_o21ai_1 _7359_ (.B1(_2081_),
    .Y(_2082_),
    .A1(_2077_),
    .A2(_2080_));
 sg13g2_nand2_1 _7360_ (.Y(_2083_),
    .A(_4329_),
    .B(_2082_));
 sg13g2_o21ai_1 _7361_ (.B1(_2083_),
    .Y(_2084_),
    .A1(_4131_),
    .A2(_2043_));
 sg13g2_nor2_1 _7362_ (.A(net245),
    .B(_4113_),
    .Y(_2085_));
 sg13g2_or2_1 _7363_ (.X(_2086_),
    .B(_2085_),
    .A(_4125_));
 sg13g2_a22oi_1 _7364_ (.Y(_2088_),
    .B1(_2086_),
    .B2(net225),
    .A2(_4255_),
    .A1(net281));
 sg13g2_o21ai_1 _7365_ (.B1(_1171_),
    .Y(_2089_),
    .A1(net286),
    .A2(_2088_));
 sg13g2_o21ai_1 _7366_ (.B1(net138),
    .Y(_2090_),
    .A1(net194),
    .A2(_4432_));
 sg13g2_a21oi_1 _7367_ (.A1(_2039_),
    .A2(_2090_),
    .Y(_2091_),
    .B1(_4267_));
 sg13g2_xnor2_1 _7368_ (.Y(_2092_),
    .A(_2089_),
    .B(_2091_));
 sg13g2_xnor2_1 _7369_ (.Y(_2093_),
    .A(_4131_),
    .B(_2043_));
 sg13g2_nand2_1 _7370_ (.Y(_2094_),
    .A(_2039_),
    .B(_2090_));
 sg13g2_xnor2_1 _7371_ (.Y(_2095_),
    .A(_4275_),
    .B(_2094_));
 sg13g2_nor2_1 _7372_ (.A(_4192_),
    .B(_2042_),
    .Y(_2096_));
 sg13g2_xnor2_1 _7373_ (.Y(_2097_),
    .A(_4305_),
    .B(_2096_));
 sg13g2_buf_1 _7374_ (.A(_0202_),
    .X(_2099_));
 sg13g2_xnor2_1 _7375_ (.Y(_2100_),
    .A(_4473_),
    .B(_2041_));
 sg13g2_o21ai_1 _7376_ (.B1(_4110_),
    .Y(_2101_),
    .A1(net239),
    .A2(net139));
 sg13g2_nor3_1 _7377_ (.A(_0230_),
    .B(net194),
    .C(_4437_),
    .Y(_2102_));
 sg13g2_a221oi_1 _7378_ (.B2(net185),
    .C1(_2102_),
    .B1(_2101_),
    .A1(net194),
    .Y(_2103_),
    .A2(_4437_));
 sg13g2_a21oi_1 _7379_ (.A1(_2099_),
    .A2(_2100_),
    .Y(_2104_),
    .B1(_2103_));
 sg13g2_nor2_1 _7380_ (.A(_2099_),
    .B(_2100_),
    .Y(_2105_));
 sg13g2_nor3_1 _7381_ (.A(_2047_),
    .B(_2104_),
    .C(_2105_),
    .Y(_2106_));
 sg13g2_xnor2_1 _7382_ (.Y(_2107_),
    .A(_4264_),
    .B(_2090_));
 sg13g2_o21ai_1 _7383_ (.B1(_2047_),
    .Y(_2108_),
    .A1(_2104_),
    .A2(_2105_));
 sg13g2_o21ai_1 _7384_ (.B1(_2108_),
    .Y(_2110_),
    .A1(_2106_),
    .A2(_2107_));
 sg13g2_o21ai_1 _7385_ (.B1(_2048_),
    .Y(_2111_),
    .A1(_2097_),
    .A2(_2110_));
 sg13g2_nand2_1 _7386_ (.Y(_2112_),
    .A(_2097_),
    .B(_2110_));
 sg13g2_a22oi_1 _7387_ (.Y(_2113_),
    .B1(_2111_),
    .B2(_2112_),
    .A2(_2095_),
    .A1(_4246_));
 sg13g2_nor2_1 _7388_ (.A(_4246_),
    .B(_2095_),
    .Y(_2114_));
 sg13g2_or2_1 _7389_ (.X(_2115_),
    .B(_2114_),
    .A(_2113_));
 sg13g2_nand2_1 _7390_ (.Y(_2116_),
    .A(_2093_),
    .B(_2115_));
 sg13g2_o21ai_1 _7391_ (.B1(_4248_),
    .Y(_2117_),
    .A1(_2093_),
    .A2(_2115_));
 sg13g2_a22oi_1 _7392_ (.Y(_2118_),
    .B1(_2116_),
    .B2(_2117_),
    .A2(_2092_),
    .A1(_4280_));
 sg13g2_nor2_1 _7393_ (.A(_4280_),
    .B(_2092_),
    .Y(_2119_));
 sg13g2_nor2_1 _7394_ (.A(_2118_),
    .B(_2119_),
    .Y(_2120_));
 sg13g2_nor2_1 _7395_ (.A(net128),
    .B(_2120_),
    .Y(_2121_));
 sg13g2_nand2_1 _7396_ (.Y(_2122_),
    .A(_4146_),
    .B(net124));
 sg13g2_nor2_1 _7397_ (.A(_2050_),
    .B(_2122_),
    .Y(_2123_));
 sg13g2_nor4_1 _7398_ (.A(_2084_),
    .B(_2089_),
    .C(_2121_),
    .D(_2123_),
    .Y(_2124_));
 sg13g2_nor2_1 _7399_ (.A(_4206_),
    .B(net127),
    .Y(_2125_));
 sg13g2_a21oi_1 _7400_ (.A1(_2048_),
    .A2(_2125_),
    .Y(_2126_),
    .B1(_2122_));
 sg13g2_nand2_2 _7401_ (.Y(_2127_),
    .A(_1531_),
    .B(_0888_));
 sg13g2_a21oi_1 _7402_ (.A1(_4321_),
    .A2(_2039_),
    .Y(_2128_),
    .B1(_4267_));
 sg13g2_or4_1 _7403_ (.A(_2127_),
    .B(net84),
    .C(_2089_),
    .D(_2128_),
    .X(_2129_));
 sg13g2_nor3_2 _7404_ (.A(_2124_),
    .B(_2126_),
    .C(_2129_),
    .Y(_2131_));
 sg13g2_nor3_1 _7405_ (.A(_2000_),
    .B(_2038_),
    .C(_2131_),
    .Y(_2132_));
 sg13g2_a21oi_1 _7406_ (.A1(_1697_),
    .A2(_1752_),
    .Y(_2133_),
    .B1(_4229_));
 sg13g2_o21ai_1 _7407_ (.B1(_0828_),
    .Y(_2134_),
    .A1(_0870_),
    .A2(_2133_));
 sg13g2_and2_1 _7408_ (.A(net188),
    .B(_2134_),
    .X(_2135_));
 sg13g2_buf_2 _7409_ (.A(_2135_),
    .X(_2136_));
 sg13g2_nor2_1 _7410_ (.A(_1002_),
    .B(_1000_),
    .Y(_2137_));
 sg13g2_a22oi_1 _7411_ (.Y(_2138_),
    .B1(_1000_),
    .B2(_4393_),
    .A2(_0869_),
    .A1(_0128_));
 sg13g2_nor2_1 _7412_ (.A(_0689_),
    .B(_2138_),
    .Y(_2139_));
 sg13g2_nor3_1 _7413_ (.A(_0128_),
    .B(net170),
    .C(net254),
    .Y(_2140_));
 sg13g2_nor2_1 _7414_ (.A(net219),
    .B(_0838_),
    .Y(_2142_));
 sg13g2_o21ai_1 _7415_ (.B1(_2142_),
    .Y(_2143_),
    .A1(net255),
    .A2(_2140_));
 sg13g2_a21o_1 _7416_ (.A2(_2143_),
    .A1(net292),
    .B1(_0392_),
    .X(_2144_));
 sg13g2_buf_1 _7417_ (.A(_2144_),
    .X(_2145_));
 sg13g2_o21ai_1 _7418_ (.B1(net81),
    .Y(_2146_),
    .A1(_2137_),
    .A2(_2139_));
 sg13g2_buf_1 _7419_ (.A(_2146_),
    .X(_2147_));
 sg13g2_nor2_1 _7420_ (.A(net88),
    .B(_0893_),
    .Y(_2148_));
 sg13g2_o21ai_1 _7421_ (.B1(_2148_),
    .Y(_2149_),
    .A1(_2136_),
    .A2(net31));
 sg13g2_nand2_1 _7422_ (.Y(_2150_),
    .A(net93),
    .B(_1551_));
 sg13g2_buf_1 _7423_ (.A(_2150_),
    .X(_2151_));
 sg13g2_nand2_1 _7424_ (.Y(_2153_),
    .A(_2272_),
    .B(_0884_));
 sg13g2_o21ai_1 _7425_ (.B1(_2153_),
    .Y(_2154_),
    .A1(_2972_),
    .A2(_0882_));
 sg13g2_buf_2 _7426_ (.A(_2154_),
    .X(_2155_));
 sg13g2_nand2_1 _7427_ (.Y(_2156_),
    .A(_2155_),
    .B(net152));
 sg13g2_buf_1 _7428_ (.A(_2156_),
    .X(_2157_));
 sg13g2_nor2_1 _7429_ (.A(_1538_),
    .B(net80),
    .Y(_2158_));
 sg13g2_nand2_1 _7430_ (.Y(_2159_),
    .A(_1564_),
    .B(net150));
 sg13g2_buf_2 _7431_ (.A(_2159_),
    .X(_2160_));
 sg13g2_nor2_1 _7432_ (.A(_2160_),
    .B(net57),
    .Y(_2161_));
 sg13g2_and2_1 _7433_ (.A(_0895_),
    .B(_1995_),
    .X(_2162_));
 sg13g2_buf_1 _7434_ (.A(_2162_),
    .X(_2164_));
 sg13g2_buf_1 _7435_ (.A(_2164_),
    .X(_2165_));
 sg13g2_buf_1 _7436_ (.A(net79),
    .X(_2166_));
 sg13g2_and2_1 _7437_ (.A(_0896_),
    .B(_1592_),
    .X(_2167_));
 sg13g2_buf_1 _7438_ (.A(_2167_),
    .X(_2168_));
 sg13g2_buf_1 _7439_ (.A(_2168_),
    .X(_2169_));
 sg13g2_a22oi_1 _7440_ (.Y(_2170_),
    .B1(_2145_),
    .B2(net47),
    .A2(_0834_),
    .A1(net115));
 sg13g2_nor2_1 _7441_ (.A(net88),
    .B(_2035_),
    .Y(_2171_));
 sg13g2_buf_2 _7442_ (.A(_2171_),
    .X(_2172_));
 sg13g2_nor3_2 _7443_ (.A(net114),
    .B(_1538_),
    .C(_0852_),
    .Y(_2173_));
 sg13g2_o21ai_1 _7444_ (.B1(net183),
    .Y(_2174_),
    .A1(_2172_),
    .A2(_2173_));
 sg13g2_o21ai_1 _7445_ (.B1(_2174_),
    .Y(_2175_),
    .A1(net119),
    .A2(_2170_));
 sg13g2_a221oi_1 _7446_ (.B2(net48),
    .C1(_2175_),
    .B1(_2161_),
    .A1(net30),
    .Y(_2176_),
    .A2(_2158_));
 sg13g2_nand2_1 _7447_ (.Y(_2177_),
    .A(net246),
    .B(_1073_));
 sg13g2_a21oi_1 _7448_ (.A1(net180),
    .A2(_0596_),
    .Y(_2178_),
    .B1(net215));
 sg13g2_nor2_1 _7449_ (.A(_1193_),
    .B(_2178_),
    .Y(_2179_));
 sg13g2_o21ai_1 _7450_ (.B1(_4116_),
    .Y(_2180_),
    .A1(_2177_),
    .A2(_2179_));
 sg13g2_nor2_1 _7451_ (.A(_0963_),
    .B(net280),
    .Y(_2181_));
 sg13g2_nand3_1 _7452_ (.B(_1147_),
    .C(_2181_),
    .A(_3406_),
    .Y(_2182_));
 sg13g2_or2_1 _7453_ (.X(_2183_),
    .B(_2182_),
    .A(_2177_));
 sg13g2_a21oi_1 _7454_ (.A1(_2180_),
    .A2(_2183_),
    .Y(_2185_),
    .B1(_3870_));
 sg13g2_nor2_1 _7455_ (.A(net229),
    .B(_2185_),
    .Y(_2186_));
 sg13g2_and2_1 _7456_ (.A(_1564_),
    .B(net150),
    .X(_2187_));
 sg13g2_buf_2 _7457_ (.A(_2187_),
    .X(_2188_));
 sg13g2_nand2_1 _7458_ (.Y(_2189_),
    .A(net52),
    .B(_2188_));
 sg13g2_inv_1 _7459_ (.Y(_2190_),
    .A(_2189_));
 sg13g2_nand2b_1 _7460_ (.Y(_2191_),
    .B(_1995_),
    .A_N(net155));
 sg13g2_buf_1 _7461_ (.A(_2191_),
    .X(_2192_));
 sg13g2_nand2_1 _7462_ (.Y(_2193_),
    .A(_1564_),
    .B(_2155_));
 sg13g2_buf_2 _7463_ (.A(_2193_),
    .X(_2194_));
 sg13g2_nor2_1 _7464_ (.A(net112),
    .B(_2194_),
    .Y(_2196_));
 sg13g2_nor3_1 _7465_ (.A(net206),
    .B(net189),
    .C(_0829_),
    .Y(_2197_));
 sg13g2_a21oi_1 _7466_ (.A1(_2197_),
    .A2(_1797_),
    .Y(_2198_),
    .B1(_1480_));
 sg13g2_nand2b_1 _7467_ (.Y(_2199_),
    .B(net292),
    .A_N(net222));
 sg13g2_nor3_1 _7468_ (.A(net256),
    .B(_0502_),
    .C(_2199_),
    .Y(_2200_));
 sg13g2_nor2_1 _7469_ (.A(_4221_),
    .B(_0991_),
    .Y(_2201_));
 sg13g2_nor2b_1 _7470_ (.A(_1763_),
    .B_N(_2200_),
    .Y(_2202_));
 sg13g2_o21ai_1 _7471_ (.B1(net207),
    .Y(_2203_),
    .A1(_2201_),
    .A2(_2202_));
 sg13g2_o21ai_1 _7472_ (.B1(_2203_),
    .Y(_2204_),
    .A1(_0991_),
    .A2(_2200_));
 sg13g2_o21ai_1 _7473_ (.B1(_2204_),
    .Y(_2205_),
    .A1(_2020_),
    .A2(_2198_));
 sg13g2_nand2_1 _7474_ (.Y(_2207_),
    .A(net188),
    .B(_2134_));
 sg13g2_buf_2 _7475_ (.A(_2207_),
    .X(_2208_));
 sg13g2_nor2b_1 _7476_ (.A(_0084_),
    .B_N(net222),
    .Y(_2209_));
 sg13g2_nand3_1 _7477_ (.B(_2209_),
    .C(_0873_),
    .A(_0840_),
    .Y(_2210_));
 sg13g2_and3_1 _7478_ (.X(_2211_),
    .A(_4066_),
    .B(_1512_),
    .C(_1422_));
 sg13g2_nand3_1 _7479_ (.B(_4168_),
    .C(_2211_),
    .A(net222),
    .Y(_2212_));
 sg13g2_nand2b_1 _7480_ (.Y(_2213_),
    .B(_2212_),
    .A_N(net175));
 sg13g2_a21o_1 _7481_ (.A2(_2210_),
    .A1(_1001_),
    .B1(_2213_),
    .X(_2214_));
 sg13g2_buf_1 _7482_ (.A(_2214_),
    .X(_2215_));
 sg13g2_nand2_2 _7483_ (.Y(_2216_),
    .A(_2208_),
    .B(_2215_));
 sg13g2_and2_1 _7484_ (.A(_1531_),
    .B(_2155_),
    .X(_2218_));
 sg13g2_buf_1 _7485_ (.A(_2218_),
    .X(_2219_));
 sg13g2_nand2_1 _7486_ (.Y(_2220_),
    .A(_1600_),
    .B(_2219_));
 sg13g2_nor2_1 _7487_ (.A(net53),
    .B(net80),
    .Y(_2221_));
 sg13g2_nand2_1 _7488_ (.Y(_2222_),
    .A(_2155_),
    .B(_0891_));
 sg13g2_buf_1 _7489_ (.A(_2222_),
    .X(_2223_));
 sg13g2_nor2_1 _7490_ (.A(net112),
    .B(net78),
    .Y(_2224_));
 sg13g2_a22oi_1 _7491_ (.Y(_2225_),
    .B1(_2224_),
    .B2(_1573_),
    .A2(_2221_),
    .A1(_2012_));
 sg13g2_o21ai_1 _7492_ (.B1(_2225_),
    .Y(_2226_),
    .A1(_2216_),
    .A2(_2220_));
 sg13g2_a221oi_1 _7493_ (.B2(_2205_),
    .C1(_2226_),
    .B1(_2196_),
    .A1(_2186_),
    .Y(_2227_),
    .A2(_2190_));
 sg13g2_nand2_1 _7494_ (.Y(_2229_),
    .A(net155),
    .B(_1995_));
 sg13g2_buf_1 _7495_ (.A(_2229_),
    .X(_2230_));
 sg13g2_nand2_1 _7496_ (.Y(_2231_),
    .A(_1531_),
    .B(_2155_));
 sg13g2_buf_2 _7497_ (.A(_2231_),
    .X(_2232_));
 sg13g2_nor2_2 _7498_ (.A(_2230_),
    .B(_2232_),
    .Y(_2233_));
 sg13g2_buf_1 _7499_ (.A(net61),
    .X(_2234_));
 sg13g2_nand2_1 _7500_ (.Y(_2235_),
    .A(net37),
    .B(_1816_));
 sg13g2_nand2b_1 _7501_ (.Y(_2236_),
    .B(_2209_),
    .A_N(_4169_));
 sg13g2_nor2_1 _7502_ (.A(_1006_),
    .B(_0866_),
    .Y(_2237_));
 sg13g2_a221oi_1 _7503_ (.B2(_4065_),
    .C1(_0849_),
    .B1(_2237_),
    .A1(_1001_),
    .Y(_2238_),
    .A2(_2236_));
 sg13g2_buf_1 _7504_ (.A(_2238_),
    .X(_2240_));
 sg13g2_buf_1 _7505_ (.A(_2240_),
    .X(_2241_));
 sg13g2_a21oi_1 _7506_ (.A1(net29),
    .A2(_2235_),
    .Y(_2242_),
    .B1(net111));
 sg13g2_and2_1 _7507_ (.A(_2155_),
    .B(_0891_),
    .X(_2243_));
 sg13g2_buf_1 _7508_ (.A(_2243_),
    .X(_2244_));
 sg13g2_nand2_1 _7509_ (.Y(_2245_),
    .A(net47),
    .B(_2244_));
 sg13g2_buf_1 _7510_ (.A(_2245_),
    .X(_2246_));
 sg13g2_buf_1 _7511_ (.A(_2215_),
    .X(_2247_));
 sg13g2_buf_1 _7512_ (.A(net46),
    .X(_2248_));
 sg13g2_nand2_1 _7513_ (.Y(_2249_),
    .A(net255),
    .B(_1697_));
 sg13g2_nor3_1 _7514_ (.A(net233),
    .B(_2249_),
    .C(_1581_),
    .Y(_2251_));
 sg13g2_or2_1 _7515_ (.X(_2252_),
    .B(_2251_),
    .A(net272));
 sg13g2_nor4_1 _7516_ (.A(net292),
    .B(_0348_),
    .C(_0524_),
    .D(_2249_),
    .Y(_2253_));
 sg13g2_nand2b_1 _7517_ (.Y(_2254_),
    .B(_2253_),
    .A_N(_0866_));
 sg13g2_nand3_1 _7518_ (.B(_2252_),
    .C(_2254_),
    .A(_0839_),
    .Y(_2255_));
 sg13g2_and2_1 _7519_ (.A(net256),
    .B(_2255_),
    .X(_2256_));
 sg13g2_buf_2 _7520_ (.A(_2256_),
    .X(_2257_));
 sg13g2_nand2_2 _7521_ (.Y(_2258_),
    .A(_2020_),
    .B(_2208_));
 sg13g2_nand2_1 _7522_ (.Y(_2259_),
    .A(_2257_),
    .B(_2258_));
 sg13g2_nand2_1 _7523_ (.Y(_2260_),
    .A(net28),
    .B(_2259_));
 sg13g2_a21oi_1 _7524_ (.A1(net258),
    .A2(_0844_),
    .Y(_2262_),
    .B1(net221));
 sg13g2_a21oi_1 _7525_ (.A1(_4068_),
    .A2(_0845_),
    .Y(_2263_),
    .B1(net97));
 sg13g2_a21oi_1 _7526_ (.A1(_4168_),
    .A2(_4093_),
    .Y(_2264_),
    .B1(_2025_));
 sg13g2_buf_1 _7527_ (.A(_2264_),
    .X(_2265_));
 sg13g2_a21oi_1 _7528_ (.A1(_2262_),
    .A2(_2263_),
    .Y(_2266_),
    .B1(net149));
 sg13g2_nor2_2 _7529_ (.A(net112),
    .B(_2160_),
    .Y(_2267_));
 sg13g2_o21ai_1 _7530_ (.B1(_2267_),
    .Y(_2268_),
    .A1(net30),
    .A2(_2266_));
 sg13g2_o21ai_1 _7531_ (.B1(_2268_),
    .Y(_2269_),
    .A1(_2246_),
    .A2(_2260_));
 sg13g2_a21oi_1 _7532_ (.A1(_2233_),
    .A2(_2242_),
    .Y(_2270_),
    .B1(_2269_));
 sg13g2_nand4_1 _7533_ (.B(_2176_),
    .C(_2227_),
    .A(_2149_),
    .Y(_2271_),
    .D(_2270_));
 sg13g2_nand2_2 _7534_ (.Y(_2273_),
    .A(net81),
    .B(_2258_));
 sg13g2_nor2_1 _7535_ (.A(_2137_),
    .B(_2139_),
    .Y(_2274_));
 sg13g2_nand2_2 _7536_ (.Y(_2275_),
    .A(_0403_),
    .B(_2255_));
 sg13g2_nand2b_1 _7537_ (.Y(_2276_),
    .B(_2275_),
    .A_N(_2274_));
 sg13g2_buf_1 _7538_ (.A(_2276_),
    .X(_2277_));
 sg13g2_nand2b_1 _7539_ (.Y(_2278_),
    .B(_2277_),
    .A_N(_2273_));
 sg13g2_nand2_1 _7540_ (.Y(_2279_),
    .A(net46),
    .B(_2278_));
 sg13g2_nor3_1 _7541_ (.A(net51),
    .B(_2232_),
    .C(_2279_),
    .Y(_2280_));
 sg13g2_a21oi_1 _7542_ (.A1(net258),
    .A2(_2143_),
    .Y(_2281_),
    .B1(_0403_));
 sg13g2_buf_1 _7543_ (.A(_2281_),
    .X(_2282_));
 sg13g2_buf_1 _7544_ (.A(_2274_),
    .X(_2284_));
 sg13g2_nand2_1 _7545_ (.Y(_2285_),
    .A(net170),
    .B(_0859_));
 sg13g2_nand2_2 _7546_ (.Y(_2286_),
    .A(net185),
    .B(net195));
 sg13g2_o21ai_1 _7547_ (.B1(_2286_),
    .Y(_2287_),
    .A1(net135),
    .A2(_2285_));
 sg13g2_or2_1 _7548_ (.X(_2288_),
    .B(net135),
    .A(_2018_));
 sg13g2_nor2_2 _7549_ (.A(_0194_),
    .B(_0859_),
    .Y(_2289_));
 sg13g2_a22oi_1 _7550_ (.Y(_2290_),
    .B1(_2288_),
    .B2(_2289_),
    .A2(_2287_),
    .A1(_2275_));
 sg13g2_nor2_1 _7551_ (.A(net91),
    .B(_2160_),
    .Y(_2291_));
 sg13g2_o21ai_1 _7552_ (.B1(_2291_),
    .Y(_2292_),
    .A1(net77),
    .A2(_2290_));
 sg13g2_nand2_1 _7553_ (.Y(_2293_),
    .A(_1544_),
    .B(_1531_));
 sg13g2_buf_1 _7554_ (.A(_2293_),
    .X(_2295_));
 sg13g2_a21o_1 _7555_ (.A2(_2223_),
    .A1(net110),
    .B1(_2029_),
    .X(_2296_));
 sg13g2_o21ai_1 _7556_ (.B1(_2296_),
    .Y(_2297_),
    .A1(net119),
    .A2(_2257_));
 sg13g2_xor2_1 _7557_ (.B(_0858_),
    .A(net170),
    .X(_2298_));
 sg13g2_buf_1 _7558_ (.A(_2298_),
    .X(_2299_));
 sg13g2_buf_1 _7559_ (.A(net134),
    .X(_2300_));
 sg13g2_buf_1 _7560_ (.A(net109),
    .X(_2301_));
 sg13g2_buf_1 _7561_ (.A(net76),
    .X(_2302_));
 sg13g2_buf_1 _7562_ (.A(net45),
    .X(_2303_));
 sg13g2_o21ai_1 _7563_ (.B1(net256),
    .Y(_2304_),
    .A1(net292),
    .A2(_2007_));
 sg13g2_buf_1 _7564_ (.A(_2304_),
    .X(_2306_));
 sg13g2_nand2_1 _7565_ (.Y(_2307_),
    .A(net116),
    .B(net133));
 sg13g2_buf_2 _7566_ (.A(_2307_),
    .X(_2308_));
 sg13g2_nand2_1 _7567_ (.Y(_2309_),
    .A(net80),
    .B(net85));
 sg13g2_a22oi_1 _7568_ (.Y(_2310_),
    .B1(_2308_),
    .B2(_2309_),
    .A2(net133),
    .A1(net83));
 sg13g2_a21oi_1 _7569_ (.A1(net27),
    .A2(net94),
    .Y(_2311_),
    .B1(_2310_));
 sg13g2_o21ai_1 _7570_ (.B1(net48),
    .Y(_2312_),
    .A1(_2297_),
    .A2(_2311_));
 sg13g2_nor2_1 _7571_ (.A(_2230_),
    .B(_2127_),
    .Y(_2313_));
 sg13g2_nand2_1 _7572_ (.Y(_2314_),
    .A(net79),
    .B(_1980_));
 sg13g2_nor2_1 _7573_ (.A(_2277_),
    .B(_2314_),
    .Y(_2315_));
 sg13g2_o21ai_1 _7574_ (.B1(net81),
    .Y(_2317_),
    .A1(_2313_),
    .A2(_2315_));
 sg13g2_nand2_2 _7575_ (.Y(_2318_),
    .A(_1544_),
    .B(net152));
 sg13g2_nor2_1 _7576_ (.A(_2192_),
    .B(_2318_),
    .Y(_2319_));
 sg13g2_buf_2 _7577_ (.A(_2319_),
    .X(_2320_));
 sg13g2_nor2_1 _7578_ (.A(_1594_),
    .B(_1989_),
    .Y(_2321_));
 sg13g2_o21ai_1 _7579_ (.B1(_1940_),
    .Y(_2322_),
    .A1(_2320_),
    .A2(_2321_));
 sg13g2_buf_1 _7580_ (.A(_1027_),
    .X(_2323_));
 sg13g2_buf_1 _7581_ (.A(_2230_),
    .X(_2324_));
 sg13g2_nor2_2 _7582_ (.A(net74),
    .B(net90),
    .Y(_2325_));
 sg13g2_o21ai_1 _7583_ (.B1(_2325_),
    .Y(_2326_),
    .A1(net29),
    .A2(net75));
 sg13g2_buf_1 _7584_ (.A(net112),
    .X(_2328_));
 sg13g2_a21oi_1 _7585_ (.A1(net110),
    .A2(net80),
    .Y(_2329_),
    .B1(net73));
 sg13g2_nand2_1 _7586_ (.Y(_2330_),
    .A(net150),
    .B(_0891_));
 sg13g2_buf_1 _7587_ (.A(_2330_),
    .X(_2331_));
 sg13g2_nor3_1 _7588_ (.A(net53),
    .B(_2331_),
    .C(net153),
    .Y(_2332_));
 sg13g2_a21oi_1 _7589_ (.A1(_1552_),
    .A2(_2329_),
    .Y(_2333_),
    .B1(_2332_));
 sg13g2_a21oi_1 _7590_ (.A1(_0095_),
    .A2(_0841_),
    .Y(_2334_),
    .B1(net189));
 sg13g2_nor2_1 _7591_ (.A(net183),
    .B(_2334_),
    .Y(_2335_));
 sg13g2_o21ai_1 _7592_ (.B1(net272),
    .Y(_2336_),
    .A1(net186),
    .A2(net187));
 sg13g2_a21oi_2 _7593_ (.B1(_1480_),
    .Y(_2337_),
    .A2(_2336_),
    .A1(_2197_));
 sg13g2_and2_1 _7594_ (.A(_1544_),
    .B(_1564_),
    .X(_2339_));
 sg13g2_buf_1 _7595_ (.A(_2339_),
    .X(_2340_));
 sg13g2_nor2_1 _7596_ (.A(net222),
    .B(_0849_),
    .Y(_2341_));
 sg13g2_or3_1 _7597_ (.A(_1914_),
    .B(_0870_),
    .C(_0873_),
    .X(_2342_));
 sg13g2_nand3_1 _7598_ (.B(_4087_),
    .C(_0846_),
    .A(_1523_),
    .Y(_2343_));
 sg13g2_nand3_1 _7599_ (.B(_2342_),
    .C(_2343_),
    .A(_2341_),
    .Y(_2344_));
 sg13g2_and3_1 _7600_ (.X(_2345_),
    .A(_1599_),
    .B(_2340_),
    .C(_2344_));
 sg13g2_buf_1 _7601_ (.A(_2345_),
    .X(_2346_));
 sg13g2_o21ai_1 _7602_ (.B1(_2346_),
    .Y(_2347_),
    .A1(_2335_),
    .A2(_2337_));
 sg13g2_nand4_1 _7603_ (.B(_2326_),
    .C(_2333_),
    .A(_2322_),
    .Y(_2348_),
    .D(_2347_));
 sg13g2_and2_1 _7604_ (.A(net152),
    .B(net150),
    .X(_2350_));
 sg13g2_buf_1 _7605_ (.A(_2350_),
    .X(_2351_));
 sg13g2_nand2_2 _7606_ (.Y(_2352_),
    .A(_2351_),
    .B(_2164_));
 sg13g2_nor2_1 _7607_ (.A(_2352_),
    .B(net196),
    .Y(_2353_));
 sg13g2_nand2_1 _7608_ (.Y(_2354_),
    .A(_2168_),
    .B(_1980_));
 sg13g2_buf_2 _7609_ (.A(_2354_),
    .X(_2355_));
 sg13g2_a21oi_1 _7610_ (.A1(net169),
    .A2(net76),
    .Y(_2356_),
    .B1(_2355_));
 sg13g2_nor3_1 _7611_ (.A(net74),
    .B(_2331_),
    .C(_2010_),
    .Y(_2357_));
 sg13g2_nor3_1 _7612_ (.A(_2353_),
    .B(_2356_),
    .C(_2357_),
    .Y(_2358_));
 sg13g2_nor2_1 _7613_ (.A(net85),
    .B(_0903_),
    .Y(_2359_));
 sg13g2_nor2_2 _7614_ (.A(net88),
    .B(_1557_),
    .Y(_2361_));
 sg13g2_nor2_1 _7615_ (.A(net73),
    .B(_2232_),
    .Y(_2362_));
 sg13g2_a221oi_1 _7616_ (.B2(_2361_),
    .C1(_2362_),
    .B1(_2335_),
    .A1(_2359_),
    .Y(_2363_),
    .A2(net86));
 sg13g2_nand2_1 _7617_ (.Y(_2364_),
    .A(_0095_),
    .B(_1583_));
 sg13g2_nor2_1 _7618_ (.A(net189),
    .B(_0535_),
    .Y(_2365_));
 sg13g2_a21oi_2 _7619_ (.B1(_2130_),
    .Y(_2366_),
    .A2(_2365_),
    .A1(_2364_));
 sg13g2_nor2_1 _7620_ (.A(net88),
    .B(_2127_),
    .Y(_2367_));
 sg13g2_and2_1 _7621_ (.A(_1564_),
    .B(_2155_),
    .X(_2368_));
 sg13g2_buf_2 _7622_ (.A(_2368_),
    .X(_2369_));
 sg13g2_nand2_1 _7623_ (.Y(_2370_),
    .A(_2369_),
    .B(net79));
 sg13g2_a221oi_1 _7624_ (.B2(net134),
    .C1(_2370_),
    .B1(_0832_),
    .A1(net258),
    .Y(_2372_),
    .A2(net221));
 sg13g2_a22oi_1 _7625_ (.Y(_2373_),
    .B1(_2372_),
    .B2(net151),
    .A2(_2367_),
    .A1(_2366_));
 sg13g2_nand3_1 _7626_ (.B(_2363_),
    .C(_2373_),
    .A(_2358_),
    .Y(_2374_));
 sg13g2_nand2_1 _7627_ (.Y(_2375_),
    .A(_1531_),
    .B(_2032_));
 sg13g2_buf_2 _7628_ (.A(_2375_),
    .X(_2376_));
 sg13g2_a21oi_1 _7629_ (.A1(net73),
    .A2(net91),
    .Y(_2377_),
    .B1(_2376_));
 sg13g2_and2_1 _7630_ (.A(net150),
    .B(_0891_),
    .X(_2378_));
 sg13g2_buf_1 _7631_ (.A(_2378_),
    .X(_2379_));
 sg13g2_o21ai_1 _7632_ (.B1(_1526_),
    .Y(_2380_),
    .A1(net108),
    .A2(_1980_));
 sg13g2_o21ai_1 _7633_ (.B1(_2380_),
    .Y(_2381_),
    .A1(_2014_),
    .A2(_2324_));
 sg13g2_nor2_1 _7634_ (.A(net110),
    .B(net91),
    .Y(_2383_));
 sg13g2_a21oi_1 _7635_ (.A1(_2035_),
    .A2(net90),
    .Y(_2384_),
    .B1(_2328_));
 sg13g2_nor4_1 _7636_ (.A(_2377_),
    .B(_2381_),
    .C(_2383_),
    .D(_2384_),
    .Y(_2385_));
 sg13g2_nand2_2 _7637_ (.Y(_2386_),
    .A(_1571_),
    .B(_2169_));
 sg13g2_and2_1 _7638_ (.A(_1531_),
    .B(net150),
    .X(_2387_));
 sg13g2_buf_2 _7639_ (.A(_2387_),
    .X(_2388_));
 sg13g2_nand2_1 _7640_ (.Y(_2389_),
    .A(_1599_),
    .B(_2388_));
 sg13g2_buf_1 _7641_ (.A(_2389_),
    .X(_2390_));
 sg13g2_a21oi_1 _7642_ (.A1(_2386_),
    .A2(_2390_),
    .Y(_2391_),
    .B1(_1987_));
 sg13g2_o21ai_1 _7643_ (.B1(net183),
    .Y(_2392_),
    .A1(_1985_),
    .A2(net134));
 sg13g2_nor2_2 _7644_ (.A(net88),
    .B(net78),
    .Y(_2394_));
 sg13g2_nor2_2 _7645_ (.A(net85),
    .B(net84),
    .Y(_2395_));
 sg13g2_nor2_1 _7646_ (.A(_2394_),
    .B(_2395_),
    .Y(_2396_));
 sg13g2_nor2_1 _7647_ (.A(_2392_),
    .B(_2396_),
    .Y(_2397_));
 sg13g2_nand2_1 _7648_ (.Y(_2398_),
    .A(net115),
    .B(net108));
 sg13g2_nor2_1 _7649_ (.A(_2136_),
    .B(_2398_),
    .Y(_2399_));
 sg13g2_nor3_1 _7650_ (.A(net88),
    .B(_2194_),
    .C(net121),
    .Y(_2400_));
 sg13g2_nor4_1 _7651_ (.A(_2391_),
    .B(_2397_),
    .C(_2399_),
    .D(_2400_),
    .Y(_2401_));
 sg13g2_nor2_2 _7652_ (.A(net74),
    .B(_2376_),
    .Y(_2402_));
 sg13g2_nand2_1 _7653_ (.Y(_2403_),
    .A(net188),
    .B(net120));
 sg13g2_nand2_1 _7654_ (.Y(_2405_),
    .A(net151),
    .B(_2403_));
 sg13g2_nor2_2 _7655_ (.A(_1538_),
    .B(_2232_),
    .Y(_2406_));
 sg13g2_and2_1 _7656_ (.A(_2155_),
    .B(_1555_),
    .X(_2407_));
 sg13g2_buf_1 _7657_ (.A(_2407_),
    .X(_2408_));
 sg13g2_o21ai_1 _7658_ (.B1(net47),
    .Y(_2409_),
    .A1(_2408_),
    .A2(net150));
 sg13g2_nand2b_1 _7659_ (.Y(_2410_),
    .B(_2409_),
    .A_N(_2406_));
 sg13g2_a21oi_1 _7660_ (.A1(_1001_),
    .A2(_2210_),
    .Y(_2411_),
    .B1(_2213_));
 sg13g2_buf_1 _7661_ (.A(_2411_),
    .X(_2412_));
 sg13g2_nor2_2 _7662_ (.A(_2136_),
    .B(net72),
    .Y(_2413_));
 sg13g2_a22oi_1 _7663_ (.Y(_2414_),
    .B1(_2410_),
    .B2(_2413_),
    .A2(_2405_),
    .A1(_2402_));
 sg13g2_nand3_1 _7664_ (.B(_2401_),
    .C(_2414_),
    .A(_2385_),
    .Y(_2416_));
 sg13g2_nand2b_1 _7665_ (.Y(_2417_),
    .B(_0850_),
    .A_N(_0844_));
 sg13g2_buf_1 _7666_ (.A(_2417_),
    .X(_2418_));
 sg13g2_o21ai_1 _7667_ (.B1(net132),
    .Y(_2419_),
    .A1(_0832_),
    .A2(net149));
 sg13g2_buf_1 _7668_ (.A(_2419_),
    .X(_2420_));
 sg13g2_nand3_1 _7669_ (.B(net92),
    .C(_2420_),
    .A(_2369_),
    .Y(_2421_));
 sg13g2_nor2_2 _7670_ (.A(net112),
    .B(net114),
    .Y(_2422_));
 sg13g2_nand2_1 _7671_ (.Y(_2423_),
    .A(_2369_),
    .B(net47));
 sg13g2_a21oi_1 _7672_ (.A1(_2323_),
    .A2(_2308_),
    .Y(_2424_),
    .B1(_2423_));
 sg13g2_a21oi_1 _7673_ (.A1(_2422_),
    .A2(net133),
    .Y(_2425_),
    .B1(_2424_));
 sg13g2_a221oi_1 _7674_ (.B2(_0645_),
    .C1(net175),
    .B1(_1583_),
    .A1(_0535_),
    .Y(_2427_),
    .A2(_0847_));
 sg13g2_buf_1 _7675_ (.A(_2427_),
    .X(_2428_));
 sg13g2_nor2_1 _7676_ (.A(net24),
    .B(_2366_),
    .Y(_2429_));
 sg13g2_nand3_1 _7677_ (.B(_4393_),
    .C(_1422_),
    .A(net219),
    .Y(_2430_));
 sg13g2_a21oi_1 _7678_ (.A1(_2016_),
    .A2(_2430_),
    .Y(_2431_),
    .B1(_1925_));
 sg13g2_nor2b_1 _7679_ (.A(_2431_),
    .B_N(_2341_),
    .Y(_2432_));
 sg13g2_nor3_1 _7680_ (.A(_1538_),
    .B(net78),
    .C(_2432_),
    .Y(_2433_));
 sg13g2_buf_2 _7681_ (.A(_2433_),
    .X(_2434_));
 sg13g2_o21ai_1 _7682_ (.B1(_2434_),
    .Y(_2435_),
    .A1(_2428_),
    .A2(_2429_));
 sg13g2_nand3_1 _7683_ (.B(_2425_),
    .C(_2435_),
    .A(_2421_),
    .Y(_2436_));
 sg13g2_nor4_1 _7684_ (.A(_2348_),
    .B(_2374_),
    .C(_2416_),
    .D(_2436_),
    .Y(_2438_));
 sg13g2_nand4_1 _7685_ (.B(_2312_),
    .C(_2317_),
    .A(_2292_),
    .Y(_2439_),
    .D(_2438_));
 sg13g2_nor3_1 _7686_ (.A(_2271_),
    .B(_2280_),
    .C(_2439_),
    .Y(_2440_));
 sg13g2_nand2_2 _7687_ (.Y(_2441_),
    .A(net115),
    .B(_1533_));
 sg13g2_a22oi_1 _7688_ (.Y(_2442_),
    .B1(net204),
    .B2(net283),
    .A2(net236),
    .A1(_3503_));
 sg13g2_or2_1 _7689_ (.X(_2443_),
    .B(net309),
    .A(net237));
 sg13g2_buf_1 _7690_ (.A(_2443_),
    .X(_2444_));
 sg13g2_nand2_1 _7691_ (.Y(_2445_),
    .A(net236),
    .B(_2444_));
 sg13g2_o21ai_1 _7692_ (.B1(_2445_),
    .Y(_2446_),
    .A1(net199),
    .A2(_2442_));
 sg13g2_a21oi_1 _7693_ (.A1(_0908_),
    .A2(_2446_),
    .Y(_2447_),
    .B1(net243));
 sg13g2_o21ai_1 _7694_ (.B1(net243),
    .Y(_2449_),
    .A1(net247),
    .A2(_2446_));
 sg13g2_o21ai_1 _7695_ (.B1(_2449_),
    .Y(_2450_),
    .A1(net191),
    .A2(_2447_));
 sg13g2_nand2_1 _7696_ (.Y(_2451_),
    .A(_0919_),
    .B(_2450_));
 sg13g2_nor2_1 _7697_ (.A(net285),
    .B(_3870_),
    .Y(_2452_));
 sg13g2_or2_1 _7698_ (.X(_2453_),
    .B(_2450_),
    .A(net247));
 sg13g2_nor2_1 _7699_ (.A(net225),
    .B(_0842_),
    .Y(_2454_));
 sg13g2_a22oi_1 _7700_ (.Y(_2455_),
    .B1(_2453_),
    .B2(_2454_),
    .A2(_2452_),
    .A1(_2451_));
 sg13g2_xnor2_1 _7701_ (.Y(_2456_),
    .A(net281),
    .B(_2455_));
 sg13g2_buf_2 _7702_ (.A(_2456_),
    .X(_2457_));
 sg13g2_inv_1 _7703_ (.Y(_2458_),
    .A(_2457_));
 sg13g2_nand2_1 _7704_ (.Y(_2460_),
    .A(_3460_),
    .B(net244));
 sg13g2_nand3_1 _7705_ (.B(net236),
    .C(net282),
    .A(_0857_),
    .Y(_2461_));
 sg13g2_a21oi_1 _7706_ (.A1(_2460_),
    .A2(_2461_),
    .Y(_2462_),
    .B1(net199));
 sg13g2_a21oi_1 _7707_ (.A1(net204),
    .A2(net282),
    .Y(_2463_),
    .B1(net283));
 sg13g2_o21ai_1 _7708_ (.B1(_0996_),
    .Y(_2464_),
    .A1(net214),
    .A2(_2463_));
 sg13g2_or2_1 _7709_ (.X(_2465_),
    .B(_2464_),
    .A(_2462_));
 sg13g2_buf_1 _7710_ (.A(_2465_),
    .X(_2466_));
 sg13g2_xnor2_1 _7711_ (.Y(_2467_),
    .A(_1095_),
    .B(net247));
 sg13g2_xnor2_1 _7712_ (.Y(_2468_),
    .A(_2466_),
    .B(_2467_));
 sg13g2_buf_2 _7713_ (.A(_2468_),
    .X(_2469_));
 sg13g2_o21ai_1 _7714_ (.B1(_1717_),
    .Y(_2470_),
    .A1(net272),
    .A2(_2469_));
 sg13g2_xnor2_1 _7715_ (.Y(_2471_),
    .A(_4126_),
    .B(_2450_));
 sg13g2_buf_1 _7716_ (.A(_2471_),
    .X(_2472_));
 sg13g2_nor2_1 _7717_ (.A(_3644_),
    .B(_0985_),
    .Y(_2473_));
 sg13g2_nor2_1 _7718_ (.A(_2181_),
    .B(_2473_),
    .Y(_2474_));
 sg13g2_xnor2_1 _7719_ (.Y(_2475_),
    .A(_2446_),
    .B(_2474_));
 sg13g2_xnor2_1 _7720_ (.Y(_2476_),
    .A(net260),
    .B(net236));
 sg13g2_nor2b_1 _7721_ (.A(net204),
    .B_N(net275),
    .Y(_2477_));
 sg13g2_a21oi_1 _7722_ (.A1(_3677_),
    .A2(_2477_),
    .Y(_2478_),
    .B1(_1151_));
 sg13g2_and2_1 _7723_ (.A(_2476_),
    .B(_2478_),
    .X(_2479_));
 sg13g2_nand2b_1 _7724_ (.Y(_2481_),
    .B(net232),
    .A_N(_1144_));
 sg13g2_nor2_1 _7725_ (.A(net199),
    .B(_0395_),
    .Y(_2482_));
 sg13g2_a221oi_1 _7726_ (.B2(_2482_),
    .C1(_2476_),
    .B1(_2481_),
    .A1(_3805_),
    .Y(_2483_),
    .A2(_2477_));
 sg13g2_nand2b_1 _7727_ (.Y(_2484_),
    .B(net237),
    .A_N(net241));
 sg13g2_a21o_1 _7728_ (.A2(_2484_),
    .A1(_3525_),
    .B1(_1248_),
    .X(_2485_));
 sg13g2_nand3_1 _7729_ (.B(_3525_),
    .C(_2484_),
    .A(_1248_),
    .Y(_2486_));
 sg13g2_a21oi_1 _7730_ (.A1(_2485_),
    .A2(_2486_),
    .Y(_2487_),
    .B1(net265));
 sg13g2_nor3_1 _7731_ (.A(_2479_),
    .B(_2483_),
    .C(_2487_),
    .Y(_2488_));
 sg13g2_a21oi_1 _7732_ (.A1(net202),
    .A2(_1391_),
    .Y(_2489_),
    .B1(net204));
 sg13g2_mux2_1 _7733_ (.A0(_0937_),
    .A1(_2489_),
    .S(net236),
    .X(_2490_));
 sg13g2_xnor2_1 _7734_ (.Y(_2492_),
    .A(_3644_),
    .B(_2490_));
 sg13g2_xnor2_1 _7735_ (.Y(_2493_),
    .A(_1686_),
    .B(_2492_));
 sg13g2_o21ai_1 _7736_ (.B1(_2487_),
    .Y(_2494_),
    .A1(_2479_),
    .A2(_2483_));
 sg13g2_o21ai_1 _7737_ (.B1(_2494_),
    .Y(_2495_),
    .A1(_2488_),
    .A2(_2493_));
 sg13g2_xor2_1 _7738_ (.B(_2475_),
    .A(net297),
    .X(_2496_));
 sg13g2_nand2b_1 _7739_ (.Y(_2497_),
    .B(_2496_),
    .A_N(_2495_));
 sg13g2_nor2_1 _7740_ (.A(_4221_),
    .B(_2492_),
    .Y(_2498_));
 sg13g2_nor2b_1 _7741_ (.A(_2496_),
    .B_N(_2495_),
    .Y(_2499_));
 sg13g2_a21oi_1 _7742_ (.A1(_2497_),
    .A2(_2498_),
    .Y(_2500_),
    .B1(_2499_));
 sg13g2_a21oi_1 _7743_ (.A1(_0051_),
    .A2(_2475_),
    .Y(_2501_),
    .B1(_2500_));
 sg13g2_inv_1 _7744_ (.Y(_2503_),
    .A(_2501_));
 sg13g2_xnor2_1 _7745_ (.Y(_2504_),
    .A(_0145_),
    .B(_2469_));
 sg13g2_and3_1 _7746_ (.X(_2505_),
    .A(_0051_),
    .B(_2475_),
    .C(_2500_));
 sg13g2_buf_1 _7747_ (.A(_2505_),
    .X(_2506_));
 sg13g2_a21oi_1 _7748_ (.A1(_2503_),
    .A2(_2504_),
    .Y(_2507_),
    .B1(_2506_));
 sg13g2_buf_2 _7749_ (.A(_2507_),
    .X(_2508_));
 sg13g2_a21oi_1 _7750_ (.A1(_0875_),
    .A2(_2466_),
    .Y(_2509_),
    .B1(net247));
 sg13g2_o21ai_1 _7751_ (.B1(_0919_),
    .Y(_2510_),
    .A1(net285),
    .A2(_2466_));
 sg13g2_o21ai_1 _7752_ (.B1(_2510_),
    .Y(_2511_),
    .A1(_1193_),
    .A2(_2509_));
 sg13g2_buf_1 _7753_ (.A(_2511_),
    .X(_2512_));
 sg13g2_nor2_1 _7754_ (.A(_2452_),
    .B(_2454_),
    .Y(_2514_));
 sg13g2_xnor2_1 _7755_ (.Y(_2515_),
    .A(_2512_),
    .B(_2514_));
 sg13g2_inv_1 _7756_ (.Y(_2516_),
    .A(_2515_));
 sg13g2_a21oi_1 _7757_ (.A1(net44),
    .A2(_2508_),
    .Y(_2517_),
    .B1(_2516_));
 sg13g2_nand3_1 _7758_ (.B(_2516_),
    .C(_2508_),
    .A(net44),
    .Y(_2518_));
 sg13g2_o21ai_1 _7759_ (.B1(_2518_),
    .Y(_2519_),
    .A1(_0868_),
    .A2(_2517_));
 sg13g2_or2_1 _7760_ (.X(_2520_),
    .B(_2508_),
    .A(net44));
 sg13g2_nor3_1 _7761_ (.A(net272),
    .B(_1080_),
    .C(_2469_),
    .Y(_2521_));
 sg13g2_o21ai_1 _7762_ (.B1(_1001_),
    .Y(_2522_),
    .A1(_2516_),
    .A2(_2521_));
 sg13g2_nand2_1 _7763_ (.Y(_2523_),
    .A(_2516_),
    .B(_2521_));
 sg13g2_nand2_1 _7764_ (.Y(_2525_),
    .A(_2522_),
    .B(_2523_));
 sg13g2_a22oi_1 _7765_ (.Y(_2526_),
    .B1(_2520_),
    .B2(_2525_),
    .A2(_2519_),
    .A1(_2470_));
 sg13g2_buf_1 _7766_ (.A(_2526_),
    .X(_2527_));
 sg13g2_buf_1 _7767_ (.A(_4066_),
    .X(_2528_));
 sg13g2_a21oi_1 _7768_ (.A1(net285),
    .A2(_2512_),
    .Y(_2529_),
    .B1(net218));
 sg13g2_or2_1 _7769_ (.X(_2530_),
    .B(_2512_),
    .A(net285));
 sg13g2_nor2_1 _7770_ (.A(_3870_),
    .B(_1149_),
    .Y(_2531_));
 sg13g2_a22oi_1 _7771_ (.Y(_2532_),
    .B1(_2530_),
    .B2(_2531_),
    .A2(_2529_),
    .A1(_3870_));
 sg13g2_xnor2_1 _7772_ (.Y(_2533_),
    .A(net262),
    .B(_2532_));
 sg13g2_a21oi_1 _7773_ (.A1(_2527_),
    .A2(_2533_),
    .Y(_2534_),
    .B1(net305));
 sg13g2_nor3_1 _7774_ (.A(net44),
    .B(_2508_),
    .C(_2470_),
    .Y(_2536_));
 sg13g2_nand3_1 _7775_ (.B(_2515_),
    .C(_2536_),
    .A(_0868_),
    .Y(_2537_));
 sg13g2_buf_1 _7776_ (.A(_2537_),
    .X(_2538_));
 sg13g2_nand2_1 _7777_ (.Y(_2539_),
    .A(_0568_),
    .B(_2538_));
 sg13g2_a21oi_1 _7778_ (.A1(net305),
    .A2(_2533_),
    .Y(_2540_),
    .B1(_2539_));
 sg13g2_or2_1 _7779_ (.X(_2541_),
    .B(_2540_),
    .A(_2534_));
 sg13g2_nand3_1 _7780_ (.B(_2457_),
    .C(_2538_),
    .A(_0315_),
    .Y(_2542_));
 sg13g2_a21oi_1 _7781_ (.A1(_2527_),
    .A2(_2542_),
    .Y(_2543_),
    .B1(_2533_));
 sg13g2_a21oi_1 _7782_ (.A1(_2458_),
    .A2(_2541_),
    .Y(_2544_),
    .B1(_2543_));
 sg13g2_a21o_1 _7783_ (.A2(_2512_),
    .A1(net262),
    .B1(net229),
    .X(_2545_));
 sg13g2_a22oi_1 _7784_ (.Y(_2547_),
    .B1(_2453_),
    .B2(_0808_),
    .A2(_2528_),
    .A1(net248));
 sg13g2_nor2_1 _7785_ (.A(_1467_),
    .B(_2547_),
    .Y(_2548_));
 sg13g2_a221oi_1 _7786_ (.B2(net248),
    .C1(_2548_),
    .B1(_2545_),
    .A1(_2528_),
    .Y(_2549_),
    .A2(_2529_));
 sg13g2_xor2_1 _7787_ (.B(_2549_),
    .A(_2544_),
    .X(_2550_));
 sg13g2_nor2_1 _7788_ (.A(net305),
    .B(_2457_),
    .Y(_2551_));
 sg13g2_a22oi_1 _7789_ (.Y(_2552_),
    .B1(_2551_),
    .B2(_2527_),
    .A2(_2538_),
    .A1(_2457_));
 sg13g2_inv_1 _7790_ (.Y(_2553_),
    .A(_2552_));
 sg13g2_a21oi_1 _7791_ (.A1(net253),
    .A2(_2538_),
    .Y(_2554_),
    .B1(_4074_));
 sg13g2_o21ai_1 _7792_ (.B1(_2527_),
    .Y(_2555_),
    .A1(_2457_),
    .A2(_2554_));
 sg13g2_nand2_1 _7793_ (.Y(_2556_),
    .A(_2538_),
    .B(_2551_));
 sg13g2_a22oi_1 _7794_ (.Y(_2558_),
    .B1(_2555_),
    .B2(_2556_),
    .A2(_2553_),
    .A1(net258));
 sg13g2_xnor2_1 _7795_ (.Y(_2559_),
    .A(_2533_),
    .B(_2558_));
 sg13g2_nor2_1 _7796_ (.A(_2550_),
    .B(_2559_),
    .Y(_2560_));
 sg13g2_nor2_1 _7797_ (.A(_4078_),
    .B(_2469_),
    .Y(_2561_));
 sg13g2_o21ai_1 _7798_ (.B1(net226),
    .Y(_2562_),
    .A1(_2561_),
    .A2(_2508_));
 sg13g2_nand2_1 _7799_ (.Y(_2563_),
    .A(_2561_),
    .B(_2508_));
 sg13g2_nand2_1 _7800_ (.Y(_2564_),
    .A(_2562_),
    .B(_2563_));
 sg13g2_a221oi_1 _7801_ (.B2(net44),
    .C1(_2536_),
    .B1(_2564_),
    .A1(_2508_),
    .Y(_2565_),
    .A2(_2521_));
 sg13g2_xnor2_1 _7802_ (.Y(_2566_),
    .A(_0868_),
    .B(_2515_));
 sg13g2_xnor2_1 _7803_ (.Y(_2567_),
    .A(_2565_),
    .B(_2566_));
 sg13g2_xor2_1 _7804_ (.B(_2498_),
    .A(_2496_),
    .X(_2569_));
 sg13g2_xnor2_1 _7805_ (.Y(_2570_),
    .A(_2495_),
    .B(_2569_));
 sg13g2_nand2b_1 _7806_ (.Y(_2571_),
    .B(_2494_),
    .A_N(_2488_));
 sg13g2_xor2_1 _7807_ (.B(_2571_),
    .A(_2493_),
    .X(_2572_));
 sg13g2_xnor2_1 _7808_ (.Y(_2573_),
    .A(_1344_),
    .B(_2561_));
 sg13g2_xnor2_1 _7809_ (.Y(_2574_),
    .A(_2472_),
    .B(_2573_));
 sg13g2_nand2_1 _7810_ (.Y(_2575_),
    .A(_2506_),
    .B(_2574_));
 sg13g2_o21ai_1 _7811_ (.B1(_2575_),
    .Y(_2576_),
    .A1(_2503_),
    .A2(_2574_));
 sg13g2_nor4_1 _7812_ (.A(_2501_),
    .B(_2506_),
    .C(_2504_),
    .D(_2574_),
    .Y(_2577_));
 sg13g2_a21oi_2 _7813_ (.B1(_2577_),
    .Y(_2578_),
    .A2(_2576_),
    .A1(_2504_));
 sg13g2_a21oi_1 _7814_ (.A1(_2570_),
    .A2(_2572_),
    .Y(_2580_),
    .B1(_2578_));
 sg13g2_nand2_1 _7815_ (.Y(_2581_),
    .A(_2527_),
    .B(_2538_));
 sg13g2_xnor2_1 _7816_ (.Y(_2582_),
    .A(_0568_),
    .B(_2457_));
 sg13g2_xnor2_1 _7817_ (.Y(_2583_),
    .A(_2581_),
    .B(_2582_));
 sg13g2_o21ai_1 _7818_ (.B1(_2583_),
    .Y(_2584_),
    .A1(_2567_),
    .A2(_2580_));
 sg13g2_and2_1 _7819_ (.A(_2560_),
    .B(_2584_),
    .X(_2585_));
 sg13g2_nand2b_1 _7820_ (.Y(_2586_),
    .B(_2585_),
    .A_N(_2441_));
 sg13g2_nand3_1 _7821_ (.B(_2440_),
    .C(_2586_),
    .A(_2132_),
    .Y(_2587_));
 sg13g2_a21oi_1 _7822_ (.A1(net52),
    .A2(_1982_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_and2_1 _7823_ (.A(_1597_),
    .B(_2588_),
    .X(_2589_));
 sg13g2_nand2_1 _7824_ (.Y(_2591_),
    .A(_3870_),
    .B(net304));
 sg13g2_a221oi_1 _7825_ (.B2(_0808_),
    .C1(_0733_),
    .B1(_2591_),
    .A1(net169),
    .Y(_2592_),
    .A2(_0645_));
 sg13g2_nor2_1 _7826_ (.A(_1602_),
    .B(_2002_),
    .Y(_2593_));
 sg13g2_or2_1 _7827_ (.X(_2594_),
    .B(_2593_),
    .A(_2313_));
 sg13g2_buf_1 _7828_ (.A(_2594_),
    .X(_2595_));
 sg13g2_nand4_1 _7829_ (.B(_2331_),
    .C(_2232_),
    .A(net80),
    .Y(_2596_),
    .D(_2160_));
 sg13g2_and2_1 _7830_ (.A(net47),
    .B(_2596_),
    .X(_2597_));
 sg13g2_nor2_1 _7831_ (.A(_2340_),
    .B(_2351_),
    .Y(_2598_));
 sg13g2_a21oi_1 _7832_ (.A1(_2598_),
    .A2(_2376_),
    .Y(_2599_),
    .B1(net84));
 sg13g2_nor3_1 _7833_ (.A(_2595_),
    .B(_2597_),
    .C(_2599_),
    .Y(_2600_));
 sg13g2_nand2_1 _7834_ (.Y(_2602_),
    .A(_1602_),
    .B(_2331_));
 sg13g2_o21ai_1 _7835_ (.B1(net115),
    .Y(_2603_),
    .A1(_2602_),
    .A2(_1533_));
 sg13g2_nor3_1 _7836_ (.A(_1566_),
    .B(_2602_),
    .C(_1533_),
    .Y(_2604_));
 sg13g2_a22oi_1 _7837_ (.Y(_2605_),
    .B1(_2598_),
    .B2(_2604_),
    .A2(_2603_),
    .A1(_1595_));
 sg13g2_nand3_1 _7838_ (.B(_2160_),
    .C(net55),
    .A(net110),
    .Y(_2606_));
 sg13g2_nor4_1 _7839_ (.A(_2602_),
    .B(_2606_),
    .C(_1980_),
    .D(_2244_),
    .Y(_2607_));
 sg13g2_buf_1 _7840_ (.A(net74),
    .X(_2608_));
 sg13g2_a21oi_1 _7841_ (.A1(_2376_),
    .A2(_2607_),
    .Y(_2609_),
    .B1(net43));
 sg13g2_nor2_1 _7842_ (.A(_2605_),
    .B(_2609_),
    .Y(_2610_));
 sg13g2_nor2_1 _7843_ (.A(net53),
    .B(_2295_),
    .Y(_2611_));
 sg13g2_o21ai_1 _7844_ (.B1(_1526_),
    .Y(_2613_),
    .A1(_2309_),
    .A2(_2351_));
 sg13g2_a22oi_1 _7845_ (.Y(_2614_),
    .B1(net43),
    .B2(net56),
    .A2(_2613_),
    .A1(_2194_));
 sg13g2_o21ai_1 _7846_ (.B1(_1997_),
    .Y(_2615_),
    .A1(_1566_),
    .A2(_2606_));
 sg13g2_nand2_1 _7847_ (.Y(_2616_),
    .A(_2309_),
    .B(_2165_));
 sg13g2_a22oi_1 _7848_ (.Y(_2617_),
    .B1(net90),
    .B2(_2616_),
    .A2(_2003_),
    .A1(_2324_));
 sg13g2_a21oi_1 _7849_ (.A1(net85),
    .A2(_2127_),
    .Y(_2618_),
    .B1(net51));
 sg13g2_a22oi_1 _7850_ (.Y(_2619_),
    .B1(_2157_),
    .B2(_2232_),
    .A2(net73),
    .A1(_1595_));
 sg13g2_a21oi_1 _7851_ (.A1(_1559_),
    .A2(net90),
    .Y(_2620_),
    .B1(net56));
 sg13g2_nor4_1 _7852_ (.A(_2617_),
    .B(_2618_),
    .C(_2619_),
    .D(_2620_),
    .Y(_2621_));
 sg13g2_a21oi_1 _7853_ (.A1(net53),
    .A2(net91),
    .Y(_2622_),
    .B1(_2160_));
 sg13g2_or3_1 _7854_ (.A(_2359_),
    .B(_2406_),
    .C(_2622_),
    .X(_2624_));
 sg13g2_nor2_1 _7855_ (.A(_2394_),
    .B(_2148_),
    .Y(_2625_));
 sg13g2_nand3_1 _7856_ (.B(_2355_),
    .C(_2625_),
    .A(_1535_),
    .Y(_2626_));
 sg13g2_nand2_1 _7857_ (.Y(_2627_),
    .A(net52),
    .B(_1980_));
 sg13g2_nand4_1 _7858_ (.B(_2246_),
    .C(_2386_),
    .A(_2627_),
    .Y(_2628_),
    .D(_0905_));
 sg13g2_nor2_1 _7859_ (.A(_2035_),
    .B(_2230_),
    .Y(_2629_));
 sg13g2_or3_1 _7860_ (.A(_2361_),
    .B(_2629_),
    .C(_2233_),
    .X(_2630_));
 sg13g2_nor4_1 _7861_ (.A(_2624_),
    .B(_2626_),
    .C(_2628_),
    .D(_2630_),
    .Y(_2631_));
 sg13g2_nand3_1 _7862_ (.B(net119),
    .C(net78),
    .A(net114),
    .Y(_2632_));
 sg13g2_nand2_1 _7863_ (.Y(_2633_),
    .A(net73),
    .B(_2423_));
 sg13g2_nand3_1 _7864_ (.B(_2318_),
    .C(net78),
    .A(_2194_),
    .Y(_2635_));
 sg13g2_o21ai_1 _7865_ (.B1(net52),
    .Y(_2636_),
    .A1(_2369_),
    .A2(_2388_));
 sg13g2_o21ai_1 _7866_ (.B1(_2636_),
    .Y(_2637_),
    .A1(net84),
    .A2(net55));
 sg13g2_a221oi_1 _7867_ (.B2(_2635_),
    .C1(_2637_),
    .B1(_2633_),
    .A1(net92),
    .Y(_2638_),
    .A2(_2632_));
 sg13g2_nand4_1 _7868_ (.B(_2621_),
    .C(_2631_),
    .A(_2615_),
    .Y(_2639_),
    .D(_2638_));
 sg13g2_nor4_1 _7869_ (.A(_2611_),
    .B(_2422_),
    .C(_2614_),
    .D(_2639_),
    .Y(_2640_));
 sg13g2_nand4_1 _7870_ (.B(_2385_),
    .C(_2610_),
    .A(_2600_),
    .Y(_2641_),
    .D(_2640_));
 sg13g2_nand2_2 _7871_ (.Y(_2642_),
    .A(_2592_),
    .B(_2641_));
 sg13g2_a21oi_1 _7872_ (.A1(_0906_),
    .A2(_2589_),
    .Y(net6),
    .B1(_2642_));
 sg13g2_nand2_1 _7873_ (.Y(_2643_),
    .A(_1997_),
    .B(_2219_));
 sg13g2_o21ai_1 _7874_ (.B1(_4146_),
    .Y(_2645_),
    .A1(net124),
    .A2(_2046_));
 sg13g2_o21ai_1 _7875_ (.B1(_0930_),
    .Y(_2646_),
    .A1(net234),
    .A2(_1106_));
 sg13g2_o21ai_1 _7876_ (.B1(_2646_),
    .Y(_2647_),
    .A1(net217),
    .A2(_0996_));
 sg13g2_a22oi_1 _7877_ (.Y(_2648_),
    .B1(_2647_),
    .B2(net216),
    .A2(_0941_),
    .A1(net248));
 sg13g2_nor2_1 _7878_ (.A(net229),
    .B(_2648_),
    .Y(_2649_));
 sg13g2_nand2_1 _7879_ (.Y(_2650_),
    .A(_2645_),
    .B(_2649_));
 sg13g2_mux2_1 _7880_ (.A0(_0826_),
    .A1(_0807_),
    .S(_0788_),
    .X(_2651_));
 sg13g2_nor2_1 _7881_ (.A(_2650_),
    .B(_2651_),
    .Y(_2652_));
 sg13g2_nor2_2 _7882_ (.A(net112),
    .B(net80),
    .Y(_2653_));
 sg13g2_o21ai_1 _7883_ (.B1(_1383_),
    .Y(_2654_),
    .A1(_2298_),
    .A2(_1551_));
 sg13g2_a21oi_1 _7884_ (.A1(_2653_),
    .A2(_2654_),
    .Y(_2656_),
    .B1(_2381_));
 sg13g2_o21ai_1 _7885_ (.B1(_2656_),
    .Y(_2657_),
    .A1(_2643_),
    .A2(_2652_));
 sg13g2_nand2_1 _7886_ (.Y(_2658_),
    .A(net52),
    .B(_1547_));
 sg13g2_nand2_1 _7887_ (.Y(_2659_),
    .A(_1884_),
    .B(_1745_));
 sg13g2_or2_1 _7888_ (.X(_2660_),
    .B(_1862_),
    .A(_1812_));
 sg13g2_buf_1 _7889_ (.A(_2660_),
    .X(_2661_));
 sg13g2_nor3_1 _7890_ (.A(net162),
    .B(net111),
    .C(_2661_),
    .Y(_2662_));
 sg13g2_nor2_1 _7891_ (.A(_2659_),
    .B(_2662_),
    .Y(_2663_));
 sg13g2_a21o_1 _7892_ (.A2(_1988_),
    .A1(_1983_),
    .B1(net55),
    .X(_2664_));
 sg13g2_a21oi_1 _7893_ (.A1(net85),
    .A2(_2664_),
    .Y(_2665_),
    .B1(_1998_));
 sg13g2_a21oi_1 _7894_ (.A1(_2196_),
    .A2(_2205_),
    .Y(_2667_),
    .B1(_2226_));
 sg13g2_a21oi_1 _7895_ (.A1(_2016_),
    .A2(_2430_),
    .Y(_2668_),
    .B1(_2033_));
 sg13g2_o21ai_1 _7896_ (.B1(_0414_),
    .Y(_2669_),
    .A1(net258),
    .A2(_2668_));
 sg13g2_nor2_1 _7897_ (.A(net153),
    .B(_2669_),
    .Y(_2670_));
 sg13g2_nor2_1 _7898_ (.A(_2428_),
    .B(_2670_),
    .Y(_2671_));
 sg13g2_o21ai_1 _7899_ (.B1(_2367_),
    .Y(_2672_),
    .A1(_2432_),
    .A2(_2671_));
 sg13g2_nand2b_1 _7900_ (.Y(_2673_),
    .B(net256),
    .A_N(_2018_));
 sg13g2_buf_2 _7901_ (.A(_2673_),
    .X(_2674_));
 sg13g2_nor2_1 _7902_ (.A(net74),
    .B(_2318_),
    .Y(_2675_));
 sg13g2_nand2_1 _7903_ (.Y(_2676_),
    .A(_2674_),
    .B(_2675_));
 sg13g2_a21oi_1 _7904_ (.A1(net45),
    .A2(net72),
    .Y(_2678_),
    .B1(_2676_));
 sg13g2_nand3_1 _7905_ (.B(net111),
    .C(_2676_),
    .A(net29),
    .Y(_2679_));
 sg13g2_o21ai_1 _7906_ (.B1(_2679_),
    .Y(_2680_),
    .A1(_2320_),
    .A2(_2678_));
 sg13g2_a21oi_2 _7907_ (.B1(net121),
    .Y(_2681_),
    .A2(net149),
    .A1(net134));
 sg13g2_nand2_1 _7908_ (.Y(_2682_),
    .A(_1996_),
    .B(_2388_));
 sg13g2_nor2_1 _7909_ (.A(net188),
    .B(_2682_),
    .Y(_2683_));
 sg13g2_a221oi_1 _7910_ (.B2(_2683_),
    .C1(_2172_),
    .B1(_2681_),
    .A1(net115),
    .Y(_2684_),
    .A2(_2188_));
 sg13g2_nand4_1 _7911_ (.B(_2672_),
    .C(_2680_),
    .A(_2667_),
    .Y(_2685_),
    .D(_2684_));
 sg13g2_nor2_1 _7912_ (.A(_2366_),
    .B(_2669_),
    .Y(_2686_));
 sg13g2_nor2_1 _7913_ (.A(_1587_),
    .B(_2686_),
    .Y(_2687_));
 sg13g2_nand2_1 _7914_ (.Y(_2689_),
    .A(net162),
    .B(_2687_));
 sg13g2_nor2_1 _7915_ (.A(_2136_),
    .B(_2275_),
    .Y(_2690_));
 sg13g2_o21ai_1 _7916_ (.B1(net46),
    .Y(_2691_),
    .A1(net77),
    .A2(_2690_));
 sg13g2_nor2_1 _7917_ (.A(_2246_),
    .B(_2691_),
    .Y(_2692_));
 sg13g2_a21oi_1 _7918_ (.A1(_2434_),
    .A2(_2689_),
    .Y(_2693_),
    .B1(_2692_));
 sg13g2_o21ai_1 _7919_ (.B1(_2693_),
    .Y(_2694_),
    .A1(_2186_),
    .A2(_2189_));
 sg13g2_nor2_1 _7920_ (.A(_2685_),
    .B(_2694_),
    .Y(_2695_));
 sg13g2_nand3_1 _7921_ (.B(net81),
    .C(_2215_),
    .A(_2674_),
    .Y(_2696_));
 sg13g2_buf_1 _7922_ (.A(_2696_),
    .X(_2697_));
 sg13g2_o21ai_1 _7923_ (.B1(net27),
    .Y(_2698_),
    .A1(net135),
    .A2(_2697_));
 sg13g2_nor2_2 _7924_ (.A(_2192_),
    .B(_2035_),
    .Y(_2699_));
 sg13g2_and2_1 _7925_ (.A(_2413_),
    .B(_2699_),
    .X(_2700_));
 sg13g2_nor3_1 _7926_ (.A(net97),
    .B(net31),
    .C(_2257_),
    .Y(_2701_));
 sg13g2_inv_1 _7927_ (.Y(_2702_),
    .A(_2701_));
 sg13g2_o21ai_1 _7928_ (.B1(_1551_),
    .Y(_2703_),
    .A1(net156),
    .A2(net57));
 sg13g2_nand2_1 _7929_ (.Y(_2704_),
    .A(net195),
    .B(_1480_));
 sg13g2_o21ai_1 _7930_ (.B1(_2704_),
    .Y(_2705_),
    .A1(net57),
    .A2(_2285_));
 sg13g2_a21o_1 _7931_ (.A2(_2703_),
    .A1(net185),
    .B1(_2705_),
    .X(_2706_));
 sg13g2_nor3_1 _7932_ (.A(_2328_),
    .B(_1558_),
    .C(_2706_),
    .Y(_2707_));
 sg13g2_a221oi_1 _7933_ (.B2(_2406_),
    .C1(_2707_),
    .B1(_2702_),
    .A1(_2698_),
    .Y(_2708_),
    .A2(_2700_));
 sg13g2_nor2_2 _7934_ (.A(_0832_),
    .B(net149),
    .Y(_2710_));
 sg13g2_o21ai_1 _7935_ (.B1(_2710_),
    .Y(_2711_),
    .A1(net169),
    .A2(net45));
 sg13g2_nor3_1 _7936_ (.A(net43),
    .B(net78),
    .C(net121),
    .Y(_2712_));
 sg13g2_a22oi_1 _7937_ (.Y(_2713_),
    .B1(_2711_),
    .B2(_2712_),
    .A2(_2681_),
    .A1(_2395_));
 sg13g2_nor2_1 _7938_ (.A(net132),
    .B(net120),
    .Y(_2714_));
 sg13g2_nor3_1 _7939_ (.A(net110),
    .B(net43),
    .C(_2714_),
    .Y(_2715_));
 sg13g2_o21ai_1 _7940_ (.B1(net183),
    .Y(_2716_),
    .A1(_2637_),
    .A2(_2715_));
 sg13g2_nor2_1 _7941_ (.A(net133),
    .B(_2337_),
    .Y(_2717_));
 sg13g2_a21oi_1 _7942_ (.A1(net255),
    .A2(_0873_),
    .Y(_2718_),
    .B1(net193));
 sg13g2_nor2b_1 _7943_ (.A(_2718_),
    .B_N(_0990_),
    .Y(_2719_));
 sg13g2_nand3_1 _7944_ (.B(_0994_),
    .C(_2211_),
    .A(net198),
    .Y(_2721_));
 sg13g2_o21ai_1 _7945_ (.B1(_2721_),
    .Y(_2722_),
    .A1(_0991_),
    .A2(_2719_));
 sg13g2_and2_1 _7946_ (.A(_1027_),
    .B(_2346_),
    .X(_2723_));
 sg13g2_buf_1 _7947_ (.A(_2723_),
    .X(_2724_));
 sg13g2_nand3b_1 _7948_ (.B(_2722_),
    .C(_2724_),
    .Y(_2725_),
    .A_N(_2717_));
 sg13g2_nand3_1 _7949_ (.B(_2716_),
    .C(_2725_),
    .A(_2713_),
    .Y(_2726_));
 sg13g2_nor2_2 _7950_ (.A(net112),
    .B(net119),
    .Y(_2727_));
 sg13g2_a21oi_1 _7951_ (.A1(_0832_),
    .A2(net45),
    .Y(_2728_),
    .B1(_2355_));
 sg13g2_a21oi_1 _7952_ (.A1(net149),
    .A2(_2727_),
    .Y(_2729_),
    .B1(_2728_));
 sg13g2_nor2_1 _7953_ (.A(net132),
    .B(net109),
    .Y(_2730_));
 sg13g2_nor2_1 _7954_ (.A(_2331_),
    .B(net116),
    .Y(_2732_));
 sg13g2_a21oi_1 _7955_ (.A1(net132),
    .A2(_2403_),
    .Y(_2733_),
    .B1(_2376_));
 sg13g2_o21ai_1 _7956_ (.B1(net48),
    .Y(_2734_),
    .A1(_2732_),
    .A2(_2733_));
 sg13g2_o21ai_1 _7957_ (.B1(_2734_),
    .Y(_2735_),
    .A1(_2729_),
    .A2(_2730_));
 sg13g2_nand2_1 _7958_ (.Y(_2736_),
    .A(_2383_),
    .B(_2420_));
 sg13g2_o21ai_1 _7959_ (.B1(_2736_),
    .Y(_2737_),
    .A1(_2600_),
    .A2(_2216_));
 sg13g2_nand2_1 _7960_ (.Y(_2738_),
    .A(net76),
    .B(_2216_));
 sg13g2_nor2_1 _7961_ (.A(_2293_),
    .B(_2191_),
    .Y(_2739_));
 sg13g2_nand2_1 _7962_ (.Y(_2740_),
    .A(net76),
    .B(net30));
 sg13g2_a22oi_1 _7963_ (.Y(_2741_),
    .B1(_2739_),
    .B2(_2740_),
    .A2(_2738_),
    .A1(_2291_));
 sg13g2_nand2_1 _7964_ (.Y(_2743_),
    .A(_2164_),
    .B(_1547_));
 sg13g2_nand2_1 _7965_ (.Y(_2744_),
    .A(_2674_),
    .B(net46));
 sg13g2_a221oi_1 _7966_ (.B2(_2743_),
    .C1(_2744_),
    .B1(_2398_),
    .A1(net45),
    .Y(_2745_),
    .A2(_2282_));
 sg13g2_nand2_1 _7967_ (.Y(_2746_),
    .A(_1526_),
    .B(_1452_));
 sg13g2_a21oi_1 _7968_ (.A1(net119),
    .A2(_1559_),
    .Y(_2747_),
    .B1(_2746_));
 sg13g2_nand2_1 _7969_ (.Y(_2748_),
    .A(_2148_),
    .B(_2215_));
 sg13g2_nand3_1 _7970_ (.B(net108),
    .C(net30),
    .A(net52),
    .Y(_2749_));
 sg13g2_o21ai_1 _7971_ (.B1(_2749_),
    .Y(_2750_),
    .A1(_2020_),
    .A2(_2748_));
 sg13g2_nor3_1 _7972_ (.A(_2745_),
    .B(_2747_),
    .C(_2750_),
    .Y(_2751_));
 sg13g2_nor2_1 _7973_ (.A(net162),
    .B(_2241_),
    .Y(_2752_));
 sg13g2_or3_1 _7974_ (.A(net310),
    .B(net311),
    .C(net312),
    .X(_2754_));
 sg13g2_buf_1 _7975_ (.A(_2754_),
    .X(_2755_));
 sg13g2_nor3_1 _7976_ (.A(_2035_),
    .B(net109),
    .C(_2755_),
    .Y(_2756_));
 sg13g2_a221oi_1 _7977_ (.B2(_2188_),
    .C1(_2756_),
    .B1(net153),
    .A1(net83),
    .Y(_2757_),
    .A2(net116));
 sg13g2_o21ai_1 _7978_ (.B1(_2344_),
    .Y(_2758_),
    .A1(net94),
    .A2(_2717_));
 sg13g2_nand2_1 _7979_ (.Y(_2759_),
    .A(_2361_),
    .B(_2758_));
 sg13g2_o21ai_1 _7980_ (.B1(_2759_),
    .Y(_2760_),
    .A1(net43),
    .A2(_2757_));
 sg13g2_a221oi_1 _7981_ (.B2(_2752_),
    .C1(_2760_),
    .B1(_2321_),
    .A1(_2617_),
    .Y(_2761_),
    .A2(_2012_));
 sg13g2_or2_1 _7982_ (.X(_2762_),
    .B(_0903_),
    .A(_1989_));
 sg13g2_nand3_1 _7983_ (.B(net281),
    .C(_1160_),
    .A(_3870_),
    .Y(_2763_));
 sg13g2_o21ai_1 _7984_ (.B1(_0820_),
    .Y(_2765_),
    .A1(_4113_),
    .A2(_2763_));
 sg13g2_buf_2 _7985_ (.A(_2765_),
    .X(_2766_));
 sg13g2_nand3_1 _7986_ (.B(_2353_),
    .C(_2766_),
    .A(net134),
    .Y(_2767_));
 sg13g2_nand2b_1 _7987_ (.Y(_2768_),
    .B(_2767_),
    .A_N(_2173_));
 sg13g2_o21ai_1 _7988_ (.B1(_2233_),
    .Y(_2769_),
    .A1(_2299_),
    .A2(_1816_));
 sg13g2_o21ai_1 _7989_ (.B1(_2769_),
    .Y(_2770_),
    .A1(_2423_),
    .A2(_2010_));
 sg13g2_nor2_1 _7990_ (.A(_1538_),
    .B(_2376_),
    .Y(_2771_));
 sg13g2_nor3_1 _7991_ (.A(_2127_),
    .B(net84),
    .C(_4512_),
    .Y(_2772_));
 sg13g2_nor4_1 _7992_ (.A(_2768_),
    .B(_2770_),
    .C(_2771_),
    .D(_2772_),
    .Y(_2773_));
 sg13g2_o21ai_1 _7993_ (.B1(_2773_),
    .Y(_2774_),
    .A1(_2762_),
    .A2(net111));
 sg13g2_nor4_1 _7994_ (.A(_2611_),
    .B(_2422_),
    .C(_2614_),
    .D(_2774_),
    .Y(_2776_));
 sg13g2_nand4_1 _7995_ (.B(_2751_),
    .C(_2761_),
    .A(_2741_),
    .Y(_2777_),
    .D(_2776_));
 sg13g2_nor4_1 _7996_ (.A(_2726_),
    .B(_2735_),
    .C(_2737_),
    .D(_2777_),
    .Y(_2778_));
 sg13g2_nand3_1 _7997_ (.B(_2708_),
    .C(_2778_),
    .A(_2695_),
    .Y(_2779_));
 sg13g2_nor2_1 _7998_ (.A(_2570_),
    .B(_2572_),
    .Y(_2780_));
 sg13g2_nor2b_1 _7999_ (.A(_2578_),
    .B_N(_2780_),
    .Y(_2781_));
 sg13g2_nor3_1 _8000_ (.A(_2583_),
    .B(_2567_),
    .C(_2781_),
    .Y(_2782_));
 sg13g2_nor2_1 _8001_ (.A(_2583_),
    .B(_2567_),
    .Y(_2783_));
 sg13g2_xor2_1 _8002_ (.B(_2574_),
    .A(_2508_),
    .X(_2784_));
 sg13g2_nand2_1 _8003_ (.Y(_2785_),
    .A(_2780_),
    .B(_2784_));
 sg13g2_nand3_1 _8004_ (.B(_2783_),
    .C(_2785_),
    .A(_2578_),
    .Y(_2787_));
 sg13g2_mux2_1 _8005_ (.A0(_2782_),
    .A1(_2787_),
    .S(_2559_),
    .X(_2788_));
 sg13g2_nor3_1 _8006_ (.A(_2441_),
    .B(_2550_),
    .C(_2788_),
    .Y(_2789_));
 sg13g2_a21oi_1 _8007_ (.A1(_0874_),
    .A2(_2252_),
    .Y(_2790_),
    .B1(_1002_));
 sg13g2_nor4_1 _8008_ (.A(_0524_),
    .B(_2249_),
    .C(_4091_),
    .D(_0866_),
    .Y(_2791_));
 sg13g2_nor4_1 _8009_ (.A(net187),
    .B(_0524_),
    .C(_4157_),
    .D(_2199_),
    .Y(_2792_));
 sg13g2_nand3_1 _8010_ (.B(_1087_),
    .C(_1581_),
    .A(net220),
    .Y(_2793_));
 sg13g2_a21oi_1 _8011_ (.A1(_0990_),
    .A2(_2793_),
    .Y(_2794_),
    .B1(_0991_));
 sg13g2_a21oi_1 _8012_ (.A1(net262),
    .A2(_2792_),
    .Y(_2795_),
    .B1(_2794_));
 sg13g2_nor4_1 _8013_ (.A(net229),
    .B(_2790_),
    .C(_2791_),
    .D(_2795_),
    .Y(_2796_));
 sg13g2_nor3_1 _8014_ (.A(_2177_),
    .B(_0934_),
    .C(_1611_),
    .Y(_2798_));
 sg13g2_nor2_1 _8015_ (.A(_1466_),
    .B(net247),
    .Y(_2799_));
 sg13g2_nor2_1 _8016_ (.A(net201),
    .B(net213),
    .Y(_2800_));
 sg13g2_nand4_1 _8017_ (.B(_3406_),
    .C(_2799_),
    .A(_1106_),
    .Y(_2801_),
    .D(_2800_));
 sg13g2_o21ai_1 _8018_ (.B1(_2801_),
    .Y(_2802_),
    .A1(net304),
    .A2(_2798_));
 sg13g2_or2_1 _8019_ (.X(_2803_),
    .B(net237),
    .A(_1358_));
 sg13g2_nand4_1 _8020_ (.B(net234),
    .C(_1007_),
    .A(_3568_),
    .Y(_2804_),
    .D(_2803_));
 sg13g2_o21ai_1 _8021_ (.B1(_2804_),
    .Y(_2805_),
    .A1(net234),
    .A2(_2802_));
 sg13g2_nor4_1 _8022_ (.A(_0722_),
    .B(_2249_),
    .C(_1581_),
    .D(_2253_),
    .Y(_2806_));
 sg13g2_nor2_1 _8023_ (.A(net206),
    .B(_2806_),
    .Y(_2807_));
 sg13g2_or2_1 _8024_ (.X(_2809_),
    .B(_0829_),
    .A(net189));
 sg13g2_o21ai_1 _8025_ (.B1(_0414_),
    .Y(_2810_),
    .A1(_2807_),
    .A2(_2809_));
 sg13g2_and2_1 _8026_ (.A(_1045_),
    .B(_1047_),
    .X(_2811_));
 sg13g2_o21ai_1 _8027_ (.B1(net180),
    .Y(_2812_),
    .A1(net160),
    .A2(net217));
 sg13g2_o21ai_1 _8028_ (.B1(net172),
    .Y(_2813_),
    .A1(net213),
    .A2(net245));
 sg13g2_a22oi_1 _8029_ (.Y(_2814_),
    .B1(_2813_),
    .B2(_2473_),
    .A2(_2812_),
    .A1(_2181_));
 sg13g2_nor4_1 _8030_ (.A(net216),
    .B(_2811_),
    .C(_1684_),
    .D(_2814_),
    .Y(_2815_));
 sg13g2_a22oi_1 _8031_ (.Y(_2816_),
    .B1(_2810_),
    .B2(_2815_),
    .A2(_2805_),
    .A1(_2796_));
 sg13g2_nor4_1 _8032_ (.A(net56),
    .B(net90),
    .C(net30),
    .D(_2816_),
    .Y(_2817_));
 sg13g2_or2_1 _8033_ (.X(_2818_),
    .B(_2817_),
    .A(_2131_));
 sg13g2_nor4_1 _8034_ (.A(_2665_),
    .B(_2779_),
    .C(_2789_),
    .D(_2818_),
    .Y(_2820_));
 sg13g2_o21ai_1 _8035_ (.B1(_2820_),
    .Y(_2821_),
    .A1(_2658_),
    .A2(_2663_));
 sg13g2_nor2_1 _8036_ (.A(net24),
    .B(_1522_),
    .Y(_2822_));
 sg13g2_and2_1 _8037_ (.A(_1477_),
    .B(_2822_),
    .X(_2823_));
 sg13g2_and2_1 _8038_ (.A(_1939_),
    .B(_1976_),
    .X(_2824_));
 sg13g2_buf_1 _8039_ (.A(_2824_),
    .X(_2825_));
 sg13g2_a21o_1 _8040_ (.A2(_2825_),
    .A1(_2752_),
    .B1(_1862_),
    .X(_2826_));
 sg13g2_nor2_1 _8041_ (.A(_0937_),
    .B(_1617_),
    .Y(_2827_));
 sg13g2_o21ai_1 _8042_ (.B1(_1718_),
    .Y(_2828_),
    .A1(_3342_),
    .A2(_3601_));
 sg13g2_a22oi_1 _8043_ (.Y(_2829_),
    .B1(_2828_),
    .B2(_1465_),
    .A2(_2827_),
    .A1(_0926_));
 sg13g2_xnor2_1 _8044_ (.Y(_2830_),
    .A(_1438_),
    .B(_2829_));
 sg13g2_buf_1 _8045_ (.A(_2830_),
    .X(_2831_));
 sg13g2_o21ai_1 _8046_ (.B1(net266),
    .Y(_2832_),
    .A1(net279),
    .A2(_0934_));
 sg13g2_nand3_1 _8047_ (.B(net276),
    .C(net278),
    .A(net277),
    .Y(_2833_));
 sg13g2_nand3_1 _8048_ (.B(net231),
    .C(_2833_),
    .A(net214),
    .Y(_2834_));
 sg13g2_a21oi_1 _8049_ (.A1(_2832_),
    .A2(_2834_),
    .Y(_2835_),
    .B1(_4440_));
 sg13g2_xor2_1 _8050_ (.B(net230),
    .A(net266),
    .X(_2836_));
 sg13g2_nor2_1 _8051_ (.A(net202),
    .B(_2836_),
    .Y(_2837_));
 sg13g2_o21ai_1 _8052_ (.B1(net284),
    .Y(_2838_),
    .A1(_0937_),
    .A2(_1611_));
 sg13g2_buf_2 _8053_ (.A(_2838_),
    .X(_2839_));
 sg13g2_nand2_2 _8054_ (.Y(_2841_),
    .A(net228),
    .B(_2839_));
 sg13g2_mux2_1 _8055_ (.A0(_2835_),
    .A1(_2837_),
    .S(_2841_),
    .X(_2842_));
 sg13g2_and3_1 _8056_ (.X(_2843_),
    .A(net203),
    .B(net131),
    .C(_2842_));
 sg13g2_buf_2 _8057_ (.A(_2843_),
    .X(_2844_));
 sg13g2_nand2_1 _8058_ (.Y(_2845_),
    .A(_0149_),
    .B(_2844_));
 sg13g2_xnor2_1 _8059_ (.Y(_2846_),
    .A(_3438_),
    .B(net270));
 sg13g2_nand2_1 _8060_ (.Y(_2847_),
    .A(_3677_),
    .B(_2846_));
 sg13g2_o21ai_1 _8061_ (.B1(_2847_),
    .Y(_2848_),
    .A1(net270),
    .A2(net194));
 sg13g2_nor2_1 _8062_ (.A(net241),
    .B(net279),
    .Y(_2849_));
 sg13g2_a21o_1 _8063_ (.A2(_2839_),
    .A1(net228),
    .B1(_2849_),
    .X(_2850_));
 sg13g2_o21ai_1 _8064_ (.B1(_2850_),
    .Y(_2852_),
    .A1(_2841_),
    .A2(_2848_));
 sg13g2_buf_1 _8065_ (.A(_2852_),
    .X(_2853_));
 sg13g2_buf_1 _8066_ (.A(_2853_),
    .X(_2854_));
 sg13g2_nand2_1 _8067_ (.Y(_2855_),
    .A(_1237_),
    .B(_2833_));
 sg13g2_nand3_1 _8068_ (.B(_2839_),
    .C(_2855_),
    .A(net228),
    .Y(_2856_));
 sg13g2_nand2b_1 _8069_ (.Y(_2857_),
    .B(net278),
    .A_N(net279));
 sg13g2_o21ai_1 _8070_ (.B1(net270),
    .Y(_2858_),
    .A1(_3794_),
    .A2(_2857_));
 sg13g2_a21o_1 _8071_ (.A2(_2839_),
    .A1(net228),
    .B1(_2858_),
    .X(_2859_));
 sg13g2_and3_1 _8072_ (.X(_2860_),
    .A(net266),
    .B(_2856_),
    .C(_2859_));
 sg13g2_buf_1 _8073_ (.A(_2860_),
    .X(_2861_));
 sg13g2_a21oi_1 _8074_ (.A1(_2856_),
    .A2(_2859_),
    .Y(_2863_),
    .B1(net266));
 sg13g2_or3_1 _8075_ (.A(_4555_),
    .B(_2861_),
    .C(_2863_),
    .X(_2864_));
 sg13g2_buf_1 _8076_ (.A(_2864_),
    .X(_2865_));
 sg13g2_buf_1 _8077_ (.A(_2865_),
    .X(_2866_));
 sg13g2_a21oi_1 _8078_ (.A1(net284),
    .A2(_1611_),
    .Y(_2867_),
    .B1(_2755_));
 sg13g2_buf_1 _8079_ (.A(_2867_),
    .X(_2868_));
 sg13g2_xnor2_1 _8080_ (.Y(_2869_),
    .A(_1281_),
    .B(_2868_));
 sg13g2_nand2_1 _8081_ (.Y(_2870_),
    .A(net240),
    .B(_1465_));
 sg13g2_a221oi_1 _8082_ (.B2(net237),
    .C1(_3794_),
    .B1(_2870_),
    .A1(_0395_),
    .Y(_2871_),
    .A2(_2868_));
 sg13g2_a21o_1 _8083_ (.A2(_2869_),
    .A1(net199),
    .B1(_2871_),
    .X(_2872_));
 sg13g2_buf_1 _8084_ (.A(_2872_),
    .X(_2874_));
 sg13g2_xnor2_1 _8085_ (.Y(_2875_),
    .A(_1237_),
    .B(_0937_));
 sg13g2_xnor2_1 _8086_ (.Y(_2876_),
    .A(_4471_),
    .B(_0934_));
 sg13g2_and3_1 _8087_ (.X(_2877_),
    .A(net228),
    .B(_2839_),
    .C(_2876_));
 sg13g2_a21oi_1 _8088_ (.A1(_2841_),
    .A2(_2875_),
    .Y(_2878_),
    .B1(_2877_));
 sg13g2_buf_1 _8089_ (.A(_2878_),
    .X(_2879_));
 sg13g2_nand2_1 _8090_ (.Y(_2880_),
    .A(_2874_),
    .B(net107));
 sg13g2_buf_2 _8091_ (.A(_2880_),
    .X(_2881_));
 sg13g2_a21oi_1 _8092_ (.A1(net71),
    .A2(net26),
    .Y(_2882_),
    .B1(_2881_));
 sg13g2_nand2_1 _8093_ (.Y(_2883_),
    .A(net122),
    .B(_2882_));
 sg13g2_nand2_1 _8094_ (.Y(_2885_),
    .A(_2845_),
    .B(_2883_));
 sg13g2_a21oi_1 _8095_ (.A1(net203),
    .A2(net131),
    .Y(_2886_),
    .B1(_2842_));
 sg13g2_buf_1 _8096_ (.A(_2886_),
    .X(_2887_));
 sg13g2_a21o_1 _8097_ (.A2(_2875_),
    .A1(_2841_),
    .B1(_2877_),
    .X(_2888_));
 sg13g2_buf_1 _8098_ (.A(_2888_),
    .X(_2889_));
 sg13g2_nand3_1 _8099_ (.B(net71),
    .C(net26),
    .A(net106),
    .Y(_2890_));
 sg13g2_a21oi_1 _8100_ (.A1(_3794_),
    .A2(_2869_),
    .Y(_2891_),
    .B1(_2871_));
 sg13g2_buf_2 _8101_ (.A(_2891_),
    .X(_2892_));
 sg13g2_o21ai_1 _8102_ (.B1(_2892_),
    .Y(_2893_),
    .A1(_2854_),
    .A2(net26));
 sg13g2_and2_1 _8103_ (.A(_2890_),
    .B(_2893_),
    .X(_2894_));
 sg13g2_inv_1 _8104_ (.Y(_2896_),
    .A(_2894_));
 sg13g2_nor2_1 _8105_ (.A(net70),
    .B(_2896_),
    .Y(_2897_));
 sg13g2_nor2_1 _8106_ (.A(net122),
    .B(_2844_),
    .Y(_2898_));
 sg13g2_nor2b_1 _8107_ (.A(_2882_),
    .B_N(net70),
    .Y(_2899_));
 sg13g2_a22oi_1 _8108_ (.Y(_2900_),
    .B1(_2899_),
    .B2(net122),
    .A2(_2898_),
    .A1(_2896_));
 sg13g2_xnor2_1 _8109_ (.Y(_2901_),
    .A(_0342_),
    .B(_0295_));
 sg13g2_buf_2 _8110_ (.A(_2901_),
    .X(_2902_));
 sg13g2_buf_1 _8111_ (.A(_0300_),
    .X(_2903_));
 sg13g2_a21oi_2 _8112_ (.B1(net69),
    .Y(_2904_),
    .A2(_0202_),
    .A1(net146));
 sg13g2_xnor2_1 _8113_ (.Y(_2905_),
    .A(_2887_),
    .B(_2904_));
 sg13g2_nor4_2 _8114_ (.A(net143),
    .B(_4201_),
    .C(_4224_),
    .Y(_2907_),
    .D(net99));
 sg13g2_xnor2_1 _8115_ (.Y(_2908_),
    .A(_2844_),
    .B(_2907_));
 sg13g2_mux2_1 _8116_ (.A0(_2905_),
    .A1(_2908_),
    .S(net122),
    .X(_2909_));
 sg13g2_xnor2_1 _8117_ (.Y(_2910_),
    .A(net64),
    .B(_2909_));
 sg13g2_xor2_1 _8118_ (.B(_2910_),
    .A(_2902_),
    .X(_2911_));
 sg13g2_a22oi_1 _8119_ (.Y(_2912_),
    .B1(_2900_),
    .B2(_2911_),
    .A2(_2897_),
    .A1(_2885_));
 sg13g2_nor2_2 _8120_ (.A(net125),
    .B(net50),
    .Y(_2913_));
 sg13g2_nor2_1 _8121_ (.A(_2861_),
    .B(_2863_),
    .Y(_2914_));
 sg13g2_buf_1 _8122_ (.A(_2914_),
    .X(_2915_));
 sg13g2_buf_1 _8123_ (.A(net107),
    .X(_2916_));
 sg13g2_nand2_1 _8124_ (.Y(_2918_),
    .A(net42),
    .B(_2916_));
 sg13g2_xnor2_1 _8125_ (.Y(_2919_),
    .A(_2913_),
    .B(_2918_));
 sg13g2_nand3_1 _8126_ (.B(net82),
    .C(net69),
    .A(net126),
    .Y(_2920_));
 sg13g2_a22oi_1 _8127_ (.Y(_2921_),
    .B1(_2904_),
    .B2(net70),
    .A2(_2920_),
    .A1(net122));
 sg13g2_o21ai_1 _8128_ (.B1(net106),
    .Y(_2922_),
    .A1(_2844_),
    .A2(_2921_));
 sg13g2_a21o_1 _8129_ (.A2(net82),
    .A1(net126),
    .B1(net69),
    .X(_2923_));
 sg13g2_a22oi_1 _8130_ (.Y(_2924_),
    .B1(_2923_),
    .B2(_0149_),
    .A2(_2907_),
    .A1(_2844_));
 sg13g2_buf_1 _8131_ (.A(_2924_),
    .X(_2925_));
 sg13g2_o21ai_1 _8132_ (.B1(net62),
    .Y(_2926_),
    .A1(net70),
    .A2(_2925_));
 sg13g2_o21ai_1 _8133_ (.B1(_2926_),
    .Y(_2927_),
    .A1(net62),
    .A2(_2922_));
 sg13g2_nor2_1 _8134_ (.A(net70),
    .B(_2925_),
    .Y(_2929_));
 sg13g2_or2_1 _8135_ (.X(_2930_),
    .B(_2921_),
    .A(_2844_));
 sg13g2_buf_1 _8136_ (.A(_2930_),
    .X(_2931_));
 sg13g2_o21ai_1 _8137_ (.B1(_2931_),
    .Y(_2932_),
    .A1(net64),
    .A2(_2929_));
 sg13g2_nor2_1 _8138_ (.A(net62),
    .B(net107),
    .Y(_2933_));
 sg13g2_a21oi_1 _8139_ (.A1(net62),
    .A2(_2931_),
    .Y(_2934_),
    .B1(_2933_));
 sg13g2_a221oi_1 _8140_ (.B2(_2934_),
    .C1(_0166_),
    .B1(_2932_),
    .A1(net32),
    .Y(_2935_),
    .A2(_2927_));
 sg13g2_o21ai_1 _8141_ (.B1(net107),
    .Y(_2936_),
    .A1(net70),
    .A2(_2925_));
 sg13g2_o21ai_1 _8142_ (.B1(_0320_),
    .Y(_2937_),
    .A1(_2844_),
    .A2(_2921_));
 sg13g2_o21ai_1 _8143_ (.B1(_2937_),
    .Y(_2938_),
    .A1(_0320_),
    .A2(_2936_));
 sg13g2_nand2_1 _8144_ (.Y(_2940_),
    .A(net62),
    .B(net107));
 sg13g2_nand2_1 _8145_ (.Y(_2941_),
    .A(net64),
    .B(net62));
 sg13g2_o21ai_1 _8146_ (.B1(_2941_),
    .Y(_2942_),
    .A1(net70),
    .A2(_2925_));
 sg13g2_and2_1 _8147_ (.A(_2940_),
    .B(_2942_),
    .X(_2943_));
 sg13g2_a221oi_1 _8148_ (.B2(_2931_),
    .C1(_0342_),
    .B1(_2943_),
    .A1(net65),
    .Y(_2944_),
    .A2(_2938_));
 sg13g2_nor2_1 _8149_ (.A(_2931_),
    .B(_2940_),
    .Y(_2945_));
 sg13g2_a21oi_1 _8150_ (.A1(_2929_),
    .A2(_2933_),
    .Y(_2946_),
    .B1(_2945_));
 sg13g2_o21ai_1 _8151_ (.B1(_2946_),
    .Y(_2947_),
    .A1(_2935_),
    .A2(_2944_));
 sg13g2_buf_2 _8152_ (.A(_2947_),
    .X(_2948_));
 sg13g2_mux2_1 _8153_ (.A0(_2912_),
    .A1(_2919_),
    .S(_2948_),
    .X(_2949_));
 sg13g2_inv_1 _8154_ (.Y(_2951_),
    .A(_2919_));
 sg13g2_mux2_1 _8155_ (.A0(_2951_),
    .A1(_2912_),
    .S(_2948_),
    .X(_2952_));
 sg13g2_a22oi_1 _8156_ (.Y(_2953_),
    .B1(net82),
    .B2(net104),
    .A2(net49),
    .A1(net126));
 sg13g2_nand4_1 _8157_ (.B(net104),
    .C(net49),
    .A(net126),
    .Y(_2954_),
    .D(net82));
 sg13g2_o21ai_1 _8158_ (.B1(_2954_),
    .Y(_2955_),
    .A1(net64),
    .A2(_2953_));
 sg13g2_buf_1 _8159_ (.A(_2955_),
    .X(_2956_));
 sg13g2_buf_1 _8160_ (.A(_2956_),
    .X(_2957_));
 sg13g2_a21oi_1 _8161_ (.A1(net240),
    .A2(_2868_),
    .Y(_2958_),
    .B1(net202));
 sg13g2_nand4_1 _8162_ (.B(net240),
    .C(net228),
    .A(net202),
    .Y(_2959_),
    .D(_2839_));
 sg13g2_nand2b_1 _8163_ (.Y(_2960_),
    .B(_2959_),
    .A_N(_2958_));
 sg13g2_buf_2 _8164_ (.A(_2960_),
    .X(_2962_));
 sg13g2_nand2_1 _8165_ (.Y(_2963_),
    .A(net131),
    .B(_2962_));
 sg13g2_buf_2 _8166_ (.A(_2963_),
    .X(_2964_));
 sg13g2_or2_1 _8167_ (.X(_2965_),
    .B(_2863_),
    .A(_2861_));
 sg13g2_buf_1 _8168_ (.A(_2965_),
    .X(_2966_));
 sg13g2_buf_1 _8169_ (.A(_2892_),
    .X(_2967_));
 sg13g2_nor2_1 _8170_ (.A(net41),
    .B(net67),
    .Y(_2968_));
 sg13g2_xnor2_1 _8171_ (.Y(_2969_),
    .A(_2964_),
    .B(_2968_));
 sg13g2_xnor2_1 _8172_ (.Y(_2970_),
    .A(net16),
    .B(_2969_));
 sg13g2_mux2_1 _8173_ (.A0(_2949_),
    .A1(_2952_),
    .S(_2970_),
    .X(_2971_));
 sg13g2_buf_1 _8174_ (.A(_2971_),
    .X(_2973_));
 sg13g2_a21oi_1 _8175_ (.A1(net64),
    .A2(net99),
    .Y(_2974_),
    .B1(net50));
 sg13g2_o21ai_1 _8176_ (.B1(_2974_),
    .Y(_2975_),
    .A1(net101),
    .A2(net98));
 sg13g2_nand2_1 _8177_ (.Y(_2976_),
    .A(net65),
    .B(net82));
 sg13g2_a21oi_1 _8178_ (.A1(net50),
    .A2(_2976_),
    .Y(_2977_),
    .B1(net125));
 sg13g2_a22oi_1 _8179_ (.Y(_2978_),
    .B1(_2975_),
    .B2(_2977_),
    .A2(net69),
    .A1(_4286_));
 sg13g2_nand3_1 _8180_ (.B(net67),
    .C(_2978_),
    .A(_2964_),
    .Y(_2979_));
 sg13g2_o21ai_1 _8181_ (.B1(net68),
    .Y(_2980_),
    .A1(_2964_),
    .A2(net67));
 sg13g2_inv_1 _8182_ (.Y(_2981_),
    .A(_2980_));
 sg13g2_nor2_1 _8183_ (.A(_2964_),
    .B(net68),
    .Y(_2982_));
 sg13g2_mux2_1 _8184_ (.A0(_2964_),
    .A1(_2982_),
    .S(_2978_),
    .X(_2984_));
 sg13g2_a22oi_1 _8185_ (.Y(_2985_),
    .B1(_2984_),
    .B2(_2874_),
    .A2(_2981_),
    .A1(_2979_));
 sg13g2_or3_1 _8186_ (.A(_2964_),
    .B(_2968_),
    .C(_2978_),
    .X(_2986_));
 sg13g2_o21ai_1 _8187_ (.B1(_2986_),
    .Y(_2987_),
    .A1(net41),
    .A2(_2985_));
 sg13g2_nor3_2 _8188_ (.A(_2964_),
    .B(net41),
    .C(net67),
    .Y(_2988_));
 sg13g2_a21o_1 _8189_ (.A2(_2988_),
    .A1(net16),
    .B1(_2913_),
    .X(_2989_));
 sg13g2_nor3_1 _8190_ (.A(_0232_),
    .B(net41),
    .C(net106),
    .Y(_2990_));
 sg13g2_o21ai_1 _8191_ (.B1(_2990_),
    .Y(_2991_),
    .A1(net16),
    .A2(_2988_));
 sg13g2_a21oi_1 _8192_ (.A1(_2989_),
    .A2(_2991_),
    .Y(_2992_),
    .B1(net131));
 sg13g2_or4_1 _8193_ (.A(_0232_),
    .B(_2956_),
    .C(_2966_),
    .D(_2988_),
    .X(_2993_));
 sg13g2_nand4_1 _8194_ (.B(net16),
    .C(net68),
    .A(_0232_),
    .Y(_2995_),
    .D(_2988_));
 sg13g2_xnor2_1 _8195_ (.Y(_2996_),
    .A(net267),
    .B(_2829_));
 sg13g2_buf_2 _8196_ (.A(_2996_),
    .X(_2997_));
 sg13g2_a21oi_1 _8197_ (.A1(_2993_),
    .A2(_2995_),
    .Y(_2998_),
    .B1(_2997_));
 sg13g2_or2_1 _8198_ (.X(_2999_),
    .B(_2988_),
    .A(net16));
 sg13g2_a21oi_1 _8199_ (.A1(_2989_),
    .A2(_2999_),
    .Y(_3000_),
    .B1(net68));
 sg13g2_nand4_1 _8200_ (.B(net16),
    .C(net131),
    .A(_2913_),
    .Y(_3001_),
    .D(net68));
 sg13g2_nand2b_1 _8201_ (.Y(_3002_),
    .B(_2997_),
    .A_N(net16));
 sg13g2_a21oi_1 _8202_ (.A1(_3001_),
    .A2(_3002_),
    .Y(_3003_),
    .B1(net42));
 sg13g2_or4_1 _8203_ (.A(_2992_),
    .B(_2998_),
    .C(_3000_),
    .D(_3003_),
    .X(_3004_));
 sg13g2_nand2_1 _8204_ (.Y(_3005_),
    .A(net101),
    .B(_4244_));
 sg13g2_inv_1 _8205_ (.Y(_3006_),
    .A(_3005_));
 sg13g2_a21oi_1 _8206_ (.A1(net67),
    .A2(_2889_),
    .Y(_3007_),
    .B1(_2997_));
 sg13g2_nand3_1 _8207_ (.B(_2881_),
    .C(_3007_),
    .A(net41),
    .Y(_3008_));
 sg13g2_o21ai_1 _8208_ (.B1(_3007_),
    .Y(_3009_),
    .A1(_2962_),
    .A2(_2881_));
 sg13g2_nand2_1 _8209_ (.Y(_3010_),
    .A(net42),
    .B(_3009_));
 sg13g2_nand2_1 _8210_ (.Y(_3011_),
    .A(_3008_),
    .B(_3010_));
 sg13g2_xnor2_1 _8211_ (.Y(_3012_),
    .A(_3006_),
    .B(_3011_));
 sg13g2_xnor2_1 _8212_ (.Y(_3013_),
    .A(_3004_),
    .B(_3012_));
 sg13g2_xnor2_1 _8213_ (.Y(_3014_),
    .A(_2987_),
    .B(_3013_));
 sg13g2_a21oi_1 _8214_ (.A1(_0166_),
    .A2(_2940_),
    .Y(_3016_),
    .B1(_2933_));
 sg13g2_nor2_1 _8215_ (.A(_2919_),
    .B(_3016_),
    .Y(_3017_));
 sg13g2_xnor2_1 _8216_ (.Y(_3018_),
    .A(net65),
    .B(_2902_));
 sg13g2_a221oi_1 _8217_ (.B2(_2931_),
    .C1(_2929_),
    .B1(_3018_),
    .A1(_2919_),
    .Y(_3019_),
    .A2(_3016_));
 sg13g2_nor2_1 _8218_ (.A(_3017_),
    .B(_3019_),
    .Y(_3020_));
 sg13g2_nor2_1 _8219_ (.A(_3014_),
    .B(_3020_),
    .Y(_3021_));
 sg13g2_nand2_1 _8220_ (.Y(_3022_),
    .A(_3014_),
    .B(_3020_));
 sg13g2_o21ai_1 _8221_ (.B1(_3022_),
    .Y(_3023_),
    .A1(_2973_),
    .A2(_3021_));
 sg13g2_buf_1 _8222_ (.A(_3023_),
    .X(_3024_));
 sg13g2_xnor2_1 _8223_ (.Y(_3025_),
    .A(_2970_),
    .B(_2912_));
 sg13g2_xor2_1 _8224_ (.B(_3025_),
    .A(_2948_),
    .X(_3027_));
 sg13g2_mux2_1 _8225_ (.A0(_2848_),
    .A1(_2849_),
    .S(_2841_),
    .X(_3028_));
 sg13g2_buf_1 _8226_ (.A(_3028_),
    .X(_3029_));
 sg13g2_o21ai_1 _8227_ (.B1(net65),
    .Y(_3030_),
    .A1(net102),
    .A2(net105));
 sg13g2_nand2_1 _8228_ (.Y(_3031_),
    .A(net143),
    .B(_3030_));
 sg13g2_o21ai_1 _8229_ (.B1(net50),
    .Y(_3032_),
    .A1(_4201_),
    .A2(net71));
 sg13g2_nand2_1 _8230_ (.Y(_3033_),
    .A(_4201_),
    .B(_2853_));
 sg13g2_nand3_1 _8231_ (.B(_3032_),
    .C(_3033_),
    .A(net101),
    .Y(_3034_));
 sg13g2_and3_1 _8232_ (.X(_3035_),
    .A(net82),
    .B(_3031_),
    .C(_3034_));
 sg13g2_nand2_1 _8233_ (.Y(_3036_),
    .A(net146),
    .B(_0202_));
 sg13g2_and3_1 _8234_ (.X(_3038_),
    .A(net49),
    .B(_3036_),
    .C(net105));
 sg13g2_buf_1 _8235_ (.A(_3038_),
    .X(_3039_));
 sg13g2_nor2_1 _8236_ (.A(_2892_),
    .B(net106),
    .Y(_3040_));
 sg13g2_buf_2 _8237_ (.A(_3040_),
    .X(_3041_));
 sg13g2_o21ai_1 _8238_ (.B1(_3041_),
    .Y(_3042_),
    .A1(_3035_),
    .A2(_3039_));
 sg13g2_buf_1 _8239_ (.A(_3042_),
    .X(_3043_));
 sg13g2_nand3_1 _8240_ (.B(_3031_),
    .C(_3034_),
    .A(net82),
    .Y(_3044_));
 sg13g2_inv_1 _8241_ (.Y(_3045_),
    .A(_3039_));
 sg13g2_nand3_1 _8242_ (.B(_3044_),
    .C(_3045_),
    .A(_2881_),
    .Y(_3046_));
 sg13g2_buf_1 _8243_ (.A(_3046_),
    .X(_3047_));
 sg13g2_xor2_1 _8244_ (.B(_0424_),
    .A(net98),
    .X(_3049_));
 sg13g2_nand2_1 _8245_ (.Y(_3050_),
    .A(net274),
    .B(_2878_));
 sg13g2_nor2_1 _8246_ (.A(net284),
    .B(_3601_),
    .Y(_3051_));
 sg13g2_a21oi_1 _8247_ (.A1(net284),
    .A2(_1611_),
    .Y(_3052_),
    .B1(_2803_));
 sg13g2_o21ai_1 _8248_ (.B1(_0911_),
    .Y(_3053_),
    .A1(_3051_),
    .A2(_3052_));
 sg13g2_nand2_1 _8249_ (.Y(_3054_),
    .A(_1358_),
    .B(_1281_));
 sg13g2_a21o_1 _8250_ (.A2(_2484_),
    .A1(_3054_),
    .B1(_2868_),
    .X(_3055_));
 sg13g2_a21oi_1 _8251_ (.A1(_3053_),
    .A2(_3055_),
    .Y(_3056_),
    .B1(_4555_));
 sg13g2_buf_1 _8252_ (.A(_3056_),
    .X(_3057_));
 sg13g2_a21oi_1 _8253_ (.A1(net223),
    .A2(net103),
    .Y(_3058_),
    .B1(_3057_));
 sg13g2_nand3_1 _8254_ (.B(net103),
    .C(_3057_),
    .A(net223),
    .Y(_3060_));
 sg13g2_o21ai_1 _8255_ (.B1(_3060_),
    .Y(_3061_),
    .A1(_3050_),
    .A2(_3058_));
 sg13g2_nand3_1 _8256_ (.B(net240),
    .C(_2868_),
    .A(net199),
    .Y(_3062_));
 sg13g2_a21o_1 _8257_ (.A2(_2868_),
    .A1(net240),
    .B1(net199),
    .X(_3063_));
 sg13g2_a21oi_1 _8258_ (.A1(_3062_),
    .A2(_3063_),
    .Y(_3064_),
    .B1(net204));
 sg13g2_xnor2_1 _8259_ (.Y(_3065_),
    .A(_0432_),
    .B(_3064_));
 sg13g2_xnor2_1 _8260_ (.Y(_3066_),
    .A(net105),
    .B(_3065_));
 sg13g2_a21o_1 _8261_ (.A2(_3061_),
    .A1(_3049_),
    .B1(_3066_),
    .X(_3067_));
 sg13g2_o21ai_1 _8262_ (.B1(_3067_),
    .Y(_3068_),
    .A1(_3049_),
    .A2(_3061_));
 sg13g2_nand3_1 _8263_ (.B(_3047_),
    .C(_3068_),
    .A(_3043_),
    .Y(_3069_));
 sg13g2_a21oi_1 _8264_ (.A1(_3044_),
    .A2(_3045_),
    .Y(_3071_),
    .B1(_2881_));
 sg13g2_nor3_1 _8265_ (.A(_3041_),
    .B(_3035_),
    .C(_3039_),
    .Y(_3072_));
 sg13g2_o21ai_1 _8266_ (.B1(_3068_),
    .Y(_3073_),
    .A1(_3071_),
    .A2(_3072_));
 sg13g2_mux2_1 _8267_ (.A0(net106),
    .A1(net105),
    .S(_2892_),
    .X(_3074_));
 sg13g2_nand2b_1 _8268_ (.Y(_3075_),
    .B(_3074_),
    .A_N(net26));
 sg13g2_nand4_1 _8269_ (.B(net107),
    .C(net71),
    .A(_2874_),
    .Y(_3076_),
    .D(_2865_));
 sg13g2_a21oi_1 _8270_ (.A1(_3075_),
    .A2(_3076_),
    .Y(_3077_),
    .B1(net122));
 sg13g2_and3_1 _8271_ (.X(_3078_),
    .A(net122),
    .B(_3075_),
    .C(_3076_));
 sg13g2_buf_1 _8272_ (.A(_3078_),
    .X(_3079_));
 sg13g2_nor2_1 _8273_ (.A(_3077_),
    .B(_3079_),
    .Y(_3080_));
 sg13g2_nor2b_1 _8274_ (.A(_2958_),
    .B_N(_2959_),
    .Y(_3082_));
 sg13g2_nor2_1 _8275_ (.A(_3082_),
    .B(_2892_),
    .Y(_3083_));
 sg13g2_nand2b_1 _8276_ (.Y(_3084_),
    .B(net106),
    .A_N(_0432_));
 sg13g2_o21ai_1 _8277_ (.B1(_3084_),
    .Y(_3085_),
    .A1(_2853_),
    .A2(_2865_));
 sg13g2_o21ai_1 _8278_ (.B1(_0432_),
    .Y(_3086_),
    .A1(net105),
    .A2(_3064_));
 sg13g2_nand3_1 _8279_ (.B(_2874_),
    .C(_2853_),
    .A(_2962_),
    .Y(_3087_));
 sg13g2_nand2_1 _8280_ (.Y(_3088_),
    .A(_3086_),
    .B(_3087_));
 sg13g2_nor4_1 _8281_ (.A(_0432_),
    .B(_2874_),
    .C(net105),
    .D(net26),
    .Y(_3089_));
 sg13g2_a221oi_1 _8282_ (.B2(net26),
    .C1(_3089_),
    .B1(_3088_),
    .A1(_3083_),
    .Y(_3090_),
    .A2(_3085_));
 sg13g2_buf_1 _8283_ (.A(_3090_),
    .X(_3091_));
 sg13g2_nor2_1 _8284_ (.A(net103),
    .B(net99),
    .Y(_3093_));
 sg13g2_nor4_1 _8285_ (.A(net195),
    .B(net142),
    .C(_2861_),
    .D(_2863_),
    .Y(_3094_));
 sg13g2_o21ai_1 _8286_ (.B1(_0432_),
    .Y(_3095_),
    .A1(_3093_),
    .A2(_3094_));
 sg13g2_nor2_1 _8287_ (.A(_1457_),
    .B(net104),
    .Y(_3096_));
 sg13g2_a221oi_1 _8288_ (.B2(_3096_),
    .C1(_2125_),
    .B1(_2866_),
    .A1(net275),
    .Y(_3097_),
    .A2(_3036_));
 sg13g2_mux2_1 _8289_ (.A0(_0149_),
    .A1(_4286_),
    .S(net26),
    .X(_3098_));
 sg13g2_a22oi_1 _8290_ (.Y(_3099_),
    .B1(_3098_),
    .B2(_3093_),
    .A2(_3097_),
    .A1(_3095_));
 sg13g2_xnor2_1 _8291_ (.Y(_3100_),
    .A(_3091_),
    .B(_3099_));
 sg13g2_xnor2_1 _8292_ (.Y(_3101_),
    .A(_3080_),
    .B(_3100_));
 sg13g2_mux2_1 _8293_ (.A0(_3069_),
    .A1(_3073_),
    .S(_3101_),
    .X(_3102_));
 sg13g2_a21oi_1 _8294_ (.A1(_3043_),
    .A2(_3047_),
    .Y(_3103_),
    .B1(net69));
 sg13g2_nand2b_1 _8295_ (.Y(_3104_),
    .B(_3103_),
    .A_N(_3101_));
 sg13g2_nand4_1 _8296_ (.B(_3101_),
    .C(_3043_),
    .A(net69),
    .Y(_3105_),
    .D(_3047_));
 sg13g2_and3_1 _8297_ (.X(_3106_),
    .A(_3102_),
    .B(_3104_),
    .C(_3105_));
 sg13g2_buf_1 _8298_ (.A(_3106_),
    .X(_3107_));
 sg13g2_nor3_1 _8299_ (.A(_3077_),
    .B(_3079_),
    .C(_3091_),
    .Y(_3108_));
 sg13g2_xnor2_1 _8300_ (.Y(_3109_),
    .A(net69),
    .B(_3099_));
 sg13g2_o21ai_1 _8301_ (.B1(_3091_),
    .Y(_3110_),
    .A1(_3077_),
    .A2(_3079_));
 sg13g2_o21ai_1 _8302_ (.B1(_3110_),
    .Y(_3111_),
    .A1(_3108_),
    .A2(_3109_));
 sg13g2_buf_1 _8303_ (.A(_3111_),
    .X(_3112_));
 sg13g2_a21oi_1 _8304_ (.A1(_0411_),
    .A2(_0413_),
    .Y(_3114_),
    .B1(_2903_));
 sg13g2_and3_1 _8305_ (.X(_3115_),
    .A(_2903_),
    .B(_0411_),
    .C(_0413_));
 sg13g2_nand2_1 _8306_ (.Y(_3116_),
    .A(_2976_),
    .B(net26));
 sg13g2_o21ai_1 _8307_ (.B1(_3116_),
    .Y(_3117_),
    .A1(_3114_),
    .A2(_3115_));
 sg13g2_nand2b_1 _8308_ (.Y(_3118_),
    .B(net98),
    .A_N(_2866_));
 sg13g2_inv_1 _8309_ (.Y(_3119_),
    .A(_0432_));
 sg13g2_a21oi_2 _8310_ (.B1(_3119_),
    .Y(_3120_),
    .A2(_3118_),
    .A1(_3117_));
 sg13g2_nor3_1 _8311_ (.A(net143),
    .B(net99),
    .C(net67),
    .Y(_3121_));
 sg13g2_nor2_1 _8312_ (.A(net69),
    .B(_3121_),
    .Y(_3122_));
 sg13g2_a21oi_1 _8313_ (.A1(_3036_),
    .A2(net67),
    .Y(_3123_),
    .B1(_3122_));
 sg13g2_nor2_1 _8314_ (.A(_2907_),
    .B(_2879_),
    .Y(_3125_));
 sg13g2_a21oi_1 _8315_ (.A1(_2879_),
    .A2(_3123_),
    .Y(_3126_),
    .B1(_3125_));
 sg13g2_xnor2_1 _8316_ (.Y(_3127_),
    .A(_3120_),
    .B(_3126_));
 sg13g2_xnor2_1 _8317_ (.Y(_3128_),
    .A(net70),
    .B(_2882_));
 sg13g2_a21oi_1 _8318_ (.A1(_2890_),
    .A2(_2893_),
    .Y(_3129_),
    .B1(_2845_));
 sg13g2_a221oi_1 _8319_ (.B2(net122),
    .C1(_3129_),
    .B1(_3128_),
    .A1(_2894_),
    .Y(_3130_),
    .A2(_2898_));
 sg13g2_xnor2_1 _8320_ (.Y(_3131_),
    .A(_2910_),
    .B(_3130_));
 sg13g2_xor2_1 _8321_ (.B(_3131_),
    .A(_3127_),
    .X(_3132_));
 sg13g2_xnor2_1 _8322_ (.Y(_3133_),
    .A(_3112_),
    .B(_3132_));
 sg13g2_nor2_1 _8323_ (.A(_2976_),
    .B(_2881_),
    .Y(_3134_));
 sg13g2_nor4_1 _8324_ (.A(_4214_),
    .B(net99),
    .C(_3041_),
    .D(net71),
    .Y(_3136_));
 sg13g2_o21ai_1 _8325_ (.B1(net101),
    .Y(_3137_),
    .A1(_3134_),
    .A2(_3136_));
 sg13g2_xnor2_1 _8326_ (.Y(_3138_),
    .A(net64),
    .B(_3041_));
 sg13g2_nand3_1 _8327_ (.B(net105),
    .C(_3138_),
    .A(net99),
    .Y(_3139_));
 sg13g2_a21oi_1 _8328_ (.A1(_3137_),
    .A2(_3139_),
    .Y(_3140_),
    .B1(net50));
 sg13g2_nor2_1 _8329_ (.A(net65),
    .B(_2854_),
    .Y(_3141_));
 sg13g2_mux2_1 _8330_ (.A0(net98),
    .A1(_3141_),
    .S(_3041_),
    .X(_3142_));
 sg13g2_nand2_1 _8331_ (.Y(_3143_),
    .A(net98),
    .B(_3029_));
 sg13g2_nor2_1 _8332_ (.A(net49),
    .B(_3143_),
    .Y(_3144_));
 sg13g2_a22oi_1 _8333_ (.Y(_3145_),
    .B1(_3144_),
    .B2(_3041_),
    .A2(_3142_),
    .A1(net49));
 sg13g2_a21oi_1 _8334_ (.A1(_2881_),
    .A2(_3144_),
    .Y(_3147_),
    .B1(net143));
 sg13g2_a21oi_1 _8335_ (.A1(net113),
    .A2(_3145_),
    .Y(_3148_),
    .B1(_3147_));
 sg13g2_nor2_2 _8336_ (.A(_3140_),
    .B(_3148_),
    .Y(_3149_));
 sg13g2_inv_1 _8337_ (.Y(_3150_),
    .A(_3149_));
 sg13g2_o21ai_1 _8338_ (.B1(_3150_),
    .Y(_3151_),
    .A1(_3107_),
    .A2(_3133_));
 sg13g2_nand2_1 _8339_ (.Y(_3152_),
    .A(_3107_),
    .B(_3133_));
 sg13g2_and2_1 _8340_ (.A(_3151_),
    .B(_3152_),
    .X(_3153_));
 sg13g2_buf_2 _8341_ (.A(_3153_),
    .X(_3154_));
 sg13g2_nor2_1 _8342_ (.A(_3027_),
    .B(_3154_),
    .Y(_3155_));
 sg13g2_or2_1 _8343_ (.X(_3156_),
    .B(_3057_),
    .A(net71));
 sg13g2_o21ai_1 _8344_ (.B1(_3156_),
    .Y(_3158_),
    .A1(net106),
    .A2(_3060_));
 sg13g2_and3_1 _8345_ (.X(_3159_),
    .A(net274),
    .B(_2962_),
    .C(_3057_));
 sg13g2_nand3b_1 _8346_ (.B(net223),
    .C(net65),
    .Y(_3160_),
    .A_N(_3057_));
 sg13g2_a21oi_1 _8347_ (.A1(net274),
    .A2(net107),
    .Y(_3161_),
    .B1(_3160_));
 sg13g2_a221oi_1 _8348_ (.B2(net106),
    .C1(_3161_),
    .B1(_3159_),
    .A1(net238),
    .Y(_3162_),
    .A2(_3158_));
 sg13g2_buf_2 _8349_ (.A(_3162_),
    .X(_3163_));
 sg13g2_xnor2_1 _8350_ (.Y(_3164_),
    .A(_3049_),
    .B(_3065_));
 sg13g2_xnor2_1 _8351_ (.Y(_3165_),
    .A(_3061_),
    .B(_3164_));
 sg13g2_buf_2 _8352_ (.A(_3165_),
    .X(_3166_));
 sg13g2_nor2_1 _8353_ (.A(_2056_),
    .B(_3093_),
    .Y(_3167_));
 sg13g2_xor2_1 _8354_ (.B(_3167_),
    .A(_3166_),
    .X(_3169_));
 sg13g2_xnor2_1 _8355_ (.Y(_3170_),
    .A(_3163_),
    .B(_3169_));
 sg13g2_o21ai_1 _8356_ (.B1(net238),
    .Y(_3171_),
    .A1(_2962_),
    .A2(net107));
 sg13g2_o21ai_1 _8357_ (.B1(_3171_),
    .Y(_3172_),
    .A1(net194),
    .A2(_0625_));
 sg13g2_o21ai_1 _8358_ (.B1(_3172_),
    .Y(_3173_),
    .A1(_3082_),
    .A2(_3050_));
 sg13g2_xor2_1 _8359_ (.B(_3173_),
    .A(_3057_),
    .X(_3174_));
 sg13g2_a21oi_1 _8360_ (.A1(_4110_),
    .A2(net49),
    .Y(_3175_),
    .B1(_2056_));
 sg13g2_nor2_1 _8361_ (.A(net190),
    .B(net194),
    .Y(_3176_));
 sg13g2_a22oi_1 _8362_ (.Y(_3177_),
    .B1(_3176_),
    .B2(net82),
    .A2(_3175_),
    .A1(net190));
 sg13g2_or2_1 _8363_ (.X(_3178_),
    .B(_3177_),
    .A(_3174_));
 sg13g2_a21o_1 _8364_ (.A2(_3178_),
    .A1(_3170_),
    .B1(_0495_),
    .X(_3180_));
 sg13g2_nand2_1 _8365_ (.Y(_3181_),
    .A(_3174_),
    .B(_3177_));
 sg13g2_nand2b_1 _8366_ (.Y(_3182_),
    .B(_3181_),
    .A_N(_3170_));
 sg13g2_nand2_1 _8367_ (.Y(_3183_),
    .A(net163),
    .B(_2916_));
 sg13g2_a21oi_1 _8368_ (.A1(_3180_),
    .A2(_3182_),
    .Y(_3184_),
    .B1(_3183_));
 sg13g2_nand2b_1 _8369_ (.Y(_3185_),
    .B(_3181_),
    .A_N(_0495_));
 sg13g2_a21oi_1 _8370_ (.A1(_3178_),
    .A2(_3185_),
    .Y(_3186_),
    .B1(_3170_));
 sg13g2_nor2_1 _8371_ (.A(_3184_),
    .B(_3186_),
    .Y(_3187_));
 sg13g2_a21o_1 _8372_ (.A2(_3047_),
    .A1(_3043_),
    .B1(_3068_),
    .X(_3188_));
 sg13g2_a21oi_1 _8373_ (.A1(_3069_),
    .A2(_3188_),
    .Y(_3189_),
    .B1(_3101_));
 sg13g2_and3_1 _8374_ (.X(_3191_),
    .A(_3101_),
    .B(_3069_),
    .C(_3188_));
 sg13g2_or2_1 _8375_ (.X(_3192_),
    .B(_3191_),
    .A(_3189_));
 sg13g2_nor2_1 _8376_ (.A(net32),
    .B(net71),
    .Y(_3193_));
 sg13g2_nor2_1 _8377_ (.A(_3033_),
    .B(_3166_),
    .Y(_3194_));
 sg13g2_a21oi_1 _8378_ (.A1(_3193_),
    .A2(_3166_),
    .Y(_3195_),
    .B1(_3194_));
 sg13g2_nor4_1 _8379_ (.A(net50),
    .B(net99),
    .C(_3163_),
    .D(_3195_),
    .Y(_3196_));
 sg13g2_nand2_1 _8380_ (.Y(_3197_),
    .A(_3192_),
    .B(_3196_));
 sg13g2_nor2_1 _8381_ (.A(_3187_),
    .B(_3197_),
    .Y(_3198_));
 sg13g2_mux2_1 _8382_ (.A0(_3163_),
    .A1(net71),
    .S(_3166_),
    .X(_3199_));
 sg13g2_mux2_1 _8383_ (.A0(_3029_),
    .A1(_3163_),
    .S(_3166_),
    .X(_3200_));
 sg13g2_mux2_1 _8384_ (.A0(_3199_),
    .A1(_3200_),
    .S(net49),
    .X(_3202_));
 sg13g2_nor2b_1 _8385_ (.A(_3163_),
    .B_N(_3166_),
    .Y(_3203_));
 sg13g2_inv_1 _8386_ (.Y(_3204_),
    .A(_3033_));
 sg13g2_o21ai_1 _8387_ (.B1(_3204_),
    .Y(_3205_),
    .A1(_3163_),
    .A2(_3166_));
 sg13g2_o21ai_1 _8388_ (.B1(_3205_),
    .Y(_3206_),
    .A1(_3143_),
    .A2(_3203_));
 sg13g2_nor2_1 _8389_ (.A(net64),
    .B(net105),
    .Y(_3207_));
 sg13g2_mux2_1 _8390_ (.A0(_3141_),
    .A1(_3207_),
    .S(_3166_),
    .X(_3208_));
 sg13g2_and2_1 _8391_ (.A(_3163_),
    .B(_3208_),
    .X(_3209_));
 sg13g2_a221oi_1 _8392_ (.B2(net50),
    .C1(_3209_),
    .B1(_3206_),
    .A1(net99),
    .Y(_3210_),
    .A2(_3202_));
 sg13g2_or3_1 _8393_ (.A(_3189_),
    .B(_3191_),
    .C(_3210_),
    .X(_3211_));
 sg13g2_o21ai_1 _8394_ (.B1(_3211_),
    .Y(_3213_),
    .A1(_3184_),
    .A2(_3186_));
 sg13g2_a21oi_1 _8395_ (.A1(_3192_),
    .A2(_3210_),
    .Y(_3214_),
    .B1(_3196_));
 sg13g2_or2_1 _8396_ (.X(_3215_),
    .B(_3149_),
    .A(_3112_));
 sg13g2_nand2_1 _8397_ (.Y(_3216_),
    .A(_3112_),
    .B(_3149_));
 sg13g2_a21oi_1 _8398_ (.A1(_3215_),
    .A2(_3216_),
    .Y(_3217_),
    .B1(_3132_));
 sg13g2_nand2b_1 _8399_ (.Y(_3218_),
    .B(_3112_),
    .A_N(_3149_));
 sg13g2_nand2b_1 _8400_ (.Y(_3219_),
    .B(_3149_),
    .A_N(_3112_));
 sg13g2_xnor2_1 _8401_ (.Y(_3220_),
    .A(_3127_),
    .B(_3131_));
 sg13g2_a21oi_1 _8402_ (.A1(_3218_),
    .A2(_3219_),
    .Y(_3221_),
    .B1(_3220_));
 sg13g2_o21ai_1 _8403_ (.B1(_3107_),
    .Y(_3222_),
    .A1(_3217_),
    .A2(_3221_));
 sg13g2_or3_1 _8404_ (.A(_3107_),
    .B(_3217_),
    .C(_3221_),
    .X(_3223_));
 sg13g2_a22oi_1 _8405_ (.Y(_3224_),
    .B1(_3222_),
    .B2(_3223_),
    .A2(_3214_),
    .A1(_3213_));
 sg13g2_buf_1 _8406_ (.A(_3224_),
    .X(_3225_));
 sg13g2_or2_1 _8407_ (.X(_3226_),
    .B(_3225_),
    .A(_3198_));
 sg13g2_buf_2 _8408_ (.A(_3226_),
    .X(_3227_));
 sg13g2_xnor2_1 _8409_ (.Y(_3228_),
    .A(_2948_),
    .B(_3025_));
 sg13g2_nand2_1 _8410_ (.Y(_3229_),
    .A(_3151_),
    .B(_3152_));
 sg13g2_or4_1 _8411_ (.A(_3228_),
    .B(_3229_),
    .C(_3198_),
    .D(_3225_),
    .X(_3230_));
 sg13g2_xnor2_1 _8412_ (.Y(_3231_),
    .A(_3014_),
    .B(_3020_));
 sg13g2_xnor2_1 _8413_ (.Y(_3232_),
    .A(_2973_),
    .B(_3231_));
 sg13g2_buf_2 _8414_ (.A(_3232_),
    .X(_3234_));
 sg13g2_inv_1 _8415_ (.Y(_3235_),
    .A(_3234_));
 sg13g2_a22oi_1 _8416_ (.Y(_3236_),
    .B1(_3230_),
    .B2(_3235_),
    .A2(_3227_),
    .A1(_3155_));
 sg13g2_nand2_1 _8417_ (.Y(_3237_),
    .A(_2907_),
    .B(_3120_));
 sg13g2_xnor2_1 _8418_ (.Y(_3238_),
    .A(net68),
    .B(_2902_));
 sg13g2_o21ai_1 _8419_ (.B1(_3238_),
    .Y(_3239_),
    .A1(_2907_),
    .A2(_3120_));
 sg13g2_nor2_1 _8420_ (.A(_2904_),
    .B(_2881_),
    .Y(_3240_));
 sg13g2_o21ai_1 _8421_ (.B1(_3240_),
    .Y(_3241_),
    .A1(_2902_),
    .A2(_3120_));
 sg13g2_nand3_1 _8422_ (.B(_3239_),
    .C(_3241_),
    .A(_3237_),
    .Y(_3242_));
 sg13g2_buf_1 _8423_ (.A(_3242_),
    .X(_3243_));
 sg13g2_and2_1 _8424_ (.A(_2902_),
    .B(_3127_),
    .X(_3245_));
 sg13g2_nor3_1 _8425_ (.A(_2902_),
    .B(_3127_),
    .C(_3131_),
    .Y(_3246_));
 sg13g2_a221oi_1 _8426_ (.B2(_3131_),
    .C1(_3246_),
    .B1(_3245_),
    .A1(_3112_),
    .Y(_3247_),
    .A2(_3132_));
 sg13g2_buf_1 _8427_ (.A(_3247_),
    .X(_3248_));
 sg13g2_nor2_1 _8428_ (.A(_3243_),
    .B(_3248_),
    .Y(_3249_));
 sg13g2_nand2_1 _8429_ (.Y(_3250_),
    .A(_3243_),
    .B(_3248_));
 sg13g2_nand2_1 _8430_ (.Y(_3251_),
    .A(_3234_),
    .B(_3250_));
 sg13g2_a22oi_1 _8431_ (.Y(_3252_),
    .B1(_3027_),
    .B2(_3154_),
    .A2(_3250_),
    .A1(_3234_));
 sg13g2_nor2_1 _8432_ (.A(_3234_),
    .B(_3250_),
    .Y(_3253_));
 sg13g2_a221oi_1 _8433_ (.B2(_3252_),
    .C1(_3253_),
    .B1(_3227_),
    .A1(_3251_),
    .Y(_3254_),
    .A2(_3155_));
 sg13g2_o21ai_1 _8434_ (.B1(_3254_),
    .Y(_3256_),
    .A1(_3236_),
    .A2(_3249_));
 sg13g2_buf_1 _8435_ (.A(_3256_),
    .X(_3257_));
 sg13g2_or2_1 _8436_ (.X(_3258_),
    .B(_3257_),
    .A(_3024_));
 sg13g2_inv_1 _8437_ (.Y(_3259_),
    .A(_3004_));
 sg13g2_nor2_1 _8438_ (.A(_2987_),
    .B(_3259_),
    .Y(_3260_));
 sg13g2_nor2_1 _8439_ (.A(_3012_),
    .B(_3260_),
    .Y(_3261_));
 sg13g2_a21oi_1 _8440_ (.A1(_2987_),
    .A2(_3259_),
    .Y(_3262_),
    .B1(_3261_));
 sg13g2_nor2_2 _8441_ (.A(_2997_),
    .B(_2918_),
    .Y(_3263_));
 sg13g2_o21ai_1 _8442_ (.B1(_3263_),
    .Y(_3264_),
    .A1(_3082_),
    .A2(_3006_));
 sg13g2_o21ai_1 _8443_ (.B1(_2997_),
    .Y(_3265_),
    .A1(net41),
    .A2(_3005_));
 sg13g2_nor2_1 _8444_ (.A(net67),
    .B(_3005_),
    .Y(_3267_));
 sg13g2_nor3_1 _8445_ (.A(net42),
    .B(net68),
    .C(_3267_),
    .Y(_3268_));
 sg13g2_a21oi_1 _8446_ (.A1(_2967_),
    .A2(_3005_),
    .Y(_3269_),
    .B1(_3268_));
 sg13g2_nand3_1 _8447_ (.B(_3265_),
    .C(_3269_),
    .A(_3264_),
    .Y(_3270_));
 sg13g2_buf_1 _8448_ (.A(_3270_),
    .X(_3271_));
 sg13g2_o21ai_1 _8449_ (.B1(_3263_),
    .Y(_3272_),
    .A1(net113),
    .A2(_2967_));
 sg13g2_nand3_1 _8450_ (.B(net63),
    .C(_3263_),
    .A(net65),
    .Y(_3273_));
 sg13g2_o21ai_1 _8451_ (.B1(_3273_),
    .Y(_3274_),
    .A1(net63),
    .A2(_3263_));
 sg13g2_a21oi_1 _8452_ (.A1(net65),
    .A2(_3263_),
    .Y(_3275_),
    .B1(net63));
 sg13g2_nor3_1 _8453_ (.A(net125),
    .B(_2997_),
    .C(_2918_),
    .Y(_3276_));
 sg13g2_nor3_1 _8454_ (.A(net113),
    .B(_3275_),
    .C(_3276_),
    .Y(_3278_));
 sg13g2_a221oi_1 _8455_ (.B2(net113),
    .C1(_3278_),
    .B1(_3274_),
    .A1(net32),
    .Y(_3279_),
    .A2(_3272_));
 sg13g2_xnor2_1 _8456_ (.Y(_3280_),
    .A(_3271_),
    .B(_3279_));
 sg13g2_o21ai_1 _8457_ (.B1(net131),
    .Y(_3281_),
    .A1(net16),
    .A2(net42));
 sg13g2_nand2_1 _8458_ (.Y(_3282_),
    .A(_2957_),
    .B(net42));
 sg13g2_a21oi_1 _8459_ (.A1(_3281_),
    .A2(_3282_),
    .Y(_3283_),
    .B1(_0232_));
 sg13g2_a22oi_1 _8460_ (.Y(_3284_),
    .B1(net42),
    .B2(_2913_),
    .A2(net131),
    .A1(_2957_));
 sg13g2_nor2b_1 _8461_ (.A(_3284_),
    .B_N(_2988_),
    .Y(_3285_));
 sg13g2_o21ai_1 _8462_ (.B1(net68),
    .Y(_3286_),
    .A1(_3283_),
    .A2(_3285_));
 sg13g2_nand2b_1 _8463_ (.Y(_3287_),
    .B(_3286_),
    .A_N(_3280_));
 sg13g2_nand2b_1 _8464_ (.Y(_3289_),
    .B(_3280_),
    .A_N(_3286_));
 sg13g2_nand2_1 _8465_ (.Y(_3290_),
    .A(_3287_),
    .B(_3289_));
 sg13g2_xor2_1 _8466_ (.B(_3290_),
    .A(_3262_),
    .X(_3291_));
 sg13g2_buf_2 _8467_ (.A(_3291_),
    .X(_3292_));
 sg13g2_a21o_1 _8468_ (.A2(_3257_),
    .A1(_3024_),
    .B1(_3292_),
    .X(_3293_));
 sg13g2_inv_1 _8469_ (.Y(_3294_),
    .A(_3287_));
 sg13g2_o21ai_1 _8470_ (.B1(_3289_),
    .Y(_3295_),
    .A1(_3262_),
    .A2(_3294_));
 sg13g2_buf_1 _8471_ (.A(_3295_),
    .X(_3296_));
 sg13g2_o21ai_1 _8472_ (.B1(_3274_),
    .Y(_3297_),
    .A1(net113),
    .A2(_3271_));
 sg13g2_nand2_1 _8473_ (.Y(_3298_),
    .A(_2874_),
    .B(_3263_));
 sg13g2_a22oi_1 _8474_ (.Y(_3300_),
    .B1(_3298_),
    .B2(net32),
    .A2(_3271_),
    .A1(net113));
 sg13g2_and2_1 _8475_ (.A(_3297_),
    .B(_3300_),
    .X(_3301_));
 sg13g2_buf_1 _8476_ (.A(_3301_),
    .X(_3302_));
 sg13g2_nor2_1 _8477_ (.A(net32),
    .B(_2889_),
    .Y(_3303_));
 sg13g2_and2_1 _8478_ (.A(net42),
    .B(_3303_),
    .X(_3304_));
 sg13g2_nor2_1 _8479_ (.A(_2915_),
    .B(_3302_),
    .Y(_3305_));
 sg13g2_a21oi_1 _8480_ (.A1(_3302_),
    .A2(_3304_),
    .Y(_3306_),
    .B1(_3305_));
 sg13g2_o21ai_1 _8481_ (.B1(_2997_),
    .Y(_3307_),
    .A1(net101),
    .A2(_3302_));
 sg13g2_o21ai_1 _8482_ (.B1(_3307_),
    .Y(_3308_),
    .A1(net113),
    .A2(_3306_));
 sg13g2_o21ai_1 _8483_ (.B1(_2915_),
    .Y(_3309_),
    .A1(_3302_),
    .A2(_3303_));
 sg13g2_nand3_1 _8484_ (.B(net63),
    .C(_3309_),
    .A(net113),
    .Y(_3311_));
 sg13g2_o21ai_1 _8485_ (.B1(_3311_),
    .Y(_3312_),
    .A1(net63),
    .A2(_3305_));
 sg13g2_a22oi_1 _8486_ (.Y(_3313_),
    .B1(_3312_),
    .B2(net131),
    .A2(_3308_),
    .A1(net63));
 sg13g2_buf_1 _8487_ (.A(_3313_),
    .X(_3314_));
 sg13g2_a21oi_1 _8488_ (.A1(net63),
    .A2(_3303_),
    .Y(_3315_),
    .B1(net41));
 sg13g2_nor2_1 _8489_ (.A(_4283_),
    .B(_3315_),
    .Y(_3316_));
 sg13g2_o21ai_1 _8490_ (.B1(_2831_),
    .Y(_3317_),
    .A1(net41),
    .A2(_3303_));
 sg13g2_a22oi_1 _8491_ (.Y(_3318_),
    .B1(_3317_),
    .B2(_4283_),
    .A2(_3316_),
    .A1(_2831_));
 sg13g2_xnor2_1 _8492_ (.Y(_3319_),
    .A(_3302_),
    .B(_3318_));
 sg13g2_nand3_1 _8493_ (.B(_3314_),
    .C(_3319_),
    .A(_3296_),
    .Y(_3320_));
 sg13g2_or3_1 _8494_ (.A(_3296_),
    .B(_3314_),
    .C(_3319_),
    .X(_3322_));
 sg13g2_a22oi_1 _8495_ (.Y(_3323_),
    .B1(_3320_),
    .B2(_3322_),
    .A2(_3293_),
    .A1(_3258_));
 sg13g2_nand2_1 _8496_ (.Y(_3324_),
    .A(_3024_),
    .B(_3257_));
 sg13g2_o21ai_1 _8497_ (.B1(_3292_),
    .Y(_3325_),
    .A1(_3024_),
    .A2(_3257_));
 sg13g2_nand3b_1 _8498_ (.B(_3314_),
    .C(_3319_),
    .Y(_3326_),
    .A_N(_3296_));
 sg13g2_nand3b_1 _8499_ (.B(_3314_),
    .C(_3296_),
    .Y(_3327_),
    .A_N(_3319_));
 sg13g2_a22oi_1 _8500_ (.Y(_3328_),
    .B1(_3326_),
    .B2(_3327_),
    .A2(_3325_),
    .A1(_3324_));
 sg13g2_nand2b_1 _8501_ (.Y(_3329_),
    .B(_3027_),
    .A_N(_3243_));
 sg13g2_nand2_1 _8502_ (.Y(_3330_),
    .A(_3243_),
    .B(_3228_));
 sg13g2_mux2_1 _8503_ (.A0(_3329_),
    .A1(_3330_),
    .S(_2973_),
    .X(_3331_));
 sg13g2_nor2_1 _8504_ (.A(_3022_),
    .B(_3292_),
    .Y(_3332_));
 sg13g2_a21oi_1 _8505_ (.A1(_3021_),
    .A2(_3292_),
    .Y(_3333_),
    .B1(_3332_));
 sg13g2_inv_1 _8506_ (.Y(_3334_),
    .A(_3329_));
 sg13g2_nand3_1 _8507_ (.B(_3292_),
    .C(_3334_),
    .A(_2973_),
    .Y(_3335_));
 sg13g2_or3_1 _8508_ (.A(_2973_),
    .B(_3292_),
    .C(_3330_),
    .X(_3336_));
 sg13g2_a21o_1 _8509_ (.A2(_3336_),
    .A1(_3335_),
    .B1(_3231_),
    .X(_3337_));
 sg13g2_o21ai_1 _8510_ (.B1(_3337_),
    .Y(_3338_),
    .A1(_3331_),
    .A2(_3333_));
 sg13g2_inv_1 _8511_ (.Y(_3339_),
    .A(_3248_));
 sg13g2_xnor2_1 _8512_ (.Y(_3340_),
    .A(_3339_),
    .B(_3154_));
 sg13g2_nand3_1 _8513_ (.B(_3154_),
    .C(_3227_),
    .A(_3339_),
    .Y(_3341_));
 sg13g2_o21ai_1 _8514_ (.B1(_3341_),
    .Y(_3343_),
    .A1(_3227_),
    .A2(_3340_));
 sg13g2_or4_1 _8515_ (.A(_3234_),
    .B(_3248_),
    .C(_3229_),
    .D(_3227_),
    .X(_3344_));
 sg13g2_and3_1 _8516_ (.X(_3345_),
    .A(_3248_),
    .B(_3154_),
    .C(_3227_));
 sg13g2_o21ai_1 _8517_ (.B1(_3339_),
    .Y(_3346_),
    .A1(_3198_),
    .A2(_3225_));
 sg13g2_or3_1 _8518_ (.A(_3339_),
    .B(_3198_),
    .C(_3225_),
    .X(_3347_));
 sg13g2_a21oi_1 _8519_ (.A1(_3346_),
    .A2(_3347_),
    .Y(_3348_),
    .B1(_3154_));
 sg13g2_o21ai_1 _8520_ (.B1(_3234_),
    .Y(_3349_),
    .A1(_3345_),
    .A2(_3348_));
 sg13g2_nand2_1 _8521_ (.Y(_3350_),
    .A(_3330_),
    .B(_3329_));
 sg13g2_a21oi_1 _8522_ (.A1(_3344_),
    .A2(_3349_),
    .Y(_3351_),
    .B1(_3350_));
 sg13g2_xor2_1 _8523_ (.B(_3292_),
    .A(_3024_),
    .X(_3352_));
 sg13g2_nand3_1 _8524_ (.B(net87),
    .C(net34),
    .A(net224),
    .Y(_3354_));
 sg13g2_a221oi_1 _8525_ (.B2(_3354_),
    .C1(net35),
    .B1(net20),
    .A1(_1106_),
    .Y(_3355_),
    .A2(_1465_));
 sg13g2_nand2b_1 _8526_ (.Y(_3356_),
    .B(_3355_),
    .A_N(_1690_));
 sg13g2_a221oi_1 _8527_ (.B2(_3352_),
    .C1(_3356_),
    .B1(_3351_),
    .A1(_3338_),
    .Y(_3357_),
    .A2(_3343_));
 sg13g2_o21ai_1 _8528_ (.B1(_3357_),
    .Y(_3358_),
    .A1(_3323_),
    .A2(_3328_));
 sg13g2_nor2b_1 _8529_ (.A(_2627_),
    .B_N(_3358_),
    .Y(_3359_));
 sg13g2_o21ai_1 _8530_ (.B1(_3359_),
    .Y(_3360_),
    .A1(_1888_),
    .A2(_2826_));
 sg13g2_o21ai_1 _8531_ (.B1(_3360_),
    .Y(_3361_),
    .A1(_1535_),
    .A2(_2823_));
 sg13g2_nand2_1 _8532_ (.Y(_3362_),
    .A(net140),
    .B(_4275_));
 sg13g2_o21ai_1 _8533_ (.B1(_4185_),
    .Y(_3363_),
    .A1(_4281_),
    .A2(_3362_));
 sg13g2_nand3b_1 _8534_ (.B(_2645_),
    .C(_3363_),
    .Y(_3365_),
    .A_N(_0826_));
 sg13g2_nor2_1 _8535_ (.A(_0788_),
    .B(_3365_),
    .Y(_3366_));
 sg13g2_nor4_1 _8536_ (.A(_2352_),
    .B(net196),
    .C(_2766_),
    .D(_3366_),
    .Y(_3367_));
 sg13g2_nor4_1 _8537_ (.A(_2657_),
    .B(_2821_),
    .C(_3361_),
    .D(_3367_),
    .Y(_3368_));
 sg13g2_nor2_1 _8538_ (.A(net169),
    .B(_0877_),
    .Y(_3369_));
 sg13g2_nand2_1 _8539_ (.Y(_3370_),
    .A(_0836_),
    .B(_3369_));
 sg13g2_a21o_1 _8540_ (.A2(_3370_),
    .A1(_0827_),
    .B1(_0905_),
    .X(_3371_));
 sg13g2_a21oi_1 _8541_ (.A1(_3368_),
    .A2(_3371_),
    .Y(net7),
    .B1(_2642_));
 sg13g2_or2_1 _8542_ (.X(_3372_),
    .B(_2651_),
    .A(_2650_));
 sg13g2_a21oi_1 _8543_ (.A1(_2717_),
    .A2(_2724_),
    .Y(_3373_),
    .B1(_2361_));
 sg13g2_a21oi_1 _8544_ (.A1(_2344_),
    .A2(_2337_),
    .Y(_3374_),
    .B1(_3373_));
 sg13g2_a22oi_1 _8545_ (.Y(_3375_),
    .B1(_2029_),
    .B2(_2244_),
    .A2(_2012_),
    .A1(_2379_));
 sg13g2_nand2b_1 _8546_ (.Y(_3376_),
    .B(_2166_),
    .A_N(_3375_));
 sg13g2_o21ai_1 _8547_ (.B1(_2295_),
    .Y(_3377_),
    .A1(net85),
    .A2(_1552_));
 sg13g2_o21ai_1 _8548_ (.B1(_2749_),
    .Y(_3378_),
    .A1(_2275_),
    .A2(_2748_));
 sg13g2_a221oi_1 _8549_ (.B2(net52),
    .C1(_3378_),
    .B1(_3377_),
    .A1(net48),
    .Y(_3379_),
    .A2(_2161_));
 sg13g2_inv_1 _8550_ (.Y(_3380_),
    .A(_2430_));
 sg13g2_nand2_1 _8551_ (.Y(_3381_),
    .A(_0874_),
    .B(_2016_));
 sg13g2_a22oi_1 _8552_ (.Y(_3382_),
    .B1(_3381_),
    .B2(_0869_),
    .A2(_3380_),
    .A1(_0874_));
 sg13g2_inv_1 _8553_ (.Y(_3383_),
    .A(_3382_));
 sg13g2_o21ai_1 _8554_ (.B1(_3383_),
    .Y(_3385_),
    .A1(_1549_),
    .A2(_1587_));
 sg13g2_nor2_1 _8555_ (.A(net24),
    .B(_3385_),
    .Y(_3386_));
 sg13g2_o21ai_1 _8556_ (.B1(_2367_),
    .Y(_3387_),
    .A1(_2432_),
    .A2(_3386_));
 sg13g2_nand3_1 _8557_ (.B(_3379_),
    .C(_3387_),
    .A(_3376_),
    .Y(_3388_));
 sg13g2_nor2_1 _8558_ (.A(net153),
    .B(_2661_),
    .Y(_3389_));
 sg13g2_nor2_1 _8559_ (.A(_2659_),
    .B(_3389_),
    .Y(_3390_));
 sg13g2_nor2_1 _8560_ (.A(_2658_),
    .B(_3390_),
    .Y(_3391_));
 sg13g2_nand2_1 _8561_ (.Y(_3392_),
    .A(_1884_),
    .B(_1887_));
 sg13g2_a21o_1 _8562_ (.A2(_2825_),
    .A1(_1481_),
    .B1(_1862_),
    .X(_3393_));
 sg13g2_o21ai_1 _8563_ (.B1(_1690_),
    .Y(_3394_),
    .A1(_3392_),
    .A2(_3393_));
 sg13g2_a21oi_1 _8564_ (.A1(_3358_),
    .A2(_3394_),
    .Y(_3396_),
    .B1(_2627_));
 sg13g2_nor4_1 _8565_ (.A(_3374_),
    .B(_3388_),
    .C(_3391_),
    .D(_3396_),
    .Y(_3397_));
 sg13g2_o21ai_1 _8566_ (.B1(_3397_),
    .Y(_3398_),
    .A1(_2643_),
    .A2(_3372_));
 sg13g2_nor2b_1 _8567_ (.A(_1535_),
    .B_N(_1477_),
    .Y(_3399_));
 sg13g2_o21ai_1 _8568_ (.B1(_2822_),
    .Y(_3400_),
    .A1(net39),
    .A2(_1481_));
 sg13g2_nand2_1 _8569_ (.Y(_3401_),
    .A(_3399_),
    .B(_3400_));
 sg13g2_a21oi_1 _8570_ (.A1(net39),
    .A2(_2323_),
    .Y(_3402_),
    .B1(net43));
 sg13g2_a22oi_1 _8571_ (.Y(_3403_),
    .B1(_3402_),
    .B2(_1580_),
    .A2(net30),
    .A1(net92));
 sg13g2_o21ai_1 _8572_ (.B1(_2684_),
    .Y(_3404_),
    .A1(net55),
    .A2(_3403_));
 sg13g2_nand2_1 _8573_ (.Y(_3405_),
    .A(net132),
    .B(net149));
 sg13g2_nor2_1 _8574_ (.A(_2194_),
    .B(_2308_),
    .Y(_3407_));
 sg13g2_a21oi_1 _8575_ (.A1(_1980_),
    .A2(_3405_),
    .Y(_3408_),
    .B1(_3407_));
 sg13g2_nand3_1 _8576_ (.B(_2248_),
    .C(_2278_),
    .A(_2351_),
    .Y(_3409_));
 sg13g2_a21oi_1 _8577_ (.A1(_3408_),
    .A2(_3409_),
    .Y(_3410_),
    .B1(net51));
 sg13g2_o21ai_1 _8578_ (.B1(net136),
    .Y(_3411_),
    .A1(_2173_),
    .A2(_2727_));
 sg13g2_o21ai_1 _8579_ (.B1(_3411_),
    .Y(_3412_),
    .A1(_2390_),
    .A2(_2405_));
 sg13g2_inv_1 _8580_ (.Y(_3413_),
    .A(_3412_));
 sg13g2_o21ai_1 _8581_ (.B1(_2595_),
    .Y(_3414_),
    .A1(net27),
    .A2(_2248_));
 sg13g2_o21ai_1 _8582_ (.B1(_2233_),
    .Y(_3415_),
    .A1(net109),
    .A2(net57));
 sg13g2_a22oi_1 _8583_ (.Y(_3416_),
    .B1(_1576_),
    .B2(net115),
    .A2(net79),
    .A1(_2340_));
 sg13g2_mux2_1 _8584_ (.A0(_2370_),
    .A1(_2386_),
    .S(net151),
    .X(_3418_));
 sg13g2_o21ai_1 _8585_ (.B1(_3418_),
    .Y(_3419_),
    .A1(net30),
    .A2(_3416_));
 sg13g2_a21oi_1 _8586_ (.A1(_2029_),
    .A2(_2402_),
    .Y(_3420_),
    .B1(_3419_));
 sg13g2_nand4_1 _8587_ (.B(_3414_),
    .C(_3415_),
    .A(_3413_),
    .Y(_3421_),
    .D(_3420_));
 sg13g2_o21ai_1 _8588_ (.B1(_2196_),
    .Y(_3422_),
    .A1(_2674_),
    .A2(_2198_));
 sg13g2_nand2b_1 _8589_ (.Y(_3423_),
    .B(_2134_),
    .A_N(_2403_));
 sg13g2_nor2_1 _8590_ (.A(net114),
    .B(_2003_),
    .Y(_3424_));
 sg13g2_nor2_1 _8591_ (.A(net80),
    .B(_2230_),
    .Y(_3425_));
 sg13g2_a221oi_1 _8592_ (.B2(_3424_),
    .C1(_3425_),
    .B1(_3423_),
    .A1(_1816_),
    .Y(_3426_),
    .A2(_2320_));
 sg13g2_a21oi_1 _8593_ (.A1(_2194_),
    .A2(_2318_),
    .Y(_3427_),
    .B1(net91));
 sg13g2_nor3_1 _8594_ (.A(_2293_),
    .B(net112),
    .C(_1480_),
    .Y(_3428_));
 sg13g2_nor3_1 _8595_ (.A(_2372_),
    .B(_3427_),
    .C(_3428_),
    .Y(_3429_));
 sg13g2_nand2_1 _8596_ (.Y(_3430_),
    .A(_3426_),
    .B(_3429_));
 sg13g2_nor4_1 _8597_ (.A(net73),
    .B(net114),
    .C(net94),
    .D(_2010_),
    .Y(_3431_));
 sg13g2_inv_1 _8598_ (.Y(_3432_),
    .A(_2325_));
 sg13g2_nand2_1 _8599_ (.Y(_3433_),
    .A(net92),
    .B(_2388_));
 sg13g2_a22oi_1 _8600_ (.Y(_3434_),
    .B1(_3432_),
    .B2(_3433_),
    .A2(_2010_),
    .A1(net29));
 sg13g2_nor4_1 _8601_ (.A(_2624_),
    .B(_3430_),
    .C(_3431_),
    .D(_3434_),
    .Y(_3435_));
 sg13g2_nand3_1 _8602_ (.B(_3422_),
    .C(_3435_),
    .A(_2225_),
    .Y(_3436_));
 sg13g2_nor3_1 _8603_ (.A(net56),
    .B(net85),
    .C(_2697_),
    .Y(_3437_));
 sg13g2_o21ai_1 _8604_ (.B1(_2400_),
    .Y(_3439_),
    .A1(net183),
    .A2(_2289_));
 sg13g2_nand3_1 _8605_ (.B(_2289_),
    .C(_2395_),
    .A(_0854_),
    .Y(_3440_));
 sg13g2_nor2_1 _8606_ (.A(net56),
    .B(net90),
    .Y(_3441_));
 sg13g2_o21ai_1 _8607_ (.B1(net24),
    .Y(_3442_),
    .A1(_2653_),
    .A2(_3441_));
 sg13g2_o21ai_1 _8608_ (.B1(net75),
    .Y(_3443_),
    .A1(net29),
    .A2(net133));
 sg13g2_nand3_1 _8609_ (.B(net48),
    .C(_3443_),
    .A(_1566_),
    .Y(_3444_));
 sg13g2_nand4_1 _8610_ (.B(_3440_),
    .C(_3442_),
    .A(_3439_),
    .Y(_3445_),
    .D(_3444_));
 sg13g2_nor4_1 _8611_ (.A(_3421_),
    .B(_3436_),
    .C(_3437_),
    .D(_3445_),
    .Y(_3446_));
 sg13g2_nor2_1 _8612_ (.A(_2608_),
    .B(_2147_),
    .Y(_3447_));
 sg13g2_a21oi_1 _8613_ (.A1(net27),
    .A2(_1482_),
    .Y(_3448_),
    .B1(net56));
 sg13g2_o21ai_1 _8614_ (.B1(_1547_),
    .Y(_3450_),
    .A1(_3447_),
    .A2(_3448_));
 sg13g2_nand3_1 _8615_ (.B(_2145_),
    .C(_2699_),
    .A(_2208_),
    .Y(_3451_));
 sg13g2_a21oi_1 _8616_ (.A1(net27),
    .A2(_2284_),
    .Y(_3452_),
    .B1(_3451_));
 sg13g2_a21oi_1 _8617_ (.A1(_2394_),
    .A2(_2681_),
    .Y(_3453_),
    .B1(_3452_));
 sg13g2_nand2_1 _8618_ (.Y(_3454_),
    .A(_2166_),
    .B(_1573_));
 sg13g2_o21ai_1 _8619_ (.B1(_3454_),
    .Y(_3455_),
    .A1(_1540_),
    .A2(_1573_));
 sg13g2_nand2_1 _8620_ (.Y(_3456_),
    .A(net134),
    .B(net77));
 sg13g2_nand2_1 _8621_ (.Y(_3457_),
    .A(_2376_),
    .B(_2223_));
 sg13g2_a221oi_1 _8622_ (.B2(net47),
    .C1(_2597_),
    .B1(_3457_),
    .A1(_2675_),
    .Y(_3458_),
    .A2(_3456_));
 sg13g2_nor2_1 _8623_ (.A(_2216_),
    .B(_3458_),
    .Y(_3459_));
 sg13g2_a21oi_1 _8624_ (.A1(_1571_),
    .A2(_3455_),
    .Y(_3461_),
    .B1(_3459_));
 sg13g2_nand4_1 _8625_ (.B(_3450_),
    .C(_3453_),
    .A(_3446_),
    .Y(_3462_),
    .D(_3461_));
 sg13g2_o21ai_1 _8626_ (.B1(_2215_),
    .Y(_3463_),
    .A1(net31),
    .A2(_2690_));
 sg13g2_buf_2 _8627_ (.A(_3463_),
    .X(_3464_));
 sg13g2_nand2_1 _8628_ (.Y(_3465_),
    .A(net92),
    .B(_2420_));
 sg13g2_o21ai_1 _8629_ (.B1(_3465_),
    .Y(_3466_),
    .A1(net73),
    .A2(_2744_));
 sg13g2_o21ai_1 _8630_ (.B1(net37),
    .Y(_3467_),
    .A1(_2687_),
    .A2(_3385_));
 sg13g2_a22oi_1 _8631_ (.Y(_3468_),
    .B1(_3467_),
    .B2(_2434_),
    .A2(_3466_),
    .A1(net108));
 sg13g2_o21ai_1 _8632_ (.B1(_3468_),
    .Y(_3469_),
    .A1(_2220_),
    .A2(_3464_));
 sg13g2_nor4_1 _8633_ (.A(_3404_),
    .B(_3410_),
    .C(_3462_),
    .D(_3469_),
    .Y(_3470_));
 sg13g2_inv_1 _8634_ (.Y(_3472_),
    .A(_2567_));
 sg13g2_nor2_1 _8635_ (.A(_3472_),
    .B(_2578_),
    .Y(_3473_));
 sg13g2_nand2b_1 _8636_ (.Y(_3474_),
    .B(_3473_),
    .A_N(_2570_));
 sg13g2_mux2_1 _8637_ (.A0(_3474_),
    .A1(_3473_),
    .S(_2583_),
    .X(_3475_));
 sg13g2_nor2b_1 _8638_ (.A(_3475_),
    .B_N(_2560_),
    .Y(_3476_));
 sg13g2_nand2b_1 _8639_ (.Y(_3477_),
    .B(_3476_),
    .A_N(_2441_));
 sg13g2_nand4_1 _8640_ (.B(_3401_),
    .C(_3470_),
    .A(_2132_),
    .Y(_3478_),
    .D(_3477_));
 sg13g2_nor2_1 _8641_ (.A(net196),
    .B(_2766_),
    .Y(_3479_));
 sg13g2_a21oi_1 _8642_ (.A1(_3366_),
    .A2(_3479_),
    .Y(_3480_),
    .B1(_2352_));
 sg13g2_nor3_1 _8643_ (.A(_3398_),
    .B(_3478_),
    .C(_3480_),
    .Y(_3481_));
 sg13g2_nand2_1 _8644_ (.Y(_3483_),
    .A(_0834_),
    .B(_0856_));
 sg13g2_a21o_1 _8645_ (.A2(_3483_),
    .A1(_0827_),
    .B1(_0905_),
    .X(_3484_));
 sg13g2_a21oi_1 _8646_ (.A1(_3481_),
    .A2(_3484_),
    .Y(net8),
    .B1(_2642_));
 sg13g2_nand2_1 _8647_ (.Y(_3485_),
    .A(_4131_),
    .B(_4108_));
 sg13g2_mux2_1 _8648_ (.A0(_3365_),
    .A1(_3485_),
    .S(_0788_),
    .X(_3486_));
 sg13g2_nor3_1 _8649_ (.A(_2352_),
    .B(_2766_),
    .C(_3486_),
    .Y(_3487_));
 sg13g2_nor2_1 _8650_ (.A(net86),
    .B(_1862_),
    .Y(_3488_));
 sg13g2_nand3_1 _8651_ (.B(_1887_),
    .C(_3488_),
    .A(_1884_),
    .Y(_3489_));
 sg13g2_a21oi_1 _8652_ (.A1(_1745_),
    .A2(_3489_),
    .Y(_3490_),
    .B1(_2658_));
 sg13g2_a22oi_1 _8653_ (.Y(_3491_),
    .B1(_1988_),
    .B2(net83),
    .A2(_2811_),
    .A1(_1566_));
 sg13g2_a21oi_1 _8654_ (.A1(_3449_),
    .A2(net283),
    .Y(_3493_),
    .B1(_3546_));
 sg13g2_a21oi_1 _8655_ (.A1(_2444_),
    .A2(_0964_),
    .Y(_3494_),
    .B1(net173));
 sg13g2_o21ai_1 _8656_ (.B1(_1062_),
    .Y(_3495_),
    .A1(_3493_),
    .A2(_3494_));
 sg13g2_o21ai_1 _8657_ (.B1(_3495_),
    .Y(_3496_),
    .A1(net243),
    .A2(_1466_));
 sg13g2_nor2_2 _8658_ (.A(_3493_),
    .B(_3494_),
    .Y(_3497_));
 sg13g2_o21ai_1 _8659_ (.B1(net247),
    .Y(_3498_),
    .A1(_1466_),
    .A2(_3497_));
 sg13g2_a221oi_1 _8660_ (.B2(net242),
    .C1(_2799_),
    .B1(_3498_),
    .A1(net191),
    .Y(_3499_),
    .A2(_3496_));
 sg13g2_buf_1 _8661_ (.A(_3499_),
    .X(_3500_));
 sg13g2_xnor2_1 _8662_ (.Y(_3501_),
    .A(_0886_),
    .B(_3500_));
 sg13g2_o21ai_1 _8663_ (.B1(_2591_),
    .Y(_3502_),
    .A1(_3870_),
    .A2(_3501_));
 sg13g2_xnor2_1 _8664_ (.Y(_3504_),
    .A(_0831_),
    .B(_3502_));
 sg13g2_xnor2_1 _8665_ (.Y(_3505_),
    .A(_0853_),
    .B(_3500_));
 sg13g2_or2_1 _8666_ (.X(_3506_),
    .B(_3505_),
    .A(net305));
 sg13g2_o21ai_1 _8667_ (.B1(_2444_),
    .Y(_3507_),
    .A1(net243),
    .A2(_0964_));
 sg13g2_o21ai_1 _8668_ (.B1(net244),
    .Y(_3508_),
    .A1(net181),
    .A2(net243));
 sg13g2_a221oi_1 _8669_ (.B2(net214),
    .C1(_1106_),
    .B1(_3508_),
    .A1(net178),
    .Y(_3509_),
    .A2(_3507_));
 sg13g2_xnor2_1 _8670_ (.Y(_3510_),
    .A(net247),
    .B(_3509_));
 sg13g2_xor2_1 _8671_ (.B(_3510_),
    .A(net171),
    .X(_3511_));
 sg13g2_o21ai_1 _8672_ (.B1(net245),
    .Y(_3512_),
    .A1(_1084_),
    .A2(_3497_));
 sg13g2_a21oi_1 _8673_ (.A1(_1084_),
    .A2(_3497_),
    .Y(_3513_),
    .B1(net245));
 sg13g2_nand2_1 _8674_ (.Y(_3515_),
    .A(net280),
    .B(_3513_));
 sg13g2_o21ai_1 _8675_ (.B1(_3515_),
    .Y(_3516_),
    .A1(net280),
    .A2(_3512_));
 sg13g2_xnor2_1 _8676_ (.Y(_3517_),
    .A(net285),
    .B(_3516_));
 sg13g2_xor2_1 _8677_ (.B(_3517_),
    .A(net257),
    .X(_3518_));
 sg13g2_nand2_1 _8678_ (.Y(_3519_),
    .A(_3511_),
    .B(_3518_));
 sg13g2_xor2_1 _8679_ (.B(_3497_),
    .A(_2474_),
    .X(_3520_));
 sg13g2_xnor2_1 _8680_ (.Y(_3521_),
    .A(net272),
    .B(_3520_));
 sg13g2_a22oi_1 _8681_ (.Y(_3522_),
    .B1(_1147_),
    .B2(net178),
    .A2(_2800_),
    .A1(_1196_));
 sg13g2_xnor2_1 _8682_ (.Y(_3523_),
    .A(net244),
    .B(_3522_));
 sg13g2_xor2_1 _8683_ (.B(_3523_),
    .A(net297),
    .X(_3524_));
 sg13g2_and2_1 _8684_ (.A(net305),
    .B(_3505_),
    .X(_3526_));
 sg13g2_nor4_1 _8685_ (.A(_3519_),
    .B(_3521_),
    .C(_3524_),
    .D(_3526_),
    .Y(_3527_));
 sg13g2_xnor2_1 _8686_ (.Y(_3528_),
    .A(net293),
    .B(net201));
 sg13g2_nand3_1 _8687_ (.B(net265),
    .C(_4110_),
    .A(net168),
    .Y(_3529_));
 sg13g2_o21ai_1 _8688_ (.B1(_3529_),
    .Y(_3530_),
    .A1(net265),
    .A2(_3054_));
 sg13g2_buf_1 _8689_ (.A(net173),
    .X(_3531_));
 sg13g2_xor2_1 _8690_ (.B(net265),
    .A(_3460_),
    .X(_3532_));
 sg13g2_nor3_1 _8691_ (.A(net174),
    .B(net168),
    .C(net265),
    .Y(_3533_));
 sg13g2_a21oi_1 _8692_ (.A1(_0857_),
    .A2(_3532_),
    .Y(_3534_),
    .B1(_3533_));
 sg13g2_nand3_1 _8693_ (.B(net168),
    .C(net265),
    .A(_1145_),
    .Y(_3535_));
 sg13g2_o21ai_1 _8694_ (.B1(_3535_),
    .Y(_3536_),
    .A1(net161),
    .A2(_3534_));
 sg13g2_nor2b_1 _8695_ (.A(_3528_),
    .B_N(_3536_),
    .Y(_3537_));
 sg13g2_a21oi_1 _8696_ (.A1(_3528_),
    .A2(_3530_),
    .Y(_3538_),
    .B1(_3537_));
 sg13g2_nor2_1 _8697_ (.A(net195),
    .B(_3538_),
    .Y(_3539_));
 sg13g2_nor2_1 _8698_ (.A(_3531_),
    .B(_2857_),
    .Y(_3540_));
 sg13g2_a21oi_1 _8699_ (.A1(net201),
    .A2(_2484_),
    .Y(_3541_),
    .B1(net254));
 sg13g2_o21ai_1 _8700_ (.B1(net163),
    .Y(_3542_),
    .A1(_3540_),
    .A2(_3541_));
 sg13g2_nand2_1 _8701_ (.Y(_3543_),
    .A(net161),
    .B(net201));
 sg13g2_o21ai_1 _8702_ (.B1(_3543_),
    .Y(_3544_),
    .A1(_3531_),
    .A2(_0964_));
 sg13g2_nand2_1 _8703_ (.Y(_3545_),
    .A(_1292_),
    .B(_3544_));
 sg13g2_nand2_1 _8704_ (.Y(_3547_),
    .A(_3816_),
    .B(net172));
 sg13g2_a21oi_1 _8705_ (.A1(net209),
    .A2(net168),
    .Y(_3548_),
    .B1(net210));
 sg13g2_a21oi_1 _8706_ (.A1(net201),
    .A2(_1196_),
    .Y(_3549_),
    .B1(_3548_));
 sg13g2_nand2_1 _8707_ (.Y(_3550_),
    .A(net163),
    .B(net214));
 sg13g2_o21ai_1 _8708_ (.B1(net254),
    .Y(_3551_),
    .A1(net161),
    .A2(_3550_));
 sg13g2_a22oi_1 _8709_ (.Y(_3552_),
    .B1(_3551_),
    .B2(net209),
    .A2(_3549_),
    .A1(_3547_));
 sg13g2_nand3_1 _8710_ (.B(_3545_),
    .C(_3552_),
    .A(_3542_),
    .Y(_3553_));
 sg13g2_a22oi_1 _8711_ (.Y(_3554_),
    .B1(_3553_),
    .B2(_3590_),
    .A2(_3539_),
    .A1(net212));
 sg13g2_nand2b_1 _8712_ (.Y(_3555_),
    .B(net161),
    .A_N(_3554_));
 sg13g2_mux2_1 _8713_ (.A0(_3539_),
    .A1(_3553_),
    .S(net212),
    .X(_3556_));
 sg13g2_a22oi_1 _8714_ (.Y(_3558_),
    .B1(_3556_),
    .B2(_3816_),
    .A2(_3553_),
    .A1(_3538_));
 sg13g2_nand3_1 _8715_ (.B(_3555_),
    .C(_3558_),
    .A(_3527_),
    .Y(_3559_));
 sg13g2_xnor2_1 _8716_ (.Y(_3560_),
    .A(net232),
    .B(_4440_));
 sg13g2_and3_1 _8717_ (.X(_3561_),
    .A(_3527_),
    .B(_3560_),
    .C(_3539_));
 sg13g2_nor2b_1 _8718_ (.A(net297),
    .B_N(_3523_),
    .Y(_3562_));
 sg13g2_nand2b_1 _8719_ (.Y(_3563_),
    .B(_3562_),
    .A_N(_3521_));
 sg13g2_o21ai_1 _8720_ (.B1(_3563_),
    .Y(_3564_),
    .A1(net193),
    .A2(_3520_));
 sg13g2_nand3_1 _8721_ (.B(_3518_),
    .C(_3564_),
    .A(_3511_),
    .Y(_3565_));
 sg13g2_xnor2_1 _8722_ (.Y(_3566_),
    .A(net242),
    .B(_3510_));
 sg13g2_nor2_1 _8723_ (.A(_1914_),
    .B(_3566_),
    .Y(_3567_));
 sg13g2_a21o_1 _8724_ (.A2(_3567_),
    .A1(_3517_),
    .B1(net222),
    .X(_3569_));
 sg13g2_o21ai_1 _8725_ (.B1(_3569_),
    .Y(_3570_),
    .A1(_3517_),
    .A2(_3567_));
 sg13g2_and2_1 _8726_ (.A(_3565_),
    .B(_3570_),
    .X(_3571_));
 sg13g2_or3_1 _8727_ (.A(_3526_),
    .B(_3561_),
    .C(_3571_),
    .X(_3572_));
 sg13g2_nand3_1 _8728_ (.B(_3559_),
    .C(_3572_),
    .A(_3506_),
    .Y(_3573_));
 sg13g2_nand2b_1 _8729_ (.Y(_3574_),
    .B(_3573_),
    .A_N(net262));
 sg13g2_nand3_1 _8730_ (.B(_3561_),
    .C(_3506_),
    .A(net262),
    .Y(_3575_));
 sg13g2_a221oi_1 _8731_ (.B2(net262),
    .C1(_3504_),
    .B1(_3573_),
    .A1(net221),
    .Y(_3576_),
    .A2(_3575_));
 sg13g2_a21o_1 _8732_ (.A2(_3574_),
    .A1(_3504_),
    .B1(_3576_),
    .X(_3577_));
 sg13g2_nor2_1 _8733_ (.A(_0886_),
    .B(_0853_),
    .Y(_3578_));
 sg13g2_nor2_1 _8734_ (.A(net246),
    .B(_3500_),
    .Y(_3580_));
 sg13g2_nor3_1 _8735_ (.A(_1762_),
    .B(_1684_),
    .C(_3580_),
    .Y(_3581_));
 sg13g2_a21oi_1 _8736_ (.A1(_1762_),
    .A2(_3578_),
    .Y(_3582_),
    .B1(_3581_));
 sg13g2_nor2_1 _8737_ (.A(_0370_),
    .B(net44),
    .Y(_3583_));
 sg13g2_inv_1 _8738_ (.Y(_3584_),
    .A(_2475_));
 sg13g2_xnor2_1 _8739_ (.Y(_3585_),
    .A(_3976_),
    .B(_2475_));
 sg13g2_nor2_1 _8740_ (.A(net297),
    .B(_2492_),
    .Y(_3586_));
 sg13g2_a22oi_1 _8741_ (.Y(_3587_),
    .B1(_3585_),
    .B2(_3586_),
    .A2(_3584_),
    .A1(_0711_));
 sg13g2_o21ai_1 _8742_ (.B1(net206),
    .Y(_3588_),
    .A1(_1344_),
    .A2(_3587_));
 sg13g2_o21ai_1 _8743_ (.B1(_2469_),
    .Y(_3589_),
    .A1(_1717_),
    .A2(_3587_));
 sg13g2_o21ai_1 _8744_ (.B1(_3589_),
    .Y(_3591_),
    .A1(_2469_),
    .A2(_3588_));
 sg13g2_nand2_1 _8745_ (.Y(_3592_),
    .A(net172),
    .B(_3054_));
 sg13g2_a22oi_1 _8746_ (.Y(_3593_),
    .B1(_3592_),
    .B2(net210),
    .A2(_1147_),
    .A1(net161));
 sg13g2_o21ai_1 _8747_ (.B1(_3547_),
    .Y(_3594_),
    .A1(net172),
    .A2(_1402_));
 sg13g2_a21oi_1 _8748_ (.A1(net209),
    .A2(_1292_),
    .Y(_3595_),
    .B1(net210));
 sg13g2_a21oi_1 _8749_ (.A1(net161),
    .A2(_3550_),
    .Y(_3596_),
    .B1(_3595_));
 sg13g2_a21oi_1 _8750_ (.A1(net201),
    .A2(_3406_),
    .Y(_3597_),
    .B1(net210));
 sg13g2_nor2_1 _8751_ (.A(net260),
    .B(_3597_),
    .Y(_3598_));
 sg13g2_a221oi_1 _8752_ (.B2(_3547_),
    .C1(_3598_),
    .B1(_3596_),
    .A1(net160),
    .Y(_3599_),
    .A2(_3594_));
 sg13g2_o21ai_1 _8753_ (.B1(_3599_),
    .Y(_3600_),
    .A1(net163),
    .A2(_3593_));
 sg13g2_nor2_1 _8754_ (.A(net168),
    .B(net269),
    .Y(_3602_));
 sg13g2_nand3_1 _8755_ (.B(net168),
    .C(net269),
    .A(net163),
    .Y(_3603_));
 sg13g2_o21ai_1 _8756_ (.B1(_3603_),
    .Y(_3604_),
    .A1(net163),
    .A2(_3532_));
 sg13g2_mux2_1 _8757_ (.A0(_3602_),
    .A1(_3604_),
    .S(net161),
    .X(_3605_));
 sg13g2_a22oi_1 _8758_ (.Y(_3606_),
    .B1(_3602_),
    .B2(_3677_),
    .A2(_1151_),
    .A1(net269));
 sg13g2_nor2_1 _8759_ (.A(_3528_),
    .B(_3606_),
    .Y(_3607_));
 sg13g2_a21oi_1 _8760_ (.A1(_3528_),
    .A2(_3605_),
    .Y(_3608_),
    .B1(_3607_));
 sg13g2_a21oi_1 _8761_ (.A1(net161),
    .A2(net212),
    .Y(_3609_),
    .B1(_3395_));
 sg13g2_nand2b_1 _8762_ (.Y(_3610_),
    .B(_3609_),
    .A_N(_3608_));
 sg13g2_xor2_1 _8763_ (.B(_2492_),
    .A(net297),
    .X(_3611_));
 sg13g2_xnor2_1 _8764_ (.Y(_3613_),
    .A(_1081_),
    .B(_2469_));
 sg13g2_xor2_1 _8765_ (.B(net44),
    .A(net222),
    .X(_3614_));
 sg13g2_nand4_1 _8766_ (.B(_3611_),
    .C(_3613_),
    .A(_3585_),
    .Y(_3615_),
    .D(_3614_));
 sg13g2_a21oi_1 _8767_ (.A1(_3600_),
    .A2(_3610_),
    .Y(_3616_),
    .B1(_3615_));
 sg13g2_a21oi_1 _8768_ (.A1(_0370_),
    .A2(net44),
    .Y(_3617_),
    .B1(_3616_));
 sg13g2_o21ai_1 _8769_ (.B1(_3617_),
    .Y(_3618_),
    .A1(_3583_),
    .A2(_3591_));
 sg13g2_nor2_1 _8770_ (.A(_2516_),
    .B(_3618_),
    .Y(_3619_));
 sg13g2_nand2_1 _8771_ (.Y(_3620_),
    .A(_2516_),
    .B(_3618_));
 sg13g2_o21ai_1 _8772_ (.B1(_3620_),
    .Y(_3621_),
    .A1(net305),
    .A2(_3619_));
 sg13g2_xor2_1 _8773_ (.B(_2457_),
    .A(net262),
    .X(_3622_));
 sg13g2_a22oi_1 _8774_ (.Y(_3624_),
    .B1(_3621_),
    .B2(_3622_),
    .A2(_2458_),
    .A1(net221));
 sg13g2_xnor2_1 _8775_ (.Y(_3625_),
    .A(net305),
    .B(_2515_));
 sg13g2_nand2_1 _8776_ (.Y(_3626_),
    .A(_3590_),
    .B(_3560_));
 sg13g2_nor4_1 _8777_ (.A(_3615_),
    .B(_3625_),
    .C(_3608_),
    .D(_3626_),
    .Y(_3627_));
 sg13g2_a221oi_1 _8778_ (.B2(_3622_),
    .C1(net229),
    .B1(_3627_),
    .A1(_0864_),
    .Y(_3628_),
    .A2(_2530_));
 sg13g2_nand2b_1 _8779_ (.Y(_3629_),
    .B(_3628_),
    .A_N(_3624_));
 sg13g2_o21ai_1 _8780_ (.B1(_3629_),
    .Y(_3630_),
    .A1(_3577_),
    .A2(_3582_));
 sg13g2_xnor2_1 _8781_ (.Y(_3631_),
    .A(net86),
    .B(_3630_));
 sg13g2_and2_1 _8782_ (.A(_2221_),
    .B(_3631_),
    .X(_3632_));
 sg13g2_nand2_1 _8783_ (.Y(_3633_),
    .A(net46),
    .B(_2273_));
 sg13g2_o21ai_1 _8784_ (.B1(_3633_),
    .Y(_3634_),
    .A1(_2351_),
    .A2(_2388_));
 sg13g2_o21ai_1 _8785_ (.B1(_3634_),
    .Y(_3635_),
    .A1(net55),
    .A2(_2029_));
 sg13g2_a21oi_1 _8786_ (.A1(_2408_),
    .A2(_3464_),
    .Y(_3636_),
    .B1(_3635_));
 sg13g2_a21oi_1 _8787_ (.A1(_1533_),
    .A2(_4512_),
    .Y(_3637_),
    .B1(_1576_));
 sg13g2_nor2_1 _8788_ (.A(net84),
    .B(_3637_),
    .Y(_3638_));
 sg13g2_nand2_1 _8789_ (.Y(_3639_),
    .A(net81),
    .B(_2196_));
 sg13g2_a21oi_1 _8790_ (.A1(_2204_),
    .A2(_2198_),
    .Y(_3640_),
    .B1(_3639_));
 sg13g2_a221oi_1 _8791_ (.B2(net86),
    .C1(_3640_),
    .B1(_3638_),
    .A1(_2224_),
    .Y(_3641_),
    .A2(_2420_));
 sg13g2_nor2b_1 _8792_ (.A(_2424_),
    .B_N(_3641_),
    .Y(_3642_));
 sg13g2_o21ai_1 _8793_ (.B1(_3642_),
    .Y(_3643_),
    .A1(net51),
    .A2(_3636_));
 sg13g2_nor3_1 _8794_ (.A(_2131_),
    .B(_3632_),
    .C(_3643_),
    .Y(_3645_));
 sg13g2_o21ai_1 _8795_ (.B1(_3645_),
    .Y(_3646_),
    .A1(_1998_),
    .A2(_3491_));
 sg13g2_nor2_1 _8796_ (.A(_2441_),
    .B(_2585_),
    .Y(_3647_));
 sg13g2_nand2_1 _8797_ (.Y(_3648_),
    .A(_2531_),
    .B(_3580_));
 sg13g2_a21o_1 _8798_ (.A2(_3395_),
    .A1(net218),
    .B1(_4438_),
    .X(_3649_));
 sg13g2_a21oi_1 _8799_ (.A1(net160),
    .A2(_3649_),
    .Y(_3650_),
    .B1(net180));
 sg13g2_o21ai_1 _8800_ (.B1(net242),
    .Y(_3651_),
    .A1(net191),
    .A2(_3650_));
 sg13g2_and2_1 _8801_ (.A(_0930_),
    .B(_3651_),
    .X(_3652_));
 sg13g2_buf_1 _8802_ (.A(_3652_),
    .X(_3653_));
 sg13g2_nand2_1 _8803_ (.Y(_3654_),
    .A(_1051_),
    .B(_3653_));
 sg13g2_o21ai_1 _8804_ (.B1(net192),
    .Y(_3656_),
    .A1(net156),
    .A2(_3654_));
 sg13g2_o21ai_1 _8805_ (.B1(_3656_),
    .Y(_3657_),
    .A1(_2234_),
    .A2(_3648_));
 sg13g2_o21ai_1 _8806_ (.B1(_0864_),
    .Y(_3658_),
    .A1(net216),
    .A2(_3653_));
 sg13g2_and2_1 _8807_ (.A(_0809_),
    .B(_3658_),
    .X(_3659_));
 sg13g2_nand3_1 _8808_ (.B(_3648_),
    .C(_3659_),
    .A(net156),
    .Y(_3660_));
 sg13g2_a21oi_1 _8809_ (.A1(_4118_),
    .A2(_3660_),
    .Y(_3661_),
    .B1(_1741_));
 sg13g2_nor2_1 _8810_ (.A(_3657_),
    .B(_3661_),
    .Y(_3662_));
 sg13g2_inv_1 _8811_ (.Y(_3663_),
    .A(_3464_));
 sg13g2_o21ai_1 _8812_ (.B1(_3663_),
    .Y(_3664_),
    .A1(_2273_),
    .A2(_3662_));
 sg13g2_a22oi_1 _8813_ (.Y(_3665_),
    .B1(_3664_),
    .B2(_2188_),
    .A2(_2691_),
    .A1(net108));
 sg13g2_nand2_1 _8814_ (.Y(_3667_),
    .A(_2208_),
    .B(_2257_));
 sg13g2_nand3b_1 _8815_ (.B(_3667_),
    .C(net45),
    .Y(_3668_),
    .A_N(net31));
 sg13g2_nand4_1 _8816_ (.B(net81),
    .C(_2258_),
    .A(_2302_),
    .Y(_3669_),
    .D(_2277_));
 sg13g2_a22oi_1 _8817_ (.Y(_3670_),
    .B1(_3669_),
    .B2(_2313_),
    .A2(_3668_),
    .A1(_2593_));
 sg13g2_nand2_1 _8818_ (.Y(_3671_),
    .A(net97),
    .B(net77));
 sg13g2_nor2b_1 _8819_ (.A(_2398_),
    .B_N(_3671_),
    .Y(_3672_));
 sg13g2_a22oi_1 _8820_ (.Y(_3673_),
    .B1(_3672_),
    .B2(_2258_),
    .A2(_2699_),
    .A1(_2674_));
 sg13g2_a21oi_1 _8821_ (.A1(_3670_),
    .A2(_3673_),
    .Y(_3674_),
    .B1(net72));
 sg13g2_a21oi_1 _8822_ (.A1(_2018_),
    .A2(_2257_),
    .Y(_3675_),
    .B1(net135));
 sg13g2_or2_1 _8823_ (.X(_3676_),
    .B(_3675_),
    .A(net77));
 sg13g2_buf_1 _8824_ (.A(_3676_),
    .X(_3678_));
 sg13g2_nor2_1 _8825_ (.A(_2232_),
    .B(_3678_),
    .Y(_3679_));
 sg13g2_a21oi_1 _8826_ (.A1(net83),
    .A2(net31),
    .Y(_3680_),
    .B1(_3679_));
 sg13g2_a21oi_1 _8827_ (.A1(net46),
    .A2(_3678_),
    .Y(_3681_),
    .B1(net29));
 sg13g2_nor4_1 _8828_ (.A(net114),
    .B(net51),
    .C(_2136_),
    .D(_3681_),
    .Y(_3682_));
 sg13g2_o21ai_1 _8829_ (.B1(_2710_),
    .Y(_3683_),
    .A1(_0612_),
    .A2(net120));
 sg13g2_nand4_1 _8830_ (.B(_1526_),
    .C(net132),
    .A(_2369_),
    .Y(_3684_),
    .D(_3683_));
 sg13g2_o21ai_1 _8831_ (.B1(net136),
    .Y(_3685_),
    .A1(_2141_),
    .A2(net97));
 sg13g2_a22oi_1 _8832_ (.Y(_3686_),
    .B1(_2402_),
    .B2(_3685_),
    .A2(_2158_),
    .A1(net162));
 sg13g2_o21ai_1 _8833_ (.B1(net79),
    .Y(_3687_),
    .A1(_2161_),
    .A2(_2732_));
 sg13g2_nand3_1 _8834_ (.B(_2219_),
    .C(_3464_),
    .A(_2169_),
    .Y(_3689_));
 sg13g2_and4_1 _8835_ (.A(_3684_),
    .B(_3686_),
    .C(_3687_),
    .D(_3689_),
    .X(_3690_));
 sg13g2_nor2b_1 _8836_ (.A(_3682_),
    .B_N(_3690_),
    .Y(_3691_));
 sg13g2_o21ai_1 _8837_ (.B1(_3691_),
    .Y(_3692_),
    .A1(net53),
    .A2(_3680_));
 sg13g2_a21o_1 _8838_ (.A2(_2275_),
    .A1(net61),
    .B1(net135),
    .X(_3693_));
 sg13g2_a21oi_1 _8839_ (.A1(_2018_),
    .A2(_2286_),
    .Y(_3694_),
    .B1(_2259_));
 sg13g2_a21oi_1 _8840_ (.A1(net135),
    .A2(_2286_),
    .Y(_3695_),
    .B1(net77));
 sg13g2_o21ai_1 _8841_ (.B1(_3695_),
    .Y(_3696_),
    .A1(_3693_),
    .A2(_3694_));
 sg13g2_nand2_1 _8842_ (.Y(_3697_),
    .A(_1527_),
    .B(_2188_));
 sg13g2_a21oi_1 _8843_ (.A1(net28),
    .A2(_3696_),
    .Y(_3698_),
    .B1(_3697_));
 sg13g2_a21oi_1 _8844_ (.A1(_2418_),
    .A2(_2683_),
    .Y(_3700_),
    .B1(_2300_));
 sg13g2_a21oi_1 _8845_ (.A1(_2208_),
    .A2(_2699_),
    .Y(_3701_),
    .B1(_2683_));
 sg13g2_a21oi_2 _8846_ (.B1(_2130_),
    .Y(_3702_),
    .A2(_0828_),
    .A1(_4078_));
 sg13g2_a21oi_1 _8847_ (.A1(_3702_),
    .A2(_2289_),
    .Y(_3703_),
    .B1(_2762_));
 sg13g2_nand3_1 _8848_ (.B(net162),
    .C(_3703_),
    .A(net57),
    .Y(_3704_));
 sg13g2_o21ai_1 _8849_ (.B1(_3704_),
    .Y(_3705_),
    .A1(_3700_),
    .A2(_3701_));
 sg13g2_a221oi_1 _8850_ (.B2(_2405_),
    .C1(_3705_),
    .B1(_2727_),
    .A1(_2337_),
    .Y(_3706_),
    .A2(_2724_));
 sg13g2_a22oi_1 _8851_ (.Y(_3707_),
    .B1(_2710_),
    .B2(_2172_),
    .A2(_2320_),
    .A1(_2235_));
 sg13g2_o21ai_1 _8852_ (.B1(_2390_),
    .Y(_3708_),
    .A1(_2355_),
    .A2(_0832_));
 sg13g2_nand2_1 _8853_ (.Y(_3709_),
    .A(_1600_),
    .B(_2244_));
 sg13g2_o21ai_1 _8854_ (.B1(_3709_),
    .Y(_3710_),
    .A1(_2355_),
    .A2(_0861_));
 sg13g2_mux2_1 _8855_ (.A0(_3708_),
    .A1(_3710_),
    .S(net169),
    .X(_3711_));
 sg13g2_a21oi_1 _8856_ (.A1(_2406_),
    .A2(_2413_),
    .Y(_3712_),
    .B1(_3711_));
 sg13g2_o21ai_1 _8857_ (.B1(net57),
    .Y(_3713_),
    .A1(_2366_),
    .A2(_3382_));
 sg13g2_nand3b_1 _8858_ (.B(_3713_),
    .C(_2434_),
    .Y(_3714_),
    .A_N(_2428_));
 sg13g2_nor2_1 _8859_ (.A(net136),
    .B(net134),
    .Y(_3715_));
 sg13g2_a22oi_1 _8860_ (.Y(_3716_),
    .B1(_3715_),
    .B2(_2394_),
    .A2(net36),
    .A1(_2422_));
 sg13g2_a21o_1 _8861_ (.A2(_2036_),
    .A1(_0612_),
    .B1(_0854_),
    .X(_3717_));
 sg13g2_o21ai_1 _8862_ (.B1(_3717_),
    .Y(_3718_),
    .A1(_2036_),
    .A2(_2172_));
 sg13g2_a21oi_1 _8863_ (.A1(net52),
    .A2(net108),
    .Y(_3719_),
    .B1(_2739_));
 sg13g2_a21oi_1 _8864_ (.A1(_2299_),
    .A2(_1480_),
    .Y(_3721_),
    .B1(_3719_));
 sg13g2_o21ai_1 _8865_ (.B1(_2755_),
    .Y(_3722_),
    .A1(net192),
    .A2(_2766_));
 sg13g2_a22oi_1 _8866_ (.Y(_3723_),
    .B1(_3722_),
    .B2(_2629_),
    .A2(_3721_),
    .A1(_1451_));
 sg13g2_nand4_1 _8867_ (.B(_3716_),
    .C(_3718_),
    .A(_3714_),
    .Y(_3724_),
    .D(_3723_));
 sg13g2_a22oi_1 _8868_ (.Y(_3725_),
    .B1(_2308_),
    .B2(_1566_),
    .A2(net133),
    .A1(net83));
 sg13g2_nand2_1 _8869_ (.Y(_3726_),
    .A(net120),
    .B(net94));
 sg13g2_nand2_1 _8870_ (.Y(_3727_),
    .A(_2165_),
    .B(_3726_));
 sg13g2_o21ai_1 _8871_ (.B1(_2020_),
    .Y(_3728_),
    .A1(_0861_),
    .A2(_2136_));
 sg13g2_nand2b_1 _8872_ (.Y(_3729_),
    .B(_3728_),
    .A_N(_2743_));
 sg13g2_nand3b_1 _8873_ (.B(_3456_),
    .C(_2247_),
    .Y(_3730_),
    .A_N(_3729_));
 sg13g2_o21ai_1 _8874_ (.B1(_3730_),
    .Y(_3732_),
    .A1(_3725_),
    .A2(_3727_));
 sg13g2_nor2_1 _8875_ (.A(_3724_),
    .B(_3732_),
    .Y(_3733_));
 sg13g2_nand4_1 _8876_ (.B(_3707_),
    .C(_3712_),
    .A(_3706_),
    .Y(_3734_),
    .D(_3733_));
 sg13g2_o21ai_1 _8877_ (.B1(net81),
    .Y(_3735_),
    .A1(_2136_),
    .A2(_2284_));
 sg13g2_a21oi_1 _8878_ (.A1(net28),
    .A2(_3735_),
    .Y(_3736_),
    .B1(_2246_));
 sg13g2_a22oi_1 _8879_ (.Y(_3737_),
    .B1(_3726_),
    .B2(_2408_),
    .A2(net149),
    .A1(_2388_));
 sg13g2_nor2_1 _8880_ (.A(net53),
    .B(_2194_),
    .Y(_3738_));
 sg13g2_o21ai_1 _8881_ (.B1(_3738_),
    .Y(_3739_),
    .A1(_2683_),
    .A2(_3405_));
 sg13g2_o21ai_1 _8882_ (.B1(_3739_),
    .Y(_3740_),
    .A1(net43),
    .A2(_3737_));
 sg13g2_a221oi_1 _8883_ (.B2(_1452_),
    .C1(_2321_),
    .B1(_3703_),
    .A1(net61),
    .Y(_3741_),
    .A2(_2320_));
 sg13g2_or2_1 _8884_ (.X(_3743_),
    .B(_2676_),
    .A(net31));
 sg13g2_o21ai_1 _8885_ (.B1(_3743_),
    .Y(_3744_),
    .A1(net86),
    .A2(_3741_));
 sg13g2_nor4_1 _8886_ (.A(_3734_),
    .B(_3736_),
    .C(_3740_),
    .D(_3744_),
    .Y(_3745_));
 sg13g2_a21oi_1 _8887_ (.A1(_1571_),
    .A2(net79),
    .Y(_3746_),
    .B1(_2173_));
 sg13g2_nand2_1 _8888_ (.Y(_3747_),
    .A(_2194_),
    .B(net78));
 sg13g2_nand3_1 _8889_ (.B(_0834_),
    .C(_3747_),
    .A(net48),
    .Y(_3748_));
 sg13g2_o21ai_1 _8890_ (.B1(_3748_),
    .Y(_3749_),
    .A1(net169),
    .A2(_3746_));
 sg13g2_a21o_1 _8891_ (.A2(_2710_),
    .A1(_2036_),
    .B1(_2172_),
    .X(_3750_));
 sg13g2_nand3_1 _8892_ (.B(_2190_),
    .C(_3654_),
    .A(net192),
    .Y(_3751_));
 sg13g2_o21ai_1 _8893_ (.B1(_2395_),
    .Y(_3752_),
    .A1(net132),
    .A2(_2286_));
 sg13g2_nand2b_1 _8894_ (.Y(_3753_),
    .B(_2681_),
    .A_N(_2392_));
 sg13g2_nand2b_1 _8895_ (.Y(_3754_),
    .B(_3753_),
    .A_N(_3752_));
 sg13g2_nand2_1 _8896_ (.Y(_3755_),
    .A(_3751_),
    .B(_3754_));
 sg13g2_a221oi_1 _8897_ (.B2(net39),
    .C1(_3755_),
    .B1(_3750_),
    .A1(_2027_),
    .Y(_3756_),
    .A2(_3749_));
 sg13g2_nand2b_1 _8898_ (.Y(_3757_),
    .B(_2233_),
    .A_N(_2242_));
 sg13g2_o21ai_1 _8899_ (.B1(net221),
    .Y(_3758_),
    .A1(_1987_),
    .A2(net76));
 sg13g2_nand3_1 _8900_ (.B(_2266_),
    .C(_3758_),
    .A(_1482_),
    .Y(_3759_));
 sg13g2_nand3_1 _8901_ (.B(net76),
    .C(net75),
    .A(net36),
    .Y(_3760_));
 sg13g2_nand2_1 _8902_ (.Y(_3761_),
    .A(_2325_),
    .B(_3760_));
 sg13g2_o21ai_1 _8903_ (.B1(net75),
    .Y(_3762_),
    .A1(_2308_),
    .A2(_2325_));
 sg13g2_a22oi_1 _8904_ (.Y(_3764_),
    .B1(_3762_),
    .B2(net29),
    .A2(_3761_),
    .A1(_3433_));
 sg13g2_a21oi_1 _8905_ (.A1(_2267_),
    .A2(_3759_),
    .Y(_3765_),
    .B1(_3764_));
 sg13g2_nand4_1 _8906_ (.B(_3756_),
    .C(_3757_),
    .A(_3745_),
    .Y(_3766_),
    .D(_3765_));
 sg13g2_nor4_1 _8907_ (.A(_3674_),
    .B(_3692_),
    .C(_3698_),
    .D(_3766_),
    .Y(_3767_));
 sg13g2_o21ai_1 _8908_ (.B1(_3767_),
    .Y(_3768_),
    .A1(net51),
    .A2(_3665_));
 sg13g2_nor4_1 _8909_ (.A(_3490_),
    .B(_3646_),
    .C(_3647_),
    .D(_3768_),
    .Y(_3769_));
 sg13g2_a21oi_1 _8910_ (.A1(_2825_),
    .A2(_3488_),
    .Y(_3770_),
    .B1(_1888_));
 sg13g2_nand2b_1 _8911_ (.Y(_3771_),
    .B(_3359_),
    .A_N(_3770_));
 sg13g2_nand3_1 _8912_ (.B(_3769_),
    .C(_3771_),
    .A(_1597_),
    .Y(_3772_));
 sg13g2_nand2_1 _8913_ (.Y(_3773_),
    .A(net121),
    .B(net39));
 sg13g2_nand3_1 _8914_ (.B(net27),
    .C(_0877_),
    .A(net132),
    .Y(_3775_));
 sg13g2_nand3_1 _8915_ (.B(_3773_),
    .C(_3775_),
    .A(net183),
    .Y(_3776_));
 sg13g2_nor2_1 _8916_ (.A(net55),
    .B(_0903_),
    .Y(_3777_));
 sg13g2_o21ai_1 _8917_ (.B1(_3777_),
    .Y(_3778_),
    .A1(_0836_),
    .A2(_0826_));
 sg13g2_a21oi_1 _8918_ (.A1(_0836_),
    .A2(_3776_),
    .Y(_3779_),
    .B1(_3778_));
 sg13g2_nor4_1 _8919_ (.A(_2657_),
    .B(_3487_),
    .C(_3772_),
    .D(_3779_),
    .Y(_3780_));
 sg13g2_nor2_1 _8920_ (.A(_2642_),
    .B(_3780_),
    .Y(net10));
 sg13g2_nor3_1 _8921_ (.A(_1814_),
    .B(net24),
    .C(_1862_),
    .Y(_3781_));
 sg13g2_and2_1 _8922_ (.A(_1884_),
    .B(_1690_),
    .X(_3782_));
 sg13g2_o21ai_1 _8923_ (.B1(_3782_),
    .Y(_3783_),
    .A1(_1812_),
    .A2(_3781_));
 sg13g2_a21oi_1 _8924_ (.A1(_1743_),
    .A2(_3783_),
    .Y(_3784_),
    .B1(_2658_));
 sg13g2_nor2_1 _8925_ (.A(_1983_),
    .B(_1999_),
    .Y(_3785_));
 sg13g2_nor2_1 _8926_ (.A(_2550_),
    .B(_2788_),
    .Y(_3786_));
 sg13g2_nor2_1 _8927_ (.A(_2441_),
    .B(_3786_),
    .Y(_3787_));
 sg13g2_nand3_1 _8928_ (.B(_2278_),
    .C(_3672_),
    .A(net28),
    .Y(_3788_));
 sg13g2_a221oi_1 _8929_ (.B2(_2020_),
    .C1(_2275_),
    .B1(_3423_),
    .A1(_2018_),
    .Y(_3789_),
    .A2(_2286_));
 sg13g2_o21ai_1 _8930_ (.B1(_3695_),
    .Y(_3790_),
    .A1(_3693_),
    .A2(_3789_));
 sg13g2_nand2_1 _8931_ (.Y(_3791_),
    .A(_2291_),
    .B(_3790_));
 sg13g2_a22oi_1 _8932_ (.Y(_3792_),
    .B1(_3788_),
    .B2(_3791_),
    .A2(net72),
    .A1(_0865_));
 sg13g2_nand2_1 _8933_ (.Y(_3793_),
    .A(net301),
    .B(net2));
 sg13g2_o21ai_1 _8934_ (.B1(_3793_),
    .Y(_3795_),
    .A1(net301),
    .A2(_2840_));
 sg13g2_nand3_1 _8935_ (.B(_3633_),
    .C(_3795_),
    .A(net152),
    .Y(_3796_));
 sg13g2_nor2_1 _8936_ (.A(_2674_),
    .B(_2136_),
    .Y(_3797_));
 sg13g2_nor2_1 _8937_ (.A(net31),
    .B(_3797_),
    .Y(_3798_));
 sg13g2_o21ai_1 _8938_ (.B1(net108),
    .Y(_3799_),
    .A1(net72),
    .A2(_3798_));
 sg13g2_a21o_1 _8939_ (.A2(_3799_),
    .A1(_3796_),
    .B1(_2004_),
    .X(_3800_));
 sg13g2_a21oi_1 _8940_ (.A1(net92),
    .A2(_1566_),
    .Y(_3801_),
    .B1(_2313_));
 sg13g2_o21ai_1 _8941_ (.B1(net47),
    .Y(_3802_),
    .A1(_2340_),
    .A2(_2388_));
 sg13g2_nand2_1 _8942_ (.Y(_3803_),
    .A(_3801_),
    .B(_3802_));
 sg13g2_a21oi_1 _8943_ (.A1(net36),
    .A2(net37),
    .Y(_3804_),
    .B1(net111));
 sg13g2_nor2_1 _8944_ (.A(_2300_),
    .B(net162),
    .Y(_3806_));
 sg13g2_o21ai_1 _8945_ (.B1(net86),
    .Y(_3807_),
    .A1(_3702_),
    .A2(_3806_));
 sg13g2_o21ai_1 _8946_ (.B1(_3807_),
    .Y(_3808_),
    .A1(net45),
    .A2(_3804_));
 sg13g2_o21ai_1 _8947_ (.B1(_0862_),
    .Y(_3809_),
    .A1(net77),
    .A2(_2257_));
 sg13g2_a21oi_1 _8948_ (.A1(_2259_),
    .A2(_3809_),
    .Y(_3810_),
    .B1(_2412_));
 sg13g2_nand2b_1 _8949_ (.Y(_3811_),
    .B(_2699_),
    .A_N(_3810_));
 sg13g2_nand3_1 _8950_ (.B(_1576_),
    .C(_2706_),
    .A(net115),
    .Y(_3812_));
 sg13g2_o21ai_1 _8951_ (.B1(_0862_),
    .Y(_3813_),
    .A1(_2282_),
    .A2(_2690_));
 sg13g2_nand2_1 _8952_ (.Y(_3814_),
    .A(_3678_),
    .B(_3813_));
 sg13g2_nor3_1 _8953_ (.A(net91),
    .B(_2318_),
    .C(net72),
    .Y(_3815_));
 sg13g2_a22oi_1 _8954_ (.Y(_3817_),
    .B1(_3814_),
    .B2(_3815_),
    .A2(_2279_),
    .A1(_2593_));
 sg13g2_nor3_1 _8955_ (.A(_0893_),
    .B(net61),
    .C(_2151_),
    .Y(_3818_));
 sg13g2_o21ai_1 _8956_ (.B1(_2331_),
    .Y(_3819_),
    .A1(_2014_),
    .A2(net136));
 sg13g2_o21ai_1 _8957_ (.B1(_1527_),
    .Y(_3820_),
    .A1(_3818_),
    .A2(_3819_));
 sg13g2_nand4_1 _8958_ (.B(_3812_),
    .C(_3817_),
    .A(_3811_),
    .Y(_3821_),
    .D(_3820_));
 sg13g2_a221oi_1 _8959_ (.B2(_2320_),
    .C1(_3821_),
    .B1(_3808_),
    .A1(_3464_),
    .Y(_3822_),
    .A2(_3803_));
 sg13g2_a21oi_1 _8960_ (.A1(_2278_),
    .A2(_3671_),
    .Y(_3823_),
    .B1(net72));
 sg13g2_nor2_1 _8961_ (.A(_2743_),
    .B(_3823_),
    .Y(_3824_));
 sg13g2_inv_1 _8962_ (.Y(_3825_),
    .A(_2220_));
 sg13g2_inv_1 _8963_ (.Y(_3826_),
    .A(_2748_));
 sg13g2_a22oi_1 _8964_ (.Y(_3828_),
    .B1(_3826_),
    .B2(net135),
    .A2(_3825_),
    .A1(_2674_));
 sg13g2_o21ai_1 _8965_ (.B1(_2403_),
    .Y(_3829_),
    .A1(net151),
    .A2(_2714_));
 sg13g2_nor3_1 _8966_ (.A(net84),
    .B(net90),
    .C(_2308_),
    .Y(_3830_));
 sg13g2_nor2_1 _8967_ (.A(_2771_),
    .B(_3830_),
    .Y(_3831_));
 sg13g2_nor2_1 _8968_ (.A(_2257_),
    .B(_2314_),
    .Y(_3832_));
 sg13g2_o21ai_1 _8969_ (.B1(_3832_),
    .Y(_3833_),
    .A1(net72),
    .A2(_3456_));
 sg13g2_nand2_1 _8970_ (.Y(_3834_),
    .A(net46),
    .B(_3832_));
 sg13g2_a22oi_1 _8971_ (.Y(_3835_),
    .B1(_3834_),
    .B2(net61),
    .A2(_3833_),
    .A1(_3831_));
 sg13g2_a221oi_1 _8972_ (.B2(_2727_),
    .C1(_3835_),
    .B1(_3829_),
    .A1(_2395_),
    .Y(_3836_),
    .A2(_3753_));
 sg13g2_o21ai_1 _8973_ (.B1(_3836_),
    .Y(_3837_),
    .A1(net77),
    .A2(_3828_));
 sg13g2_o21ai_1 _8974_ (.B1(net36),
    .Y(_3839_),
    .A1(net76),
    .A2(net24));
 sg13g2_nor2b_1 _8975_ (.A(_2432_),
    .B_N(_2367_),
    .Y(_3840_));
 sg13g2_a21oi_1 _8976_ (.A1(_1587_),
    .A2(_3840_),
    .Y(_3841_),
    .B1(_3428_));
 sg13g2_nor4_1 _8977_ (.A(net74),
    .B(net78),
    .C(net120),
    .D(_2029_),
    .Y(_3842_));
 sg13g2_a21oi_1 _8978_ (.A1(_2372_),
    .A2(_2681_),
    .Y(_3843_),
    .B1(_3842_));
 sg13g2_o21ai_1 _8979_ (.B1(_3843_),
    .Y(_3844_),
    .A1(net24),
    .A2(_3841_));
 sg13g2_a21oi_1 _8980_ (.A1(_3703_),
    .A2(_3839_),
    .Y(_3845_),
    .B1(_3844_));
 sg13g2_inv_1 _8981_ (.Y(_3846_),
    .A(_3831_));
 sg13g2_a21oi_1 _8982_ (.A1(net97),
    .A2(_3702_),
    .Y(_3847_),
    .B1(net153));
 sg13g2_nor3_1 _8983_ (.A(net111),
    .B(_3415_),
    .C(_3847_),
    .Y(_3848_));
 sg13g2_a21oi_1 _8984_ (.A1(net133),
    .A2(_3846_),
    .Y(_3850_),
    .B1(_3848_));
 sg13g2_nand3_1 _8985_ (.B(_3845_),
    .C(_3850_),
    .A(_2425_),
    .Y(_3851_));
 sg13g2_nor4_1 _8986_ (.A(net169),
    .B(net110),
    .C(net74),
    .D(_2730_),
    .Y(_3852_));
 sg13g2_o21ai_1 _8987_ (.B1(net136),
    .Y(_3853_),
    .A1(_2400_),
    .A2(_3852_));
 sg13g2_nor3_1 _8988_ (.A(net74),
    .B(_0893_),
    .C(net94),
    .Y(_3854_));
 sg13g2_xnor2_1 _8989_ (.Y(_3855_),
    .A(net120),
    .B(net133));
 sg13g2_nand2_1 _8990_ (.Y(_3856_),
    .A(net116),
    .B(_3855_));
 sg13g2_nor3_1 _8991_ (.A(_2355_),
    .B(_2392_),
    .C(_2714_),
    .Y(_3857_));
 sg13g2_a221oi_1 _8992_ (.B2(_3856_),
    .C1(_3857_),
    .B1(_3854_),
    .A1(_2359_),
    .Y(_3858_),
    .A2(net111));
 sg13g2_and2_1 _8993_ (.A(_2012_),
    .B(_3425_),
    .X(_3859_));
 sg13g2_a22oi_1 _8994_ (.Y(_3860_),
    .B1(net109),
    .B2(_1571_),
    .A2(_0834_),
    .A1(_2388_));
 sg13g2_a22oi_1 _8995_ (.Y(_3861_),
    .B1(_2010_),
    .B2(_1576_),
    .A2(_1551_),
    .A1(_2340_));
 sg13g2_nand2b_1 _8996_ (.Y(_3862_),
    .B(net79),
    .A_N(_3861_));
 sg13g2_o21ai_1 _8997_ (.B1(_3862_),
    .Y(_3863_),
    .A1(net73),
    .A2(_3860_));
 sg13g2_nand4_1 _8998_ (.B(net83),
    .C(_1986_),
    .A(net47),
    .Y(_3864_),
    .D(_1573_));
 sg13g2_o21ai_1 _8999_ (.B1(_3864_),
    .Y(_3865_),
    .A1(_2246_),
    .A2(_2413_));
 sg13g2_a22oi_1 _9000_ (.Y(_3866_),
    .B1(_2386_),
    .B2(net88),
    .A2(_2035_),
    .A1(net110));
 sg13g2_nor2_1 _9001_ (.A(_2224_),
    .B(_3866_),
    .Y(_3867_));
 sg13g2_nand3_1 _9002_ (.B(_1451_),
    .C(_2321_),
    .A(net36),
    .Y(_3868_));
 sg13g2_o21ai_1 _9003_ (.B1(_3868_),
    .Y(_3869_),
    .A1(_2029_),
    .A2(_3867_));
 sg13g2_nor4_1 _9004_ (.A(_3859_),
    .B(_3863_),
    .C(_3865_),
    .D(_3869_),
    .Y(_3871_));
 sg13g2_o21ai_1 _9005_ (.B1(_1813_),
    .Y(_3872_),
    .A1(net120),
    .A2(_2010_));
 sg13g2_nand2_1 _9006_ (.Y(_3873_),
    .A(_1579_),
    .B(net134));
 sg13g2_nand3_1 _9007_ (.B(net79),
    .C(net75),
    .A(_1566_),
    .Y(_3874_));
 sg13g2_a21oi_1 _9008_ (.A1(_3872_),
    .A2(_3873_),
    .Y(_3875_),
    .B1(_3874_));
 sg13g2_o21ai_1 _9009_ (.B1(net57),
    .Y(_3876_),
    .A1(_1551_),
    .A2(_3702_));
 sg13g2_nand3b_1 _9010_ (.B(_2267_),
    .C(_3876_),
    .Y(_3877_),
    .A_N(_2240_));
 sg13g2_a21oi_1 _9011_ (.A1(_1813_),
    .A2(_2337_),
    .Y(_3878_),
    .B1(net94));
 sg13g2_nand2b_1 _9012_ (.Y(_3879_),
    .B(_2346_),
    .A_N(_3878_));
 sg13g2_nand4_1 _9013_ (.B(_1579_),
    .C(net75),
    .A(_2361_),
    .Y(_3880_),
    .D(_2722_));
 sg13g2_nor3_1 _9014_ (.A(_1538_),
    .B(net119),
    .C(_2298_),
    .Y(_3882_));
 sg13g2_nor2_1 _9015_ (.A(_2653_),
    .B(_3882_),
    .Y(_3883_));
 sg13g2_or2_1 _9016_ (.X(_3884_),
    .B(_3883_),
    .A(_2654_));
 sg13g2_nand4_1 _9017_ (.B(_3879_),
    .C(_3880_),
    .A(_3877_),
    .Y(_3885_),
    .D(_3884_));
 sg13g2_nor4_1 _9018_ (.A(net91),
    .B(net80),
    .C(net109),
    .D(net37),
    .Y(_3886_));
 sg13g2_nor4_1 _9019_ (.A(_3640_),
    .B(_3875_),
    .C(_3885_),
    .D(_3886_),
    .Y(_3887_));
 sg13g2_nand4_1 _9020_ (.B(_3858_),
    .C(_3871_),
    .A(_3853_),
    .Y(_3888_),
    .D(_3887_));
 sg13g2_nor4_1 _9021_ (.A(_3824_),
    .B(_3837_),
    .C(_3851_),
    .D(_3888_),
    .Y(_3889_));
 sg13g2_nand3_1 _9022_ (.B(_2027_),
    .C(_2036_),
    .A(_2141_),
    .Y(_3890_));
 sg13g2_o21ai_1 _9023_ (.B1(_3890_),
    .Y(_3891_),
    .A1(net121),
    .A2(_2390_));
 sg13g2_nor3_1 _9024_ (.A(net121),
    .B(_2265_),
    .C(_2390_),
    .Y(_3893_));
 sg13g2_a21o_1 _9025_ (.A2(_3891_),
    .A1(net29),
    .B1(_3893_),
    .X(_3894_));
 sg13g2_nor2_1 _9026_ (.A(_2670_),
    .B(_3806_),
    .Y(_3895_));
 sg13g2_o21ai_1 _9027_ (.B1(net37),
    .Y(_3896_),
    .A1(_1587_),
    .A2(_3895_));
 sg13g2_nand2b_1 _9028_ (.Y(_3897_),
    .B(_3896_),
    .A_N(_2428_));
 sg13g2_a21oi_1 _9029_ (.A1(net61),
    .A2(_2273_),
    .Y(_3898_),
    .B1(_2701_));
 sg13g2_nand2_1 _9030_ (.Y(_3899_),
    .A(_2406_),
    .B(net46));
 sg13g2_o21ai_1 _9031_ (.B1(_3690_),
    .Y(_3900_),
    .A1(_3898_),
    .A2(_3899_));
 sg13g2_a221oi_1 _9032_ (.B2(_2434_),
    .C1(_3900_),
    .B1(_3897_),
    .A1(_1986_),
    .Y(_3901_),
    .A2(_3894_));
 sg13g2_nand4_1 _9033_ (.B(_3822_),
    .C(_3889_),
    .A(_3800_),
    .Y(_3902_),
    .D(_3901_));
 sg13g2_a21oi_1 _9034_ (.A1(net192),
    .A2(_3580_),
    .Y(_3904_),
    .B1(_2273_));
 sg13g2_nor2b_1 _9035_ (.A(_3500_),
    .B_N(_3578_),
    .Y(_3905_));
 sg13g2_nand2b_1 _9036_ (.Y(_3906_),
    .B(_1149_),
    .A_N(_0831_));
 sg13g2_nor3_1 _9037_ (.A(net156),
    .B(_3905_),
    .C(_3906_),
    .Y(_3907_));
 sg13g2_a21oi_1 _9038_ (.A1(net156),
    .A2(net196),
    .Y(_3908_),
    .B1(_3907_));
 sg13g2_nand2_1 _9039_ (.Y(_3909_),
    .A(net245),
    .B(_2182_));
 sg13g2_o21ai_1 _9040_ (.B1(net216),
    .Y(_3910_),
    .A1(_2179_),
    .A2(_3909_));
 sg13g2_o21ai_1 _9041_ (.B1(net230),
    .Y(_3911_),
    .A1(_4110_),
    .A2(_2857_));
 sg13g2_a21o_1 _9042_ (.A2(_3911_),
    .A1(_2473_),
    .B1(_1438_),
    .X(_3912_));
 sg13g2_nand4_1 _9043_ (.B(net281),
    .C(_3578_),
    .A(net217),
    .Y(_3913_),
    .D(_3912_));
 sg13g2_nand3_1 _9044_ (.B(_4114_),
    .C(_3913_),
    .A(net170),
    .Y(_3914_));
 sg13g2_o21ai_1 _9045_ (.B1(_3914_),
    .Y(_3915_),
    .A1(_1040_),
    .A2(_3500_));
 sg13g2_a21oi_1 _9046_ (.A1(_3881_),
    .A2(_3915_),
    .Y(_3916_),
    .B1(_3906_));
 sg13g2_a21o_1 _9047_ (.A2(_3910_),
    .A1(net192),
    .B1(_3916_),
    .X(_3917_));
 sg13g2_nor2_1 _9048_ (.A(_1183_),
    .B(net196),
    .Y(_3918_));
 sg13g2_nand2_1 _9049_ (.Y(_3919_),
    .A(net156),
    .B(_3653_));
 sg13g2_a22oi_1 _9050_ (.Y(_3920_),
    .B1(_3919_),
    .B2(_0912_),
    .A2(_3918_),
    .A1(_3917_));
 sg13g2_mux2_1 _9051_ (.A0(_3908_),
    .A1(_3920_),
    .S(_0194_),
    .X(_3921_));
 sg13g2_a21oi_1 _9052_ (.A1(_3904_),
    .A2(_3921_),
    .Y(_3922_),
    .B1(_3464_));
 sg13g2_nor3_1 _9053_ (.A(net51),
    .B(_2160_),
    .C(_3922_),
    .Y(_3923_));
 sg13g2_mux2_1 _9054_ (.A0(net86),
    .A1(_2308_),
    .S(_3630_),
    .X(_3925_));
 sg13g2_nor4_1 _9055_ (.A(net53),
    .B(_2157_),
    .C(_1168_),
    .D(_3925_),
    .Y(_3926_));
 sg13g2_nor4_1 _9056_ (.A(_3792_),
    .B(_3902_),
    .C(_3923_),
    .D(_3926_),
    .Y(_3927_));
 sg13g2_nand2b_1 _9057_ (.Y(_3928_),
    .B(_3927_),
    .A_N(_2818_));
 sg13g2_nor4_1 _9058_ (.A(_3784_),
    .B(_3785_),
    .C(_3787_),
    .D(_3928_),
    .Y(_3929_));
 sg13g2_nand3_1 _9059_ (.B(net37),
    .C(_1976_),
    .A(net36),
    .Y(_3930_));
 sg13g2_a21oi_1 _9060_ (.A1(_1939_),
    .A2(_3930_),
    .Y(_3931_),
    .B1(_2661_));
 sg13g2_nand2b_1 _9061_ (.Y(_3932_),
    .B(_3782_),
    .A_N(_3931_));
 sg13g2_a22oi_1 _9062_ (.Y(_3933_),
    .B1(_3932_),
    .B2(_3359_),
    .A2(_3399_),
    .A1(_1522_));
 sg13g2_nand2_1 _9063_ (.Y(_3934_),
    .A(_3929_),
    .B(_3933_));
 sg13g2_nand3_1 _9064_ (.B(net136),
    .C(_0855_),
    .A(_0836_),
    .Y(_3936_));
 sg13g2_a21oi_1 _9065_ (.A1(_0827_),
    .A2(_3936_),
    .Y(_3937_),
    .B1(_0905_));
 sg13g2_nor2_1 _9066_ (.A(_3934_),
    .B(_3937_),
    .Y(_3938_));
 sg13g2_inv_1 _9067_ (.Y(_3939_),
    .A(_0727_));
 sg13g2_o21ai_1 _9068_ (.B1(_3939_),
    .Y(_3940_),
    .A1(_0824_),
    .A2(net14));
 sg13g2_a221oi_1 _9069_ (.B2(_0782_),
    .C1(_0766_),
    .B1(_3940_),
    .A1(_0727_),
    .Y(_3941_),
    .A2(_0784_));
 sg13g2_xor2_1 _9070_ (.B(_3941_),
    .A(_4387_),
    .X(_3942_));
 sg13g2_a21oi_1 _9071_ (.A1(net27),
    .A2(_2766_),
    .Y(_3943_),
    .B1(_1365_));
 sg13g2_o21ai_1 _9072_ (.B1(_3943_),
    .Y(_3944_),
    .A1(_3365_),
    .A2(_3942_));
 sg13g2_nor2_1 _9073_ (.A(_0824_),
    .B(_0758_),
    .Y(_3945_));
 sg13g2_a21oi_1 _9074_ (.A1(_0824_),
    .A2(_0801_),
    .Y(_3946_),
    .B1(_0736_));
 sg13g2_o21ai_1 _9075_ (.B1(_0781_),
    .Y(_3947_),
    .A1(_3939_),
    .A2(_0779_));
 sg13g2_nor3_1 _9076_ (.A(_3945_),
    .B(_3946_),
    .C(_3947_),
    .Y(_3948_));
 sg13g2_xnor2_1 _9077_ (.Y(_3949_),
    .A(_4387_),
    .B(_3948_));
 sg13g2_or3_1 _9078_ (.A(_2766_),
    .B(_3485_),
    .C(_3949_),
    .X(_3950_));
 sg13g2_nand2_1 _9079_ (.Y(_3951_),
    .A(net39),
    .B(_2766_));
 sg13g2_nand4_1 _9080_ (.B(_3944_),
    .C(_3950_),
    .A(_2755_),
    .Y(_3952_),
    .D(_3951_));
 sg13g2_a21oi_1 _9081_ (.A1(net39),
    .A2(_0912_),
    .Y(_3953_),
    .B1(_2352_));
 sg13g2_nor2_1 _9082_ (.A(net39),
    .B(_2643_),
    .Y(_3954_));
 sg13g2_a22oi_1 _9083_ (.Y(_3955_),
    .B1(_3954_),
    .B2(_3372_),
    .A2(_3953_),
    .A1(_3952_));
 sg13g2_a21oi_1 _9084_ (.A1(_3938_),
    .A2(_3955_),
    .Y(net11),
    .B1(_2642_));
 sg13g2_nand3_1 _9085_ (.B(net286),
    .C(_3653_),
    .A(net246),
    .Y(_3956_));
 sg13g2_o21ai_1 _9086_ (.B1(net156),
    .Y(_3957_),
    .A1(_2186_),
    .A2(_3956_));
 sg13g2_nand2_1 _9087_ (.Y(_3958_),
    .A(_2285_),
    .B(_3956_));
 sg13g2_o21ai_1 _9088_ (.B1(_3958_),
    .Y(_3959_),
    .A1(_1183_),
    .A2(_3956_));
 sg13g2_a21oi_1 _9089_ (.A1(_0809_),
    .A2(_3959_),
    .Y(_3960_),
    .B1(_2186_));
 sg13g2_a21oi_1 _9090_ (.A1(_1741_),
    .A2(_3957_),
    .Y(_3961_),
    .B1(_3960_));
 sg13g2_o21ai_1 _9091_ (.B1(_4114_),
    .Y(_3962_),
    .A1(_2177_),
    .A2(_4113_));
 sg13g2_a21oi_1 _9092_ (.A1(net248),
    .A2(_3962_),
    .Y(_3963_),
    .B1(net229));
 sg13g2_nor4_1 _9093_ (.A(_2273_),
    .B(_3659_),
    .C(_3961_),
    .D(_3963_),
    .Y(_3964_));
 sg13g2_o21ai_1 _9094_ (.B1(_2188_),
    .Y(_3966_),
    .A1(_3464_),
    .A2(_3964_));
 sg13g2_a22oi_1 _9095_ (.Y(_3967_),
    .B1(_3633_),
    .B2(_2219_),
    .A2(_2260_),
    .A1(net108));
 sg13g2_a21oi_1 _9096_ (.A1(_3966_),
    .A2(_3967_),
    .Y(_3968_),
    .B1(net51));
 sg13g2_a21oi_1 _9097_ (.A1(_0865_),
    .A2(net135),
    .Y(_3969_),
    .B1(_2257_));
 sg13g2_o21ai_1 _9098_ (.B1(net81),
    .Y(_3970_),
    .A1(_3797_),
    .A2(_3969_));
 sg13g2_a21oi_1 _9099_ (.A1(net28),
    .A2(_3970_),
    .Y(_3971_),
    .B1(_2398_));
 sg13g2_inv_1 _9100_ (.Y(_3972_),
    .A(_2172_));
 sg13g2_o21ai_1 _9101_ (.B1(_3405_),
    .Y(_3973_),
    .A1(_0834_),
    .A2(_0863_));
 sg13g2_a21oi_1 _9102_ (.A1(_2029_),
    .A2(_2172_),
    .Y(_3974_),
    .B1(_2402_));
 sg13g2_a21oi_1 _9103_ (.A1(_3972_),
    .A2(_3973_),
    .Y(_3975_),
    .B1(_3974_));
 sg13g2_nor3_1 _9104_ (.A(net119),
    .B(_2746_),
    .C(_3806_),
    .Y(_3977_));
 sg13g2_a21oi_1 _9105_ (.A1(_2306_),
    .A2(_3425_),
    .Y(_3978_),
    .B1(_3977_));
 sg13g2_a21oi_1 _9106_ (.A1(net27),
    .A2(_1168_),
    .Y(_3979_),
    .B1(_3978_));
 sg13g2_nand3_1 _9107_ (.B(net48),
    .C(_1482_),
    .A(_2340_),
    .Y(_3980_));
 sg13g2_nand3_1 _9108_ (.B(net36),
    .C(net75),
    .A(_2422_),
    .Y(_3981_));
 sg13g2_a22oi_1 _9109_ (.Y(_3982_),
    .B1(net97),
    .B2(_2653_),
    .A2(net83),
    .A1(_1526_));
 sg13g2_o21ai_1 _9110_ (.B1(_2771_),
    .Y(_3983_),
    .A1(net109),
    .A2(net75));
 sg13g2_o21ai_1 _9111_ (.B1(_3983_),
    .Y(_3984_),
    .A1(net153),
    .A2(_3982_));
 sg13g2_a21oi_1 _9112_ (.A1(_2012_),
    .A2(_2325_),
    .Y(_3985_),
    .B1(_3984_));
 sg13g2_nand4_1 _9113_ (.B(_3980_),
    .C(_3981_),
    .A(_3752_),
    .Y(_3986_),
    .D(_3985_));
 sg13g2_o21ai_1 _9114_ (.B1(_2413_),
    .Y(_3988_),
    .A1(_2595_),
    .A2(_3424_));
 sg13g2_nor3_1 _9115_ (.A(_0623_),
    .B(net56),
    .C(_2301_),
    .Y(_3989_));
 sg13g2_nand3_1 _9116_ (.B(_2710_),
    .C(_3989_),
    .A(_2379_),
    .Y(_3990_));
 sg13g2_nand3b_1 _9117_ (.B(net92),
    .C(_2369_),
    .Y(_3991_),
    .A_N(_1573_));
 sg13g2_nand3_1 _9118_ (.B(_1573_),
    .C(_2727_),
    .A(net136),
    .Y(_3992_));
 sg13g2_nand4_1 _9119_ (.B(_3990_),
    .C(_3991_),
    .A(_3988_),
    .Y(_3993_),
    .D(_3992_));
 sg13g2_nor4_1 _9120_ (.A(_3975_),
    .B(_3979_),
    .C(_3986_),
    .D(_3993_),
    .Y(_3994_));
 sg13g2_o21ai_1 _9121_ (.B1(_1548_),
    .Y(_3995_),
    .A1(_2408_),
    .A2(_1576_));
 sg13g2_a21oi_1 _9122_ (.A1(_1991_),
    .A2(_3995_),
    .Y(_3996_),
    .B1(_1540_));
 sg13g2_nor2_1 _9123_ (.A(_1991_),
    .B(_2012_),
    .Y(_3997_));
 sg13g2_a21oi_1 _9124_ (.A1(net83),
    .A2(_1580_),
    .Y(_3999_),
    .B1(_3997_));
 sg13g2_nor3_1 _9125_ (.A(_2608_),
    .B(_2303_),
    .C(_3999_),
    .Y(_4000_));
 sg13g2_nor2_1 _9126_ (.A(_2220_),
    .B(_2697_),
    .Y(_4001_));
 sg13g2_nor2_1 _9127_ (.A(_3709_),
    .B(_2681_),
    .Y(_4002_));
 sg13g2_nor4_1 _9128_ (.A(_3996_),
    .B(_4000_),
    .C(_4001_),
    .D(_4002_),
    .Y(_4003_));
 sg13g2_nor2_1 _9129_ (.A(net114),
    .B(_1539_),
    .Y(_4004_));
 sg13g2_a22oi_1 _9130_ (.Y(_4005_),
    .B1(_2682_),
    .B2(_2355_),
    .A2(_0863_),
    .A1(_0832_));
 sg13g2_a21oi_1 _9131_ (.A1(_0623_),
    .A2(_2301_),
    .Y(_4006_),
    .B1(_2390_));
 sg13g2_nor4_1 _9132_ (.A(_2265_),
    .B(_4004_),
    .C(_4005_),
    .D(_4006_),
    .Y(_4007_));
 sg13g2_a21oi_1 _9133_ (.A1(_2386_),
    .A2(net149),
    .Y(_4008_),
    .B1(_4007_));
 sg13g2_a22oi_1 _9134_ (.Y(_4010_),
    .B1(net151),
    .B2(_1571_),
    .A2(_0834_),
    .A1(_2369_));
 sg13g2_nor2_1 _9135_ (.A(net43),
    .B(_4010_),
    .Y(_4011_));
 sg13g2_a22oi_1 _9136_ (.Y(_4012_),
    .B1(_2320_),
    .B2(_3873_),
    .A2(net153),
    .A1(_2359_));
 sg13g2_nor2_1 _9137_ (.A(_2241_),
    .B(_4012_),
    .Y(_4013_));
 sg13g2_nor2_1 _9138_ (.A(net31),
    .B(_3729_),
    .Y(_4014_));
 sg13g2_nor4_1 _9139_ (.A(_4008_),
    .B(_4011_),
    .C(_4013_),
    .D(_4014_),
    .Y(_4015_));
 sg13g2_a221oi_1 _9140_ (.B2(_3424_),
    .C1(_2036_),
    .B1(_2247_),
    .A1(_2595_),
    .Y(_4016_),
    .A2(_2208_));
 sg13g2_o21ai_1 _9141_ (.B1(_1558_),
    .Y(_4017_),
    .A1(net110),
    .A2(_2418_));
 sg13g2_nand2_1 _9142_ (.Y(_4018_),
    .A(net48),
    .B(_4017_));
 sg13g2_a22oi_1 _9143_ (.Y(_4019_),
    .B1(_4016_),
    .B2(_4018_),
    .A2(_2037_),
    .A1(net45));
 sg13g2_a21oi_1 _9144_ (.A1(_1365_),
    .A2(_3654_),
    .Y(_4021_),
    .B1(_2189_));
 sg13g2_a21oi_1 _9145_ (.A1(net151),
    .A2(_2289_),
    .Y(_4022_),
    .B1(_2420_));
 sg13g2_nor2b_1 _9146_ (.A(_4022_),
    .B_N(_3738_),
    .Y(_4023_));
 sg13g2_nand2_1 _9147_ (.Y(_4024_),
    .A(net76),
    .B(_2697_));
 sg13g2_nor3_1 _9148_ (.A(net91),
    .B(_2318_),
    .C(_2216_),
    .Y(_4025_));
 sg13g2_o21ai_1 _9149_ (.B1(net109),
    .Y(_4026_),
    .A1(net262),
    .A2(_2262_));
 sg13g2_nand3_1 _9150_ (.B(net151),
    .C(_4026_),
    .A(_1482_),
    .Y(_4027_));
 sg13g2_a22oi_1 _9151_ (.Y(_4028_),
    .B1(_4027_),
    .B2(_2267_),
    .A2(_4025_),
    .A1(_4024_));
 sg13g2_o21ai_1 _9152_ (.B1(net97),
    .Y(_4029_),
    .A1(net116),
    .A2(_1342_));
 sg13g2_o21ai_1 _9153_ (.B1(_4029_),
    .Y(_4030_),
    .A1(net61),
    .A2(net111));
 sg13g2_nand2_1 _9154_ (.Y(_4032_),
    .A(_2233_),
    .B(_4030_));
 sg13g2_nand3_1 _9155_ (.B(_4028_),
    .C(_4032_),
    .A(_2741_),
    .Y(_4033_));
 sg13g2_nor4_1 _9156_ (.A(_4019_),
    .B(_4021_),
    .C(_4023_),
    .D(_4033_),
    .Y(_4034_));
 sg13g2_nand4_1 _9157_ (.B(_4003_),
    .C(_4015_),
    .A(_3994_),
    .Y(_4035_),
    .D(_4034_));
 sg13g2_o21ai_1 _9158_ (.B1(net28),
    .Y(_4036_),
    .A1(_2314_),
    .A2(_3456_));
 sg13g2_o21ai_1 _9159_ (.B1(_2675_),
    .Y(_4037_),
    .A1(_2234_),
    .A2(net28));
 sg13g2_nand2_1 _9160_ (.Y(_4038_),
    .A(_2246_),
    .B(_4037_));
 sg13g2_o21ai_1 _9161_ (.B1(_4038_),
    .Y(_4039_),
    .A1(_3798_),
    .A2(_4036_));
 sg13g2_a21oi_1 _9162_ (.A1(_2302_),
    .A2(_2674_),
    .Y(_4040_),
    .B1(_3667_));
 sg13g2_o21ai_1 _9163_ (.B1(_3671_),
    .Y(_4041_),
    .A1(_2147_),
    .A2(_4040_));
 sg13g2_nand3_1 _9164_ (.B(_2699_),
    .C(_4041_),
    .A(net28),
    .Y(_4043_));
 sg13g2_a21o_1 _9165_ (.A2(_2277_),
    .A1(_2303_),
    .B1(_2697_),
    .X(_4044_));
 sg13g2_a21oi_1 _9166_ (.A1(net162),
    .A2(_2669_),
    .Y(_4045_),
    .B1(_1587_));
 sg13g2_o21ai_1 _9167_ (.B1(net37),
    .Y(_4046_),
    .A1(_3382_),
    .A2(_4045_));
 sg13g2_a22oi_1 _9168_ (.Y(_4047_),
    .B1(_4046_),
    .B2(_2434_),
    .A2(_4044_),
    .A1(_2406_));
 sg13g2_nand3_1 _9169_ (.B(_4043_),
    .C(_4047_),
    .A(_4039_),
    .Y(_4048_));
 sg13g2_nor4_1 _9170_ (.A(_3968_),
    .B(_3971_),
    .C(_4035_),
    .D(_4048_),
    .Y(_4049_));
 sg13g2_o21ai_1 _9171_ (.B1(_4049_),
    .Y(_4050_),
    .A1(_2441_),
    .A2(_3476_));
 sg13g2_nor2_1 _9172_ (.A(_3646_),
    .B(_4050_),
    .Y(_4051_));
 sg13g2_o21ai_1 _9173_ (.B1(_3399_),
    .Y(_4052_),
    .A1(net30),
    .A2(_1522_));
 sg13g2_nand2_1 _9174_ (.Y(_4054_),
    .A(_4051_),
    .B(_4052_));
 sg13g2_nor3_1 _9175_ (.A(_0812_),
    .B(net121),
    .C(_3369_),
    .Y(_4055_));
 sg13g2_nor2_1 _9176_ (.A(_3778_),
    .B(_4055_),
    .Y(_4056_));
 sg13g2_nor3_1 _9177_ (.A(_3398_),
    .B(_4054_),
    .C(_4056_),
    .Y(_4057_));
 sg13g2_nand2_1 _9178_ (.Y(_4058_),
    .A(_3950_),
    .B(_3951_));
 sg13g2_nor2b_1 _9179_ (.A(_3944_),
    .B_N(_3963_),
    .Y(_4059_));
 sg13g2_o21ai_1 _9180_ (.B1(_2353_),
    .Y(_4060_),
    .A1(_4058_),
    .A2(_4059_));
 sg13g2_a21oi_1 _9181_ (.A1(_4057_),
    .A2(_4060_),
    .Y(net12),
    .B1(_2642_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \counter[0]$_SDFFE_PP0P__333  (.L_HI(net333));
 sg13g2_buf_1 _9184_ (.A(net317),
    .X(uio_oe[0]));
 sg13g2_buf_1 _9185_ (.A(net318),
    .X(uio_oe[1]));
 sg13g2_buf_1 _9186_ (.A(net319),
    .X(uio_oe[2]));
 sg13g2_buf_1 _9187_ (.A(net320),
    .X(uio_oe[3]));
 sg13g2_buf_1 _9188_ (.A(net321),
    .X(uio_oe[4]));
 sg13g2_buf_1 _9189_ (.A(net322),
    .X(uio_oe[5]));
 sg13g2_buf_1 _9190_ (.A(net323),
    .X(uio_oe[6]));
 sg13g2_buf_1 _9191_ (.A(net324),
    .X(uio_oe[7]));
 sg13g2_buf_1 _9192_ (.A(net325),
    .X(uio_out[0]));
 sg13g2_buf_1 _9193_ (.A(net326),
    .X(uio_out[1]));
 sg13g2_buf_1 _9194_ (.A(net327),
    .X(uio_out[2]));
 sg13g2_buf_1 _9195_ (.A(net328),
    .X(uio_out[3]));
 sg13g2_buf_1 _9196_ (.A(net329),
    .X(uio_out[4]));
 sg13g2_buf_1 _9197_ (.A(net330),
    .X(uio_out[5]));
 sg13g2_buf_1 _9198_ (.A(net331),
    .X(uio_out[6]));
 sg13g2_buf_1 _9199_ (.A(net332),
    .X(uio_out[7]));
 sg13g2_buf_1 _9200_ (.A(\hvsync_gen.vsync ),
    .X(net9));
 sg13g2_buf_1 _9201_ (.A(hsync),
    .X(net13));
 sg13g2_dfrbp_1 \counter[0]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net333),
    .D(_0024_),
    .Q_N(_4599_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net334),
    .D(_0025_),
    .Q_N(_4598_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net335),
    .D(_0026_),
    .Q_N(_0019_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net336),
    .D(_0027_),
    .Q_N(_0020_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net337),
    .D(_0028_),
    .Q_N(_4597_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net338),
    .D(_0029_),
    .Q_N(_0021_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFFE_PP0P_  (.CLK(counter_clk),
    .RESET_B(net339),
    .D(_0030_),
    .Q_N(_4596_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net340),
    .D(_0031_),
    .Q_N(_0023_),
    .Q(\flag.flag_abrosexual_inst.pix_x[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net341),
    .D(_0032_),
    .Q_N(_0018_),
    .Q(\flag.flag_abrosexual_inst.pix_x[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net342),
    .D(_0033_),
    .Q_N(_0017_),
    .Q(\flag.flag_abrosexual_inst.pix_x[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net343),
    .D(_0034_),
    .Q_N(_0016_),
    .Q(\flag.flag_abrosexual_inst.pix_x[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net344),
    .D(_0035_),
    .Q_N(_0014_),
    .Q(\flag.flag_abrosexual_inst.pix_x[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net345),
    .D(_0036_),
    .Q_N(_0013_),
    .Q(\flag.flag_abrosexual_inst.pix_x[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net346),
    .D(_0037_),
    .Q_N(_0012_),
    .Q(\flag.flag_abrosexual_inst.pix_x[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net347),
    .D(_0038_),
    .Q_N(_0011_),
    .Q(\flag.flag_abrosexual_inst.pix_x[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net348),
    .D(_0039_),
    .Q_N(_0007_),
    .Q(\flag.flag_abrosexual_inst.pix_x[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net349),
    .D(_0040_),
    .Q_N(_0004_),
    .Q(\flag.flag_abrosexual_inst.pix_x[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net350),
    .D(_0000_),
    .Q_N(_4595_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net351),
    .D(_0041_),
    .Q_N(_0022_),
    .Q(\flag.flag_abrosexual_inst.pix_y[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net352),
    .D(_0042_),
    .Q_N(_0015_),
    .Q(\flag.flag_abrosexual_inst.pix_y[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net353),
    .D(_0043_),
    .Q_N(_0008_),
    .Q(\flag.flag_abrosexual_inst.pix_y[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net354),
    .D(_0044_),
    .Q_N(_0002_),
    .Q(\flag.flag_abrosexual_inst.pix_y[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net355),
    .D(_0045_),
    .Q_N(_0009_),
    .Q(\flag.flag_abrosexual_inst.pix_y[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net356),
    .D(_0046_),
    .Q_N(_0003_),
    .Q(\flag.flag_abrosexual_inst.pix_y[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net357),
    .D(_0047_),
    .Q_N(_0006_),
    .Q(\flag.flag_abrosexual_inst.pix_y[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net358),
    .D(_0048_),
    .Q_N(_0010_),
    .Q(\flag.flag_abrosexual_inst.pix_y[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net359),
    .D(_0049_),
    .Q_N(_0005_),
    .Q(\flag.flag_abrosexual_inst.pix_y[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net360),
    .D(_0050_),
    .Q_N(_4600_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net361),
    .D(_0001_),
    .Q_N(_4594_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_buf_1 input1 (.A(uio_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(uio_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(uio_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(uio_in[6]),
    .X(net5));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[0]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[1]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[2]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[3]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[4]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[5]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[6]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout14 (.A(_0734_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1175_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_2957_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1103_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_1100_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_1064_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1756_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1061_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1020_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1678_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1548_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1015_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_2866_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2303_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2248_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_2234_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2151_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2147_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2048_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1637_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1635_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1608_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1580_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1452_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1342_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0865_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1643_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2966_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_2915_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2608_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2472_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2302_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2247_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2169_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2166_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2060_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2047_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2004_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_1600_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1595_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1579_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1559_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1540_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1451_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1341_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1016_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0943_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0863_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0295_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_4350_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_4244_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_4214_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2666_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2967_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_2916_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2903_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_2887_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_2854_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_2412_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_2328_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2324_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2323_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_2301_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_2282_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_2223_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_2165_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_2157_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_2145_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2099_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2006_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2003_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1991_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_1814_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_1631_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_1594_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_1577_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1558_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1539_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1527_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1383_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1168_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0971_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0958_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0862_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_0420_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_0173_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_4399_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_4246_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_4235_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_4213_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_4175_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_3029_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_2889_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_2879_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2379_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2300_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_2295_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_2241_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2192_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2045_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_2014_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_1997_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_1813_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1658_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1630_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1602_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0861_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0854_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0141_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_4557_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_4280_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_4248_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_4206_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_4174_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_4146_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_4142_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_4097_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_2831_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_2418_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_2306_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_2299_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_2284_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_1986_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_1603_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_4473_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_4432_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_4264_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_4261_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_4219_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_4217_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_4208_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_4192_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_4154_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_4145_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_4096_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_2265_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_2032_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_2027_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_1555_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_1552_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_0932_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_0896_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_0859_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_4191_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_4153_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_4072_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_3482_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_3531_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_1481_),
    .X(net162));
 sg13g2_buf_2 fanout163 (.A(_0858_),
    .X(net163));
 sg13g2_buf_2 fanout164 (.A(_4512_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_4402_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_4136_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_4071_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_3471_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_0623_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_0194_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_1495_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_1420_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_1145_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0857_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_0849_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_4228_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_4162_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_3816_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_3731_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_3568_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_3460_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_2250_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_2141_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_2033_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_1741_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_0722_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_0689_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_0612_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_0370_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_0183_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_1407_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_1365_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_1357_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_1196_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_1183_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_0912_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_4134_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_4087_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_3805_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_3720_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_3557_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_3514_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_3503_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_3449_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_2184_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_1925_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_1806_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_1730_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_1708_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_1697_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_1512_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_1479_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_1292_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_1248_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_1204_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_1051_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_0930_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_0809_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_0711_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_0458_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_0414_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_0359_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_0172_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_0095_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_1467_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_1344_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_0922_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_0911_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_0808_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_0592_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_0441_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_0230_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_0145_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_3881_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_3590_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_3546_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_3438_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_3364_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_1468_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_1391_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_1358_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_1193_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_1095_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_1084_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_1073_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_1040_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_0919_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_0864_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_0798_),
    .X(net249));
 sg13g2_buf_4 fanout250 (.X(net250),
    .A(_0700_));
 sg13g2_buf_2 fanout251 (.A(_0667_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_0590_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_0568_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_0447_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_0436_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_0403_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_0348_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_0315_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_0161_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_0128_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_0084_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_2528_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_1717_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_1437_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_0608_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_0394_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_4527_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_4525_),
    .X(net268));
 sg13g2_buf_2 fanout269 (.A(_4389_),
    .X(net269));
 sg13g2_buf_2 fanout270 (.A(_4315_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_4221_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_4078_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_3579_),
    .X(net273));
 sg13g2_buf_2 fanout274 (.A(_3353_),
    .X(net274));
 sg13g2_buf_2 fanout275 (.A(_1457_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_1380_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_1347_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_1270_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_1226_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_1182_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_1149_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_0985_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_0963_),
    .X(net283));
 sg13g2_buf_2 fanout284 (.A(_0908_),
    .X(net284));
 sg13g2_buf_2 fanout285 (.A(_0886_),
    .X(net285));
 sg13g2_buf_2 fanout286 (.A(_0853_),
    .X(net286));
 sg13g2_buf_2 fanout287 (.A(_0831_),
    .X(net287));
 sg13g2_buf_2 fanout288 (.A(_0656_),
    .X(net288));
 sg13g2_buf_2 fanout289 (.A(_0480_),
    .X(net289));
 sg13g2_buf_2 fanout290 (.A(_0392_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_0337_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_0304_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_0227_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_0150_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_0117_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_0073_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0051_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_1483_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_1080_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_0883_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_0881_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_4423_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_4388_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_4114_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_4073_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_1446_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_1369_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_0974_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_0952_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0875_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_0842_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_0776_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_0381_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_0293_),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(_0062_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_4583_),
    .X(net316));
 sg13g2_tielo _9184__317 (.L_LO(net317));
 sg13g2_tielo _9185__318 (.L_LO(net318));
 sg13g2_tielo _9186__319 (.L_LO(net319));
 sg13g2_tielo _9187__320 (.L_LO(net320));
 sg13g2_tielo _9188__321 (.L_LO(net321));
 sg13g2_tielo _9189__322 (.L_LO(net322));
 sg13g2_tielo _9190__323 (.L_LO(net323));
 sg13g2_tielo _9191__324 (.L_LO(net324));
 sg13g2_tielo _9192__325 (.L_LO(net325));
 sg13g2_tielo _9193__326 (.L_LO(net326));
 sg13g2_tielo _9194__327 (.L_LO(net327));
 sg13g2_tielo _9195__328 (.L_LO(net328));
 sg13g2_tielo _9196__329 (.L_LO(net329));
 sg13g2_tielo _9197__330 (.L_LO(net330));
 sg13g2_tielo _9198__331 (.L_LO(net331));
 sg13g2_tielo _9199__332 (.L_LO(net332));
 sg13g2_tiehi \counter[1]$_SDFFE_PP0P__334  (.L_HI(net334));
 sg13g2_tiehi \counter[2]$_SDFFE_PP0P__335  (.L_HI(net335));
 sg13g2_tiehi \counter[3]$_SDFFE_PP0P__336  (.L_HI(net336));
 sg13g2_tiehi \counter[4]$_SDFFE_PP0P__337  (.L_HI(net337));
 sg13g2_tiehi \counter[5]$_SDFFE_PP0P__338  (.L_HI(net338));
 sg13g2_tiehi \counter[6]$_SDFFE_PP0P__339  (.L_HI(net339));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__340  (.L_HI(net340));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__341  (.L_HI(net341));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__342  (.L_HI(net342));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__343  (.L_HI(net343));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__344  (.L_HI(net344));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__345  (.L_HI(net345));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__346  (.L_HI(net346));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__347  (.L_HI(net347));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__348  (.L_HI(net348));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__349  (.L_HI(net349));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__350  (.L_HI(net350));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__351  (.L_HI(net351));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__352  (.L_HI(net352));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__353  (.L_HI(net353));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__354  (.L_HI(net354));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__355  (.L_HI(net355));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__356  (.L_HI(net356));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__357  (.L_HI(net357));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__358  (.L_HI(net358));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__359  (.L_HI(net359));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__360  (.L_HI(net360));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__361  (.L_HI(net361));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_3356_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(_3356_));
 sg13g2_antennanp ANTENNA_4 (.A(clk));
 sg13g2_antennanp ANTENNA_5 (.A(_3356_));
 sg13g2_antennanp ANTENNA_6 (.A(clk));
 sg13g2_antennanp ANTENNA_7 (.A(_3356_));
 sg13g2_antennanp ANTENNA_8 (.A(clk));
 sg13g2_antennanp ANTENNA_9 (.A(_3356_));
 sg13g2_antennanp ANTENNA_10 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_fill_2 FILLER_0_133 ();
 sg13g2_fill_1 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_148 ();
 sg13g2_fill_2 FILLER_0_155 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_191 ();
 sg13g2_fill_2 FILLER_0_198 ();
 sg13g2_fill_1 FILLER_0_200 ();
 sg13g2_fill_1 FILLER_0_218 ();
 sg13g2_fill_1 FILLER_0_223 ();
 sg13g2_fill_2 FILLER_0_242 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_279 ();
 sg13g2_fill_1 FILLER_0_289 ();
 sg13g2_fill_1 FILLER_0_314 ();
 sg13g2_fill_1 FILLER_0_366 ();
 sg13g2_fill_1 FILLER_0_379 ();
 sg13g2_fill_2 FILLER_0_385 ();
 sg13g2_fill_2 FILLER_0_397 ();
 sg13g2_fill_1 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_153 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_fill_1 FILLER_1_163 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_4 FILLER_1_189 ();
 sg13g2_fill_1 FILLER_1_232 ();
 sg13g2_decap_4 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_262 ();
 sg13g2_fill_1 FILLER_1_278 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_289 ();
 sg13g2_fill_1 FILLER_1_302 ();
 sg13g2_fill_2 FILLER_1_359 ();
 sg13g2_fill_1 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_395 ();
 sg13g2_fill_1 FILLER_1_411 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_fill_2 FILLER_2_98 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_fill_1 FILLER_2_119 ();
 sg13g2_fill_2 FILLER_2_128 ();
 sg13g2_fill_1 FILLER_2_130 ();
 sg13g2_fill_1 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_204 ();
 sg13g2_fill_1 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_233 ();
 sg13g2_fill_2 FILLER_2_247 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_fill_1 FILLER_2_315 ();
 sg13g2_fill_1 FILLER_2_327 ();
 sg13g2_fill_2 FILLER_2_368 ();
 sg13g2_fill_1 FILLER_2_380 ();
 sg13g2_fill_1 FILLER_2_402 ();
 sg13g2_fill_1 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_2_414 ();
 sg13g2_decap_8 FILLER_2_418 ();
 sg13g2_decap_4 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_fill_2 FILLER_3_63 ();
 sg13g2_fill_1 FILLER_3_65 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_118 ();
 sg13g2_fill_2 FILLER_3_127 ();
 sg13g2_fill_1 FILLER_3_129 ();
 sg13g2_fill_1 FILLER_3_147 ();
 sg13g2_fill_1 FILLER_3_207 ();
 sg13g2_fill_1 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_237 ();
 sg13g2_fill_1 FILLER_3_239 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_274 ();
 sg13g2_fill_1 FILLER_3_317 ();
 sg13g2_fill_1 FILLER_3_324 ();
 sg13g2_fill_2 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_163 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_fill_1 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_fill_2 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_303 ();
 sg13g2_fill_2 FILLER_4_314 ();
 sg13g2_fill_1 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_1 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_62 ();
 sg13g2_fill_2 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_112 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_fill_2 FILLER_5_179 ();
 sg13g2_fill_1 FILLER_5_196 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_220 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_fill_1 FILLER_5_237 ();
 sg13g2_decap_4 FILLER_5_248 ();
 sg13g2_fill_2 FILLER_5_310 ();
 sg13g2_fill_1 FILLER_5_312 ();
 sg13g2_fill_1 FILLER_5_322 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_fill_2 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_418 ();
 sg13g2_decap_4 FILLER_5_425 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_4 FILLER_6_42 ();
 sg13g2_fill_1 FILLER_6_46 ();
 sg13g2_fill_1 FILLER_6_69 ();
 sg13g2_fill_1 FILLER_6_85 ();
 sg13g2_fill_2 FILLER_6_122 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_fill_2 FILLER_6_190 ();
 sg13g2_fill_2 FILLER_6_197 ();
 sg13g2_fill_1 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_263 ();
 sg13g2_fill_1 FILLER_6_270 ();
 sg13g2_fill_1 FILLER_6_276 ();
 sg13g2_fill_1 FILLER_6_303 ();
 sg13g2_fill_1 FILLER_6_309 ();
 sg13g2_fill_1 FILLER_6_322 ();
 sg13g2_fill_2 FILLER_6_351 ();
 sg13g2_fill_1 FILLER_6_353 ();
 sg13g2_fill_2 FILLER_6_370 ();
 sg13g2_fill_1 FILLER_6_372 ();
 sg13g2_fill_1 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_decap_4 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_fill_1 FILLER_7_80 ();
 sg13g2_decap_4 FILLER_7_93 ();
 sg13g2_fill_1 FILLER_7_97 ();
 sg13g2_fill_1 FILLER_7_107 ();
 sg13g2_fill_2 FILLER_7_113 ();
 sg13g2_fill_1 FILLER_7_122 ();
 sg13g2_fill_1 FILLER_7_198 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_fill_1 FILLER_7_410 ();
 sg13g2_decap_8 FILLER_7_416 ();
 sg13g2_decap_8 FILLER_7_423 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_4 FILLER_8_42 ();
 sg13g2_fill_2 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_65 ();
 sg13g2_fill_1 FILLER_8_71 ();
 sg13g2_fill_1 FILLER_8_78 ();
 sg13g2_fill_2 FILLER_8_87 ();
 sg13g2_fill_1 FILLER_8_110 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_fill_1 FILLER_8_229 ();
 sg13g2_decap_4 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_245 ();
 sg13g2_fill_1 FILLER_8_250 ();
 sg13g2_fill_1 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_263 ();
 sg13g2_fill_1 FILLER_8_268 ();
 sg13g2_fill_1 FILLER_8_279 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_decap_4 FILLER_8_299 ();
 sg13g2_fill_1 FILLER_8_303 ();
 sg13g2_fill_1 FILLER_8_312 ();
 sg13g2_fill_1 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_1 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_fill_2 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_89 ();
 sg13g2_fill_1 FILLER_9_99 ();
 sg13g2_fill_1 FILLER_9_136 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_172 ();
 sg13g2_fill_1 FILLER_9_211 ();
 sg13g2_fill_2 FILLER_9_247 ();
 sg13g2_fill_1 FILLER_9_255 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_fill_1 FILLER_9_324 ();
 sg13g2_fill_2 FILLER_9_335 ();
 sg13g2_fill_1 FILLER_9_337 ();
 sg13g2_fill_1 FILLER_9_348 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_409 ();
 sg13g2_fill_1 FILLER_9_411 ();
 sg13g2_decap_8 FILLER_9_416 ();
 sg13g2_decap_8 FILLER_9_423 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_48 ();
 sg13g2_fill_1 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_91 ();
 sg13g2_fill_1 FILLER_10_97 ();
 sg13g2_fill_1 FILLER_10_108 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_fill_1 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_146 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_167 ();
 sg13g2_fill_1 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_fill_2 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_fill_2 FILLER_10_230 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_321 ();
 sg13g2_fill_2 FILLER_10_330 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_fill_1 FILLER_10_382 ();
 sg13g2_fill_2 FILLER_10_390 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_fill_2 FILLER_10_428 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_58 ();
 sg13g2_fill_2 FILLER_11_91 ();
 sg13g2_fill_2 FILLER_11_98 ();
 sg13g2_fill_2 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_111 ();
 sg13g2_fill_1 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_138 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_fill_1 FILLER_11_163 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_2 FILLER_11_259 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_320 ();
 sg13g2_fill_1 FILLER_11_336 ();
 sg13g2_fill_1 FILLER_11_342 ();
 sg13g2_fill_2 FILLER_11_372 ();
 sg13g2_fill_1 FILLER_11_374 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_32 ();
 sg13g2_fill_2 FILLER_12_57 ();
 sg13g2_fill_1 FILLER_12_81 ();
 sg13g2_fill_2 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_fill_1 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_160 ();
 sg13g2_decap_4 FILLER_12_210 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_fill_2 FILLER_12_342 ();
 sg13g2_fill_1 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_fill_1 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_12_414 ();
 sg13g2_decap_8 FILLER_12_421 ();
 sg13g2_fill_2 FILLER_12_428 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_77 ();
 sg13g2_fill_1 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_2 FILLER_13_129 ();
 sg13g2_fill_1 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_169 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_fill_1 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_372 ();
 sg13g2_fill_1 FILLER_13_381 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_225 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_fill_1 FILLER_14_251 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_fill_1 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_267 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_fill_2 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_298 ();
 sg13g2_fill_1 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_352 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_2 FILLER_14_388 ();
 sg13g2_fill_1 FILLER_14_394 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_fill_2 FILLER_14_427 ();
 sg13g2_fill_1 FILLER_14_429 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_28 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_fill_1 FILLER_15_122 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_160 ();
 sg13g2_fill_1 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_decap_4 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_15_188 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_289 ();
 sg13g2_fill_2 FILLER_15_340 ();
 sg13g2_fill_1 FILLER_15_342 ();
 sg13g2_fill_2 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_280 ();
 sg13g2_fill_2 FILLER_16_329 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_fill_2 FILLER_16_384 ();
 sg13g2_fill_1 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_28 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_fill_1 FILLER_17_122 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_142 ();
 sg13g2_fill_1 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_188 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_fill_1 FILLER_17_237 ();
 sg13g2_fill_1 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_fill_2 FILLER_17_384 ();
 sg13g2_fill_2 FILLER_17_401 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_4 FILLER_17_424 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_fill_1 FILLER_18_101 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_2 FILLER_18_123 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_18_211 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_252 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_276 ();
 sg13g2_fill_2 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_1 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_363 ();
 sg13g2_fill_1 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_186 ();
 sg13g2_fill_1 FILLER_19_192 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_fill_2 FILLER_19_233 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_291 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_330 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_decap_4 FILLER_19_388 ();
 sg13g2_fill_2 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_fill_2 FILLER_19_427 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_decap_4 FILLER_20_35 ();
 sg13g2_fill_1 FILLER_20_53 ();
 sg13g2_fill_2 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_107 ();
 sg13g2_fill_1 FILLER_20_114 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_fill_1 FILLER_20_131 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_229 ();
 sg13g2_decap_4 FILLER_20_242 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_1 FILLER_20_251 ();
 sg13g2_fill_1 FILLER_20_279 ();
 sg13g2_fill_1 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_decap_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_20_383 ();
 sg13g2_fill_1 FILLER_20_392 ();
 sg13g2_fill_2 FILLER_20_397 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_fill_2 FILLER_20_427 ();
 sg13g2_fill_1 FILLER_20_429 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_4 FILLER_21_21 ();
 sg13g2_fill_2 FILLER_21_25 ();
 sg13g2_fill_1 FILLER_21_128 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_192 ();
 sg13g2_fill_2 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_2 FILLER_21_217 ();
 sg13g2_fill_1 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_233 ();
 sg13g2_fill_2 FILLER_21_238 ();
 sg13g2_fill_1 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_258 ();
 sg13g2_fill_1 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_380 ();
 sg13g2_fill_1 FILLER_21_401 ();
 sg13g2_decap_8 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_416 ();
 sg13g2_decap_8 FILLER_21_423 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_56 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_fill_2 FILLER_22_105 ();
 sg13g2_fill_2 FILLER_22_127 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_175 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_2 FILLER_22_196 ();
 sg13g2_fill_2 FILLER_22_203 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_248 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_261 ();
 sg13g2_decap_4 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_280 ();
 sg13g2_fill_1 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_297 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_2 FILLER_22_345 ();
 sg13g2_fill_1 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_fill_1 FILLER_22_390 ();
 sg13g2_fill_2 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_415 ();
 sg13g2_decap_8 FILLER_22_422 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_51 ();
 sg13g2_fill_1 FILLER_23_64 ();
 sg13g2_fill_1 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_fill_2 FILLER_23_341 ();
 sg13g2_decap_4 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_4 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_1 FILLER_24_24 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_fill_1 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_81 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_2 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_235 ();
 sg13g2_fill_2 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_4 FILLER_24_275 ();
 sg13g2_fill_2 FILLER_24_279 ();
 sg13g2_fill_1 FILLER_24_287 ();
 sg13g2_fill_1 FILLER_24_292 ();
 sg13g2_fill_2 FILLER_24_297 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_2 FILLER_24_358 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_decap_4 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_414 ();
 sg13g2_decap_8 FILLER_24_421 ();
 sg13g2_fill_2 FILLER_24_428 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_18 ();
 sg13g2_fill_2 FILLER_25_46 ();
 sg13g2_fill_1 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_54 ();
 sg13g2_fill_1 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_68 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_97 ();
 sg13g2_fill_1 FILLER_25_160 ();
 sg13g2_fill_2 FILLER_25_165 ();
 sg13g2_fill_1 FILLER_25_175 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_289 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_327 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_341 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_354 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_2 FILLER_25_397 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_418 ();
 sg13g2_decap_4 FILLER_25_425 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_31 ();
 sg13g2_fill_1 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_50 ();
 sg13g2_fill_1 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_170 ();
 sg13g2_decap_4 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_202 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_223 ();
 sg13g2_fill_1 FILLER_26_239 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_303 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_343 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_4 FILLER_26_424 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_23 ();
 sg13g2_fill_2 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_157 ();
 sg13g2_fill_2 FILLER_27_169 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_232 ();
 sg13g2_fill_2 FILLER_27_237 ();
 sg13g2_fill_1 FILLER_27_239 ();
 sg13g2_fill_2 FILLER_27_244 ();
 sg13g2_decap_4 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_303 ();
 sg13g2_fill_1 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_320 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_fill_1 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_355 ();
 sg13g2_fill_2 FILLER_27_367 ();
 sg13g2_fill_1 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_378 ();
 sg13g2_fill_1 FILLER_27_384 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_fill_2 FILLER_27_404 ();
 sg13g2_decap_8 FILLER_27_412 ();
 sg13g2_decap_8 FILLER_27_419 ();
 sg13g2_decap_4 FILLER_27_426 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_fill_2 FILLER_28_78 ();
 sg13g2_fill_1 FILLER_28_80 ();
 sg13g2_fill_2 FILLER_28_115 ();
 sg13g2_decap_4 FILLER_28_122 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_1 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_1 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_113 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_237 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_decap_4 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_2 FILLER_29_300 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_145 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_173 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_291 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_1 FILLER_30_323 ();
 sg13g2_fill_2 FILLER_30_333 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_2 FILLER_30_403 ();
 sg13g2_fill_1 FILLER_30_412 ();
 sg13g2_decap_8 FILLER_30_416 ();
 sg13g2_decap_8 FILLER_30_423 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_1 FILLER_31_36 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_66 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_decap_4 FILLER_31_89 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_136 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_fill_2 FILLER_31_192 ();
 sg13g2_fill_1 FILLER_31_194 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_262 ();
 sg13g2_fill_1 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_294 ();
 sg13g2_fill_1 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_312 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_1 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_1 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_71 ();
 sg13g2_fill_1 FILLER_32_82 ();
 sg13g2_fill_1 FILLER_32_92 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_123 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_2 FILLER_32_167 ();
 sg13g2_fill_1 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_217 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_decap_4 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_418 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_2 FILLER_33_14 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_fill_1 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_136 ();
 sg13g2_fill_2 FILLER_33_203 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_262 ();
 sg13g2_fill_1 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_284 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_decap_4 FILLER_33_304 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_1 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_386 ();
 sg13g2_decap_4 FILLER_33_396 ();
 sg13g2_fill_2 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_412 ();
 sg13g2_decap_8 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_2 FILLER_34_37 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_162 ();
 sg13g2_fill_1 FILLER_34_171 ();
 sg13g2_fill_2 FILLER_34_186 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_248 ();
 sg13g2_fill_2 FILLER_34_264 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_422 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_decap_4 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_47 ();
 sg13g2_fill_1 FILLER_35_61 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_117 ();
 sg13g2_fill_1 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_170 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_1 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_1 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_333 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_385 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_414 ();
 sg13g2_decap_8 FILLER_35_421 ();
 sg13g2_fill_2 FILLER_35_428 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_227 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_fill_1 FILLER_36_277 ();
 sg13g2_decap_4 FILLER_36_283 ();
 sg13g2_decap_4 FILLER_36_291 ();
 sg13g2_fill_1 FILLER_36_299 ();
 sg13g2_fill_1 FILLER_36_324 ();
 sg13g2_fill_2 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_4 FILLER_36_424 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_4 FILLER_37_42 ();
 sg13g2_fill_1 FILLER_37_46 ();
 sg13g2_fill_1 FILLER_37_71 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_288 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_342 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_410 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_159 ();
 sg13g2_fill_2 FILLER_38_183 ();
 sg13g2_fill_1 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_fill_2 FILLER_38_241 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_fill_2 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_298 ();
 sg13g2_fill_2 FILLER_38_310 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_decap_4 FILLER_38_400 ();
 sg13g2_fill_1 FILLER_38_404 ();
 sg13g2_decap_4 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_4 FILLER_38_424 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_44 ();
 sg13g2_fill_1 FILLER_39_50 ();
 sg13g2_fill_1 FILLER_39_55 ();
 sg13g2_fill_1 FILLER_39_60 ();
 sg13g2_fill_1 FILLER_39_65 ();
 sg13g2_fill_2 FILLER_39_83 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_fill_1 FILLER_39_120 ();
 sg13g2_fill_1 FILLER_39_125 ();
 sg13g2_fill_1 FILLER_39_160 ();
 sg13g2_fill_2 FILLER_39_183 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_285 ();
 sg13g2_fill_1 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_321 ();
 sg13g2_fill_1 FILLER_39_350 ();
 sg13g2_fill_1 FILLER_39_367 ();
 sg13g2_fill_2 FILLER_39_376 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_390 ();
 sg13g2_decap_4 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_415 ();
 sg13g2_decap_8 FILLER_39_422 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_4 FILLER_40_42 ();
 sg13g2_fill_1 FILLER_40_46 ();
 sg13g2_fill_2 FILLER_40_60 ();
 sg13g2_fill_2 FILLER_40_68 ();
 sg13g2_fill_1 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_2 FILLER_40_113 ();
 sg13g2_fill_1 FILLER_40_115 ();
 sg13g2_fill_1 FILLER_40_134 ();
 sg13g2_fill_2 FILLER_40_151 ();
 sg13g2_fill_2 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_227 ();
 sg13g2_fill_2 FILLER_40_234 ();
 sg13g2_fill_2 FILLER_40_267 ();
 sg13g2_fill_1 FILLER_40_269 ();
 sg13g2_fill_2 FILLER_40_307 ();
 sg13g2_fill_2 FILLER_40_313 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_fill_1 FILLER_40_332 ();
 sg13g2_fill_2 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_fill_2 FILLER_40_365 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_fill_1 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_fill_2 FILLER_41_42 ();
 sg13g2_fill_1 FILLER_41_48 ();
 sg13g2_fill_1 FILLER_41_54 ();
 sg13g2_fill_1 FILLER_41_67 ();
 sg13g2_fill_1 FILLER_41_73 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_1 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_115 ();
 sg13g2_fill_1 FILLER_41_137 ();
 sg13g2_fill_1 FILLER_41_162 ();
 sg13g2_fill_1 FILLER_41_167 ();
 sg13g2_fill_2 FILLER_41_180 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_fill_2 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_236 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_decap_4 FILLER_41_263 ();
 sg13g2_fill_2 FILLER_41_275 ();
 sg13g2_fill_1 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_314 ();
 sg13g2_fill_1 FILLER_41_326 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_348 ();
 sg13g2_fill_1 FILLER_41_358 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_41_414 ();
 sg13g2_decap_8 FILLER_41_421 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_53 ();
 sg13g2_fill_2 FILLER_42_78 ();
 sg13g2_fill_1 FILLER_42_80 ();
 sg13g2_fill_1 FILLER_42_103 ();
 sg13g2_fill_2 FILLER_42_135 ();
 sg13g2_fill_2 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_171 ();
 sg13g2_fill_1 FILLER_42_207 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_284 ();
 sg13g2_fill_1 FILLER_42_291 ();
 sg13g2_fill_1 FILLER_42_297 ();
 sg13g2_fill_2 FILLER_42_313 ();
 sg13g2_fill_1 FILLER_42_339 ();
 sg13g2_decap_4 FILLER_42_347 ();
 sg13g2_fill_1 FILLER_42_351 ();
 sg13g2_fill_1 FILLER_42_362 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_fill_1 FILLER_42_400 ();
 sg13g2_decap_8 FILLER_42_411 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_decap_4 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_4 FILLER_43_42 ();
 sg13g2_fill_1 FILLER_43_46 ();
 sg13g2_fill_1 FILLER_43_52 ();
 sg13g2_fill_2 FILLER_43_59 ();
 sg13g2_fill_1 FILLER_43_66 ();
 sg13g2_fill_2 FILLER_43_73 ();
 sg13g2_fill_1 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_140 ();
 sg13g2_fill_1 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_158 ();
 sg13g2_fill_2 FILLER_43_168 ();
 sg13g2_fill_2 FILLER_43_186 ();
 sg13g2_fill_1 FILLER_43_202 ();
 sg13g2_fill_1 FILLER_43_207 ();
 sg13g2_fill_1 FILLER_43_215 ();
 sg13g2_fill_1 FILLER_43_220 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_247 ();
 sg13g2_fill_1 FILLER_43_258 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_295 ();
 sg13g2_fill_1 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_340 ();
 sg13g2_fill_2 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_388 ();
 sg13g2_decap_8 FILLER_43_421 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_2 FILLER_44_59 ();
 sg13g2_fill_1 FILLER_44_61 ();
 sg13g2_fill_1 FILLER_44_94 ();
 sg13g2_fill_1 FILLER_44_107 ();
 sg13g2_fill_2 FILLER_44_154 ();
 sg13g2_fill_1 FILLER_44_164 ();
 sg13g2_fill_2 FILLER_44_180 ();
 sg13g2_fill_2 FILLER_44_192 ();
 sg13g2_fill_1 FILLER_44_194 ();
 sg13g2_fill_1 FILLER_44_206 ();
 sg13g2_fill_1 FILLER_44_212 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_decap_4 FILLER_44_246 ();
 sg13g2_fill_1 FILLER_44_250 ();
 sg13g2_fill_2 FILLER_44_263 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_274 ();
 sg13g2_fill_2 FILLER_44_304 ();
 sg13g2_fill_1 FILLER_44_306 ();
 sg13g2_fill_1 FILLER_44_326 ();
 sg13g2_fill_1 FILLER_44_352 ();
 sg13g2_decap_4 FILLER_44_357 ();
 sg13g2_fill_2 FILLER_44_361 ();
 sg13g2_fill_2 FILLER_44_378 ();
 sg13g2_fill_2 FILLER_44_412 ();
 sg13g2_decap_8 FILLER_44_418 ();
 sg13g2_decap_4 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_fill_2 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_104 ();
 sg13g2_fill_1 FILLER_45_118 ();
 sg13g2_fill_1 FILLER_45_142 ();
 sg13g2_fill_1 FILLER_45_147 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_fill_1 FILLER_45_194 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_fill_2 FILLER_45_228 ();
 sg13g2_fill_2 FILLER_45_234 ();
 sg13g2_fill_2 FILLER_45_245 ();
 sg13g2_fill_2 FILLER_45_276 ();
 sg13g2_fill_1 FILLER_45_278 ();
 sg13g2_fill_1 FILLER_45_294 ();
 sg13g2_fill_1 FILLER_45_327 ();
 sg13g2_fill_1 FILLER_45_343 ();
 sg13g2_fill_2 FILLER_45_352 ();
 sg13g2_fill_1 FILLER_45_354 ();
 sg13g2_fill_2 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_416 ();
 sg13g2_decap_8 FILLER_45_423 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_1 FILLER_46_83 ();
 sg13g2_fill_2 FILLER_46_97 ();
 sg13g2_fill_1 FILLER_46_109 ();
 sg13g2_fill_1 FILLER_46_118 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_fill_1 FILLER_46_189 ();
 sg13g2_fill_1 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_254 ();
 sg13g2_fill_2 FILLER_46_276 ();
 sg13g2_decap_4 FILLER_46_288 ();
 sg13g2_fill_2 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_345 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_decap_4 FILLER_46_372 ();
 sg13g2_fill_1 FILLER_46_379 ();
 sg13g2_fill_2 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_fill_2 FILLER_46_427 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_4 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_39 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_fill_1 FILLER_47_59 ();
 sg13g2_fill_1 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_74 ();
 sg13g2_fill_2 FILLER_47_79 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_1 FILLER_47_153 ();
 sg13g2_decap_4 FILLER_47_158 ();
 sg13g2_fill_1 FILLER_47_162 ();
 sg13g2_fill_1 FILLER_47_184 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_fill_2 FILLER_47_257 ();
 sg13g2_fill_2 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_decap_8 FILLER_47_409 ();
 sg13g2_decap_8 FILLER_47_416 ();
 sg13g2_decap_8 FILLER_47_423 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_37 ();
 sg13g2_fill_1 FILLER_48_48 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_114 ();
 sg13g2_fill_1 FILLER_48_121 ();
 sg13g2_decap_4 FILLER_48_132 ();
 sg13g2_fill_1 FILLER_48_141 ();
 sg13g2_fill_1 FILLER_48_152 ();
 sg13g2_fill_1 FILLER_48_157 ();
 sg13g2_fill_2 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_fill_1 FILLER_48_170 ();
 sg13g2_fill_1 FILLER_48_175 ();
 sg13g2_fill_2 FILLER_48_186 ();
 sg13g2_fill_1 FILLER_48_188 ();
 sg13g2_fill_2 FILLER_48_224 ();
 sg13g2_fill_1 FILLER_48_263 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_fill_1 FILLER_48_315 ();
 sg13g2_decap_4 FILLER_48_324 ();
 sg13g2_fill_2 FILLER_48_340 ();
 sg13g2_fill_1 FILLER_48_342 ();
 sg13g2_fill_2 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_349 ();
 sg13g2_fill_2 FILLER_48_380 ();
 sg13g2_fill_1 FILLER_48_389 ();
 sg13g2_fill_2 FILLER_48_398 ();
 sg13g2_decap_8 FILLER_48_408 ();
 sg13g2_decap_8 FILLER_48_415 ();
 sg13g2_decap_8 FILLER_48_422 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_64 ();
 sg13g2_fill_1 FILLER_49_71 ();
 sg13g2_fill_1 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_fill_1 FILLER_49_114 ();
 sg13g2_fill_2 FILLER_49_144 ();
 sg13g2_fill_1 FILLER_49_146 ();
 sg13g2_fill_2 FILLER_49_152 ();
 sg13g2_fill_1 FILLER_49_217 ();
 sg13g2_fill_1 FILLER_49_228 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_246 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_287 ();
 sg13g2_fill_1 FILLER_49_289 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_2 FILLER_49_324 ();
 sg13g2_fill_2 FILLER_49_339 ();
 sg13g2_fill_1 FILLER_49_350 ();
 sg13g2_decap_4 FILLER_49_375 ();
 sg13g2_fill_2 FILLER_49_384 ();
 sg13g2_fill_1 FILLER_49_389 ();
 sg13g2_fill_1 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_405 ();
 sg13g2_decap_8 FILLER_49_412 ();
 sg13g2_decap_8 FILLER_49_419 ();
 sg13g2_decap_4 FILLER_49_426 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_37 ();
 sg13g2_fill_1 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_decap_4 FILLER_50_68 ();
 sg13g2_fill_2 FILLER_50_126 ();
 sg13g2_fill_1 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_161 ();
 sg13g2_fill_2 FILLER_50_168 ();
 sg13g2_fill_1 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_181 ();
 sg13g2_fill_1 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_2 FILLER_50_231 ();
 sg13g2_fill_2 FILLER_50_242 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_353 ();
 sg13g2_fill_1 FILLER_50_359 ();
 sg13g2_decap_8 FILLER_50_365 ();
 sg13g2_decap_8 FILLER_50_372 ();
 sg13g2_decap_8 FILLER_50_379 ();
 sg13g2_decap_8 FILLER_50_386 ();
 sg13g2_decap_8 FILLER_50_393 ();
 sg13g2_decap_8 FILLER_50_400 ();
 sg13g2_decap_8 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_50_414 ();
 sg13g2_decap_8 FILLER_50_421 ();
 sg13g2_fill_2 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_4 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_39 ();
 sg13g2_fill_2 FILLER_51_99 ();
 sg13g2_fill_1 FILLER_51_106 ();
 sg13g2_fill_1 FILLER_51_115 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_134 ();
 sg13g2_fill_2 FILLER_51_146 ();
 sg13g2_fill_1 FILLER_51_148 ();
 sg13g2_fill_1 FILLER_51_196 ();
 sg13g2_decap_4 FILLER_51_203 ();
 sg13g2_fill_1 FILLER_51_207 ();
 sg13g2_fill_1 FILLER_51_220 ();
 sg13g2_decap_4 FILLER_51_246 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_1 FILLER_51_257 ();
 sg13g2_fill_2 FILLER_51_353 ();
 sg13g2_fill_2 FILLER_51_359 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_decap_8 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_51_414 ();
 sg13g2_decap_8 FILLER_51_421 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_4 FILLER_52_28 ();
 sg13g2_fill_2 FILLER_52_32 ();
 sg13g2_fill_2 FILLER_52_57 ();
 sg13g2_fill_1 FILLER_52_64 ();
 sg13g2_fill_2 FILLER_52_110 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_124 ();
 sg13g2_fill_1 FILLER_52_166 ();
 sg13g2_fill_2 FILLER_52_171 ();
 sg13g2_fill_1 FILLER_52_206 ();
 sg13g2_fill_1 FILLER_52_212 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_258 ();
 sg13g2_decap_4 FILLER_52_274 ();
 sg13g2_fill_1 FILLER_52_278 ();
 sg13g2_fill_2 FILLER_52_293 ();
 sg13g2_decap_4 FILLER_52_321 ();
 sg13g2_fill_1 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_365 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_fill_2 FILLER_52_427 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_4 FILLER_53_28 ();
 sg13g2_fill_2 FILLER_53_32 ();
 sg13g2_fill_1 FILLER_53_57 ();
 sg13g2_fill_1 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_75 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_1 FILLER_53_141 ();
 sg13g2_fill_1 FILLER_53_161 ();
 sg13g2_fill_1 FILLER_53_166 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_fill_1 FILLER_53_234 ();
 sg13g2_fill_1 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_267 ();
 sg13g2_fill_2 FILLER_53_328 ();
 sg13g2_fill_2 FILLER_53_362 ();
 sg13g2_fill_1 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_376 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_decap_8 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_397 ();
 sg13g2_decap_8 FILLER_53_404 ();
 sg13g2_decap_8 FILLER_53_411 ();
 sg13g2_decap_8 FILLER_53_418 ();
 sg13g2_decap_4 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_fill_2 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_fill_1 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_1 FILLER_54_104 ();
 sg13g2_fill_1 FILLER_54_182 ();
 sg13g2_fill_2 FILLER_54_194 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_229 ();
 sg13g2_fill_2 FILLER_54_235 ();
 sg13g2_fill_1 FILLER_54_264 ();
 sg13g2_fill_2 FILLER_54_348 ();
 sg13g2_fill_1 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_369 ();
 sg13g2_decap_8 FILLER_54_376 ();
 sg13g2_decap_8 FILLER_54_383 ();
 sg13g2_decap_8 FILLER_54_390 ();
 sg13g2_decap_8 FILLER_54_397 ();
 sg13g2_decap_8 FILLER_54_404 ();
 sg13g2_decap_8 FILLER_54_411 ();
 sg13g2_decap_8 FILLER_54_418 ();
 sg13g2_decap_4 FILLER_54_425 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_fill_2 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_fill_1 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_61 ();
 sg13g2_fill_1 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_fill_1 FILLER_55_120 ();
 sg13g2_fill_2 FILLER_55_126 ();
 sg13g2_fill_1 FILLER_55_136 ();
 sg13g2_fill_1 FILLER_55_142 ();
 sg13g2_fill_1 FILLER_55_148 ();
 sg13g2_fill_1 FILLER_55_159 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_fill_1 FILLER_55_176 ();
 sg13g2_fill_1 FILLER_55_217 ();
 sg13g2_fill_1 FILLER_55_222 ();
 sg13g2_fill_1 FILLER_55_228 ();
 sg13g2_fill_1 FILLER_55_234 ();
 sg13g2_fill_1 FILLER_55_239 ();
 sg13g2_fill_2 FILLER_55_245 ();
 sg13g2_fill_2 FILLER_55_256 ();
 sg13g2_fill_1 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_347 ();
 sg13g2_decap_8 FILLER_55_372 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_55_414 ();
 sg13g2_decap_8 FILLER_55_421 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_decap_4 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_96 ();
 sg13g2_fill_1 FILLER_56_109 ();
 sg13g2_fill_2 FILLER_56_118 ();
 sg13g2_fill_2 FILLER_56_133 ();
 sg13g2_fill_1 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_148 ();
 sg13g2_fill_2 FILLER_56_172 ();
 sg13g2_fill_1 FILLER_56_182 ();
 sg13g2_fill_1 FILLER_56_197 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_212 ();
 sg13g2_fill_1 FILLER_56_229 ();
 sg13g2_fill_2 FILLER_56_235 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_1 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_300 ();
 sg13g2_fill_2 FILLER_56_361 ();
 sg13g2_fill_1 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_376 ();
 sg13g2_decap_8 FILLER_56_383 ();
 sg13g2_decap_8 FILLER_56_390 ();
 sg13g2_decap_8 FILLER_56_397 ();
 sg13g2_decap_8 FILLER_56_404 ();
 sg13g2_decap_8 FILLER_56_411 ();
 sg13g2_decap_8 FILLER_56_418 ();
 sg13g2_decap_4 FILLER_56_425 ();
 sg13g2_fill_1 FILLER_56_429 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_4 FILLER_57_35 ();
 sg13g2_fill_1 FILLER_57_100 ();
 sg13g2_fill_1 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_172 ();
 sg13g2_fill_2 FILLER_57_219 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_fill_1 FILLER_57_238 ();
 sg13g2_fill_1 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_fill_2 FILLER_57_264 ();
 sg13g2_fill_2 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_308 ();
 sg13g2_fill_1 FILLER_57_315 ();
 sg13g2_fill_2 FILLER_57_321 ();
 sg13g2_fill_1 FILLER_57_323 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_fill_2 FILLER_57_427 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_4 FILLER_58_35 ();
 sg13g2_fill_1 FILLER_58_78 ();
 sg13g2_fill_2 FILLER_58_94 ();
 sg13g2_fill_1 FILLER_58_96 ();
 sg13g2_fill_2 FILLER_58_148 ();
 sg13g2_fill_1 FILLER_58_150 ();
 sg13g2_fill_2 FILLER_58_156 ();
 sg13g2_fill_1 FILLER_58_168 ();
 sg13g2_decap_4 FILLER_58_173 ();
 sg13g2_fill_2 FILLER_58_229 ();
 sg13g2_fill_1 FILLER_58_235 ();
 sg13g2_decap_8 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_401 ();
 sg13g2_decap_8 FILLER_58_408 ();
 sg13g2_decap_8 FILLER_58_415 ();
 sg13g2_decap_8 FILLER_58_422 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_fill_2 FILLER_59_35 ();
 sg13g2_fill_1 FILLER_59_37 ();
 sg13g2_fill_1 FILLER_59_90 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_104 ();
 sg13g2_fill_2 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_131 ();
 sg13g2_fill_1 FILLER_59_138 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_1 FILLER_59_158 ();
 sg13g2_fill_1 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_220 ();
 sg13g2_fill_2 FILLER_59_230 ();
 sg13g2_fill_1 FILLER_59_241 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_fill_1 FILLER_59_276 ();
 sg13g2_fill_1 FILLER_59_282 ();
 sg13g2_fill_2 FILLER_59_288 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_314 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_fill_2 FILLER_59_396 ();
 sg13g2_fill_2 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_59_412 ();
 sg13g2_decap_8 FILLER_59_419 ();
 sg13g2_decap_4 FILLER_59_426 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_35 ();
 sg13g2_decap_4 FILLER_60_41 ();
 sg13g2_fill_1 FILLER_60_49 ();
 sg13g2_fill_2 FILLER_60_102 ();
 sg13g2_fill_1 FILLER_60_108 ();
 sg13g2_fill_1 FILLER_60_138 ();
 sg13g2_fill_1 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_167 ();
 sg13g2_fill_2 FILLER_60_173 ();
 sg13g2_fill_1 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_261 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_fill_1 FILLER_60_291 ();
 sg13g2_fill_2 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_312 ();
 sg13g2_fill_2 FILLER_60_319 ();
 sg13g2_fill_2 FILLER_60_395 ();
 sg13g2_fill_2 FILLER_60_401 ();
 sg13g2_decap_8 FILLER_60_415 ();
 sg13g2_decap_8 FILLER_60_422 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_fill_2 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_127 ();
 sg13g2_fill_1 FILLER_61_129 ();
 sg13g2_fill_1 FILLER_61_234 ();
 sg13g2_fill_1 FILLER_61_240 ();
 sg13g2_fill_1 FILLER_61_245 ();
 sg13g2_fill_1 FILLER_61_274 ();
 sg13g2_fill_2 FILLER_61_304 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_fill_2 FILLER_61_351 ();
 sg13g2_fill_1 FILLER_61_353 ();
 sg13g2_fill_1 FILLER_61_382 ();
 sg13g2_fill_1 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_397 ();
 sg13g2_fill_2 FILLER_61_411 ();
 sg13g2_fill_1 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_fill_2 FILLER_62_42 ();
 sg13g2_fill_2 FILLER_62_114 ();
 sg13g2_fill_2 FILLER_62_120 ();
 sg13g2_fill_1 FILLER_62_122 ();
 sg13g2_fill_1 FILLER_62_132 ();
 sg13g2_fill_1 FILLER_62_148 ();
 sg13g2_fill_1 FILLER_62_162 ();
 sg13g2_fill_1 FILLER_62_172 ();
 sg13g2_fill_1 FILLER_62_197 ();
 sg13g2_fill_2 FILLER_62_206 ();
 sg13g2_fill_1 FILLER_62_214 ();
 sg13g2_fill_2 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_264 ();
 sg13g2_fill_2 FILLER_62_273 ();
 sg13g2_fill_2 FILLER_62_300 ();
 sg13g2_fill_1 FILLER_62_324 ();
 sg13g2_fill_1 FILLER_62_356 ();
 sg13g2_fill_1 FILLER_62_362 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_2 FILLER_62_377 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_2 FILLER_62_423 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_fill_2 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_fill_1 FILLER_63_162 ();
 sg13g2_fill_2 FILLER_63_171 ();
 sg13g2_fill_1 FILLER_63_173 ();
 sg13g2_fill_1 FILLER_63_203 ();
 sg13g2_fill_2 FILLER_63_223 ();
 sg13g2_fill_1 FILLER_63_260 ();
 sg13g2_fill_1 FILLER_63_271 ();
 sg13g2_fill_2 FILLER_63_362 ();
 sg13g2_fill_2 FILLER_63_373 ();
 sg13g2_fill_1 FILLER_63_380 ();
 sg13g2_fill_2 FILLER_63_423 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_fill_2 FILLER_64_42 ();
 sg13g2_fill_1 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_88 ();
 sg13g2_fill_1 FILLER_64_172 ();
 sg13g2_fill_2 FILLER_64_178 ();
 sg13g2_fill_1 FILLER_64_186 ();
 sg13g2_fill_1 FILLER_64_191 ();
 sg13g2_fill_2 FILLER_64_210 ();
 sg13g2_fill_1 FILLER_64_212 ();
 sg13g2_fill_2 FILLER_64_228 ();
 sg13g2_fill_1 FILLER_64_245 ();
 sg13g2_fill_1 FILLER_64_251 ();
 sg13g2_fill_1 FILLER_64_262 ();
 sg13g2_fill_1 FILLER_64_274 ();
 sg13g2_fill_1 FILLER_64_296 ();
 sg13g2_fill_2 FILLER_64_309 ();
 sg13g2_fill_1 FILLER_64_344 ();
 sg13g2_fill_2 FILLER_64_350 ();
 sg13g2_fill_1 FILLER_64_352 ();
 sg13g2_fill_2 FILLER_64_363 ();
 sg13g2_fill_2 FILLER_64_413 ();
 sg13g2_fill_2 FILLER_64_427 ();
 sg13g2_fill_1 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_fill_2 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_44 ();
 sg13g2_fill_1 FILLER_65_64 ();
 sg13g2_fill_1 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_169 ();
 sg13g2_fill_1 FILLER_65_184 ();
 sg13g2_fill_2 FILLER_65_189 ();
 sg13g2_fill_1 FILLER_65_191 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_1 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_276 ();
 sg13g2_fill_2 FILLER_65_318 ();
 sg13g2_fill_1 FILLER_65_320 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_373 ();
 sg13g2_fill_1 FILLER_65_379 ();
 sg13g2_fill_2 FILLER_65_421 ();
 sg13g2_fill_2 FILLER_65_427 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_4 FILLER_66_42 ();
 sg13g2_fill_1 FILLER_66_58 ();
 sg13g2_fill_2 FILLER_66_64 ();
 sg13g2_fill_1 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_158 ();
 sg13g2_fill_2 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_211 ();
 sg13g2_fill_1 FILLER_66_218 ();
 sg13g2_fill_2 FILLER_66_228 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_1 FILLER_66_346 ();
 sg13g2_fill_2 FILLER_66_356 ();
 sg13g2_decap_4 FILLER_66_363 ();
 sg13g2_fill_1 FILLER_66_367 ();
 sg13g2_fill_1 FILLER_66_392 ();
 sg13g2_fill_2 FILLER_66_416 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_2 FILLER_67_71 ();
 sg13g2_fill_1 FILLER_67_73 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_1 FILLER_67_100 ();
 sg13g2_fill_2 FILLER_67_111 ();
 sg13g2_fill_1 FILLER_67_122 ();
 sg13g2_fill_2 FILLER_67_153 ();
 sg13g2_fill_1 FILLER_67_155 ();
 sg13g2_fill_1 FILLER_67_165 ();
 sg13g2_fill_1 FILLER_67_183 ();
 sg13g2_fill_1 FILLER_67_194 ();
 sg13g2_fill_1 FILLER_67_203 ();
 sg13g2_fill_2 FILLER_67_234 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_273 ();
 sg13g2_fill_2 FILLER_67_283 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_fill_1 FILLER_67_347 ();
 sg13g2_fill_2 FILLER_67_367 ();
 sg13g2_fill_2 FILLER_67_375 ();
 sg13g2_fill_1 FILLER_67_404 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_4 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_60 ();
 sg13g2_decap_4 FILLER_68_69 ();
 sg13g2_fill_2 FILLER_68_107 ();
 sg13g2_fill_1 FILLER_68_124 ();
 sg13g2_fill_2 FILLER_68_134 ();
 sg13g2_fill_1 FILLER_68_150 ();
 sg13g2_fill_1 FILLER_68_217 ();
 sg13g2_fill_1 FILLER_68_255 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_302 ();
 sg13g2_fill_1 FILLER_68_304 ();
 sg13g2_fill_1 FILLER_68_345 ();
 sg13g2_fill_2 FILLER_68_350 ();
 sg13g2_fill_1 FILLER_68_352 ();
 sg13g2_decap_4 FILLER_68_362 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_2 FILLER_68_385 ();
 sg13g2_fill_2 FILLER_68_414 ();
 sg13g2_decap_4 FILLER_68_419 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_77 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_fill_1 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_129 ();
 sg13g2_fill_2 FILLER_69_170 ();
 sg13g2_fill_1 FILLER_69_184 ();
 sg13g2_fill_1 FILLER_69_202 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_375 ();
 sg13g2_decap_4 FILLER_69_386 ();
 sg13g2_fill_1 FILLER_69_390 ();
 sg13g2_fill_2 FILLER_69_396 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_86 ();
 sg13g2_fill_2 FILLER_70_96 ();
 sg13g2_fill_2 FILLER_70_102 ();
 sg13g2_fill_1 FILLER_70_109 ();
 sg13g2_fill_1 FILLER_70_127 ();
 sg13g2_fill_2 FILLER_70_137 ();
 sg13g2_fill_2 FILLER_70_190 ();
 sg13g2_fill_1 FILLER_70_205 ();
 sg13g2_fill_1 FILLER_70_211 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_fill_1 FILLER_70_222 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_261 ();
 sg13g2_fill_1 FILLER_70_300 ();
 sg13g2_fill_2 FILLER_70_317 ();
 sg13g2_fill_1 FILLER_70_325 ();
 sg13g2_fill_1 FILLER_70_331 ();
 sg13g2_fill_1 FILLER_70_336 ();
 sg13g2_fill_1 FILLER_70_342 ();
 sg13g2_fill_1 FILLER_70_349 ();
 sg13g2_fill_1 FILLER_70_354 ();
 sg13g2_decap_4 FILLER_70_360 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_fill_1 FILLER_70_396 ();
 sg13g2_fill_2 FILLER_70_405 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_fill_2 FILLER_71_91 ();
 sg13g2_fill_1 FILLER_71_149 ();
 sg13g2_fill_2 FILLER_71_176 ();
 sg13g2_fill_1 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_187 ();
 sg13g2_fill_1 FILLER_71_212 ();
 sg13g2_decap_4 FILLER_71_244 ();
 sg13g2_fill_1 FILLER_71_248 ();
 sg13g2_fill_1 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_294 ();
 sg13g2_fill_1 FILLER_71_303 ();
 sg13g2_fill_1 FILLER_71_308 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_2 FILLER_71_368 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_380 ();
 sg13g2_fill_2 FILLER_71_396 ();
 sg13g2_fill_1 FILLER_71_398 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_fill_2 FILLER_72_98 ();
 sg13g2_fill_1 FILLER_72_100 ();
 sg13g2_fill_2 FILLER_72_194 ();
 sg13g2_fill_1 FILLER_72_204 ();
 sg13g2_fill_1 FILLER_72_246 ();
 sg13g2_fill_1 FILLER_72_257 ();
 sg13g2_fill_1 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_288 ();
 sg13g2_fill_1 FILLER_72_290 ();
 sg13g2_fill_2 FILLER_72_296 ();
 sg13g2_fill_1 FILLER_72_355 ();
 sg13g2_fill_1 FILLER_72_360 ();
 sg13g2_fill_2 FILLER_72_365 ();
 sg13g2_fill_1 FILLER_72_367 ();
 sg13g2_fill_1 FILLER_72_385 ();
 sg13g2_decap_4 FILLER_72_426 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_4 FILLER_73_105 ();
 sg13g2_fill_1 FILLER_73_123 ();
 sg13g2_fill_2 FILLER_73_179 ();
 sg13g2_fill_1 FILLER_73_181 ();
 sg13g2_fill_1 FILLER_73_186 ();
 sg13g2_fill_2 FILLER_73_207 ();
 sg13g2_fill_1 FILLER_73_213 ();
 sg13g2_fill_1 FILLER_73_218 ();
 sg13g2_fill_2 FILLER_73_240 ();
 sg13g2_fill_1 FILLER_73_242 ();
 sg13g2_fill_1 FILLER_73_248 ();
 sg13g2_fill_1 FILLER_73_290 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_1 FILLER_73_301 ();
 sg13g2_fill_1 FILLER_73_313 ();
 sg13g2_fill_1 FILLER_73_319 ();
 sg13g2_decap_4 FILLER_73_358 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_368 ();
 sg13g2_fill_2 FILLER_73_395 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_2 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_211 ();
 sg13g2_fill_1 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_243 ();
 sg13g2_fill_1 FILLER_74_250 ();
 sg13g2_fill_2 FILLER_74_262 ();
 sg13g2_fill_1 FILLER_74_269 ();
 sg13g2_fill_1 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_285 ();
 sg13g2_fill_1 FILLER_74_292 ();
 sg13g2_fill_1 FILLER_74_305 ();
 sg13g2_fill_2 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_354 ();
 sg13g2_fill_1 FILLER_74_356 ();
 sg13g2_fill_1 FILLER_74_379 ();
 sg13g2_fill_1 FILLER_74_390 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_fill_1 FILLER_75_112 ();
 sg13g2_decap_4 FILLER_75_134 ();
 sg13g2_fill_1 FILLER_75_141 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_1 FILLER_75_206 ();
 sg13g2_fill_1 FILLER_75_211 ();
 sg13g2_fill_1 FILLER_75_221 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_2 FILLER_75_245 ();
 sg13g2_fill_1 FILLER_75_247 ();
 sg13g2_fill_1 FILLER_75_260 ();
 sg13g2_fill_1 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_278 ();
 sg13g2_fill_1 FILLER_75_340 ();
 sg13g2_fill_2 FILLER_75_388 ();
 sg13g2_fill_1 FILLER_75_409 ();
 sg13g2_decap_4 FILLER_75_426 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_4 FILLER_76_119 ();
 sg13g2_fill_1 FILLER_76_123 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_167 ();
 sg13g2_fill_1 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_208 ();
 sg13g2_fill_1 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_267 ();
 sg13g2_fill_2 FILLER_76_273 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_fill_2 FILLER_76_287 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_fill_2 FILLER_76_352 ();
 sg13g2_fill_1 FILLER_76_362 ();
 sg13g2_fill_1 FILLER_76_368 ();
 sg13g2_fill_1 FILLER_76_399 ();
 sg13g2_fill_2 FILLER_76_419 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_4 FILLER_77_126 ();
 sg13g2_fill_2 FILLER_77_219 ();
 sg13g2_decap_4 FILLER_77_240 ();
 sg13g2_fill_1 FILLER_77_249 ();
 sg13g2_fill_2 FILLER_77_270 ();
 sg13g2_fill_1 FILLER_77_277 ();
 sg13g2_fill_1 FILLER_77_301 ();
 sg13g2_fill_2 FILLER_77_317 ();
 sg13g2_fill_2 FILLER_77_334 ();
 sg13g2_fill_1 FILLER_77_341 ();
 sg13g2_fill_1 FILLER_77_355 ();
 sg13g2_fill_1 FILLER_77_385 ();
 sg13g2_fill_1 FILLER_77_410 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_fill_2 FILLER_78_147 ();
 sg13g2_fill_1 FILLER_78_149 ();
 sg13g2_fill_1 FILLER_78_180 ();
 sg13g2_fill_1 FILLER_78_185 ();
 sg13g2_fill_1 FILLER_78_190 ();
 sg13g2_fill_2 FILLER_78_195 ();
 sg13g2_fill_1 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_207 ();
 sg13g2_fill_1 FILLER_78_213 ();
 sg13g2_fill_1 FILLER_78_218 ();
 sg13g2_fill_2 FILLER_78_223 ();
 sg13g2_fill_1 FILLER_78_229 ();
 sg13g2_fill_1 FILLER_78_235 ();
 sg13g2_fill_1 FILLER_78_269 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_fill_1 FILLER_78_311 ();
 sg13g2_fill_2 FILLER_78_339 ();
 sg13g2_fill_2 FILLER_78_366 ();
 sg13g2_fill_1 FILLER_78_368 ();
 sg13g2_fill_2 FILLER_78_377 ();
 sg13g2_fill_2 FILLER_78_393 ();
 sg13g2_fill_1 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_fill_2 FILLER_79_147 ();
 sg13g2_fill_1 FILLER_79_169 ();
 sg13g2_fill_1 FILLER_79_174 ();
 sg13g2_fill_1 FILLER_79_205 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_217 ();
 sg13g2_fill_1 FILLER_79_223 ();
 sg13g2_fill_1 FILLER_79_229 ();
 sg13g2_fill_1 FILLER_79_254 ();
 sg13g2_fill_1 FILLER_79_285 ();
 sg13g2_fill_2 FILLER_79_291 ();
 sg13g2_fill_1 FILLER_79_314 ();
 sg13g2_fill_1 FILLER_79_324 ();
 sg13g2_fill_2 FILLER_79_370 ();
 sg13g2_fill_1 FILLER_79_372 ();
 sg13g2_fill_2 FILLER_79_378 ();
 sg13g2_fill_1 FILLER_79_380 ();
 sg13g2_fill_2 FILLER_79_402 ();
 sg13g2_decap_4 FILLER_79_415 ();
 sg13g2_fill_1 FILLER_79_419 ();
 sg13g2_decap_4 FILLER_79_425 ();
 sg13g2_fill_1 FILLER_79_429 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_1 FILLER_80_210 ();
 sg13g2_fill_1 FILLER_80_224 ();
 sg13g2_fill_2 FILLER_80_250 ();
 sg13g2_fill_1 FILLER_80_272 ();
 sg13g2_fill_1 FILLER_80_278 ();
 sg13g2_fill_1 FILLER_80_307 ();
 sg13g2_fill_1 FILLER_80_317 ();
 sg13g2_fill_1 FILLER_80_332 ();
 sg13g2_fill_2 FILLER_80_384 ();
 sg13g2_fill_1 FILLER_80_386 ();
 sg13g2_fill_2 FILLER_80_395 ();
 sg13g2_fill_1 FILLER_80_397 ();
 sg13g2_fill_1 FILLER_80_429 ();
endmodule
